module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 ;
  wire n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 ;
  assign n130 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n131 = ( ~x0 & x1 ) | ( ~x0 & n130 ) | ( x1 & n130 ) ;
  assign n132 = ( ~x2 & n130 ) | ( ~x2 & n131 ) | ( n130 & n131 ) ;
  assign n133 = ( x0 & x1 ) | ( x0 & x2 ) | ( x1 & x2 ) ;
  assign n134 = ( x3 & ~x4 ) | ( x3 & n133 ) | ( ~x4 & n133 ) ;
  assign n135 = ( ~x3 & x4 ) | ( ~x3 & n134 ) | ( x4 & n134 ) ;
  assign n136 = ( ~n133 & n134 ) | ( ~n133 & n135 ) | ( n134 & n135 ) ;
  assign n137 = ( x3 & x4 ) | ( x3 & n133 ) | ( x4 & n133 ) ;
  assign n138 = ( x5 & ~x6 ) | ( x5 & n137 ) | ( ~x6 & n137 ) ;
  assign n139 = ( ~x5 & x6 ) | ( ~x5 & n138 ) | ( x6 & n138 ) ;
  assign n140 = ( ~n137 & n138 ) | ( ~n137 & n139 ) | ( n138 & n139 ) ;
  assign n141 = ( x5 & x6 ) | ( x5 & n137 ) | ( x6 & n137 ) ;
  assign n142 = ( x7 & ~x8 ) | ( x7 & n141 ) | ( ~x8 & n141 ) ;
  assign n143 = ( ~x7 & x8 ) | ( ~x7 & n142 ) | ( x8 & n142 ) ;
  assign n144 = ( ~n141 & n142 ) | ( ~n141 & n143 ) | ( n142 & n143 ) ;
  assign n145 = ( x7 & x8 ) | ( x7 & n141 ) | ( x8 & n141 ) ;
  assign n146 = ( x9 & ~x10 ) | ( x9 & n145 ) | ( ~x10 & n145 ) ;
  assign n147 = ( ~x9 & x10 ) | ( ~x9 & n146 ) | ( x10 & n146 ) ;
  assign n148 = ( ~n145 & n146 ) | ( ~n145 & n147 ) | ( n146 & n147 ) ;
  assign n149 = ( x9 & x10 ) | ( x9 & n145 ) | ( x10 & n145 ) ;
  assign n150 = ( x11 & ~x12 ) | ( x11 & n149 ) | ( ~x12 & n149 ) ;
  assign n151 = ( ~x11 & x12 ) | ( ~x11 & n150 ) | ( x12 & n150 ) ;
  assign n152 = ( ~n149 & n150 ) | ( ~n149 & n151 ) | ( n150 & n151 ) ;
  assign n153 = ( x11 & x12 ) | ( x11 & n149 ) | ( x12 & n149 ) ;
  assign n154 = ( x13 & ~x14 ) | ( x13 & n153 ) | ( ~x14 & n153 ) ;
  assign n155 = ( ~x13 & x14 ) | ( ~x13 & n154 ) | ( x14 & n154 ) ;
  assign n156 = ( ~n153 & n154 ) | ( ~n153 & n155 ) | ( n154 & n155 ) ;
  assign n157 = ( x13 & x14 ) | ( x13 & n153 ) | ( x14 & n153 ) ;
  assign n158 = ( x15 & ~x16 ) | ( x15 & n157 ) | ( ~x16 & n157 ) ;
  assign n159 = ( ~x15 & x16 ) | ( ~x15 & n158 ) | ( x16 & n158 ) ;
  assign n160 = ( ~n157 & n158 ) | ( ~n157 & n159 ) | ( n158 & n159 ) ;
  assign n161 = ( x15 & x16 ) | ( x15 & n157 ) | ( x16 & n157 ) ;
  assign n162 = ( x17 & ~x18 ) | ( x17 & n161 ) | ( ~x18 & n161 ) ;
  assign n163 = ( ~x17 & x18 ) | ( ~x17 & n162 ) | ( x18 & n162 ) ;
  assign n164 = ( ~n161 & n162 ) | ( ~n161 & n163 ) | ( n162 & n163 ) ;
  assign n165 = ( x17 & x18 ) | ( x17 & n161 ) | ( x18 & n161 ) ;
  assign n166 = ( x19 & ~x20 ) | ( x19 & n165 ) | ( ~x20 & n165 ) ;
  assign n167 = ( ~x19 & x20 ) | ( ~x19 & n166 ) | ( x20 & n166 ) ;
  assign n168 = ( ~n165 & n166 ) | ( ~n165 & n167 ) | ( n166 & n167 ) ;
  assign n169 = ( x19 & x20 ) | ( x19 & n165 ) | ( x20 & n165 ) ;
  assign n170 = ( x21 & ~x22 ) | ( x21 & n169 ) | ( ~x22 & n169 ) ;
  assign n171 = ( ~x21 & x22 ) | ( ~x21 & n170 ) | ( x22 & n170 ) ;
  assign n172 = ( ~n169 & n170 ) | ( ~n169 & n171 ) | ( n170 & n171 ) ;
  assign n173 = ( x21 & x22 ) | ( x21 & n169 ) | ( x22 & n169 ) ;
  assign n174 = ( x23 & ~x24 ) | ( x23 & n173 ) | ( ~x24 & n173 ) ;
  assign n175 = ( ~x23 & x24 ) | ( ~x23 & n174 ) | ( x24 & n174 ) ;
  assign n176 = ( ~n173 & n174 ) | ( ~n173 & n175 ) | ( n174 & n175 ) ;
  assign n177 = ( x23 & x24 ) | ( x23 & n173 ) | ( x24 & n173 ) ;
  assign n178 = ( x25 & ~x26 ) | ( x25 & n177 ) | ( ~x26 & n177 ) ;
  assign n179 = ( ~x25 & x26 ) | ( ~x25 & n178 ) | ( x26 & n178 ) ;
  assign n180 = ( ~n177 & n178 ) | ( ~n177 & n179 ) | ( n178 & n179 ) ;
  assign n181 = ( x25 & x26 ) | ( x25 & n177 ) | ( x26 & n177 ) ;
  assign n182 = ( x27 & ~x28 ) | ( x27 & n181 ) | ( ~x28 & n181 ) ;
  assign n183 = ( ~x27 & x28 ) | ( ~x27 & n182 ) | ( x28 & n182 ) ;
  assign n184 = ( ~n181 & n182 ) | ( ~n181 & n183 ) | ( n182 & n183 ) ;
  assign n185 = ( x27 & x28 ) | ( x27 & n181 ) | ( x28 & n181 ) ;
  assign n186 = ( x29 & ~x30 ) | ( x29 & n185 ) | ( ~x30 & n185 ) ;
  assign n187 = ( ~x29 & x30 ) | ( ~x29 & n186 ) | ( x30 & n186 ) ;
  assign n188 = ( ~n185 & n186 ) | ( ~n185 & n187 ) | ( n186 & n187 ) ;
  assign n189 = ( x29 & x30 ) | ( x29 & n185 ) | ( x30 & n185 ) ;
  assign n190 = ( x31 & ~x32 ) | ( x31 & n189 ) | ( ~x32 & n189 ) ;
  assign n191 = ( ~x31 & x32 ) | ( ~x31 & n190 ) | ( x32 & n190 ) ;
  assign n192 = ( ~n189 & n190 ) | ( ~n189 & n191 ) | ( n190 & n191 ) ;
  assign n193 = ( x31 & x32 ) | ( x31 & n189 ) | ( x32 & n189 ) ;
  assign n194 = ( x33 & ~x34 ) | ( x33 & n193 ) | ( ~x34 & n193 ) ;
  assign n195 = ( ~x33 & x34 ) | ( ~x33 & n194 ) | ( x34 & n194 ) ;
  assign n196 = ( ~n193 & n194 ) | ( ~n193 & n195 ) | ( n194 & n195 ) ;
  assign n197 = ( x33 & x34 ) | ( x33 & n193 ) | ( x34 & n193 ) ;
  assign n198 = ( x35 & ~x36 ) | ( x35 & n197 ) | ( ~x36 & n197 ) ;
  assign n199 = ( ~x35 & x36 ) | ( ~x35 & n198 ) | ( x36 & n198 ) ;
  assign n200 = ( ~n197 & n198 ) | ( ~n197 & n199 ) | ( n198 & n199 ) ;
  assign n201 = ( x35 & x36 ) | ( x35 & n197 ) | ( x36 & n197 ) ;
  assign n202 = ( x37 & ~x38 ) | ( x37 & n201 ) | ( ~x38 & n201 ) ;
  assign n203 = ( ~x37 & x38 ) | ( ~x37 & n202 ) | ( x38 & n202 ) ;
  assign n204 = ( ~n201 & n202 ) | ( ~n201 & n203 ) | ( n202 & n203 ) ;
  assign n205 = ( x37 & x38 ) | ( x37 & n201 ) | ( x38 & n201 ) ;
  assign n206 = ( x39 & ~x40 ) | ( x39 & n205 ) | ( ~x40 & n205 ) ;
  assign n207 = ( ~x39 & x40 ) | ( ~x39 & n206 ) | ( x40 & n206 ) ;
  assign n208 = ( ~n205 & n206 ) | ( ~n205 & n207 ) | ( n206 & n207 ) ;
  assign n209 = ( x39 & x40 ) | ( x39 & n205 ) | ( x40 & n205 ) ;
  assign n210 = ( x41 & ~x42 ) | ( x41 & n209 ) | ( ~x42 & n209 ) ;
  assign n211 = ( ~x41 & x42 ) | ( ~x41 & n210 ) | ( x42 & n210 ) ;
  assign n212 = ( ~n209 & n210 ) | ( ~n209 & n211 ) | ( n210 & n211 ) ;
  assign n213 = ( x41 & x42 ) | ( x41 & n209 ) | ( x42 & n209 ) ;
  assign n214 = ( x43 & ~x44 ) | ( x43 & n213 ) | ( ~x44 & n213 ) ;
  assign n215 = ( ~x43 & x44 ) | ( ~x43 & n214 ) | ( x44 & n214 ) ;
  assign n216 = ( ~n213 & n214 ) | ( ~n213 & n215 ) | ( n214 & n215 ) ;
  assign n217 = ( x43 & x44 ) | ( x43 & n213 ) | ( x44 & n213 ) ;
  assign n218 = ( x45 & ~x46 ) | ( x45 & n217 ) | ( ~x46 & n217 ) ;
  assign n219 = ( ~x45 & x46 ) | ( ~x45 & n218 ) | ( x46 & n218 ) ;
  assign n220 = ( ~n217 & n218 ) | ( ~n217 & n219 ) | ( n218 & n219 ) ;
  assign n221 = ( x45 & x46 ) | ( x45 & n217 ) | ( x46 & n217 ) ;
  assign n222 = ( x47 & ~x48 ) | ( x47 & n221 ) | ( ~x48 & n221 ) ;
  assign n223 = ( ~x47 & x48 ) | ( ~x47 & n222 ) | ( x48 & n222 ) ;
  assign n224 = ( ~n221 & n222 ) | ( ~n221 & n223 ) | ( n222 & n223 ) ;
  assign n225 = ( x47 & x48 ) | ( x47 & n221 ) | ( x48 & n221 ) ;
  assign n226 = ( x49 & ~x50 ) | ( x49 & n225 ) | ( ~x50 & n225 ) ;
  assign n227 = ( ~x49 & x50 ) | ( ~x49 & n226 ) | ( x50 & n226 ) ;
  assign n228 = ( ~n225 & n226 ) | ( ~n225 & n227 ) | ( n226 & n227 ) ;
  assign n229 = ( x49 & x50 ) | ( x49 & n225 ) | ( x50 & n225 ) ;
  assign n230 = ( x51 & ~x52 ) | ( x51 & n229 ) | ( ~x52 & n229 ) ;
  assign n231 = ( ~x51 & x52 ) | ( ~x51 & n230 ) | ( x52 & n230 ) ;
  assign n232 = ( ~n229 & n230 ) | ( ~n229 & n231 ) | ( n230 & n231 ) ;
  assign n233 = ( x51 & x52 ) | ( x51 & n229 ) | ( x52 & n229 ) ;
  assign n234 = ( x53 & ~x54 ) | ( x53 & n233 ) | ( ~x54 & n233 ) ;
  assign n235 = ( ~x53 & x54 ) | ( ~x53 & n234 ) | ( x54 & n234 ) ;
  assign n236 = ( ~n233 & n234 ) | ( ~n233 & n235 ) | ( n234 & n235 ) ;
  assign n237 = ( x53 & x54 ) | ( x53 & n233 ) | ( x54 & n233 ) ;
  assign n238 = ( x55 & ~x56 ) | ( x55 & n237 ) | ( ~x56 & n237 ) ;
  assign n239 = ( ~x55 & x56 ) | ( ~x55 & n238 ) | ( x56 & n238 ) ;
  assign n240 = ( ~n237 & n238 ) | ( ~n237 & n239 ) | ( n238 & n239 ) ;
  assign n241 = ( x55 & x56 ) | ( x55 & n237 ) | ( x56 & n237 ) ;
  assign n242 = ( x57 & ~x58 ) | ( x57 & n241 ) | ( ~x58 & n241 ) ;
  assign n243 = ( ~x57 & x58 ) | ( ~x57 & n242 ) | ( x58 & n242 ) ;
  assign n244 = ( ~n241 & n242 ) | ( ~n241 & n243 ) | ( n242 & n243 ) ;
  assign n245 = ( x57 & x58 ) | ( x57 & n241 ) | ( x58 & n241 ) ;
  assign n246 = ( x59 & ~x60 ) | ( x59 & n245 ) | ( ~x60 & n245 ) ;
  assign n247 = ( ~x59 & x60 ) | ( ~x59 & n246 ) | ( x60 & n246 ) ;
  assign n248 = ( ~n245 & n246 ) | ( ~n245 & n247 ) | ( n246 & n247 ) ;
  assign n249 = ( x59 & x60 ) | ( x59 & n245 ) | ( x60 & n245 ) ;
  assign n250 = ( x61 & ~x62 ) | ( x61 & n249 ) | ( ~x62 & n249 ) ;
  assign n251 = ( ~x61 & x62 ) | ( ~x61 & n250 ) | ( x62 & n250 ) ;
  assign n252 = ( ~n249 & n250 ) | ( ~n249 & n251 ) | ( n250 & n251 ) ;
  assign n253 = ( x61 & x62 ) | ( x61 & n249 ) | ( x62 & n249 ) ;
  assign n254 = ( x63 & ~x64 ) | ( x63 & n253 ) | ( ~x64 & n253 ) ;
  assign n255 = ( ~x63 & x64 ) | ( ~x63 & n254 ) | ( x64 & n254 ) ;
  assign n256 = ( ~n253 & n254 ) | ( ~n253 & n255 ) | ( n254 & n255 ) ;
  assign n257 = ( x63 & x64 ) | ( x63 & n253 ) | ( x64 & n253 ) ;
  assign n258 = ( x65 & ~x66 ) | ( x65 & n257 ) | ( ~x66 & n257 ) ;
  assign n259 = ( ~x65 & x66 ) | ( ~x65 & n258 ) | ( x66 & n258 ) ;
  assign n260 = ( ~n257 & n258 ) | ( ~n257 & n259 ) | ( n258 & n259 ) ;
  assign n261 = ( x65 & x66 ) | ( x65 & n257 ) | ( x66 & n257 ) ;
  assign n262 = ( x67 & ~x68 ) | ( x67 & n261 ) | ( ~x68 & n261 ) ;
  assign n263 = ( ~x67 & x68 ) | ( ~x67 & n262 ) | ( x68 & n262 ) ;
  assign n264 = ( ~n261 & n262 ) | ( ~n261 & n263 ) | ( n262 & n263 ) ;
  assign n265 = ( x67 & x68 ) | ( x67 & n261 ) | ( x68 & n261 ) ;
  assign n266 = ( x69 & ~x70 ) | ( x69 & n265 ) | ( ~x70 & n265 ) ;
  assign n267 = ( ~x69 & x70 ) | ( ~x69 & n266 ) | ( x70 & n266 ) ;
  assign n268 = ( ~n265 & n266 ) | ( ~n265 & n267 ) | ( n266 & n267 ) ;
  assign n269 = ( x69 & x70 ) | ( x69 & n265 ) | ( x70 & n265 ) ;
  assign n270 = ( x71 & ~x72 ) | ( x71 & n269 ) | ( ~x72 & n269 ) ;
  assign n271 = ( ~x71 & x72 ) | ( ~x71 & n270 ) | ( x72 & n270 ) ;
  assign n272 = ( ~n269 & n270 ) | ( ~n269 & n271 ) | ( n270 & n271 ) ;
  assign n273 = ( x71 & x72 ) | ( x71 & n269 ) | ( x72 & n269 ) ;
  assign n274 = ( x73 & ~x74 ) | ( x73 & n273 ) | ( ~x74 & n273 ) ;
  assign n275 = ( ~x73 & x74 ) | ( ~x73 & n274 ) | ( x74 & n274 ) ;
  assign n276 = ( ~n273 & n274 ) | ( ~n273 & n275 ) | ( n274 & n275 ) ;
  assign n277 = ( x73 & x74 ) | ( x73 & n273 ) | ( x74 & n273 ) ;
  assign n278 = ( x75 & ~x76 ) | ( x75 & n277 ) | ( ~x76 & n277 ) ;
  assign n279 = ( ~x75 & x76 ) | ( ~x75 & n278 ) | ( x76 & n278 ) ;
  assign n280 = ( ~n277 & n278 ) | ( ~n277 & n279 ) | ( n278 & n279 ) ;
  assign n281 = ( x75 & x76 ) | ( x75 & n277 ) | ( x76 & n277 ) ;
  assign n282 = ( x77 & ~x78 ) | ( x77 & n281 ) | ( ~x78 & n281 ) ;
  assign n283 = ( ~x77 & x78 ) | ( ~x77 & n282 ) | ( x78 & n282 ) ;
  assign n284 = ( ~n281 & n282 ) | ( ~n281 & n283 ) | ( n282 & n283 ) ;
  assign n285 = ( x77 & x78 ) | ( x77 & n281 ) | ( x78 & n281 ) ;
  assign n286 = ( x79 & ~x80 ) | ( x79 & n285 ) | ( ~x80 & n285 ) ;
  assign n287 = ( ~x79 & x80 ) | ( ~x79 & n286 ) | ( x80 & n286 ) ;
  assign n288 = ( ~n285 & n286 ) | ( ~n285 & n287 ) | ( n286 & n287 ) ;
  assign n289 = ( x79 & x80 ) | ( x79 & n285 ) | ( x80 & n285 ) ;
  assign n290 = ( x81 & ~x82 ) | ( x81 & n289 ) | ( ~x82 & n289 ) ;
  assign n291 = ( ~x81 & x82 ) | ( ~x81 & n290 ) | ( x82 & n290 ) ;
  assign n292 = ( ~n289 & n290 ) | ( ~n289 & n291 ) | ( n290 & n291 ) ;
  assign n293 = ( x81 & x82 ) | ( x81 & n289 ) | ( x82 & n289 ) ;
  assign n294 = ( x83 & ~x84 ) | ( x83 & n293 ) | ( ~x84 & n293 ) ;
  assign n295 = ( ~x83 & x84 ) | ( ~x83 & n294 ) | ( x84 & n294 ) ;
  assign n296 = ( ~n293 & n294 ) | ( ~n293 & n295 ) | ( n294 & n295 ) ;
  assign n297 = ( x83 & x84 ) | ( x83 & n293 ) | ( x84 & n293 ) ;
  assign n298 = ( x85 & ~x86 ) | ( x85 & n297 ) | ( ~x86 & n297 ) ;
  assign n299 = ( ~x85 & x86 ) | ( ~x85 & n298 ) | ( x86 & n298 ) ;
  assign n300 = ( ~n297 & n298 ) | ( ~n297 & n299 ) | ( n298 & n299 ) ;
  assign n301 = ( x85 & x86 ) | ( x85 & n297 ) | ( x86 & n297 ) ;
  assign n302 = ( x87 & ~x88 ) | ( x87 & n301 ) | ( ~x88 & n301 ) ;
  assign n303 = ( ~x87 & x88 ) | ( ~x87 & n302 ) | ( x88 & n302 ) ;
  assign n304 = ( ~n301 & n302 ) | ( ~n301 & n303 ) | ( n302 & n303 ) ;
  assign n305 = ( x87 & x88 ) | ( x87 & n301 ) | ( x88 & n301 ) ;
  assign n306 = ( x89 & ~x90 ) | ( x89 & n305 ) | ( ~x90 & n305 ) ;
  assign n307 = ( ~x89 & x90 ) | ( ~x89 & n306 ) | ( x90 & n306 ) ;
  assign n308 = ( ~n305 & n306 ) | ( ~n305 & n307 ) | ( n306 & n307 ) ;
  assign n309 = ( x89 & x90 ) | ( x89 & n305 ) | ( x90 & n305 ) ;
  assign n310 = ( x91 & ~x92 ) | ( x91 & n309 ) | ( ~x92 & n309 ) ;
  assign n311 = ( ~x91 & x92 ) | ( ~x91 & n310 ) | ( x92 & n310 ) ;
  assign n312 = ( ~n309 & n310 ) | ( ~n309 & n311 ) | ( n310 & n311 ) ;
  assign n313 = ( x91 & x92 ) | ( x91 & n309 ) | ( x92 & n309 ) ;
  assign n314 = ( x93 & ~x94 ) | ( x93 & n313 ) | ( ~x94 & n313 ) ;
  assign n315 = ( ~x93 & x94 ) | ( ~x93 & n314 ) | ( x94 & n314 ) ;
  assign n316 = ( ~n313 & n314 ) | ( ~n313 & n315 ) | ( n314 & n315 ) ;
  assign n317 = ( x93 & x94 ) | ( x93 & n313 ) | ( x94 & n313 ) ;
  assign n318 = ( x95 & ~x96 ) | ( x95 & n317 ) | ( ~x96 & n317 ) ;
  assign n319 = ( ~x95 & x96 ) | ( ~x95 & n318 ) | ( x96 & n318 ) ;
  assign n320 = ( ~n317 & n318 ) | ( ~n317 & n319 ) | ( n318 & n319 ) ;
  assign n321 = ( x95 & x96 ) | ( x95 & n317 ) | ( x96 & n317 ) ;
  assign n322 = ( x97 & ~x98 ) | ( x97 & n321 ) | ( ~x98 & n321 ) ;
  assign n323 = ( ~x97 & x98 ) | ( ~x97 & n322 ) | ( x98 & n322 ) ;
  assign n324 = ( ~n321 & n322 ) | ( ~n321 & n323 ) | ( n322 & n323 ) ;
  assign n325 = ( x97 & x98 ) | ( x97 & n321 ) | ( x98 & n321 ) ;
  assign n326 = ( x99 & ~x100 ) | ( x99 & n325 ) | ( ~x100 & n325 ) ;
  assign n327 = ( ~x99 & x100 ) | ( ~x99 & n326 ) | ( x100 & n326 ) ;
  assign n328 = ( ~n325 & n326 ) | ( ~n325 & n327 ) | ( n326 & n327 ) ;
  assign n329 = ( x99 & x100 ) | ( x99 & n325 ) | ( x100 & n325 ) ;
  assign n330 = ( x101 & ~x102 ) | ( x101 & n329 ) | ( ~x102 & n329 ) ;
  assign n331 = ( ~x101 & x102 ) | ( ~x101 & n330 ) | ( x102 & n330 ) ;
  assign n332 = ( ~n329 & n330 ) | ( ~n329 & n331 ) | ( n330 & n331 ) ;
  assign n333 = ( x101 & x102 ) | ( x101 & n329 ) | ( x102 & n329 ) ;
  assign n334 = ( x103 & ~x104 ) | ( x103 & n333 ) | ( ~x104 & n333 ) ;
  assign n335 = ( ~x103 & x104 ) | ( ~x103 & n334 ) | ( x104 & n334 ) ;
  assign n336 = ( ~n333 & n334 ) | ( ~n333 & n335 ) | ( n334 & n335 ) ;
  assign n337 = ( x103 & x104 ) | ( x103 & n333 ) | ( x104 & n333 ) ;
  assign n338 = ( x105 & ~x106 ) | ( x105 & n337 ) | ( ~x106 & n337 ) ;
  assign n339 = ( ~x105 & x106 ) | ( ~x105 & n338 ) | ( x106 & n338 ) ;
  assign n340 = ( ~n337 & n338 ) | ( ~n337 & n339 ) | ( n338 & n339 ) ;
  assign n341 = ( x105 & x106 ) | ( x105 & n337 ) | ( x106 & n337 ) ;
  assign n342 = ( x107 & ~x108 ) | ( x107 & n341 ) | ( ~x108 & n341 ) ;
  assign n343 = ( ~x107 & x108 ) | ( ~x107 & n342 ) | ( x108 & n342 ) ;
  assign n344 = ( ~n341 & n342 ) | ( ~n341 & n343 ) | ( n342 & n343 ) ;
  assign n345 = ( x107 & x108 ) | ( x107 & n341 ) | ( x108 & n341 ) ;
  assign n346 = ( x109 & ~x110 ) | ( x109 & n345 ) | ( ~x110 & n345 ) ;
  assign n347 = ( ~x109 & x110 ) | ( ~x109 & n346 ) | ( x110 & n346 ) ;
  assign n348 = ( ~n345 & n346 ) | ( ~n345 & n347 ) | ( n346 & n347 ) ;
  assign n349 = ( x109 & x110 ) | ( x109 & n345 ) | ( x110 & n345 ) ;
  assign n350 = ( x111 & ~x112 ) | ( x111 & n349 ) | ( ~x112 & n349 ) ;
  assign n351 = ( ~x111 & x112 ) | ( ~x111 & n350 ) | ( x112 & n350 ) ;
  assign n352 = ( ~n349 & n350 ) | ( ~n349 & n351 ) | ( n350 & n351 ) ;
  assign n353 = ( x111 & x112 ) | ( x111 & n349 ) | ( x112 & n349 ) ;
  assign n354 = ( x113 & ~x114 ) | ( x113 & n353 ) | ( ~x114 & n353 ) ;
  assign n355 = ( ~x113 & x114 ) | ( ~x113 & n354 ) | ( x114 & n354 ) ;
  assign n356 = ( ~n353 & n354 ) | ( ~n353 & n355 ) | ( n354 & n355 ) ;
  assign n357 = ( x113 & x114 ) | ( x113 & n353 ) | ( x114 & n353 ) ;
  assign n358 = ( x115 & ~x116 ) | ( x115 & n357 ) | ( ~x116 & n357 ) ;
  assign n359 = ( ~x115 & x116 ) | ( ~x115 & n358 ) | ( x116 & n358 ) ;
  assign n360 = ( ~n357 & n358 ) | ( ~n357 & n359 ) | ( n358 & n359 ) ;
  assign n361 = ( x115 & x116 ) | ( x115 & n357 ) | ( x116 & n357 ) ;
  assign n362 = ( x117 & ~x118 ) | ( x117 & n361 ) | ( ~x118 & n361 ) ;
  assign n363 = ( ~x117 & x118 ) | ( ~x117 & n362 ) | ( x118 & n362 ) ;
  assign n364 = ( ~n361 & n362 ) | ( ~n361 & n363 ) | ( n362 & n363 ) ;
  assign n365 = ( x117 & x118 ) | ( x117 & n361 ) | ( x118 & n361 ) ;
  assign n366 = ( x119 & ~x120 ) | ( x119 & n365 ) | ( ~x120 & n365 ) ;
  assign n367 = ( ~x119 & x120 ) | ( ~x119 & n366 ) | ( x120 & n366 ) ;
  assign n368 = ( ~n365 & n366 ) | ( ~n365 & n367 ) | ( n366 & n367 ) ;
  assign n369 = ( x119 & x120 ) | ( x119 & n365 ) | ( x120 & n365 ) ;
  assign n370 = ( x121 & ~x122 ) | ( x121 & n369 ) | ( ~x122 & n369 ) ;
  assign n371 = ( ~x121 & x122 ) | ( ~x121 & n370 ) | ( x122 & n370 ) ;
  assign n372 = ( ~n369 & n370 ) | ( ~n369 & n371 ) | ( n370 & n371 ) ;
  assign n373 = ( x121 & x122 ) | ( x121 & n369 ) | ( x122 & n369 ) ;
  assign n374 = ( x123 & ~x124 ) | ( x123 & n373 ) | ( ~x124 & n373 ) ;
  assign n375 = ( ~x123 & x124 ) | ( ~x123 & n374 ) | ( x124 & n374 ) ;
  assign n376 = ( ~n373 & n374 ) | ( ~n373 & n375 ) | ( n374 & n375 ) ;
  assign n377 = ( x123 & x124 ) | ( x123 & n373 ) | ( x124 & n373 ) ;
  assign n378 = ( x125 & ~x126 ) | ( x125 & n377 ) | ( ~x126 & n377 ) ;
  assign n379 = ( ~x125 & x126 ) | ( ~x125 & n378 ) | ( x126 & n378 ) ;
  assign n380 = ( ~n377 & n378 ) | ( ~n377 & n379 ) | ( n378 & n379 ) ;
  assign n381 = ( x125 & x126 ) | ( x125 & n377 ) | ( x126 & n377 ) ;
  assign n382 = ( x127 & ~x128 ) | ( x127 & n381 ) | ( ~x128 & n381 ) ;
  assign n383 = ( ~x127 & x128 ) | ( ~x127 & n382 ) | ( x128 & n382 ) ;
  assign n384 = ( ~n381 & n382 ) | ( ~n381 & n383 ) | ( n382 & n383 ) ;
  assign n385 = ( x127 & x128 ) | ( x127 & n381 ) | ( x128 & n381 ) ;
  assign y0 = n132 ;
  assign y1 = n136 ;
  assign y2 = n140 ;
  assign y3 = n144 ;
  assign y4 = n148 ;
  assign y5 = n152 ;
  assign y6 = n156 ;
  assign y7 = n160 ;
  assign y8 = n164 ;
  assign y9 = n168 ;
  assign y10 = n172 ;
  assign y11 = n176 ;
  assign y12 = n180 ;
  assign y13 = n184 ;
  assign y14 = n188 ;
  assign y15 = n192 ;
  assign y16 = n196 ;
  assign y17 = n200 ;
  assign y18 = n204 ;
  assign y19 = n208 ;
  assign y20 = n212 ;
  assign y21 = n216 ;
  assign y22 = n220 ;
  assign y23 = n224 ;
  assign y24 = n228 ;
  assign y25 = n232 ;
  assign y26 = n236 ;
  assign y27 = n240 ;
  assign y28 = n244 ;
  assign y29 = n248 ;
  assign y30 = n252 ;
  assign y31 = n256 ;
  assign y32 = n260 ;
  assign y33 = n264 ;
  assign y34 = n268 ;
  assign y35 = n272 ;
  assign y36 = n276 ;
  assign y37 = n280 ;
  assign y38 = n284 ;
  assign y39 = n288 ;
  assign y40 = n292 ;
  assign y41 = n296 ;
  assign y42 = n300 ;
  assign y43 = n304 ;
  assign y44 = n308 ;
  assign y45 = n312 ;
  assign y46 = n316 ;
  assign y47 = n320 ;
  assign y48 = n324 ;
  assign y49 = n328 ;
  assign y50 = n332 ;
  assign y51 = n336 ;
  assign y52 = n340 ;
  assign y53 = n344 ;
  assign y54 = n348 ;
  assign y55 = n352 ;
  assign y56 = n356 ;
  assign y57 = n360 ;
  assign y58 = n364 ;
  assign y59 = n368 ;
  assign y60 = n372 ;
  assign y61 = n376 ;
  assign y62 = n380 ;
  assign y63 = n384 ;
  assign y64 = n385 ;
endmodule
