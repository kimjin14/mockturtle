module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 ;
  wire n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 ;
  assign n148 = x13 | x14 ;
  assign n149 = x6 | x7 ;
  assign n150 = n148 | n149 ;
  assign n151 = x17 | x21 ;
  assign n152 = x8 | x12 ;
  assign n153 = n151 | n152 ;
  assign n154 = n150 | n153 ;
  assign n155 = x18 | x19 ;
  assign n156 = x4 | x16 ;
  assign n157 = n155 | n156 ;
  assign n158 = x5 | x22 ;
  assign n159 = x9 | x11 ;
  assign n160 = n158 | n159 ;
  assign n161 = n157 | n160 ;
  assign n162 = n154 | n161 ;
  assign n163 = x0 | x54 ;
  assign n164 = ( x0 & n162 ) | ( x0 & n163 ) | ( n162 & n163 ) ;
  assign n165 = ~x54 & n164 ;
  assign n166 = ~x56 & n158 ;
  assign n167 = x6 | x12 ;
  assign n168 = x17 | n157 ;
  assign n169 = n167 | n168 ;
  assign n170 = x8 | x21 ;
  assign n171 = x7 | n170 ;
  assign n172 = x10 & ~n148 ;
  assign n173 = ~n171 & n172 ;
  assign n174 = ~x13 & x14 ;
  assign n175 = ~n171 & n174 ;
  assign n176 = x14 & ~n175 ;
  assign n177 = x8 & x21 ;
  assign n178 = ( x7 & n170 ) | ( x7 & ~n177 ) | ( n170 & ~n177 ) ;
  assign n179 = ( x7 & x13 ) | ( x7 & n170 ) | ( x13 & n170 ) ;
  assign n180 = x13 & ~n178 ;
  assign n181 = ( n178 & ~n179 ) | ( n178 & n180 ) | ( ~n179 & n180 ) ;
  assign n182 = ( n175 & ~n176 ) | ( n175 & n181 ) | ( ~n176 & n181 ) ;
  assign n183 = ~x10 & n182 ;
  assign n184 = ( ~n158 & n173 ) | ( ~n158 & n183 ) | ( n173 & n183 ) ;
  assign n185 = ~n169 & n184 ;
  assign n186 = ( ~n159 & n166 ) | ( ~n159 & n185 ) | ( n166 & n185 ) ;
  assign n187 = ~n158 & n159 ;
  assign n188 = ( n164 & n165 ) | ( n164 & ~n187 ) | ( n165 & ~n187 ) ;
  assign n189 = ( x56 & n164 ) | ( x56 & n188 ) | ( n164 & n188 ) ;
  assign n190 = ( n165 & ~n186 ) | ( n165 & n189 ) | ( ~n186 & n189 ) ;
  assign n191 = x129 | n190 ;
  assign n192 = x3 | n191 ;
  assign n193 = x11 | x12 ;
  assign n194 = n170 | n193 ;
  assign n195 = n157 | n194 ;
  assign n196 = x7 | x13 ;
  assign n197 = x5 | x6 ;
  assign n198 = n196 | n197 ;
  assign n199 = x10 | x22 ;
  assign n200 = n148 | n199 ;
  assign n201 = ( ~x13 & n198 ) | ( ~x13 & n200 ) | ( n198 & n200 ) ;
  assign n202 = n195 | n201 ;
  assign n203 = ~x17 & x54 ;
  assign n204 = n202 & n203 ;
  assign n205 = x1 | n204 ;
  assign n206 = ~x14 & x54 ;
  assign n207 = x8 | x11 ;
  assign n208 = n151 | n207 ;
  assign n209 = x6 & x12 ;
  assign n210 = ( x5 & n167 ) | ( x5 & ~n209 ) | ( n167 & ~n209 ) ;
  assign n211 = ( x5 & x7 ) | ( x5 & n167 ) | ( x7 & n167 ) ;
  assign n212 = x7 & ~n210 ;
  assign n213 = ( n210 & ~n211 ) | ( n210 & n212 ) | ( ~n211 & n212 ) ;
  assign n214 = ~x13 & n213 ;
  assign n215 = ~x7 & x13 ;
  assign n216 = x5 | n167 ;
  assign n217 = n215 & ~n216 ;
  assign n218 = n214 | n217 ;
  assign n219 = ( x9 & ~n157 ) | ( x9 & n218 ) | ( ~n157 & n218 ) ;
  assign n220 = n196 | n216 ;
  assign n221 = ( x9 & n157 ) | ( x9 & n220 ) | ( n157 & n220 ) ;
  assign n222 = n219 & ~n221 ;
  assign n223 = ~n208 & n222 ;
  assign n224 = n206 & n223 ;
  assign n225 = ~n199 & n224 ;
  assign n226 = n205 & ~n225 ;
  assign n227 = x129 | n226 ;
  assign n228 = x3 | n227 ;
  assign n229 = x122 & x127 ;
  assign n230 = x41 | x46 ;
  assign n231 = x38 | x50 ;
  assign n232 = n230 | n231 ;
  assign n233 = x42 | x44 ;
  assign n234 = x40 | n233 ;
  assign n235 = x2 | n234 ;
  assign n236 = n232 | n235 ;
  assign n237 = x15 | x20 ;
  assign n238 = x24 | x49 ;
  assign n239 = n237 | n238 ;
  assign n240 = x45 | n238 ;
  assign n241 = x43 | x47 ;
  assign n242 = x48 | n241 ;
  assign n243 = n240 | n242 ;
  assign n244 = n239 | n243 ;
  assign n245 = n236 | n244 ;
  assign n246 = x82 & n245 ;
  assign n247 = n229 | n246 ;
  assign n248 = x65 | n247 ;
  assign n249 = x38 | x40 ;
  assign n250 = n233 | n249 ;
  assign n251 = x46 | x50 ;
  assign n252 = x41 | n251 ;
  assign n253 = n250 | n252 ;
  assign n254 = x43 | n253 ;
  assign n255 = x47 | x48 ;
  assign n256 = x45 | n255 ;
  assign n257 = x24 | x45 ;
  assign n258 = x49 | n237 ;
  assign n259 = n257 | n258 ;
  assign n260 = ( ~x45 & n256 ) | ( ~x45 & n259 ) | ( n256 & n259 ) ;
  assign n261 = n254 | n260 ;
  assign n262 = x82 & n261 ;
  assign n263 = ~x82 & n229 ;
  assign n264 = n262 | n263 ;
  assign n265 = x2 & n264 ;
  assign n266 = n248 & ~n265 ;
  assign n267 = x129 | n266 ;
  assign n268 = x9 | x14 ;
  assign n269 = n199 | n268 ;
  assign n270 = n198 | n269 ;
  assign n271 = x17 | n195 ;
  assign n272 = n270 | n271 ;
  assign n273 = x61 | x118 ;
  assign n274 = n272 & ~n273 ;
  assign n275 = x0 & ~x123 ;
  assign n276 = ~x113 & n275 ;
  assign n277 = n274 | n276 ;
  assign n278 = ~x129 & n277 ;
  assign n279 = x10 & ~x22 ;
  assign n280 = ~n268 & n279 ;
  assign n281 = ~n220 & n280 ;
  assign n282 = ~x16 & x54 ;
  assign n283 = x4 | n155 ;
  assign n284 = n282 & ~n283 ;
  assign n285 = ~n208 & n284 ;
  assign n286 = n281 & n285 ;
  assign n287 = x4 & ~x54 ;
  assign n288 = n286 | n287 ;
  assign n289 = ~x129 & n288 ;
  assign n290 = ~x3 & n289 ;
  assign n291 = x5 & ~x54 ;
  assign n292 = x7 | n167 ;
  assign n293 = x25 | x29 ;
  assign n294 = x28 & ~n293 ;
  assign n295 = ~n292 & n294 ;
  assign n296 = x13 | n269 ;
  assign n297 = n295 & ~n296 ;
  assign n298 = x59 | n208 ;
  assign n299 = ( ~x5 & n284 ) | ( ~x5 & n291 ) | ( n284 & n291 ) ;
  assign n300 = ~n298 & n299 ;
  assign n301 = n297 & n300 ;
  assign n302 = n291 | n301 ;
  assign n303 = ~x129 & n302 ;
  assign n304 = ~x3 & n303 ;
  assign n305 = x6 & ~x54 ;
  assign n306 = x5 | x7 ;
  assign n307 = x25 & ~x29 ;
  assign n308 = ~x28 & n307 ;
  assign n309 = ~x12 & n308 ;
  assign n310 = ~n306 & n309 ;
  assign n311 = ~n296 & n310 ;
  assign n312 = ( ~x6 & n284 ) | ( ~x6 & n305 ) | ( n284 & n305 ) ;
  assign n313 = ~n298 & n312 ;
  assign n314 = n311 & n313 ;
  assign n315 = n305 | n314 ;
  assign n316 = ~x129 & n315 ;
  assign n317 = ~x3 & n316 ;
  assign n318 = x7 & ~x54 ;
  assign n319 = x18 | x21 ;
  assign n320 = x8 & ~x17 ;
  assign n321 = ~n319 & n320 ;
  assign n322 = x4 | x19 ;
  assign n323 = x7 | n322 ;
  assign n324 = n282 & ~n323 ;
  assign n325 = n321 & n324 ;
  assign n326 = x6 | n193 ;
  assign n327 = x5 | n326 ;
  assign n328 = n296 | n327 ;
  assign n329 = n325 & ~n328 ;
  assign n330 = n318 | n329 ;
  assign n331 = ~x129 & n330 ;
  assign n332 = ~x3 & n331 ;
  assign n333 = x8 & ~x54 ;
  assign n334 = n220 | n269 ;
  assign n335 = x17 | x18 ;
  assign n336 = ~x11 & x21 ;
  assign n337 = ~n335 & n336 ;
  assign n338 = x8 | n322 ;
  assign n339 = n282 & ~n338 ;
  assign n340 = n337 & n339 ;
  assign n341 = ~n334 & n340 ;
  assign n342 = n333 | n341 ;
  assign n343 = ~x129 & n342 ;
  assign n344 = ~x3 & n343 ;
  assign n345 = x9 & ~x54 ;
  assign n346 = x11 & ~n306 ;
  assign n347 = ~n167 & n346 ;
  assign n348 = ~n200 & n347 ;
  assign n349 = x9 | n322 ;
  assign n350 = n282 & ~n349 ;
  assign n351 = x8 | n151 ;
  assign n352 = n319 | n351 ;
  assign n353 = n350 & ~n352 ;
  assign n354 = n348 & n353 ;
  assign n355 = n345 | n354 ;
  assign n356 = ~x129 & n355 ;
  assign n357 = ~x3 & n356 ;
  assign n358 = x10 & ~x54 ;
  assign n359 = x10 | n322 ;
  assign n360 = n282 & ~n359 ;
  assign n361 = ~n352 & n360 ;
  assign n362 = n306 | n326 ;
  assign n363 = x9 | x22 ;
  assign n364 = n174 & ~n363 ;
  assign n365 = ~n362 & n364 ;
  assign n366 = n361 & n365 ;
  assign n367 = n358 | n366 ;
  assign n368 = ~x129 & n367 ;
  assign n369 = ~x3 & n368 ;
  assign n370 = x11 & ~x54 ;
  assign n371 = x11 | n322 ;
  assign n372 = n282 & ~n371 ;
  assign n373 = ~n352 & n372 ;
  assign n374 = ~x10 & x22 ;
  assign n375 = ~n268 & n374 ;
  assign n376 = ~n220 & n375 ;
  assign n377 = n373 & n376 ;
  assign n378 = n370 | n377 ;
  assign n379 = ~x129 & n378 ;
  assign n380 = ~x3 & n379 ;
  assign n381 = x12 & ~x54 ;
  assign n382 = x12 | n322 ;
  assign n383 = n282 & ~n382 ;
  assign n384 = x18 & ~n351 ;
  assign n385 = n383 & n384 ;
  assign n386 = x11 | n270 ;
  assign n387 = n385 & ~n386 ;
  assign n388 = n381 | n387 ;
  assign n389 = ~x129 & n388 ;
  assign n390 = ~x3 & n389 ;
  assign n391 = x13 & ~x54 ;
  assign n392 = ( ~x13 & n284 ) | ( ~x13 & n391 ) | ( n284 & n391 ) ;
  assign n393 = ~n298 & n392 ;
  assign n394 = x25 | x28 ;
  assign n395 = ( n293 & n294 ) | ( n293 & ~n394 ) | ( n294 & ~n394 ) ;
  assign n396 = ~n216 & n395 ;
  assign n397 = x7 | n269 ;
  assign n398 = n396 & ~n397 ;
  assign n399 = n393 & n398 ;
  assign n400 = n391 | n399 ;
  assign n401 = ~x129 & n400 ;
  assign n402 = ~x3 & n401 ;
  assign n403 = x14 & ~x54 ;
  assign n404 = ~x16 & n206 ;
  assign n405 = ~n322 & n404 ;
  assign n406 = ~n352 & n405 ;
  assign n407 = ~x9 & x13 ;
  assign n408 = ~n199 & n407 ;
  assign n409 = ~n362 & n408 ;
  assign n410 = n406 & n409 ;
  assign n411 = n403 | n410 ;
  assign n412 = ~x129 & n411 ;
  assign n413 = ~x3 & n412 ;
  assign n414 = x45 | x48 ;
  assign n415 = x41 | x43 ;
  assign n416 = x47 | n415 ;
  assign n417 = n414 | n416 ;
  assign n418 = n240 | n417 ;
  assign n419 = x15 | n418 ;
  assign n420 = x46 | n231 ;
  assign n421 = x82 & n234 ;
  assign n422 = ( x82 & n420 ) | ( x82 & n421 ) | ( n420 & n421 ) ;
  assign n423 = ( x82 & n419 ) | ( x82 & n422 ) | ( n419 & n422 ) ;
  assign n424 = n229 | n423 ;
  assign n425 = x70 | n424 ;
  assign n426 = n243 | n253 ;
  assign n427 = x15 & n426 ;
  assign n428 = x2 | x20 ;
  assign n429 = ~x15 & n428 ;
  assign n430 = ~n254 & n429 ;
  assign n431 = ~n238 & n430 ;
  assign n432 = ~n256 & n431 ;
  assign n433 = n427 | n432 ;
  assign n434 = x82 & n433 ;
  assign n435 = x15 & n263 ;
  assign n436 = n434 | n435 ;
  assign n437 = n425 & ~n436 ;
  assign n438 = x129 | n437 ;
  assign n439 = x16 & ~x54 ;
  assign n440 = ( x6 & n214 ) | ( x6 & n217 ) | ( n214 & n217 ) ;
  assign n441 = ~n269 & n440 ;
  assign n442 = n285 & n441 ;
  assign n443 = n439 | n442 ;
  assign n444 = ~x129 & n443 ;
  assign n445 = ~x3 & n444 ;
  assign n446 = x17 & ~x54 ;
  assign n447 = x7 | n197 ;
  assign n448 = x12 | n394 ;
  assign n449 = n447 | n448 ;
  assign n450 = n296 | n449 ;
  assign n451 = x11 | n170 ;
  assign n452 = ~x29 & x59 ;
  assign n453 = ~n451 & n452 ;
  assign n454 = ( n203 & n284 ) | ( n203 & n439 ) | ( n284 & n439 ) ;
  assign n455 = n453 & n454 ;
  assign n456 = ~n450 & n455 ;
  assign n457 = n446 | n456 ;
  assign n458 = ~x129 & n457 ;
  assign n459 = ~x3 & n458 ;
  assign n460 = x18 & ~x54 ;
  assign n461 = x16 & x54 ;
  assign n462 = ~n283 & n461 ;
  assign n463 = ~n208 & n462 ;
  assign n464 = ~n334 & n463 ;
  assign n465 = n460 | n464 ;
  assign n466 = ~x129 & n465 ;
  assign n467 = ~x3 & n466 ;
  assign n468 = x19 & ~x54 ;
  assign n469 = x17 & ~n451 ;
  assign n470 = n284 & n469 ;
  assign n471 = ~n334 & n470 ;
  assign n472 = n468 | n471 ;
  assign n473 = ~x129 & n472 ;
  assign n474 = ~x3 & n473 ;
  assign n475 = x40 | x42 ;
  assign n476 = n231 | n475 ;
  assign n477 = x44 | n258 ;
  assign n478 = n476 | n477 ;
  assign n479 = x43 | n230 ;
  assign n480 = n256 | n479 ;
  assign n481 = ( ~x45 & n257 ) | ( ~x45 & n480 ) | ( n257 & n480 ) ;
  assign n482 = n478 | n481 ;
  assign n483 = x82 & n482 ;
  assign n484 = n229 | n483 ;
  assign n485 = x71 | n484 ;
  assign n486 = x50 | n249 ;
  assign n487 = x15 | x49 ;
  assign n488 = n233 | n487 ;
  assign n489 = n486 | n488 ;
  assign n490 = n481 | n489 ;
  assign n491 = x20 & n490 ;
  assign n492 = x2 & ~n482 ;
  assign n493 = n491 | n492 ;
  assign n494 = x82 & n493 ;
  assign n495 = x20 & n263 ;
  assign n496 = n494 | n495 ;
  assign n497 = n485 & ~n496 ;
  assign n498 = x129 | n497 ;
  assign n499 = x21 & ~x54 ;
  assign n500 = n207 | n335 ;
  assign n501 = ~x21 & x54 ;
  assign n502 = x19 & n501 ;
  assign n503 = ~n156 & n502 ;
  assign n504 = ~n500 & n503 ;
  assign n505 = ~n334 & n504 ;
  assign n506 = n499 | n505 ;
  assign n507 = ~x129 & n506 ;
  assign n508 = ~x3 & n507 ;
  assign n509 = x22 & ~x54 ;
  assign n510 = x22 | n322 ;
  assign n511 = n282 & ~n510 ;
  assign n512 = ~n352 & n511 ;
  assign n513 = x9 | x10 ;
  assign n514 = n148 | n513 ;
  assign n515 = x5 & ~x7 ;
  assign n516 = ~n326 & n515 ;
  assign n517 = ~n514 & n516 ;
  assign n518 = n512 & n517 ;
  assign n519 = n509 | n518 ;
  assign n520 = ~x129 & n519 ;
  assign n521 = ~x3 & n520 ;
  assign n522 = ~x23 & x55 ;
  assign n523 = x129 | n522 ;
  assign n524 = x61 & ~n523 ;
  assign n525 = n428 | n487 ;
  assign n526 = x82 & n525 ;
  assign n527 = n229 & ~n526 ;
  assign n528 = ( x82 & n417 ) | ( x82 & n422 ) | ( n417 & n422 ) ;
  assign n529 = n527 | n528 ;
  assign n530 = ~x24 & n529 ;
  assign n531 = x2 | x45 ;
  assign n532 = n255 | n531 ;
  assign n533 = n258 | n532 ;
  assign n534 = x82 & n254 ;
  assign n535 = ( x82 & n533 ) | ( x82 & n534 ) | ( n533 & n534 ) ;
  assign n536 = n229 | n535 ;
  assign n537 = x63 & ~n536 ;
  assign n538 = x24 & x82 ;
  assign n539 = ~n233 & n538 ;
  assign n540 = ~n486 & n539 ;
  assign n541 = ~n480 & n540 ;
  assign n542 = x129 | n541 ;
  assign n543 = n537 | n542 ;
  assign n544 = n530 | n543 ;
  assign n545 = x25 & ~x116 ;
  assign n546 = x26 & n545 ;
  assign n547 = x39 | x52 ;
  assign n548 = x51 | n547 ;
  assign n549 = n546 | n548 ;
  assign n550 = x26 & x116 ;
  assign n551 = x95 | x100 ;
  assign n552 = x97 & ~x110 ;
  assign n553 = ( ~x110 & n551 ) | ( ~x110 & n552 ) | ( n551 & n552 ) ;
  assign n554 = x25 & ~n553 ;
  assign n555 = n550 | n554 ;
  assign n556 = ( n546 & n549 ) | ( n546 & n555 ) | ( n549 & n555 ) ;
  assign n557 = ~x85 & n556 ;
  assign n558 = x26 | x27 ;
  assign n559 = x85 & n545 ;
  assign n560 = x85 | x110 ;
  assign n561 = x96 | n560 ;
  assign n562 = x85 & x116 ;
  assign n563 = ( x100 & ~n561 ) | ( x100 & n562 ) | ( ~n561 & n562 ) ;
  assign n564 = ( ~n558 & n559 ) | ( ~n558 & n563 ) | ( n559 & n563 ) ;
  assign n565 = ~n558 & n564 ;
  assign n566 = ( ~x27 & n557 ) | ( ~x27 & n565 ) | ( n557 & n565 ) ;
  assign n567 = ~n548 & n554 ;
  assign n568 = x26 | x85 ;
  assign n569 = ~x51 & x116 ;
  assign n570 = ~n547 & n569 ;
  assign n571 = ( x27 & n545 ) | ( x27 & n570 ) | ( n545 & n570 ) ;
  assign n572 = ~n568 & n571 ;
  assign n573 = ( n567 & ~n568 ) | ( n567 & n572 ) | ( ~n568 & n572 ) ;
  assign n574 = ~x53 & n573 ;
  assign n575 = ( ~x53 & n566 ) | ( ~x53 & n574 ) | ( n566 & n574 ) ;
  assign n576 = x27 | x85 ;
  assign n577 = ~x53 & x58 ;
  assign n578 = ~n576 & n577 ;
  assign n579 = ( ~x26 & n545 ) | ( ~x26 & n550 ) | ( n545 & n550 ) ;
  assign n580 = n578 & n579 ;
  assign n581 = x58 & ~n580 ;
  assign n582 = x53 & ~x85 ;
  assign n583 = ~x27 & n582 ;
  assign n584 = n579 & n583 ;
  assign n585 = ( n580 & ~n581 ) | ( n580 & n584 ) | ( ~n581 & n584 ) ;
  assign n586 = ( n575 & ~n581 ) | ( n575 & n585 ) | ( ~n581 & n585 ) ;
  assign n587 = ~x129 & n586 ;
  assign n588 = ~x3 & n587 ;
  assign n589 = x85 & ~x116 ;
  assign n590 = x110 | n589 ;
  assign n591 = n550 | n590 ;
  assign n592 = x96 | n591 ;
  assign n593 = ~x26 & n562 ;
  assign n594 = n592 & ~n593 ;
  assign n595 = x100 & ~n594 ;
  assign n596 = x85 | n570 ;
  assign n597 = x26 & ~n596 ;
  assign n598 = n595 | n597 ;
  assign n599 = ~x129 & n598 ;
  assign n600 = ~x3 & n599 ;
  assign n601 = x27 | x53 ;
  assign n602 = x58 | n601 ;
  assign n603 = n600 & ~n602 ;
  assign n604 = x95 & ~x96 ;
  assign n605 = x27 & x116 ;
  assign n606 = n590 | n605 ;
  assign n607 = n604 & ~n606 ;
  assign n608 = ~x27 & n562 ;
  assign n609 = n607 | n608 ;
  assign n610 = ~x100 & n609 ;
  assign n611 = x27 & ~n596 ;
  assign n612 = n610 | n611 ;
  assign n613 = ~x129 & n612 ;
  assign n614 = ~x3 & n613 ;
  assign n615 = x53 | x58 ;
  assign n616 = x26 | n615 ;
  assign n617 = n614 & ~n616 ;
  assign n618 = ~x26 & n548 ;
  assign n619 = x27 | n548 ;
  assign n620 = ~n618 & n619 ;
  assign n621 = n553 | n620 ;
  assign n622 = x26 & ~x27 ;
  assign n623 = ~x26 & x27 ;
  assign n624 = n622 | n623 ;
  assign n625 = ~x116 & n624 ;
  assign n626 = n621 & ~n625 ;
  assign n627 = x28 & ~n626 ;
  assign n628 = x26 | x100 ;
  assign n629 = x110 | n628 ;
  assign n630 = n604 & ~n629 ;
  assign n631 = ~n548 & n550 ;
  assign n632 = n630 | n631 ;
  assign n633 = ~x27 & n632 ;
  assign n634 = n605 & n618 ;
  assign n635 = n633 | n634 ;
  assign n636 = n627 | n635 ;
  assign n637 = ~x85 & n636 ;
  assign n638 = ( ~x85 & x100 ) | ( ~x85 & x116 ) | ( x100 & x116 ) ;
  assign n639 = ( x28 & x85 ) | ( x28 & x116 ) | ( x85 & x116 ) ;
  assign n640 = ~n638 & n639 ;
  assign n641 = ~n558 & n640 ;
  assign n642 = n637 | n641 ;
  assign n643 = ~x53 & n642 ;
  assign n644 = ~x26 & n582 ;
  assign n645 = x28 & ~x116 ;
  assign n646 = ~x27 & n645 ;
  assign n647 = n644 & n646 ;
  assign n648 = n643 | n647 ;
  assign n649 = ~x58 & n648 ;
  assign n650 = ~n568 & n577 ;
  assign n651 = n646 & n650 ;
  assign n652 = n649 | n651 ;
  assign n653 = ~x129 & n652 ;
  assign n654 = ~x3 & n653 ;
  assign n655 = x29 & ~x116 ;
  assign n656 = n576 | n615 ;
  assign n657 = x26 & ~n656 ;
  assign n658 = ( n605 & n655 ) | ( n605 & n657 ) | ( n655 & n657 ) ;
  assign n659 = ~x96 & n552 ;
  assign n660 = x97 | n551 ;
  assign n661 = x29 & ~n660 ;
  assign n662 = ( ~n551 & n659 ) | ( ~n551 & n661 ) | ( n659 & n661 ) ;
  assign n663 = x29 & x110 ;
  assign n664 = ~x58 & n663 ;
  assign n665 = ( ~x58 & n662 ) | ( ~x58 & n664 ) | ( n662 & n664 ) ;
  assign n666 = x97 & x116 ;
  assign n667 = ( n577 & n655 ) | ( n577 & n666 ) | ( n655 & n666 ) ;
  assign n668 = n577 & n667 ;
  assign n669 = ( ~x53 & n665 ) | ( ~x53 & n668 ) | ( n665 & n668 ) ;
  assign n670 = x27 & n655 ;
  assign n671 = ~n615 & n670 ;
  assign n672 = x27 & ~n671 ;
  assign n673 = x53 & ~x58 ;
  assign n674 = n655 & n673 ;
  assign n675 = ( n671 & ~n672 ) | ( n671 & n674 ) | ( ~n672 & n674 ) ;
  assign n676 = ( n669 & ~n672 ) | ( n669 & n675 ) | ( ~n672 & n675 ) ;
  assign n677 = ~x85 & n676 ;
  assign n678 = x85 & ~n615 ;
  assign n679 = ~n601 & n678 ;
  assign n680 = n655 & n679 ;
  assign n681 = x26 | n680 ;
  assign n682 = n677 | n681 ;
  assign n683 = ( ~x26 & n658 ) | ( ~x26 & n682 ) | ( n658 & n682 ) ;
  assign n684 = ~x129 & n683 ;
  assign n685 = ~x3 & n684 ;
  assign n686 = x88 & x106 ;
  assign n687 = ( ~x60 & x106 ) | ( ~x60 & x109 ) | ( x106 & x109 ) ;
  assign n688 = ( x30 & ~x106 ) | ( x30 & x109 ) | ( ~x106 & x109 ) ;
  assign n689 = ~n687 & n688 ;
  assign n690 = n686 | n689 ;
  assign n691 = ~x129 & n690 ;
  assign n692 = x89 & x106 ;
  assign n693 = ( ~x30 & x106 ) | ( ~x30 & x109 ) | ( x106 & x109 ) ;
  assign n694 = ( x31 & ~x106 ) | ( x31 & x109 ) | ( ~x106 & x109 ) ;
  assign n695 = ~n693 & n694 ;
  assign n696 = n692 | n695 ;
  assign n697 = ~x129 & n696 ;
  assign n698 = x99 & x106 ;
  assign n699 = ( ~x31 & x106 ) | ( ~x31 & x109 ) | ( x106 & x109 ) ;
  assign n700 = ( x32 & ~x106 ) | ( x32 & x109 ) | ( ~x106 & x109 ) ;
  assign n701 = ~n699 & n700 ;
  assign n702 = n698 | n701 ;
  assign n703 = ~x129 & n702 ;
  assign n704 = x90 & x106 ;
  assign n705 = ( ~x32 & x106 ) | ( ~x32 & x109 ) | ( x106 & x109 ) ;
  assign n706 = ( x33 & ~x106 ) | ( x33 & x109 ) | ( ~x106 & x109 ) ;
  assign n707 = ~n705 & n706 ;
  assign n708 = n704 | n707 ;
  assign n709 = ~x129 & n708 ;
  assign n710 = x91 & x106 ;
  assign n711 = ( ~x33 & x106 ) | ( ~x33 & x109 ) | ( x106 & x109 ) ;
  assign n712 = ( x34 & ~x106 ) | ( x34 & x109 ) | ( ~x106 & x109 ) ;
  assign n713 = ~n711 & n712 ;
  assign n714 = n710 | n713 ;
  assign n715 = ~x129 & n714 ;
  assign n716 = x92 & x106 ;
  assign n717 = ( ~x34 & x106 ) | ( ~x34 & x109 ) | ( x106 & x109 ) ;
  assign n718 = ( x35 & ~x106 ) | ( x35 & x109 ) | ( ~x106 & x109 ) ;
  assign n719 = ~n717 & n718 ;
  assign n720 = n716 | n719 ;
  assign n721 = ~x129 & n720 ;
  assign n722 = x98 & x106 ;
  assign n723 = ( ~x35 & x106 ) | ( ~x35 & x109 ) | ( x106 & x109 ) ;
  assign n724 = ( x36 & ~x106 ) | ( x36 & x109 ) | ( ~x106 & x109 ) ;
  assign n725 = ~n723 & n724 ;
  assign n726 = n722 | n725 ;
  assign n727 = ~x129 & n726 ;
  assign n728 = x93 & x106 ;
  assign n729 = ( ~x36 & x106 ) | ( ~x36 & x109 ) | ( x106 & x109 ) ;
  assign n730 = ( x37 & ~x106 ) | ( x37 & x109 ) | ( ~x106 & x109 ) ;
  assign n731 = ~n729 & n730 ;
  assign n732 = n728 | n731 ;
  assign n733 = ~x129 & n732 ;
  assign n734 = n239 | n531 ;
  assign n735 = x82 & n734 ;
  assign n736 = n229 & ~n735 ;
  assign n737 = ( ~x48 & n263 ) | ( ~x48 & n736 ) | ( n263 & n736 ) ;
  assign n738 = ( ~n241 & n263 ) | ( ~n241 & n737 ) | ( n263 & n737 ) ;
  assign n739 = ( ~n252 & n263 ) | ( ~n252 & n738 ) | ( n263 & n738 ) ;
  assign n740 = n421 | n739 ;
  assign n741 = ~x38 & n740 ;
  assign n742 = n230 | n241 ;
  assign n743 = x50 | n234 ;
  assign n744 = n742 | n743 ;
  assign n745 = ( ~x45 & n414 ) | ( ~x45 & n734 ) | ( n414 & n734 ) ;
  assign n746 = n744 | n745 ;
  assign n747 = x82 & n746 ;
  assign n748 = n229 | n747 ;
  assign n749 = x74 & ~n748 ;
  assign n750 = x82 & n250 ;
  assign n751 = ( x129 & ~n421 ) | ( x129 & n750 ) | ( ~n421 & n750 ) ;
  assign n752 = ( x38 & x129 ) | ( x38 & n751 ) | ( x129 & n751 ) ;
  assign n753 = n749 | n752 ;
  assign n754 = n741 | n753 ;
  assign n755 = ~x51 & x109 ;
  assign n756 = ~n547 & n755 ;
  assign n757 = x106 | n756 ;
  assign n758 = x52 & ~n755 ;
  assign n759 = ( ~x52 & n755 ) | ( ~x52 & n758 ) | ( n755 & n758 ) ;
  assign n760 = x39 & ~n759 ;
  assign n761 = n757 | n760 ;
  assign n762 = ~x129 & n761 ;
  assign n763 = x82 & n233 ;
  assign n764 = ( ~n232 & n263 ) | ( ~n232 & n738 ) | ( n263 & n738 ) ;
  assign n765 = n763 | n764 ;
  assign n766 = ~x40 & n765 ;
  assign n767 = n231 | n233 ;
  assign n768 = n742 | n767 ;
  assign n769 = n745 | n768 ;
  assign n770 = x82 & n769 ;
  assign n771 = n229 | n770 ;
  assign n772 = x73 & ~n771 ;
  assign n773 = ~n233 & n421 ;
  assign n774 = x129 | n773 ;
  assign n775 = n772 | n774 ;
  assign n776 = n766 | n775 ;
  assign n777 = n422 | n738 ;
  assign n778 = ~x41 & n777 ;
  assign n779 = n241 | n251 ;
  assign n780 = n745 | n779 ;
  assign n781 = ( x82 & n750 ) | ( x82 & n780 ) | ( n750 & n780 ) ;
  assign n782 = n229 | n781 ;
  assign n783 = x76 & ~n782 ;
  assign n784 = n249 | n251 ;
  assign n785 = x41 & x82 ;
  assign n786 = ~n233 & n785 ;
  assign n787 = ~n784 & n786 ;
  assign n788 = x129 | n787 ;
  assign n789 = n783 | n788 ;
  assign n790 = n778 | n789 ;
  assign n791 = x44 & x82 ;
  assign n792 = ( n263 & ~n416 ) | ( n263 & n737 ) | ( ~n416 & n737 ) ;
  assign n793 = ( n263 & ~n784 ) | ( n263 & n792 ) | ( ~n784 & n792 ) ;
  assign n794 = n791 | n793 ;
  assign n795 = ~x42 & n794 ;
  assign n796 = x44 | n486 ;
  assign n797 = n742 | n796 ;
  assign n798 = n745 | n797 ;
  assign n799 = x82 & n798 ;
  assign n800 = n229 | n799 ;
  assign n801 = x72 & ~n800 ;
  assign n802 = ~x44 & x82 ;
  assign n803 = x42 & n802 ;
  assign n804 = x129 | n803 ;
  assign n805 = n801 | n804 ;
  assign n806 = n795 | n805 ;
  assign n807 = x82 & n253 ;
  assign n808 = ( ~n255 & n263 ) | ( ~n255 & n736 ) | ( n263 & n736 ) ;
  assign n809 = n807 | n808 ;
  assign n810 = ~x43 & n809 ;
  assign n811 = n239 | n532 ;
  assign n812 = ( x82 & n807 ) | ( x82 & n811 ) | ( n807 & n811 ) ;
  assign n813 = n229 | n812 ;
  assign n814 = x77 & ~n813 ;
  assign n815 = x43 & ~n475 ;
  assign n816 = n802 & n815 ;
  assign n817 = ~n232 & n816 ;
  assign n818 = x129 | n817 ;
  assign n819 = n814 | n818 ;
  assign n820 = n810 | n819 ;
  assign n821 = x129 | n791 ;
  assign n822 = n742 | n745 ;
  assign n823 = n476 | n822 ;
  assign n824 = x82 & n823 ;
  assign n825 = ( x44 & n229 ) | ( x44 & n824 ) | ( n229 & n824 ) ;
  assign n826 = ( x67 & n229 ) | ( x67 & ~n824 ) | ( n229 & ~n824 ) ;
  assign n827 = ~n825 & n826 ;
  assign n828 = n821 | n827 ;
  assign n829 = ( x82 & n241 ) | ( x82 & n807 ) | ( n241 & n807 ) ;
  assign n830 = ( x48 & x82 ) | ( x48 & n829 ) | ( x82 & n829 ) ;
  assign n831 = ( ~x24 & n263 ) | ( ~x24 & n527 ) | ( n263 & n527 ) ;
  assign n832 = n830 | n831 ;
  assign n833 = ~x45 & n832 ;
  assign n834 = x2 | n255 ;
  assign n835 = n239 | n834 ;
  assign n836 = n254 | n835 ;
  assign n837 = x82 & n836 ;
  assign n838 = n229 | n837 ;
  assign n839 = x68 & ~n838 ;
  assign n840 = n242 | n252 ;
  assign n841 = x38 | n475 ;
  assign n842 = x45 & ~n841 ;
  assign n843 = n802 & n842 ;
  assign n844 = ~n840 & n843 ;
  assign n845 = x129 | n844 ;
  assign n846 = n839 | n845 ;
  assign n847 = n833 | n846 ;
  assign n848 = x50 | n250 ;
  assign n849 = n416 | n745 ;
  assign n850 = n848 | n849 ;
  assign n851 = x82 & n850 ;
  assign n852 = n229 | n851 ;
  assign n853 = ( n792 & n848 ) | ( n792 & n852 ) | ( n848 & n852 ) ;
  assign n854 = ~x46 & n853 ;
  assign n855 = x75 & ~n852 ;
  assign n856 = n422 & ~n848 ;
  assign n857 = x129 | n856 ;
  assign n858 = n855 | n857 ;
  assign n859 = n854 | n858 ;
  assign n860 = ( x82 & n534 ) | ( x82 & n745 ) | ( n534 & n745 ) ;
  assign n861 = n229 | n860 ;
  assign n862 = x64 & ~n861 ;
  assign n863 = n415 | n420 ;
  assign n864 = x47 & ~n475 ;
  assign n865 = n802 & n864 ;
  assign n866 = ~n863 & n865 ;
  assign n867 = x129 | n866 ;
  assign n868 = n862 | n867 ;
  assign n869 = ( ~x47 & n534 ) | ( ~x47 & n808 ) | ( n534 & n808 ) ;
  assign n870 = n868 | n869 ;
  assign n871 = x2 | x47 ;
  assign n872 = n259 | n871 ;
  assign n873 = ( x82 & n534 ) | ( x82 & n872 ) | ( n534 & n872 ) ;
  assign n874 = n229 | n873 ;
  assign n875 = x62 & ~n874 ;
  assign n876 = n241 | n252 ;
  assign n877 = x48 & ~n841 ;
  assign n878 = n802 & n877 ;
  assign n879 = ~n876 & n878 ;
  assign n880 = x129 | n879 ;
  assign n881 = n875 | n880 ;
  assign n882 = ( ~x48 & n737 ) | ( ~x48 & n829 ) | ( n737 & n829 ) ;
  assign n883 = n881 | n882 ;
  assign n884 = n238 | n848 ;
  assign n885 = n480 | n884 ;
  assign n886 = x82 & n885 ;
  assign n887 = n229 | n886 ;
  assign n888 = x69 | n887 ;
  assign n889 = x24 | x42 ;
  assign n890 = n796 | n889 ;
  assign n891 = n480 | n890 ;
  assign n892 = x49 & n891 ;
  assign n893 = x2 | n237 ;
  assign n894 = ~n884 & n893 ;
  assign n895 = ~n742 & n894 ;
  assign n896 = ~n414 & n895 ;
  assign n897 = n892 | n896 ;
  assign n898 = x82 & n897 ;
  assign n899 = x49 & n263 ;
  assign n900 = n898 | n899 ;
  assign n901 = n888 & ~n900 ;
  assign n902 = x129 | n901 ;
  assign n903 = n479 | n834 ;
  assign n904 = n259 | n903 ;
  assign n905 = x82 & n904 ;
  assign n906 = n229 & ~n905 ;
  assign n907 = n750 | n906 ;
  assign n908 = ~x50 & n907 ;
  assign n909 = ( x82 & n750 ) | ( x82 & n822 ) | ( n750 & n822 ) ;
  assign n910 = n229 | n909 ;
  assign n911 = x66 & ~n910 ;
  assign n912 = x50 & ~n841 ;
  assign n913 = n802 & n912 ;
  assign n914 = x129 | n913 ;
  assign n915 = n911 | n914 ;
  assign n916 = n908 | n915 ;
  assign n917 = x51 & ~x109 ;
  assign n918 = ( ~x51 & x106 ) | ( ~x51 & x109 ) | ( x106 & x109 ) ;
  assign n919 = ( ~x129 & n917 ) | ( ~x129 & n918 ) | ( n917 & n918 ) ;
  assign n920 = ( ~x52 & x106 ) | ( ~x52 & n755 ) | ( x106 & n755 ) ;
  assign n921 = ( ~x129 & n758 ) | ( ~x129 & n920 ) | ( n758 & n920 ) ;
  assign n922 = x58 & x116 ;
  assign n923 = x58 | x110 ;
  assign n924 = x96 | n923 ;
  assign n925 = n551 | n924 ;
  assign n926 = ~n922 & n925 ;
  assign n927 = x53 | n926 ;
  assign n928 = x97 & ~n927 ;
  assign n929 = ~x116 & n673 ;
  assign n930 = n928 | n929 ;
  assign n931 = ~x129 & n930 ;
  assign n932 = ~x3 & n931 ;
  assign n933 = ~n576 & n932 ;
  assign n934 = ~x26 & n933 ;
  assign n935 = ( n534 & ~n807 ) | ( n534 & n813 ) | ( ~n807 & n813 ) ;
  assign n936 = ~x129 & n935 ;
  assign n937 = x123 | x129 ;
  assign n938 = x114 & ~x122 ;
  assign n939 = ~n937 & n938 ;
  assign n940 = x58 & ~x116 ;
  assign n941 = ~x26 & x58 ;
  assign n942 = x37 & ~x116 ;
  assign n943 = n941 | n942 ;
  assign n944 = ~n940 & n943 ;
  assign n945 = ( x58 & x94 ) | ( x58 & n550 ) | ( x94 & n550 ) ;
  assign n946 = ( ~x58 & n941 ) | ( ~x58 & n945 ) | ( n941 & n945 ) ;
  assign n947 = n944 | n946 ;
  assign n948 = ~x53 & n947 ;
  assign n949 = ~x26 & x37 ;
  assign n950 = ~x58 & n949 ;
  assign n951 = n948 | n950 ;
  assign n952 = ~x85 & n951 ;
  assign n953 = ~n615 & n949 ;
  assign n954 = n952 | n953 ;
  assign n955 = ~x27 & n954 ;
  assign n956 = x85 | n615 ;
  assign n957 = n949 & ~n956 ;
  assign n958 = n955 | n957 ;
  assign n959 = ~x129 & n958 ;
  assign n960 = ~x3 & n959 ;
  assign n961 = x26 | x53 ;
  assign n962 = x85 | n961 ;
  assign n963 = x116 | n962 ;
  assign n964 = ( x26 & x53 ) | ( x26 & x85 ) | ( x53 & x85 ) ;
  assign n965 = x58 | n964 ;
  assign n966 = n963 & n965 ;
  assign n967 = x57 & ~n966 ;
  assign n968 = x60 & n922 ;
  assign n969 = ~n962 & n968 ;
  assign n970 = n967 | n969 ;
  assign n971 = ~x27 & n970 ;
  assign n972 = x57 & ~x58 ;
  assign n973 = ~n962 & n972 ;
  assign n974 = n971 | n973 ;
  assign n975 = ~x129 & n974 ;
  assign n976 = ~x3 & n975 ;
  assign n977 = ~n558 & n940 ;
  assign n978 = x116 & n624 ;
  assign n979 = ~x58 & n978 ;
  assign n980 = ~n548 & n979 ;
  assign n981 = n977 | n980 ;
  assign n982 = ~x129 & n981 ;
  assign n983 = ~x3 & n982 ;
  assign n984 = ~x53 & n983 ;
  assign n985 = ~x85 & n984 ;
  assign n986 = ( x53 & x58 ) | ( x53 & x116 ) | ( x58 & x116 ) ;
  assign n987 = n553 & ~n615 ;
  assign n988 = n986 | n987 ;
  assign n989 = x59 & ~n988 ;
  assign n990 = x96 & n987 ;
  assign n991 = n989 | n990 ;
  assign n992 = ~x85 & n991 ;
  assign n993 = x59 & ~x116 ;
  assign n994 = n678 & n993 ;
  assign n995 = n992 | n994 ;
  assign n996 = ~x27 & n995 ;
  assign n997 = x27 & ~n956 ;
  assign n998 = n993 & n997 ;
  assign n999 = n996 | n998 ;
  assign n1000 = ~x26 & n999 ;
  assign n1001 = n657 & n993 ;
  assign n1002 = n1000 | n1001 ;
  assign n1003 = ~x129 & n1002 ;
  assign n1004 = ~x3 & n1003 ;
  assign n1005 = x117 | x122 ;
  assign n1006 = x60 & n1005 ;
  assign n1007 = x123 & ~n1005 ;
  assign n1008 = n1006 | n1007 ;
  assign n1009 = ~x114 & x123 ;
  assign n1010 = ~x122 & n1009 ;
  assign n1011 = ~x129 & n1010 ;
  assign n1012 = x136 & ~x137 ;
  assign n1013 = x132 & x133 ;
  assign n1014 = x131 & n1013 ;
  assign n1015 = ~x138 & n1014 ;
  assign n1016 = n1012 & n1015 ;
  assign n1017 = x62 & ~n1016 ;
  assign n1018 = ~x136 & x140 ;
  assign n1019 = ( ~x140 & n1016 ) | ( ~x140 & n1018 ) | ( n1016 & n1018 ) ;
  assign n1020 = n1017 | n1019 ;
  assign n1021 = ~x129 & n1020 ;
  assign n1022 = x63 & ~n1016 ;
  assign n1023 = ~x142 & n1016 ;
  assign n1024 = n1022 | n1023 ;
  assign n1025 = ~x129 & n1024 ;
  assign n1026 = x64 & ~n1016 ;
  assign n1027 = ~x136 & x139 ;
  assign n1028 = ( ~x139 & n1016 ) | ( ~x139 & n1027 ) | ( n1016 & n1027 ) ;
  assign n1029 = n1026 | n1028 ;
  assign n1030 = ~x129 & n1029 ;
  assign n1031 = x65 & ~n1016 ;
  assign n1032 = ~x146 & n1016 ;
  assign n1033 = n1031 | n1032 ;
  assign n1034 = ~x129 & n1033 ;
  assign n1035 = x136 | x137 ;
  assign n1036 = n1015 & ~n1035 ;
  assign n1037 = ( x129 & x143 ) | ( x129 & n1036 ) | ( x143 & n1036 ) ;
  assign n1038 = ( x66 & ~x129 ) | ( x66 & n1036 ) | ( ~x129 & n1036 ) ;
  assign n1039 = ~n1037 & n1038 ;
  assign n1040 = ( x129 & x139 ) | ( x129 & n1036 ) | ( x139 & n1036 ) ;
  assign n1041 = ( x67 & ~x129 ) | ( x67 & n1036 ) | ( ~x129 & n1036 ) ;
  assign n1042 = ~n1040 & n1041 ;
  assign n1043 = x68 & ~n1016 ;
  assign n1044 = ~x136 & x141 ;
  assign n1045 = ( ~x141 & n1016 ) | ( ~x141 & n1044 ) | ( n1016 & n1044 ) ;
  assign n1046 = n1043 | n1045 ;
  assign n1047 = ~x129 & n1046 ;
  assign n1048 = x69 & ~n1016 ;
  assign n1049 = ~x143 & n1016 ;
  assign n1050 = n1048 | n1049 ;
  assign n1051 = ~x129 & n1050 ;
  assign n1052 = x70 & ~n1016 ;
  assign n1053 = ~x144 & n1016 ;
  assign n1054 = n1052 | n1053 ;
  assign n1055 = ~x129 & n1054 ;
  assign n1056 = x71 & ~n1016 ;
  assign n1057 = ~x145 & n1016 ;
  assign n1058 = n1056 | n1057 ;
  assign n1059 = ~x129 & n1058 ;
  assign n1060 = ( x129 & x140 ) | ( x129 & n1036 ) | ( x140 & n1036 ) ;
  assign n1061 = ( x72 & ~x129 ) | ( x72 & n1036 ) | ( ~x129 & n1036 ) ;
  assign n1062 = ~n1060 & n1061 ;
  assign n1063 = ( x129 & x141 ) | ( x129 & n1036 ) | ( x141 & n1036 ) ;
  assign n1064 = ( x73 & ~x129 ) | ( x73 & n1036 ) | ( ~x129 & n1036 ) ;
  assign n1065 = ~n1063 & n1064 ;
  assign n1066 = ( x129 & x142 ) | ( x129 & n1036 ) | ( x142 & n1036 ) ;
  assign n1067 = ( x74 & ~x129 ) | ( x74 & n1036 ) | ( ~x129 & n1036 ) ;
  assign n1068 = ~n1066 & n1067 ;
  assign n1069 = ( x129 & x144 ) | ( x129 & n1036 ) | ( x144 & n1036 ) ;
  assign n1070 = ( x75 & ~x129 ) | ( x75 & n1036 ) | ( ~x129 & n1036 ) ;
  assign n1071 = ~n1069 & n1070 ;
  assign n1072 = ( x129 & x145 ) | ( x129 & n1036 ) | ( x145 & n1036 ) ;
  assign n1073 = ( x76 & ~x129 ) | ( x76 & n1036 ) | ( ~x129 & n1036 ) ;
  assign n1074 = ~n1072 & n1073 ;
  assign n1075 = ( x129 & x146 ) | ( x129 & n1036 ) | ( x146 & n1036 ) ;
  assign n1076 = ( x77 & ~x129 ) | ( x77 & n1036 ) | ( ~x129 & n1036 ) ;
  assign n1077 = ~n1075 & n1076 ;
  assign n1078 = ~x136 & x137 ;
  assign n1079 = n1015 & n1078 ;
  assign n1080 = ( x129 & ~x142 ) | ( x129 & n1079 ) | ( ~x142 & n1079 ) ;
  assign n1081 = ( x78 & ~x129 ) | ( x78 & n1079 ) | ( ~x129 & n1079 ) ;
  assign n1082 = ~n1080 & n1081 ;
  assign n1083 = ( x129 & ~x143 ) | ( x129 & n1079 ) | ( ~x143 & n1079 ) ;
  assign n1084 = ( x79 & ~x129 ) | ( x79 & n1079 ) | ( ~x129 & n1079 ) ;
  assign n1085 = ~n1083 & n1084 ;
  assign n1086 = ( x129 & ~x144 ) | ( x129 & n1079 ) | ( ~x144 & n1079 ) ;
  assign n1087 = ( x80 & ~x129 ) | ( x80 & n1079 ) | ( ~x129 & n1079 ) ;
  assign n1088 = ~n1086 & n1087 ;
  assign n1089 = ( x129 & ~x145 ) | ( x129 & n1079 ) | ( ~x145 & n1079 ) ;
  assign n1090 = ( x81 & ~x129 ) | ( x81 & n1079 ) | ( ~x129 & n1079 ) ;
  assign n1091 = ~n1089 & n1090 ;
  assign n1092 = ( x129 & ~x146 ) | ( x129 & n1079 ) | ( ~x146 & n1079 ) ;
  assign n1093 = ( x82 & ~x129 ) | ( x82 & n1079 ) | ( ~x129 & n1079 ) ;
  assign n1094 = ~n1092 & n1093 ;
  assign n1095 = ( x89 & x136 ) | ( x89 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1096 = ( ~x62 & x136 ) | ( ~x62 & x138 ) | ( x136 & x138 ) ;
  assign n1097 = n1095 & n1096 ;
  assign n1098 = ( ~x119 & x136 ) | ( ~x119 & x138 ) | ( x136 & x138 ) ;
  assign n1099 = ( x72 & x136 ) | ( x72 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1100 = n1098 | n1099 ;
  assign n1101 = ~n1097 & n1100 ;
  assign n1102 = x137 | n1101 ;
  assign n1103 = x136 & ~x138 ;
  assign n1104 = x31 & n1103 ;
  assign n1105 = ( x115 & x136 ) | ( x115 & x138 ) | ( x136 & x138 ) ;
  assign n1106 = ( x87 & ~x136 ) | ( x87 & x138 ) | ( ~x136 & x138 ) ;
  assign n1107 = ~n1105 & n1106 ;
  assign n1108 = n1104 | n1107 ;
  assign n1109 = x137 & n1108 ;
  assign n1110 = n1102 & ~n1109 ;
  assign n1111 = ( x129 & ~x141 ) | ( x129 & n1079 ) | ( ~x141 & n1079 ) ;
  assign n1112 = ( x84 & ~x129 ) | ( x84 & n1079 ) | ( ~x129 & n1079 ) ;
  assign n1113 = ~n1111 & n1112 ;
  assign n1114 = ~n560 & n660 ;
  assign n1115 = ( n561 & n589 ) | ( n561 & n1114 ) | ( n589 & n1114 ) ;
  assign n1116 = ~x129 & n1115 ;
  assign n1117 = ~x3 & n1116 ;
  assign n1118 = ~n602 & n1117 ;
  assign n1119 = ~x26 & n1118 ;
  assign n1120 = ( x129 & ~x139 ) | ( x129 & n1079 ) | ( ~x139 & n1079 ) ;
  assign n1121 = ( x86 & ~x129 ) | ( x86 & n1079 ) | ( ~x129 & n1079 ) ;
  assign n1122 = ~n1120 & n1121 ;
  assign n1123 = ( x129 & ~x140 ) | ( x129 & n1079 ) | ( ~x140 & n1079 ) ;
  assign n1124 = ( x87 & ~x129 ) | ( x87 & n1079 ) | ( ~x129 & n1079 ) ;
  assign n1125 = ~n1123 & n1124 ;
  assign n1126 = x136 & x137 ;
  assign n1127 = n1015 & n1126 ;
  assign n1128 = ( x129 & ~x139 ) | ( x129 & n1127 ) | ( ~x139 & n1127 ) ;
  assign n1129 = ( x88 & ~x129 ) | ( x88 & n1127 ) | ( ~x129 & n1127 ) ;
  assign n1130 = ~n1128 & n1129 ;
  assign n1131 = ( x129 & ~x140 ) | ( x129 & n1127 ) | ( ~x140 & n1127 ) ;
  assign n1132 = ( x89 & ~x129 ) | ( x89 & n1127 ) | ( ~x129 & n1127 ) ;
  assign n1133 = ~n1131 & n1132 ;
  assign n1134 = ( x129 & ~x142 ) | ( x129 & n1127 ) | ( ~x142 & n1127 ) ;
  assign n1135 = ( x90 & ~x129 ) | ( x90 & n1127 ) | ( ~x129 & n1127 ) ;
  assign n1136 = ~n1134 & n1135 ;
  assign n1137 = ( x129 & ~x143 ) | ( x129 & n1127 ) | ( ~x143 & n1127 ) ;
  assign n1138 = ( x91 & ~x129 ) | ( x91 & n1127 ) | ( ~x129 & n1127 ) ;
  assign n1139 = ~n1137 & n1138 ;
  assign n1140 = ( x129 & ~x144 ) | ( x129 & n1127 ) | ( ~x144 & n1127 ) ;
  assign n1141 = ( x92 & ~x129 ) | ( x92 & n1127 ) | ( ~x129 & n1127 ) ;
  assign n1142 = ~n1140 & n1141 ;
  assign n1143 = ( x129 & ~x146 ) | ( x129 & n1127 ) | ( ~x146 & n1127 ) ;
  assign n1144 = ( x93 & ~x129 ) | ( x93 & n1127 ) | ( ~x129 & n1127 ) ;
  assign n1145 = ~n1143 & n1144 ;
  assign n1146 = x138 & n1014 ;
  assign n1147 = x82 & ~n1035 ;
  assign n1148 = n1146 & n1147 ;
  assign n1149 = ( x129 & ~x142 ) | ( x129 & n1148 ) | ( ~x142 & n1148 ) ;
  assign n1150 = ( x94 & ~x129 ) | ( x94 & n1148 ) | ( ~x129 & n1148 ) ;
  assign n1151 = ~n1149 & n1150 ;
  assign n1152 = x3 | n1014 ;
  assign n1153 = x110 | n1152 ;
  assign n1154 = x138 & n1147 ;
  assign n1155 = n1014 & ~n1154 ;
  assign n1156 = n1153 & ~n1155 ;
  assign n1157 = x95 & ~n1156 ;
  assign n1158 = x143 & n1148 ;
  assign n1159 = n1157 | n1158 ;
  assign n1160 = ~x129 & n1159 ;
  assign n1161 = x96 & ~n1156 ;
  assign n1162 = x146 & n1148 ;
  assign n1163 = n1161 | n1162 ;
  assign n1164 = ~x129 & n1163 ;
  assign n1165 = x97 & ~n1156 ;
  assign n1166 = x145 & n1148 ;
  assign n1167 = n1165 | n1166 ;
  assign n1168 = ~x129 & n1167 ;
  assign n1169 = ( x129 & ~x145 ) | ( x129 & n1127 ) | ( ~x145 & n1127 ) ;
  assign n1170 = ( x98 & ~x129 ) | ( x98 & n1127 ) | ( ~x129 & n1127 ) ;
  assign n1171 = ~n1169 & n1170 ;
  assign n1172 = ( x129 & ~x141 ) | ( x129 & n1127 ) | ( ~x141 & n1127 ) ;
  assign n1173 = ( x99 & ~x129 ) | ( x99 & n1127 ) | ( ~x129 & n1127 ) ;
  assign n1174 = ~n1172 & n1173 ;
  assign n1175 = x100 & ~n1156 ;
  assign n1176 = x144 & n1148 ;
  assign n1177 = n1175 | n1176 ;
  assign n1178 = ~x129 & n1177 ;
  assign n1179 = ( ~x124 & x136 ) | ( ~x124 & x138 ) | ( x136 & x138 ) ;
  assign n1180 = ( x77 & x136 ) | ( x77 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1181 = n1179 | n1180 ;
  assign n1182 = ( x93 & x136 ) | ( x93 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1183 = ( ~x65 & x136 ) | ( ~x65 & x138 ) | ( x136 & x138 ) ;
  assign n1184 = n1182 & n1183 ;
  assign n1185 = n1181 & ~n1184 ;
  assign n1186 = x137 | n1185 ;
  assign n1187 = x37 & n1103 ;
  assign n1188 = ( ~x96 & x136 ) | ( ~x96 & x138 ) | ( x136 & x138 ) ;
  assign n1189 = ( x82 & ~x136 ) | ( x82 & x138 ) | ( ~x136 & x138 ) ;
  assign n1190 = ~n1188 & n1189 ;
  assign n1191 = n1187 | n1190 ;
  assign n1192 = x137 & n1191 ;
  assign n1193 = n1186 & ~n1192 ;
  assign n1194 = x91 & n1012 ;
  assign n1195 = x95 & n1078 ;
  assign n1196 = n1194 | n1195 ;
  assign n1197 = x138 & n1196 ;
  assign n1198 = ( x79 & x136 ) | ( x79 & x137 ) | ( x136 & x137 ) ;
  assign n1199 = ( x34 & ~x136 ) | ( x34 & x137 ) | ( ~x136 & x137 ) ;
  assign n1200 = n1198 & n1199 ;
  assign n1201 = ( x69 & x136 ) | ( x69 & x137 ) | ( x136 & x137 ) ;
  assign n1202 = ( x66 & ~x136 ) | ( x66 & x137 ) | ( ~x136 & x137 ) ;
  assign n1203 = n1201 | n1202 ;
  assign n1204 = ~n1200 & n1203 ;
  assign n1205 = x138 | n1204 ;
  assign n1206 = ~n1197 & n1205 ;
  assign n1207 = x90 & n1012 ;
  assign n1208 = x94 & n1078 ;
  assign n1209 = n1207 | n1208 ;
  assign n1210 = x138 & n1209 ;
  assign n1211 = ( x78 & x136 ) | ( x78 & x137 ) | ( x136 & x137 ) ;
  assign n1212 = ( x33 & ~x136 ) | ( x33 & x137 ) | ( ~x136 & x137 ) ;
  assign n1213 = n1211 & n1212 ;
  assign n1214 = ( x63 & x136 ) | ( x63 & x137 ) | ( x136 & x137 ) ;
  assign n1215 = ( x74 & ~x136 ) | ( x74 & x137 ) | ( ~x136 & x137 ) ;
  assign n1216 = n1214 | n1215 ;
  assign n1217 = ~n1213 & n1216 ;
  assign n1218 = x138 | n1217 ;
  assign n1219 = ~n1210 & n1218 ;
  assign n1220 = x99 & n1012 ;
  assign n1221 = ~x112 & n1078 ;
  assign n1222 = n1220 | n1221 ;
  assign n1223 = x138 & n1222 ;
  assign n1224 = ( x68 & x136 ) | ( x68 & x137 ) | ( x136 & x137 ) ;
  assign n1225 = ( x73 & ~x136 ) | ( x73 & x137 ) | ( ~x136 & x137 ) ;
  assign n1226 = n1224 | n1225 ;
  assign n1227 = ( x84 & x136 ) | ( x84 & x137 ) | ( x136 & x137 ) ;
  assign n1228 = ( x32 & ~x136 ) | ( x32 & x137 ) | ( ~x136 & x137 ) ;
  assign n1229 = n1227 & n1228 ;
  assign n1230 = n1226 & ~n1229 ;
  assign n1231 = x138 | n1230 ;
  assign n1232 = ~n1223 & n1231 ;
  assign n1233 = ( x92 & x136 ) | ( x92 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1234 = ( ~x70 & x136 ) | ( ~x70 & x138 ) | ( x136 & x138 ) ;
  assign n1235 = n1233 & n1234 ;
  assign n1236 = ( ~x125 & x136 ) | ( ~x125 & x138 ) | ( x136 & x138 ) ;
  assign n1237 = ( x75 & x136 ) | ( x75 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1238 = n1236 | n1237 ;
  assign n1239 = ~n1235 & n1238 ;
  assign n1240 = x137 | n1239 ;
  assign n1241 = x35 & n1103 ;
  assign n1242 = ( ~x100 & x136 ) | ( ~x100 & x138 ) | ( x136 & x138 ) ;
  assign n1243 = ( x80 & ~x136 ) | ( x80 & x138 ) | ( ~x136 & x138 ) ;
  assign n1244 = ~n1242 & n1243 ;
  assign n1245 = n1241 | n1244 ;
  assign n1246 = x137 & n1245 ;
  assign n1247 = n1240 & ~n1246 ;
  assign n1248 = ~n616 & n1114 ;
  assign n1249 = ~x27 & n1248 ;
  assign n1250 = n562 | n1249 ;
  assign n1251 = ~x129 & n1250 ;
  assign n1252 = ~x3 & n1251 ;
  assign n1253 = ( x98 & x136 ) | ( x98 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1254 = ( ~x71 & x136 ) | ( ~x71 & x138 ) | ( x136 & x138 ) ;
  assign n1255 = n1253 & n1254 ;
  assign n1256 = ( ~x23 & x136 ) | ( ~x23 & x138 ) | ( x136 & x138 ) ;
  assign n1257 = ( x76 & x136 ) | ( x76 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1258 = n1256 | n1257 ;
  assign n1259 = ~n1255 & n1258 ;
  assign n1260 = x137 | n1259 ;
  assign n1261 = x36 & n1103 ;
  assign n1262 = ( ~x97 & x136 ) | ( ~x97 & x138 ) | ( x136 & x138 ) ;
  assign n1263 = ( x81 & ~x136 ) | ( x81 & x138 ) | ( ~x136 & x138 ) ;
  assign n1264 = ~n1262 & n1263 ;
  assign n1265 = n1261 | n1264 ;
  assign n1266 = x137 & n1265 ;
  assign n1267 = n1260 & ~n1266 ;
  assign n1268 = ( x88 & x136 ) | ( x88 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1269 = ( ~x64 & x136 ) | ( ~x64 & x138 ) | ( x136 & x138 ) ;
  assign n1270 = n1268 & n1269 ;
  assign n1271 = ( ~x120 & x136 ) | ( ~x120 & x138 ) | ( x136 & x138 ) ;
  assign n1272 = ( x67 & x136 ) | ( x67 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1273 = n1271 | n1272 ;
  assign n1274 = ~n1270 & n1273 ;
  assign n1275 = x137 | n1274 ;
  assign n1276 = x30 & n1103 ;
  assign n1277 = ( ~x111 & x136 ) | ( ~x111 & x138 ) | ( x136 & x138 ) ;
  assign n1278 = ( x86 & ~x136 ) | ( x86 & x138 ) | ( ~x136 & x138 ) ;
  assign n1279 = ~n1277 & n1278 ;
  assign n1280 = n1276 | n1279 ;
  assign n1281 = x137 & n1280 ;
  assign n1282 = n1275 & ~n1281 ;
  assign n1283 = ( x26 & n618 ) | ( x26 & n624 ) | ( n618 & n624 ) ;
  assign n1284 = ~x129 & n1283 ;
  assign n1285 = ~x3 & n1284 ;
  assign n1286 = x116 & n1285 ;
  assign n1287 = ~x97 & n577 ;
  assign n1288 = n673 | n1287 ;
  assign n1289 = ~x129 & n1288 ;
  assign n1290 = ~x3 & n1289 ;
  assign n1291 = x116 & n1290 ;
  assign n1292 = x111 & ~n1154 ;
  assign n1293 = ~x137 & x138 ;
  assign n1294 = x82 & n1293 ;
  assign n1295 = n1027 & n1294 ;
  assign n1296 = n1292 | n1295 ;
  assign n1297 = n1014 & n1296 ;
  assign n1298 = ~x129 & n1297 ;
  assign n1299 = n1044 & n1294 ;
  assign n1300 = x112 | n1154 ;
  assign n1301 = ~n1299 & n1300 ;
  assign n1302 = n1014 & ~n1301 ;
  assign n1303 = ~x129 & n1302 ;
  assign n1304 = ( ~x54 & x113 ) | ( ~x54 & x129 ) | ( x113 & x129 ) ;
  assign n1305 = x11 | x22 ;
  assign n1306 = ( x54 & x129 ) | ( x54 & ~n1305 ) | ( x129 & ~n1305 ) ;
  assign n1307 = n1304 | n1306 ;
  assign n1308 = x3 | n1307 ;
  assign n1309 = n1018 & n1294 ;
  assign n1310 = x115 | n1154 ;
  assign n1311 = ~n1309 & n1310 ;
  assign n1312 = n1014 & ~n1311 ;
  assign n1313 = ~x129 & n1312 ;
  assign n1314 = x4 | x12 ;
  assign n1315 = x7 | x9 ;
  assign n1316 = n1314 | n1315 ;
  assign n1317 = ~x129 & n1316 ;
  assign n1318 = ~x3 & n1317 ;
  assign n1319 = x54 & n1318 ;
  assign n1320 = x122 & ~x129 ;
  assign n1321 = ~x54 & x118 ;
  assign n1322 = x54 & ~x59 ;
  assign n1323 = n395 & n1322 ;
  assign n1324 = n1321 | n1323 ;
  assign n1325 = ~x129 & n1324 ;
  assign n1326 = ~x129 & n551 ;
  assign n1327 = x110 | x120 ;
  assign n1328 = x3 | n1327 ;
  assign n1329 = ~x129 & n1328 ;
  assign n1330 = ~x111 & n1329 ;
  assign n1331 = x81 & x120 ;
  assign n1332 = ~x129 & n1331 ;
  assign n1333 = x129 | x134 ;
  assign n1334 = x129 | x135 ;
  assign n1335 = x57 & ~x129 ;
  assign n1336 = ~x96 & x125 ;
  assign n1337 = x3 | n1336 ;
  assign n1338 = ~x129 & n1337 ;
  assign n1339 = ~x126 & n1013 ;
  assign y0 = x108 ;
  assign y1 = x83 ;
  assign y2 = x104 ;
  assign y3 = x103 ;
  assign y4 = x102 ;
  assign y5 = x105 ;
  assign y6 = x107 ;
  assign y7 = x101 ;
  assign y8 = x126 ;
  assign y9 = x121 ;
  assign y10 = x1 ;
  assign y11 = x0 ;
  assign y12 = ~1'b0 ;
  assign y13 = x130 ;
  assign y14 = x128 ;
  assign y15 = n192 ;
  assign y16 = n228 ;
  assign y17 = ~n267 ;
  assign y18 = n278 ;
  assign y19 = n290 ;
  assign y20 = n304 ;
  assign y21 = n317 ;
  assign y22 = n332 ;
  assign y23 = n344 ;
  assign y24 = n357 ;
  assign y25 = n369 ;
  assign y26 = n380 ;
  assign y27 = n390 ;
  assign y28 = n402 ;
  assign y29 = n413 ;
  assign y30 = ~n438 ;
  assign y31 = n445 ;
  assign y32 = n459 ;
  assign y33 = n467 ;
  assign y34 = n474 ;
  assign y35 = ~n498 ;
  assign y36 = n508 ;
  assign y37 = n521 ;
  assign y38 = n524 ;
  assign y39 = ~n544 ;
  assign y40 = n588 ;
  assign y41 = n603 ;
  assign y42 = n617 ;
  assign y43 = n654 ;
  assign y44 = n685 ;
  assign y45 = n691 ;
  assign y46 = n697 ;
  assign y47 = n703 ;
  assign y48 = n709 ;
  assign y49 = n715 ;
  assign y50 = n721 ;
  assign y51 = n727 ;
  assign y52 = n733 ;
  assign y53 = ~n754 ;
  assign y54 = n762 ;
  assign y55 = ~n776 ;
  assign y56 = ~n790 ;
  assign y57 = ~n806 ;
  assign y58 = ~n820 ;
  assign y59 = ~n828 ;
  assign y60 = ~n847 ;
  assign y61 = ~n859 ;
  assign y62 = ~n870 ;
  assign y63 = ~n883 ;
  assign y64 = ~n902 ;
  assign y65 = ~n916 ;
  assign y66 = n919 ;
  assign y67 = n921 ;
  assign y68 = n934 ;
  assign y69 = ~n936 ;
  assign y70 = n939 ;
  assign y71 = n960 ;
  assign y72 = n976 ;
  assign y73 = n985 ;
  assign y74 = n1004 ;
  assign y75 = n1008 ;
  assign y76 = n1011 ;
  assign y77 = ~n1021 ;
  assign y78 = ~n1025 ;
  assign y79 = ~n1030 ;
  assign y80 = ~n1034 ;
  assign y81 = ~n1039 ;
  assign y82 = ~n1042 ;
  assign y83 = ~n1047 ;
  assign y84 = ~n1051 ;
  assign y85 = ~n1055 ;
  assign y86 = ~n1059 ;
  assign y87 = ~n1062 ;
  assign y88 = ~n1065 ;
  assign y89 = ~n1068 ;
  assign y90 = ~n1071 ;
  assign y91 = ~n1074 ;
  assign y92 = ~n1077 ;
  assign y93 = n1082 ;
  assign y94 = n1085 ;
  assign y95 = n1088 ;
  assign y96 = n1091 ;
  assign y97 = n1094 ;
  assign y98 = ~n1110 ;
  assign y99 = n1113 ;
  assign y100 = n1119 ;
  assign y101 = n1122 ;
  assign y102 = n1125 ;
  assign y103 = n1130 ;
  assign y104 = n1133 ;
  assign y105 = n1136 ;
  assign y106 = n1139 ;
  assign y107 = n1142 ;
  assign y108 = n1145 ;
  assign y109 = n1151 ;
  assign y110 = n1160 ;
  assign y111 = n1164 ;
  assign y112 = n1168 ;
  assign y113 = n1171 ;
  assign y114 = n1174 ;
  assign y115 = n1178 ;
  assign y116 = ~n1193 ;
  assign y117 = ~n1206 ;
  assign y118 = ~n1219 ;
  assign y119 = ~n1232 ;
  assign y120 = ~n1247 ;
  assign y121 = n1252 ;
  assign y122 = ~n1267 ;
  assign y123 = ~n1282 ;
  assign y124 = n1286 ;
  assign y125 = n1291 ;
  assign y126 = n1298 ;
  assign y127 = n1303 ;
  assign y128 = ~n1308 ;
  assign y129 = n937 ;
  assign y130 = n1313 ;
  assign y131 = n1319 ;
  assign y132 = ~n1320 ;
  assign y133 = n1325 ;
  assign y134 = n1326 ;
  assign y135 = n1330 ;
  assign y136 = n1332 ;
  assign y137 = n1333 ;
  assign y138 = n1334 ;
  assign y139 = n1335 ;
  assign y140 = n1338 ;
  assign y141 = n1339 ;
endmodule
