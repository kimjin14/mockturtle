module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 ;
  assign n513 = ~x259 & x387 ;
  assign n514 = x259 & ~x387 ;
  assign n515 = n513 & ~n514 ;
  assign n516 = x260 & ~x388 ;
  assign n517 = ( x388 & n515 ) | ( x388 & ~n516 ) | ( n515 & ~n516 ) ;
  assign n518 = ( ~x388 & n514 ) | ( ~x388 & n516 ) | ( n514 & n516 ) ;
  assign n519 = x256 & ~x384 ;
  assign n520 = x257 | n519 ;
  assign n521 = ~x257 & x385 ;
  assign n522 = ( x385 & ~n519 ) | ( x385 & n521 ) | ( ~n519 & n521 ) ;
  assign n523 = n520 & ~n522 ;
  assign n524 = ( x258 & ~x386 ) | ( x258 & n523 ) | ( ~x386 & n523 ) ;
  assign n525 = ( ~n517 & n518 ) | ( ~n517 & n524 ) | ( n518 & n524 ) ;
  assign n526 = ~x263 & x391 ;
  assign n527 = x262 & ~x390 ;
  assign n528 = ~n526 & n527 ;
  assign n529 = x263 & ~x391 ;
  assign n530 = x264 | n529 ;
  assign n531 = n528 | n530 ;
  assign n532 = ~x392 & n531 ;
  assign n533 = x264 & ~x392 ;
  assign n534 = ~x262 & x390 ;
  assign n535 = ( ~x263 & x391 ) | ( ~x263 & n534 ) | ( x391 & n534 ) ;
  assign n536 = ( x392 & ~n533 ) | ( x392 & n535 ) | ( ~n533 & n535 ) ;
  assign n537 = ( ~x259 & x386 ) | ( ~x259 & x387 ) | ( x386 & x387 ) ;
  assign n538 = ( x260 & x261 ) | ( x260 & ~x389 ) | ( x261 & ~x389 ) ;
  assign n539 = x261 & ~x389 ;
  assign n540 = ( ~n537 & n538 ) | ( ~n537 & n539 ) | ( n538 & n539 ) ;
  assign n541 = ( x258 & x259 ) | ( x258 & ~x387 ) | ( x259 & ~x387 ) ;
  assign n542 = ( n538 & n539 ) | ( n538 & n541 ) | ( n539 & n541 ) ;
  assign n543 = ( n523 & n540 ) | ( n523 & n542 ) | ( n540 & n542 ) ;
  assign n544 = ( n532 & ~n536 ) | ( n532 & n543 ) | ( ~n536 & n543 ) ;
  assign n545 = ~x261 & x389 ;
  assign n546 = ( ~n532 & n536 ) | ( ~n532 & n545 ) | ( n536 & n545 ) ;
  assign n547 = ( n525 & n544 ) | ( n525 & ~n546 ) | ( n544 & ~n546 ) ;
  assign n548 = x264 & n529 ;
  assign n549 = ( x264 & n528 ) | ( x264 & n548 ) | ( n528 & n548 ) ;
  assign n550 = x264 & ~x391 ;
  assign n551 = x263 & x264 ;
  assign n552 = ( ~n534 & n550 ) | ( ~n534 & n551 ) | ( n550 & n551 ) ;
  assign n553 = ( n543 & n549 ) | ( n543 & n552 ) | ( n549 & n552 ) ;
  assign n554 = ( ~n545 & n549 ) | ( ~n545 & n552 ) | ( n549 & n552 ) ;
  assign n555 = ( n525 & n553 ) | ( n525 & n554 ) | ( n553 & n554 ) ;
  assign n556 = n547 | n555 ;
  assign n557 = ~x271 & x399 ;
  assign n558 = x270 & ~x398 ;
  assign n559 = ~n557 & n558 ;
  assign n560 = x271 & ~x399 ;
  assign n561 = x272 & n560 ;
  assign n562 = ( x272 & n559 ) | ( x272 & n561 ) | ( n559 & n561 ) ;
  assign n563 = ~x270 & x398 ;
  assign n564 = x272 & ~x399 ;
  assign n565 = x271 & x272 ;
  assign n566 = ( ~n563 & n564 ) | ( ~n563 & n565 ) | ( n564 & n565 ) ;
  assign n567 = ~x268 & x396 ;
  assign n568 = x266 & ~x394 ;
  assign n569 = ~x267 & x395 ;
  assign n570 = n568 & ~n569 ;
  assign n571 = x267 & ~x395 ;
  assign n572 = ~n567 & n571 ;
  assign n573 = ( ~n567 & n570 ) | ( ~n567 & n572 ) | ( n570 & n572 ) ;
  assign n574 = ~x269 & x397 ;
  assign n575 = x268 & ~x396 ;
  assign n576 = ~n574 & n575 ;
  assign n577 = x269 & ~x397 ;
  assign n578 = n576 | n577 ;
  assign n579 = n574 & ~n577 ;
  assign n580 = ( n573 & n578 ) | ( n573 & ~n579 ) | ( n578 & ~n579 ) ;
  assign n581 = ( n562 & n566 ) | ( n562 & n580 ) | ( n566 & n580 ) ;
  assign n582 = ~n563 & n577 ;
  assign n583 = ( ~n557 & n559 ) | ( ~n557 & n582 ) | ( n559 & n582 ) ;
  assign n584 = n560 | n583 ;
  assign n585 = ~x266 & x394 ;
  assign n586 = ( ~x267 & x395 ) | ( ~x267 & n585 ) | ( x395 & n585 ) ;
  assign n587 = n567 | n574 ;
  assign n588 = ( ~n576 & n586 ) | ( ~n576 & n587 ) | ( n586 & n587 ) ;
  assign n589 = x272 & ~n588 ;
  assign n590 = ( n566 & n584 ) | ( n566 & n589 ) | ( n584 & n589 ) ;
  assign n591 = ( ~x393 & n581 ) | ( ~x393 & n590 ) | ( n581 & n590 ) ;
  assign n592 = ( x265 & n581 ) | ( x265 & n590 ) | ( n581 & n590 ) ;
  assign n593 = ( n556 & n591 ) | ( n556 & n592 ) | ( n591 & n592 ) ;
  assign n594 = ( ~x271 & x399 ) | ( ~x271 & n563 ) | ( x399 & n563 ) ;
  assign n595 = x272 & ~x400 ;
  assign n596 = ( x400 & n594 ) | ( x400 & ~n595 ) | ( n594 & ~n595 ) ;
  assign n597 = ( ~x400 & n560 ) | ( ~x400 & n595 ) | ( n560 & n595 ) ;
  assign n598 = ( ~x400 & n559 ) | ( ~x400 & n597 ) | ( n559 & n597 ) ;
  assign n599 = ( n580 & ~n596 ) | ( n580 & n598 ) | ( ~n596 & n598 ) ;
  assign n600 = ( x400 & n588 ) | ( x400 & ~n595 ) | ( n588 & ~n595 ) ;
  assign n601 = ( ~n584 & n596 ) | ( ~n584 & n600 ) | ( n596 & n600 ) ;
  assign n602 = ( x393 & ~n599 ) | ( x393 & n601 ) | ( ~n599 & n601 ) ;
  assign n603 = ( x265 & n599 ) | ( x265 & ~n601 ) | ( n599 & ~n601 ) ;
  assign n604 = ( n556 & ~n602 ) | ( n556 & n603 ) | ( ~n602 & n603 ) ;
  assign n605 = n593 | n604 ;
  assign n606 = ~x277 & x405 ;
  assign n607 = x276 & ~x404 ;
  assign n608 = ~n606 & n607 ;
  assign n609 = ~x274 & x402 ;
  assign n610 = ( ~x275 & x403 ) | ( ~x275 & n609 ) | ( x403 & n609 ) ;
  assign n611 = ~x276 & x404 ;
  assign n612 = n606 | n611 ;
  assign n613 = ( ~n608 & n610 ) | ( ~n608 & n612 ) | ( n610 & n612 ) ;
  assign n614 = ~x279 & x407 ;
  assign n615 = ~x278 & x406 ;
  assign n616 = x277 & ~x405 ;
  assign n617 = ~n615 & n616 ;
  assign n618 = x278 & ~x406 ;
  assign n619 = ~n614 & n618 ;
  assign n620 = ( ~n614 & n617 ) | ( ~n614 & n619 ) | ( n617 & n619 ) ;
  assign n621 = x279 & ~x407 ;
  assign n622 = x280 & ~x408 ;
  assign n623 = ( ~x408 & n621 ) | ( ~x408 & n622 ) | ( n621 & n622 ) ;
  assign n624 = ( ~x408 & n620 ) | ( ~x408 & n623 ) | ( n620 & n623 ) ;
  assign n625 = n615 & ~n618 ;
  assign n626 = n614 | n625 ;
  assign n627 = ( x408 & ~n623 ) | ( x408 & n626 ) | ( ~n623 & n626 ) ;
  assign n628 = ( n613 & ~n624 ) | ( n613 & n627 ) | ( ~n624 & n627 ) ;
  assign n629 = n614 & ~n621 ;
  assign n630 = ( ~n621 & n625 ) | ( ~n621 & n629 ) | ( n625 & n629 ) ;
  assign n631 = ( x408 & ~n622 ) | ( x408 & n630 ) | ( ~n622 & n630 ) ;
  assign n632 = ( ~x408 & n619 ) | ( ~x408 & n623 ) | ( n619 & n623 ) ;
  assign n633 = x274 & ~x402 ;
  assign n634 = ~x275 & x403 ;
  assign n635 = n633 & ~n634 ;
  assign n636 = x275 & ~x403 ;
  assign n637 = ~n611 & n636 ;
  assign n638 = ( ~n611 & n635 ) | ( ~n611 & n637 ) | ( n635 & n637 ) ;
  assign n639 = n608 | n616 ;
  assign n640 = n606 & ~n616 ;
  assign n641 = ( n638 & n639 ) | ( n638 & ~n640 ) | ( n639 & ~n640 ) ;
  assign n642 = ( ~n631 & n632 ) | ( ~n631 & n641 ) | ( n632 & n641 ) ;
  assign n643 = ( x401 & n628 ) | ( x401 & ~n642 ) | ( n628 & ~n642 ) ;
  assign n644 = ( x273 & ~n628 ) | ( x273 & n642 ) | ( ~n628 & n642 ) ;
  assign n645 = ( n605 & ~n643 ) | ( n605 & n644 ) | ( ~n643 & n644 ) ;
  assign n646 = x280 & ~n630 ;
  assign n647 = x280 & n621 ;
  assign n648 = ( x280 & n619 ) | ( x280 & n647 ) | ( n619 & n647 ) ;
  assign n649 = ( n641 & n646 ) | ( n641 & n648 ) | ( n646 & n648 ) ;
  assign n650 = ( x280 & n620 ) | ( x280 & n647 ) | ( n620 & n647 ) ;
  assign n651 = ( x280 & ~n626 ) | ( x280 & n647 ) | ( ~n626 & n647 ) ;
  assign n652 = ( ~n613 & n650 ) | ( ~n613 & n651 ) | ( n650 & n651 ) ;
  assign n653 = ( ~x401 & n649 ) | ( ~x401 & n652 ) | ( n649 & n652 ) ;
  assign n654 = ( x273 & n649 ) | ( x273 & n652 ) | ( n649 & n652 ) ;
  assign n655 = ( n605 & n653 ) | ( n605 & n654 ) | ( n653 & n654 ) ;
  assign n656 = n645 | n655 ;
  assign n657 = ~x304 & x432 ;
  assign n658 = ~x311 & x439 ;
  assign n659 = ~x310 & x438 ;
  assign n660 = n658 | n659 ;
  assign n661 = ~x309 & x437 ;
  assign n662 = ~x308 & x436 ;
  assign n663 = n661 | n662 ;
  assign n664 = n660 | n663 ;
  assign n665 = ~x305 & x433 ;
  assign n666 = ~x307 & x435 ;
  assign n667 = ~x306 & x434 ;
  assign n668 = n666 | n667 ;
  assign n669 = n665 | n668 ;
  assign n670 = n664 | n669 ;
  assign n671 = n657 | n670 ;
  assign n672 = ~x303 & x431 ;
  assign n673 = ~x302 & x430 ;
  assign n674 = n672 | n673 ;
  assign n675 = ~x300 & x428 ;
  assign n676 = ~x301 & x429 ;
  assign n677 = n675 | n676 ;
  assign n678 = n674 | n677 ;
  assign n679 = ~x299 & x427 ;
  assign n680 = ~x298 & x426 ;
  assign n681 = n679 | n680 ;
  assign n682 = ~x297 & x425 ;
  assign n683 = ~x296 & x424 ;
  assign n684 = n682 | n683 ;
  assign n685 = n681 | n684 ;
  assign n686 = n678 | n685 ;
  assign n687 = ~x288 & x416 ;
  assign n688 = ~x295 & x423 ;
  assign n689 = ~x294 & x422 ;
  assign n690 = n688 | n689 ;
  assign n691 = ~x292 & x420 ;
  assign n692 = ~x293 & x421 ;
  assign n693 = n691 | n692 ;
  assign n694 = n690 | n693 ;
  assign n695 = ~x289 & x417 ;
  assign n696 = ~x291 & x419 ;
  assign n697 = ~x290 & x418 ;
  assign n698 = n696 | n697 ;
  assign n699 = n695 | n698 ;
  assign n700 = n694 | n699 ;
  assign n701 = n687 | n700 ;
  assign n702 = ~x285 & x413 ;
  assign n703 = x284 & ~x412 ;
  assign n704 = ~n702 & n703 ;
  assign n705 = ~x282 & x410 ;
  assign n706 = ( ~x283 & x411 ) | ( ~x283 & n705 ) | ( x411 & n705 ) ;
  assign n707 = ~x284 & x412 ;
  assign n708 = n702 | n707 ;
  assign n709 = ( ~n704 & n706 ) | ( ~n704 & n708 ) | ( n706 & n708 ) ;
  assign n710 = ~x287 & x415 ;
  assign n711 = ~x286 & x414 ;
  assign n712 = x286 & ~x414 ;
  assign n713 = n711 & ~n712 ;
  assign n714 = n710 | n713 ;
  assign n715 = x285 & ~x413 ;
  assign n716 = ~n711 & n715 ;
  assign n717 = ~n710 & n712 ;
  assign n718 = ( ~n710 & n716 ) | ( ~n710 & n717 ) | ( n716 & n717 ) ;
  assign n719 = ( n709 & n714 ) | ( n709 & ~n718 ) | ( n714 & ~n718 ) ;
  assign n720 = x287 & ~x415 ;
  assign n721 = ( n701 & n719 ) | ( n701 & ~n720 ) | ( n719 & ~n720 ) ;
  assign n722 = n701 | n721 ;
  assign n723 = x294 & ~x422 ;
  assign n724 = ~n688 & n723 ;
  assign n725 = n694 & ~n724 ;
  assign n726 = x288 & ~x416 ;
  assign n727 = ( x289 & ~x417 ) | ( x289 & n726 ) | ( ~x417 & n726 ) ;
  assign n728 = x290 & ~x418 ;
  assign n729 = ~n697 & n728 ;
  assign n730 = ( ~n697 & n727 ) | ( ~n697 & n729 ) | ( n727 & n729 ) ;
  assign n731 = ( x291 & ~x419 ) | ( x291 & n730 ) | ( ~x419 & n730 ) ;
  assign n732 = ( n724 & ~n725 ) | ( n724 & n731 ) | ( ~n725 & n731 ) ;
  assign n733 = x292 & ~x420 ;
  assign n734 = ( x293 & ~x421 ) | ( x293 & n733 ) | ( ~x421 & n733 ) ;
  assign n735 = ( ~x295 & x423 ) | ( ~x295 & n689 ) | ( x423 & n689 ) ;
  assign n736 = x295 & ~x423 ;
  assign n737 = ( n734 & ~n735 ) | ( n734 & n736 ) | ( ~n735 & n736 ) ;
  assign n738 = ~n686 & n737 ;
  assign n739 = ( ~n686 & n732 ) | ( ~n686 & n738 ) | ( n732 & n738 ) ;
  assign n740 = ( n686 & n722 ) | ( n686 & ~n739 ) | ( n722 & ~n739 ) ;
  assign n741 = x296 & ~x424 ;
  assign n742 = ( x297 & ~x425 ) | ( x297 & n741 ) | ( ~x425 & n741 ) ;
  assign n743 = x298 & ~x426 ;
  assign n744 = ~n680 & n743 ;
  assign n745 = ( ~n680 & n742 ) | ( ~n680 & n744 ) | ( n742 & n744 ) ;
  assign n746 = ( x299 & ~x427 ) | ( x299 & n745 ) | ( ~x427 & n745 ) ;
  assign n747 = ~n678 & n746 ;
  assign n748 = x300 & ~x428 ;
  assign n749 = ( x301 & ~x429 ) | ( x301 & n748 ) | ( ~x429 & n748 ) ;
  assign n750 = ~n674 & n749 ;
  assign n751 = x303 & ~x431 ;
  assign n752 = x302 & ~x430 ;
  assign n753 = ~n672 & n752 ;
  assign n754 = n751 | n753 ;
  assign n755 = n750 | n754 ;
  assign n756 = n747 | n755 ;
  assign n757 = ~n671 & n756 ;
  assign n758 = ( n671 & n740 ) | ( n671 & ~n757 ) | ( n740 & ~n757 ) ;
  assign n759 = ~x319 & x447 ;
  assign n760 = ~x318 & x446 ;
  assign n761 = n759 | n760 ;
  assign n762 = ~x317 & x445 ;
  assign n763 = ~x316 & x444 ;
  assign n764 = n762 | n763 ;
  assign n765 = n761 | n764 ;
  assign n766 = ~x315 & x443 ;
  assign n767 = ~x314 & x442 ;
  assign n768 = n766 | n767 ;
  assign n769 = ~x313 & x441 ;
  assign n770 = ~x312 & x440 ;
  assign n771 = n769 | n770 ;
  assign n772 = n768 | n771 ;
  assign n773 = n765 | n772 ;
  assign n774 = x316 & ~x444 ;
  assign n775 = ( x317 & ~x445 ) | ( x317 & n774 ) | ( ~x445 & n774 ) ;
  assign n776 = ~n761 & n775 ;
  assign n777 = x318 & ~x446 ;
  assign n778 = ~n759 & n777 ;
  assign n779 = n776 | n778 ;
  assign n780 = n773 & ~n779 ;
  assign n781 = x319 & ~x447 ;
  assign n782 = x312 & ~x440 ;
  assign n783 = ( x313 & ~x441 ) | ( x313 & n782 ) | ( ~x441 & n782 ) ;
  assign n784 = x314 & ~x442 ;
  assign n785 = ~n767 & n784 ;
  assign n786 = ( ~n767 & n783 ) | ( ~n767 & n785 ) | ( n783 & n785 ) ;
  assign n787 = ( x315 & ~x443 ) | ( x315 & n786 ) | ( ~x443 & n786 ) ;
  assign n788 = n765 & ~n781 ;
  assign n789 = ( n781 & n787 ) | ( n781 & ~n788 ) | ( n787 & ~n788 ) ;
  assign n790 = n780 & ~n789 ;
  assign n791 = ~x327 & x455 ;
  assign n792 = x326 & ~x454 ;
  assign n793 = ~n791 & n792 ;
  assign n794 = ~x326 & x454 ;
  assign n795 = n791 | n794 ;
  assign n796 = ~x325 & x453 ;
  assign n797 = ~x324 & x452 ;
  assign n798 = n796 | n797 ;
  assign n799 = n795 | n798 ;
  assign n800 = ~x323 & x451 ;
  assign n801 = ~x322 & x450 ;
  assign n802 = n800 | n801 ;
  assign n803 = ~x321 & x449 ;
  assign n804 = ~x320 & x448 ;
  assign n805 = n803 | n804 ;
  assign n806 = n802 | n805 ;
  assign n807 = n799 | n806 ;
  assign n808 = x320 & ~x448 ;
  assign n809 = ( x321 & ~x449 ) | ( x321 & n808 ) | ( ~x449 & n808 ) ;
  assign n810 = x322 & ~x450 ;
  assign n811 = ~n801 & n810 ;
  assign n812 = ( ~n801 & n809 ) | ( ~n801 & n811 ) | ( n809 & n811 ) ;
  assign n813 = ( x323 & ~x451 ) | ( x323 & n812 ) | ( ~x451 & n812 ) ;
  assign n814 = ( n799 & n807 ) | ( n799 & ~n813 ) | ( n807 & ~n813 ) ;
  assign n815 = ~n793 & n814 ;
  assign n816 = ~x335 & x463 ;
  assign n817 = ~x334 & x462 ;
  assign n818 = n816 | n817 ;
  assign n819 = ~x333 & x461 ;
  assign n820 = ~x332 & x460 ;
  assign n821 = n819 | n820 ;
  assign n822 = n818 | n821 ;
  assign n823 = ~x331 & x459 ;
  assign n824 = ~x330 & x458 ;
  assign n825 = n823 | n824 ;
  assign n826 = ~x329 & x457 ;
  assign n827 = ~x328 & x456 ;
  assign n828 = n826 | n827 ;
  assign n829 = n825 | n828 ;
  assign n830 = x324 & ~x452 ;
  assign n831 = ( x325 & ~x453 ) | ( x325 & n830 ) | ( ~x453 & n830 ) ;
  assign n832 = ( ~x327 & x455 ) | ( ~x327 & n794 ) | ( x455 & n794 ) ;
  assign n833 = x327 & ~x455 ;
  assign n834 = ( n831 & ~n832 ) | ( n831 & n833 ) | ( ~n832 & n833 ) ;
  assign n835 = ~n829 & n834 ;
  assign n836 = x328 & ~x456 ;
  assign n837 = ( x329 & ~x457 ) | ( x329 & n836 ) | ( ~x457 & n836 ) ;
  assign n838 = x330 & ~x458 ;
  assign n839 = ~n824 & n838 ;
  assign n840 = ( ~n824 & n837 ) | ( ~n824 & n839 ) | ( n837 & n839 ) ;
  assign n841 = ( x331 & ~x459 ) | ( x331 & n840 ) | ( ~x459 & n840 ) ;
  assign n842 = ~n822 & n841 ;
  assign n843 = ( ~n822 & n835 ) | ( ~n822 & n842 ) | ( n835 & n842 ) ;
  assign n844 = n822 | n829 ;
  assign n845 = ( n822 & ~n841 ) | ( n822 & n844 ) | ( ~n841 & n844 ) ;
  assign n846 = ( n815 & ~n843 ) | ( n815 & n845 ) | ( ~n843 & n845 ) ;
  assign n847 = ~n793 & n799 ;
  assign n848 = ( n793 & n813 ) | ( n793 & ~n847 ) | ( n813 & ~n847 ) ;
  assign n849 = ( n843 & ~n845 ) | ( n843 & n848 ) | ( ~n845 & n848 ) ;
  assign n850 = ( n790 & n846 ) | ( n790 & ~n849 ) | ( n846 & ~n849 ) ;
  assign n851 = ~x343 & x471 ;
  assign n852 = ~x342 & x470 ;
  assign n853 = n851 | n852 ;
  assign n854 = ~x341 & x469 ;
  assign n855 = ~x340 & x468 ;
  assign n856 = n854 | n855 ;
  assign n857 = n853 | n856 ;
  assign n858 = ~x336 & x464 ;
  assign n859 = ~x339 & x467 ;
  assign n860 = ~x338 & x466 ;
  assign n861 = n859 | n860 ;
  assign n862 = ~x337 & x465 ;
  assign n863 = x335 & ~x463 ;
  assign n864 = ~n862 & n863 ;
  assign n865 = ~n861 & n864 ;
  assign n866 = ~n858 & n865 ;
  assign n867 = n858 | n862 ;
  assign n868 = n861 | n867 ;
  assign n869 = x332 & ~x460 ;
  assign n870 = ( ~x334 & x461 ) | ( ~x334 & x462 ) | ( x461 & x462 ) ;
  assign n871 = ( x333 & x334 ) | ( x333 & ~x462 ) | ( x334 & ~x462 ) ;
  assign n872 = ( n869 & ~n870 ) | ( n869 & n871 ) | ( ~n870 & n871 ) ;
  assign n873 = ~n816 & n872 ;
  assign n874 = ( n866 & ~n868 ) | ( n866 & n873 ) | ( ~n868 & n873 ) ;
  assign n875 = x336 & ~x464 ;
  assign n876 = ( x337 & ~x465 ) | ( x337 & n875 ) | ( ~x465 & n875 ) ;
  assign n877 = x338 & ~x466 ;
  assign n878 = ~n860 & n877 ;
  assign n879 = ( ~n860 & n876 ) | ( ~n860 & n878 ) | ( n876 & n878 ) ;
  assign n880 = ( x339 & ~x467 ) | ( x339 & n879 ) | ( ~x467 & n879 ) ;
  assign n881 = ~n857 & n880 ;
  assign n882 = ( ~n857 & n874 ) | ( ~n857 & n881 ) | ( n874 & n881 ) ;
  assign n883 = x343 & ~x471 ;
  assign n884 = x340 & ~x468 ;
  assign n885 = ( ~x342 & x469 ) | ( ~x342 & x470 ) | ( x469 & x470 ) ;
  assign n886 = ( x341 & x342 ) | ( x341 & ~x470 ) | ( x342 & ~x470 ) ;
  assign n887 = ( n884 & ~n885 ) | ( n884 & n886 ) | ( ~n885 & n886 ) ;
  assign n888 = n851 & ~n883 ;
  assign n889 = ( n883 & n887 ) | ( n883 & ~n888 ) | ( n887 & ~n888 ) ;
  assign n890 = n882 | n889 ;
  assign n891 = ~x351 & x479 ;
  assign n892 = x350 & ~x478 ;
  assign n893 = ~n891 & n892 ;
  assign n894 = ~x350 & x478 ;
  assign n895 = n891 | n894 ;
  assign n896 = ~x349 & x477 ;
  assign n897 = ~x348 & x476 ;
  assign n898 = n896 | n897 ;
  assign n899 = n895 | n898 ;
  assign n900 = ~x347 & x475 ;
  assign n901 = ~x346 & x474 ;
  assign n902 = n900 | n901 ;
  assign n903 = ~x345 & x473 ;
  assign n904 = ~x344 & x472 ;
  assign n905 = n903 | n904 ;
  assign n906 = n902 | n905 ;
  assign n907 = n899 | n906 ;
  assign n908 = x344 & ~x472 ;
  assign n909 = ( x345 & ~x473 ) | ( x345 & n908 ) | ( ~x473 & n908 ) ;
  assign n910 = x346 & ~x474 ;
  assign n911 = ~n901 & n910 ;
  assign n912 = ( ~n901 & n909 ) | ( ~n901 & n911 ) | ( n909 & n911 ) ;
  assign n913 = ( x347 & ~x475 ) | ( x347 & n912 ) | ( ~x475 & n912 ) ;
  assign n914 = ( n899 & n907 ) | ( n899 & ~n913 ) | ( n907 & ~n913 ) ;
  assign n915 = ~n893 & n914 ;
  assign n916 = ~x355 & x483 ;
  assign n917 = ~x354 & x482 ;
  assign n918 = n916 | n917 ;
  assign n919 = ~x352 & x480 ;
  assign n920 = ~x353 & x481 ;
  assign n921 = n919 | n920 ;
  assign n922 = n918 | n921 ;
  assign n923 = x351 & ~x479 ;
  assign n924 = n895 & ~n923 ;
  assign n925 = x348 & ~x476 ;
  assign n926 = ( x349 & ~x477 ) | ( x349 & n925 ) | ( ~x477 & n925 ) ;
  assign n927 = ( n923 & ~n924 ) | ( n923 & n926 ) | ( ~n924 & n926 ) ;
  assign n928 = ~n922 & n927 ;
  assign n929 = ( n915 & n922 ) | ( n915 & ~n928 ) | ( n922 & ~n928 ) ;
  assign n930 = ~n893 & n899 ;
  assign n931 = ( n893 & n913 ) | ( n893 & ~n930 ) | ( n913 & ~n930 ) ;
  assign n932 = ( ~n922 & n928 ) | ( ~n922 & n931 ) | ( n928 & n931 ) ;
  assign n933 = ( n890 & ~n929 ) | ( n890 & n932 ) | ( ~n929 & n932 ) ;
  assign n934 = ~n851 & n887 ;
  assign n935 = n857 | n868 ;
  assign n936 = ( n857 & ~n880 ) | ( n857 & n935 ) | ( ~n880 & n935 ) ;
  assign n937 = ~n934 & n936 ;
  assign n938 = n883 & ~n906 ;
  assign n939 = n913 | n938 ;
  assign n940 = ~n899 & n939 ;
  assign n941 = ( n914 & n937 ) | ( n914 & ~n940 ) | ( n937 & ~n940 ) ;
  assign n942 = ~n893 & n895 ;
  assign n943 = ( n893 & n926 ) | ( n893 & ~n942 ) | ( n926 & ~n942 ) ;
  assign n944 = n918 | n919 ;
  assign n945 = ~n920 & n923 ;
  assign n946 = ~n944 & n945 ;
  assign n947 = ( ~n922 & n943 ) | ( ~n922 & n946 ) | ( n943 & n946 ) ;
  assign n948 = ( n922 & n941 ) | ( n922 & ~n947 ) | ( n941 & ~n947 ) ;
  assign n949 = ( n850 & ~n933 ) | ( n850 & n948 ) | ( ~n933 & n948 ) ;
  assign n950 = x304 & ~x432 ;
  assign n951 = ( x305 & ~x433 ) | ( x305 & n950 ) | ( ~x433 & n950 ) ;
  assign n952 = x306 & ~x434 ;
  assign n953 = ~n667 & n952 ;
  assign n954 = ( ~n667 & n951 ) | ( ~n667 & n953 ) | ( n951 & n953 ) ;
  assign n955 = ( x307 & ~x435 ) | ( x307 & n954 ) | ( ~x435 & n954 ) ;
  assign n956 = ~n664 & n955 ;
  assign n957 = x308 & ~x436 ;
  assign n958 = ( x309 & ~x437 ) | ( x309 & n957 ) | ( ~x437 & n957 ) ;
  assign n959 = x310 & ~x438 ;
  assign n960 = ~n659 & n959 ;
  assign n961 = ( ~n659 & n958 ) | ( ~n659 & n960 ) | ( n958 & n960 ) ;
  assign n962 = ( x311 & ~x439 ) | ( x311 & n961 ) | ( ~x439 & n961 ) ;
  assign n963 = ~n773 & n962 ;
  assign n964 = ( ~n773 & n956 ) | ( ~n773 & n963 ) | ( n956 & n963 ) ;
  assign n965 = ~n765 & n787 ;
  assign n966 = n779 | n965 ;
  assign n967 = n964 | n966 ;
  assign n968 = n781 & ~n805 ;
  assign n969 = ~n802 & n968 ;
  assign n970 = n813 | n969 ;
  assign n971 = ( n793 & ~n847 ) | ( n793 & n970 ) | ( ~n847 & n970 ) ;
  assign n972 = ( n843 & ~n845 ) | ( n843 & n971 ) | ( ~n845 & n971 ) ;
  assign n973 = ( ~n846 & n967 ) | ( ~n846 & n972 ) | ( n967 & n972 ) ;
  assign n974 = ( n933 & ~n948 ) | ( n933 & n973 ) | ( ~n948 & n973 ) ;
  assign n975 = ( n758 & n949 ) | ( n758 & ~n974 ) | ( n949 & ~n974 ) ;
  assign n976 = x383 & ~x511 ;
  assign n977 = x382 & ~x510 ;
  assign n978 = ~n976 & n977 ;
  assign n979 = ~x382 & x510 ;
  assign n980 = x380 & ~x508 ;
  assign n981 = ( x381 & ~x509 ) | ( x381 & n980 ) | ( ~x509 & n980 ) ;
  assign n982 = ~n979 & n981 ;
  assign n983 = ( ~n976 & n978 ) | ( ~n976 & n982 ) | ( n978 & n982 ) ;
  assign n984 = ~x383 & x511 ;
  assign n985 = ~x381 & x509 ;
  assign n986 = n979 | n985 ;
  assign n987 = ~x380 & x508 ;
  assign n988 = n976 | n987 ;
  assign n989 = n986 | n988 ;
  assign n990 = ~n984 & n989 ;
  assign n991 = ~n983 & n990 ;
  assign n992 = x384 & n991 ;
  assign n993 = n978 | n984 ;
  assign n994 = n976 & ~n984 ;
  assign n995 = ( n982 & n993 ) | ( n982 & ~n994 ) | ( n993 & ~n994 ) ;
  assign n996 = x384 & ~n995 ;
  assign n997 = ~x359 & x487 ;
  assign n998 = x358 & ~x486 ;
  assign n999 = ~n997 & n998 ;
  assign n1000 = ~x358 & x486 ;
  assign n1001 = n997 | n1000 ;
  assign n1002 = ~x357 & x485 ;
  assign n1003 = ~x356 & x484 ;
  assign n1004 = n1002 | n1003 ;
  assign n1005 = n1001 | n1004 ;
  assign n1006 = ~n999 & n1005 ;
  assign n1007 = x352 & ~x480 ;
  assign n1008 = ( x353 & ~x481 ) | ( x353 & n1007 ) | ( ~x481 & n1007 ) ;
  assign n1009 = x354 & ~x482 ;
  assign n1010 = ~n917 & n1009 ;
  assign n1011 = ( ~n917 & n1008 ) | ( ~n917 & n1010 ) | ( n1008 & n1010 ) ;
  assign n1012 = ( x355 & ~x483 ) | ( x355 & n1011 ) | ( ~x483 & n1011 ) ;
  assign n1013 = ( n999 & ~n1006 ) | ( n999 & n1012 ) | ( ~n1006 & n1012 ) ;
  assign n1014 = x356 & ~x484 ;
  assign n1015 = ( x357 & ~x485 ) | ( x357 & n1014 ) | ( ~x485 & n1014 ) ;
  assign n1016 = ~n1001 & n1015 ;
  assign n1017 = x359 & ~x487 ;
  assign n1018 = n1016 | n1017 ;
  assign n1019 = n1013 | n1018 ;
  assign n1020 = ~x369 & x497 ;
  assign n1021 = ~x367 & x495 ;
  assign n1022 = ~x366 & x494 ;
  assign n1023 = n1021 | n1022 ;
  assign n1024 = x364 & ~x492 ;
  assign n1025 = ( x365 & ~x493 ) | ( x365 & n1024 ) | ( ~x493 & n1024 ) ;
  assign n1026 = ~n1023 & n1025 ;
  assign n1027 = x367 & ~x495 ;
  assign n1028 = x366 & ~x494 ;
  assign n1029 = ~n1021 & n1028 ;
  assign n1030 = n1027 | n1029 ;
  assign n1031 = n1026 | n1030 ;
  assign n1032 = ~n1020 & n1031 ;
  assign n1033 = ~x362 & x490 ;
  assign n1034 = x360 & ~x488 ;
  assign n1035 = ( x361 & ~x489 ) | ( x361 & n1034 ) | ( ~x489 & n1034 ) ;
  assign n1036 = x362 & ~x490 ;
  assign n1037 = ~n1033 & n1036 ;
  assign n1038 = ( ~n1033 & n1035 ) | ( ~n1033 & n1037 ) | ( n1035 & n1037 ) ;
  assign n1039 = ( x363 & ~x491 ) | ( x363 & n1038 ) | ( ~x491 & n1038 ) ;
  assign n1040 = ~x365 & x493 ;
  assign n1041 = ~x364 & x492 ;
  assign n1042 = n1040 | n1041 ;
  assign n1043 = n1023 | n1042 ;
  assign n1044 = ~x363 & x491 ;
  assign n1045 = n1033 | n1044 ;
  assign n1046 = ~x361 & x489 ;
  assign n1047 = ~x360 & x488 ;
  assign n1048 = n1046 | n1047 ;
  assign n1049 = n1045 | n1048 ;
  assign n1050 = n1043 | n1049 ;
  assign n1051 = ( ~n1039 & n1043 ) | ( ~n1039 & n1050 ) | ( n1043 & n1050 ) ;
  assign n1052 = ( n1020 & ~n1032 ) | ( n1020 & n1051 ) | ( ~n1032 & n1051 ) ;
  assign n1053 = n1039 & ~n1043 ;
  assign n1054 = ( ~n1020 & n1032 ) | ( ~n1020 & n1053 ) | ( n1032 & n1053 ) ;
  assign n1055 = ( n1019 & ~n1052 ) | ( n1019 & n1054 ) | ( ~n1052 & n1054 ) ;
  assign n1056 = ~x379 & x507 ;
  assign n1057 = ~x378 & x506 ;
  assign n1058 = n1056 | n1057 ;
  assign n1059 = ~x377 & x505 ;
  assign n1060 = ~x376 & x504 ;
  assign n1061 = n1059 | n1060 ;
  assign n1062 = n1058 | n1061 ;
  assign n1063 = x376 & ~x504 ;
  assign n1064 = ( x377 & ~x505 ) | ( x377 & n1063 ) | ( ~x505 & n1063 ) ;
  assign n1065 = x378 & ~x506 ;
  assign n1066 = ~n1057 & n1065 ;
  assign n1067 = ( ~n1057 & n1064 ) | ( ~n1057 & n1066 ) | ( n1064 & n1066 ) ;
  assign n1068 = ( x379 & ~x507 ) | ( x379 & n1067 ) | ( ~x507 & n1067 ) ;
  assign n1069 = n1062 & ~n1068 ;
  assign n1070 = ~x375 & x503 ;
  assign n1071 = ~x374 & x502 ;
  assign n1072 = n1070 | n1071 ;
  assign n1073 = ~x373 & x501 ;
  assign n1074 = ~x372 & x500 ;
  assign n1075 = n1073 | n1074 ;
  assign n1076 = n1072 | n1075 ;
  assign n1077 = ~x370 & x498 ;
  assign n1078 = x368 & ~x496 ;
  assign n1079 = ( x369 & ~x497 ) | ( x369 & n1078 ) | ( ~x497 & n1078 ) ;
  assign n1080 = x370 & ~x498 ;
  assign n1081 = ~n1077 & n1080 ;
  assign n1082 = ( ~n1077 & n1079 ) | ( ~n1077 & n1081 ) | ( n1079 & n1081 ) ;
  assign n1083 = ( x371 & ~x499 ) | ( x371 & n1082 ) | ( ~x499 & n1082 ) ;
  assign n1084 = ~x371 & x499 ;
  assign n1085 = n1077 | n1084 ;
  assign n1086 = ~x368 & x496 ;
  assign n1087 = n1085 | n1086 ;
  assign n1088 = n1076 | n1087 ;
  assign n1089 = ( n1076 & ~n1083 ) | ( n1076 & n1088 ) | ( ~n1083 & n1088 ) ;
  assign n1090 = x374 & ~x502 ;
  assign n1091 = ~n1070 & n1090 ;
  assign n1092 = x372 & ~x500 ;
  assign n1093 = ( x373 & ~x501 ) | ( x373 & n1092 ) | ( ~x501 & n1092 ) ;
  assign n1094 = ~n1072 & n1093 ;
  assign n1095 = n1091 | n1094 ;
  assign n1096 = n1089 & ~n1095 ;
  assign n1097 = x375 & ~x503 ;
  assign n1098 = ( n1068 & ~n1069 ) | ( n1068 & n1097 ) | ( ~n1069 & n1097 ) ;
  assign n1099 = ( n1069 & n1096 ) | ( n1069 & ~n1098 ) | ( n1096 & ~n1098 ) ;
  assign n1100 = n1076 & ~n1091 ;
  assign n1101 = ( n1083 & n1091 ) | ( n1083 & ~n1100 ) | ( n1091 & ~n1100 ) ;
  assign n1102 = n1094 | n1101 ;
  assign n1103 = ( ~n1069 & n1098 ) | ( ~n1069 & n1102 ) | ( n1098 & n1102 ) ;
  assign n1104 = ( n1055 & ~n1099 ) | ( n1055 & n1103 ) | ( ~n1099 & n1103 ) ;
  assign n1105 = ( n992 & n996 ) | ( n992 & ~n1104 ) | ( n996 & ~n1104 ) ;
  assign n1106 = ~n1039 & n1049 ;
  assign n1107 = ( n1017 & n1039 ) | ( n1017 & ~n1106 ) | ( n1039 & ~n1106 ) ;
  assign n1108 = ~n1029 & n1043 ;
  assign n1109 = ~n1026 & n1108 ;
  assign n1110 = n1026 | n1029 ;
  assign n1111 = ( n1106 & n1109 ) | ( n1106 & ~n1110 ) | ( n1109 & ~n1110 ) ;
  assign n1112 = n1006 & ~n1016 ;
  assign n1113 = ( n1109 & ~n1110 ) | ( n1109 & n1112 ) | ( ~n1110 & n1112 ) ;
  assign n1114 = ( ~n1107 & n1111 ) | ( ~n1107 & n1113 ) | ( n1111 & n1113 ) ;
  assign n1115 = ~n1027 & n1114 ;
  assign n1116 = n1094 | n1097 ;
  assign n1117 = ~n1062 & n1116 ;
  assign n1118 = n1068 | n1117 ;
  assign n1119 = ( ~n1069 & n1101 ) | ( ~n1069 & n1118 ) | ( n1101 & n1118 ) ;
  assign n1120 = ( n992 & n996 ) | ( n992 & ~n1119 ) | ( n996 & ~n1119 ) ;
  assign n1121 = n1020 | n1086 ;
  assign n1122 = n1085 | n1121 ;
  assign n1123 = n1076 | n1122 ;
  assign n1124 = ( n1076 & ~n1083 ) | ( n1076 & n1123 ) | ( ~n1083 & n1123 ) ;
  assign n1125 = ~n1091 & n1124 ;
  assign n1126 = ( n1069 & ~n1118 ) | ( n1069 & n1125 ) | ( ~n1118 & n1125 ) ;
  assign n1127 = ( n992 & n996 ) | ( n992 & n1126 ) | ( n996 & n1126 ) ;
  assign n1128 = ( n1115 & n1120 ) | ( n1115 & n1127 ) | ( n1120 & n1127 ) ;
  assign n1129 = ( n975 & n1105 ) | ( n975 & n1128 ) | ( n1105 & n1128 ) ;
  assign n1130 = n732 | n737 ;
  assign n1131 = n717 | n720 ;
  assign n1132 = x282 & ~x410 ;
  assign n1133 = ~x283 & x411 ;
  assign n1134 = n1132 & ~n1133 ;
  assign n1135 = x283 & ~x411 ;
  assign n1136 = ~n707 & n1135 ;
  assign n1137 = ( ~n707 & n1134 ) | ( ~n707 & n1136 ) | ( n1134 & n1136 ) ;
  assign n1138 = n704 | n715 ;
  assign n1139 = n702 & ~n715 ;
  assign n1140 = ( n1137 & n1138 ) | ( n1137 & ~n1139 ) | ( n1138 & ~n1139 ) ;
  assign n1141 = n710 & ~n720 ;
  assign n1142 = ( n713 & ~n720 ) | ( n713 & n1141 ) | ( ~n720 & n1141 ) ;
  assign n1143 = ( n1131 & n1140 ) | ( n1131 & ~n1142 ) | ( n1140 & ~n1142 ) ;
  assign n1144 = ~n701 & n1143 ;
  assign n1145 = n1130 | n1144 ;
  assign n1146 = n750 | n753 ;
  assign n1147 = n747 | n1146 ;
  assign n1148 = ( ~n671 & n751 ) | ( ~n671 & n1147 ) | ( n751 & n1147 ) ;
  assign n1149 = n686 & ~n1146 ;
  assign n1150 = ~n747 & n1149 ;
  assign n1151 = ( n671 & ~n751 ) | ( n671 & n1150 ) | ( ~n751 & n1150 ) ;
  assign n1152 = ( n1145 & n1148 ) | ( n1145 & ~n1151 ) | ( n1148 & ~n1151 ) ;
  assign n1153 = ~n671 & n1152 ;
  assign n1154 = ( ~n949 & n974 ) | ( ~n949 & n1153 ) | ( n974 & n1153 ) ;
  assign n1155 = ( n1105 & n1128 ) | ( n1105 & ~n1154 ) | ( n1128 & ~n1154 ) ;
  assign n1156 = ( x409 & n1129 ) | ( x409 & n1155 ) | ( n1129 & n1155 ) ;
  assign n1157 = ( ~x281 & n1129 ) | ( ~x281 & n1155 ) | ( n1129 & n1155 ) ;
  assign n1158 = ( ~n656 & n1156 ) | ( ~n656 & n1157 ) | ( n1156 & n1157 ) ;
  assign n1159 = x256 & ~n991 ;
  assign n1160 = x256 & n995 ;
  assign n1161 = ( n1104 & n1159 ) | ( n1104 & n1160 ) | ( n1159 & n1160 ) ;
  assign n1162 = ( n1119 & n1159 ) | ( n1119 & n1160 ) | ( n1159 & n1160 ) ;
  assign n1163 = ( ~n1126 & n1159 ) | ( ~n1126 & n1160 ) | ( n1159 & n1160 ) ;
  assign n1164 = ( ~n1115 & n1162 ) | ( ~n1115 & n1163 ) | ( n1162 & n1163 ) ;
  assign n1165 = ( ~n975 & n1161 ) | ( ~n975 & n1164 ) | ( n1161 & n1164 ) ;
  assign n1166 = ( n1154 & n1161 ) | ( n1154 & n1164 ) | ( n1161 & n1164 ) ;
  assign n1167 = ( ~x409 & n1165 ) | ( ~x409 & n1166 ) | ( n1165 & n1166 ) ;
  assign n1168 = ( x281 & n1165 ) | ( x281 & n1166 ) | ( n1165 & n1166 ) ;
  assign n1169 = ( n656 & n1167 ) | ( n656 & n1168 ) | ( n1167 & n1168 ) ;
  assign n1170 = n1158 | n1169 ;
  assign n1171 = x385 & n991 ;
  assign n1172 = x385 & ~n995 ;
  assign n1173 = ( ~n1104 & n1171 ) | ( ~n1104 & n1172 ) | ( n1171 & n1172 ) ;
  assign n1174 = ( ~n1119 & n1171 ) | ( ~n1119 & n1172 ) | ( n1171 & n1172 ) ;
  assign n1175 = ( n1126 & n1171 ) | ( n1126 & n1172 ) | ( n1171 & n1172 ) ;
  assign n1176 = ( n1115 & n1174 ) | ( n1115 & n1175 ) | ( n1174 & n1175 ) ;
  assign n1177 = ( n975 & n1173 ) | ( n975 & n1176 ) | ( n1173 & n1176 ) ;
  assign n1178 = ( ~n1154 & n1173 ) | ( ~n1154 & n1176 ) | ( n1173 & n1176 ) ;
  assign n1179 = ( x409 & n1177 ) | ( x409 & n1178 ) | ( n1177 & n1178 ) ;
  assign n1180 = ( ~x281 & n1177 ) | ( ~x281 & n1178 ) | ( n1177 & n1178 ) ;
  assign n1181 = ( ~n656 & n1179 ) | ( ~n656 & n1180 ) | ( n1179 & n1180 ) ;
  assign n1182 = x257 & ~n991 ;
  assign n1183 = x257 & n995 ;
  assign n1184 = ( n1104 & n1182 ) | ( n1104 & n1183 ) | ( n1182 & n1183 ) ;
  assign n1185 = ( n1119 & n1182 ) | ( n1119 & n1183 ) | ( n1182 & n1183 ) ;
  assign n1186 = ( ~n1126 & n1182 ) | ( ~n1126 & n1183 ) | ( n1182 & n1183 ) ;
  assign n1187 = ( ~n1115 & n1185 ) | ( ~n1115 & n1186 ) | ( n1185 & n1186 ) ;
  assign n1188 = ( ~n975 & n1184 ) | ( ~n975 & n1187 ) | ( n1184 & n1187 ) ;
  assign n1189 = ( n1154 & n1184 ) | ( n1154 & n1187 ) | ( n1184 & n1187 ) ;
  assign n1190 = ( ~x409 & n1188 ) | ( ~x409 & n1189 ) | ( n1188 & n1189 ) ;
  assign n1191 = ( x281 & n1188 ) | ( x281 & n1189 ) | ( n1188 & n1189 ) ;
  assign n1192 = ( n656 & n1190 ) | ( n656 & n1191 ) | ( n1190 & n1191 ) ;
  assign n1193 = n1181 | n1192 ;
  assign n1194 = ~x7 & x135 ;
  assign n1195 = x6 & ~x134 ;
  assign n1196 = ~n1194 & n1195 ;
  assign n1197 = x7 & ~x135 ;
  assign n1198 = x8 | n1197 ;
  assign n1199 = n1196 | n1198 ;
  assign n1200 = ~x136 & n1199 ;
  assign n1201 = x8 & ~x136 ;
  assign n1202 = ~x6 & x134 ;
  assign n1203 = ( ~x7 & x135 ) | ( ~x7 & n1202 ) | ( x135 & n1202 ) ;
  assign n1204 = ( x136 & ~n1201 ) | ( x136 & n1203 ) | ( ~n1201 & n1203 ) ;
  assign n1205 = x2 & ~x130 ;
  assign n1206 = x0 & ~x128 ;
  assign n1207 = ( x1 & ~x129 ) | ( x1 & n1206 ) | ( ~x129 & n1206 ) ;
  assign n1208 = ~x2 & x130 ;
  assign n1209 = ~n1205 & n1208 ;
  assign n1210 = ( n1205 & n1207 ) | ( n1205 & ~n1209 ) | ( n1207 & ~n1209 ) ;
  assign n1211 = ( x3 & x4 ) | ( x3 & ~x132 ) | ( x4 & ~x132 ) ;
  assign n1212 = ( x5 & ~x133 ) | ( x5 & n1211 ) | ( ~x133 & n1211 ) ;
  assign n1213 = ( ~x4 & x131 ) | ( ~x4 & x132 ) | ( x131 & x132 ) ;
  assign n1214 = ( ~x5 & x133 ) | ( ~x5 & n1213 ) | ( x133 & n1213 ) ;
  assign n1215 = ( n1210 & n1212 ) | ( n1210 & ~n1214 ) | ( n1212 & ~n1214 ) ;
  assign n1216 = ( n1200 & ~n1204 ) | ( n1200 & n1215 ) | ( ~n1204 & n1215 ) ;
  assign n1217 = x8 & n1197 ;
  assign n1218 = ( x8 & n1196 ) | ( x8 & n1217 ) | ( n1196 & n1217 ) ;
  assign n1219 = x8 & ~x135 ;
  assign n1220 = x7 & x8 ;
  assign n1221 = ( ~n1202 & n1219 ) | ( ~n1202 & n1220 ) | ( n1219 & n1220 ) ;
  assign n1222 = ( n1215 & n1218 ) | ( n1215 & n1221 ) | ( n1218 & n1221 ) ;
  assign n1223 = n1216 | n1222 ;
  assign n1224 = ~x15 & x143 ;
  assign n1225 = x14 & ~x142 ;
  assign n1226 = ~n1224 & n1225 ;
  assign n1227 = x15 & ~x143 ;
  assign n1228 = x16 & n1227 ;
  assign n1229 = ( x16 & n1226 ) | ( x16 & n1228 ) | ( n1226 & n1228 ) ;
  assign n1230 = ~x14 & x142 ;
  assign n1231 = x16 & ~x143 ;
  assign n1232 = x15 & x16 ;
  assign n1233 = ( ~n1230 & n1231 ) | ( ~n1230 & n1232 ) | ( n1231 & n1232 ) ;
  assign n1234 = ~x12 & x140 ;
  assign n1235 = x10 & ~x138 ;
  assign n1236 = ~x11 & x139 ;
  assign n1237 = n1235 & ~n1236 ;
  assign n1238 = x11 & ~x139 ;
  assign n1239 = ~n1234 & n1238 ;
  assign n1240 = ( ~n1234 & n1237 ) | ( ~n1234 & n1239 ) | ( n1237 & n1239 ) ;
  assign n1241 = ~x13 & x141 ;
  assign n1242 = x12 & ~x140 ;
  assign n1243 = ~n1241 & n1242 ;
  assign n1244 = x13 & ~x141 ;
  assign n1245 = n1243 | n1244 ;
  assign n1246 = n1241 & ~n1244 ;
  assign n1247 = ( n1240 & n1245 ) | ( n1240 & ~n1246 ) | ( n1245 & ~n1246 ) ;
  assign n1248 = ( n1229 & n1233 ) | ( n1229 & n1247 ) | ( n1233 & n1247 ) ;
  assign n1249 = ~n1230 & n1244 ;
  assign n1250 = ( ~n1224 & n1226 ) | ( ~n1224 & n1249 ) | ( n1226 & n1249 ) ;
  assign n1251 = n1227 | n1250 ;
  assign n1252 = ~x10 & x138 ;
  assign n1253 = ( ~x11 & x139 ) | ( ~x11 & n1252 ) | ( x139 & n1252 ) ;
  assign n1254 = n1234 | n1241 ;
  assign n1255 = ( ~n1243 & n1253 ) | ( ~n1243 & n1254 ) | ( n1253 & n1254 ) ;
  assign n1256 = x16 & ~n1255 ;
  assign n1257 = ( n1233 & n1251 ) | ( n1233 & n1256 ) | ( n1251 & n1256 ) ;
  assign n1258 = ( ~x137 & n1248 ) | ( ~x137 & n1257 ) | ( n1248 & n1257 ) ;
  assign n1259 = ( x9 & n1248 ) | ( x9 & n1257 ) | ( n1248 & n1257 ) ;
  assign n1260 = ( n1223 & n1258 ) | ( n1223 & n1259 ) | ( n1258 & n1259 ) ;
  assign n1261 = ( ~x15 & x143 ) | ( ~x15 & n1230 ) | ( x143 & n1230 ) ;
  assign n1262 = x16 & ~x144 ;
  assign n1263 = ( x144 & n1261 ) | ( x144 & ~n1262 ) | ( n1261 & ~n1262 ) ;
  assign n1264 = ( ~x144 & n1227 ) | ( ~x144 & n1262 ) | ( n1227 & n1262 ) ;
  assign n1265 = ( ~x144 & n1226 ) | ( ~x144 & n1264 ) | ( n1226 & n1264 ) ;
  assign n1266 = ( n1247 & ~n1263 ) | ( n1247 & n1265 ) | ( ~n1263 & n1265 ) ;
  assign n1267 = ( x144 & n1255 ) | ( x144 & ~n1262 ) | ( n1255 & ~n1262 ) ;
  assign n1268 = ( ~n1251 & n1263 ) | ( ~n1251 & n1267 ) | ( n1263 & n1267 ) ;
  assign n1269 = ( x137 & ~n1266 ) | ( x137 & n1268 ) | ( ~n1266 & n1268 ) ;
  assign n1270 = ( x9 & n1266 ) | ( x9 & ~n1268 ) | ( n1266 & ~n1268 ) ;
  assign n1271 = ( n1223 & ~n1269 ) | ( n1223 & n1270 ) | ( ~n1269 & n1270 ) ;
  assign n1272 = n1260 | n1271 ;
  assign n1273 = ~x21 & x149 ;
  assign n1274 = x20 & ~x148 ;
  assign n1275 = ~n1273 & n1274 ;
  assign n1276 = ~x18 & x146 ;
  assign n1277 = ( ~x19 & x147 ) | ( ~x19 & n1276 ) | ( x147 & n1276 ) ;
  assign n1278 = ~x20 & x148 ;
  assign n1279 = n1273 | n1278 ;
  assign n1280 = ( ~n1275 & n1277 ) | ( ~n1275 & n1279 ) | ( n1277 & n1279 ) ;
  assign n1281 = ~x23 & x151 ;
  assign n1282 = ~x22 & x150 ;
  assign n1283 = x21 & ~x149 ;
  assign n1284 = ~n1282 & n1283 ;
  assign n1285 = x22 & ~x150 ;
  assign n1286 = ~n1281 & n1285 ;
  assign n1287 = ( ~n1281 & n1284 ) | ( ~n1281 & n1286 ) | ( n1284 & n1286 ) ;
  assign n1288 = x23 & ~x151 ;
  assign n1289 = x24 & ~x152 ;
  assign n1290 = ( ~x152 & n1288 ) | ( ~x152 & n1289 ) | ( n1288 & n1289 ) ;
  assign n1291 = ( ~x152 & n1287 ) | ( ~x152 & n1290 ) | ( n1287 & n1290 ) ;
  assign n1292 = n1282 & ~n1285 ;
  assign n1293 = n1281 | n1292 ;
  assign n1294 = ( x152 & ~n1290 ) | ( x152 & n1293 ) | ( ~n1290 & n1293 ) ;
  assign n1295 = ( n1280 & ~n1291 ) | ( n1280 & n1294 ) | ( ~n1291 & n1294 ) ;
  assign n1296 = n1281 & ~n1288 ;
  assign n1297 = ( ~n1288 & n1292 ) | ( ~n1288 & n1296 ) | ( n1292 & n1296 ) ;
  assign n1298 = ( x152 & ~n1289 ) | ( x152 & n1297 ) | ( ~n1289 & n1297 ) ;
  assign n1299 = ( ~x152 & n1286 ) | ( ~x152 & n1290 ) | ( n1286 & n1290 ) ;
  assign n1300 = x18 & ~x146 ;
  assign n1301 = ~x19 & x147 ;
  assign n1302 = n1300 & ~n1301 ;
  assign n1303 = x19 & ~x147 ;
  assign n1304 = ~n1278 & n1303 ;
  assign n1305 = ( ~n1278 & n1302 ) | ( ~n1278 & n1304 ) | ( n1302 & n1304 ) ;
  assign n1306 = n1275 | n1283 ;
  assign n1307 = n1273 & ~n1283 ;
  assign n1308 = ( n1305 & n1306 ) | ( n1305 & ~n1307 ) | ( n1306 & ~n1307 ) ;
  assign n1309 = ( ~n1298 & n1299 ) | ( ~n1298 & n1308 ) | ( n1299 & n1308 ) ;
  assign n1310 = ( x145 & n1295 ) | ( x145 & ~n1309 ) | ( n1295 & ~n1309 ) ;
  assign n1311 = ( x17 & ~n1295 ) | ( x17 & n1309 ) | ( ~n1295 & n1309 ) ;
  assign n1312 = ( n1272 & ~n1310 ) | ( n1272 & n1311 ) | ( ~n1310 & n1311 ) ;
  assign n1313 = x24 & ~n1297 ;
  assign n1314 = x24 & n1288 ;
  assign n1315 = ( x24 & n1286 ) | ( x24 & n1314 ) | ( n1286 & n1314 ) ;
  assign n1316 = ( n1308 & n1313 ) | ( n1308 & n1315 ) | ( n1313 & n1315 ) ;
  assign n1317 = ( x24 & n1287 ) | ( x24 & n1314 ) | ( n1287 & n1314 ) ;
  assign n1318 = ( x24 & ~n1293 ) | ( x24 & n1314 ) | ( ~n1293 & n1314 ) ;
  assign n1319 = ( ~n1280 & n1317 ) | ( ~n1280 & n1318 ) | ( n1317 & n1318 ) ;
  assign n1320 = ( ~x145 & n1316 ) | ( ~x145 & n1319 ) | ( n1316 & n1319 ) ;
  assign n1321 = ( x17 & n1316 ) | ( x17 & n1319 ) | ( n1316 & n1319 ) ;
  assign n1322 = ( n1272 & n1320 ) | ( n1272 & n1321 ) | ( n1320 & n1321 ) ;
  assign n1323 = n1312 | n1322 ;
  assign n1324 = ( x25 & ~x153 ) | ( x25 & n1323 ) | ( ~x153 & n1323 ) ;
  assign n1325 = ~x48 & x176 ;
  assign n1326 = ~x55 & x183 ;
  assign n1327 = ~x54 & x182 ;
  assign n1328 = n1326 | n1327 ;
  assign n1329 = ~x53 & x181 ;
  assign n1330 = ~x52 & x180 ;
  assign n1331 = n1329 | n1330 ;
  assign n1332 = n1328 | n1331 ;
  assign n1333 = ~x49 & x177 ;
  assign n1334 = ~x51 & x179 ;
  assign n1335 = ~x50 & x178 ;
  assign n1336 = n1334 | n1335 ;
  assign n1337 = n1333 | n1336 ;
  assign n1338 = n1332 | n1337 ;
  assign n1339 = n1325 | n1338 ;
  assign n1340 = ~x47 & x175 ;
  assign n1341 = ~x46 & x174 ;
  assign n1342 = n1340 | n1341 ;
  assign n1343 = ~x44 & x172 ;
  assign n1344 = ~x45 & x173 ;
  assign n1345 = n1343 | n1344 ;
  assign n1346 = n1342 | n1345 ;
  assign n1347 = ~x43 & x171 ;
  assign n1348 = ~x42 & x170 ;
  assign n1349 = n1347 | n1348 ;
  assign n1350 = ~x41 & x169 ;
  assign n1351 = ~x40 & x168 ;
  assign n1352 = n1350 | n1351 ;
  assign n1353 = n1349 | n1352 ;
  assign n1354 = n1346 | n1353 ;
  assign n1355 = ~x32 & x160 ;
  assign n1356 = ~x39 & x167 ;
  assign n1357 = ~x38 & x166 ;
  assign n1358 = n1356 | n1357 ;
  assign n1359 = ~x36 & x164 ;
  assign n1360 = ~x37 & x165 ;
  assign n1361 = n1359 | n1360 ;
  assign n1362 = n1358 | n1361 ;
  assign n1363 = ~x33 & x161 ;
  assign n1364 = ~x35 & x163 ;
  assign n1365 = ~x34 & x162 ;
  assign n1366 = n1364 | n1365 ;
  assign n1367 = n1363 | n1366 ;
  assign n1368 = n1362 | n1367 ;
  assign n1369 = n1355 | n1368 ;
  assign n1370 = ~x29 & x157 ;
  assign n1371 = x28 & ~x156 ;
  assign n1372 = ~n1370 & n1371 ;
  assign n1373 = ~x26 & x154 ;
  assign n1374 = ( ~x27 & x155 ) | ( ~x27 & n1373 ) | ( x155 & n1373 ) ;
  assign n1375 = ~x28 & x156 ;
  assign n1376 = n1370 | n1375 ;
  assign n1377 = ( ~n1372 & n1374 ) | ( ~n1372 & n1376 ) | ( n1374 & n1376 ) ;
  assign n1378 = ~x31 & x159 ;
  assign n1379 = ~x30 & x158 ;
  assign n1380 = x30 & ~x158 ;
  assign n1381 = n1379 & ~n1380 ;
  assign n1382 = n1378 | n1381 ;
  assign n1383 = x29 & ~x157 ;
  assign n1384 = ~n1379 & n1383 ;
  assign n1385 = ~n1378 & n1380 ;
  assign n1386 = ( ~n1378 & n1384 ) | ( ~n1378 & n1385 ) | ( n1384 & n1385 ) ;
  assign n1387 = ( n1377 & n1382 ) | ( n1377 & ~n1386 ) | ( n1382 & ~n1386 ) ;
  assign n1388 = x31 & ~x159 ;
  assign n1389 = ( n1369 & n1387 ) | ( n1369 & ~n1388 ) | ( n1387 & ~n1388 ) ;
  assign n1390 = n1369 | n1389 ;
  assign n1391 = x38 & ~x166 ;
  assign n1392 = ~n1356 & n1391 ;
  assign n1393 = n1362 & ~n1392 ;
  assign n1394 = x32 & ~x160 ;
  assign n1395 = ( x33 & ~x161 ) | ( x33 & n1394 ) | ( ~x161 & n1394 ) ;
  assign n1396 = x34 & ~x162 ;
  assign n1397 = ~n1365 & n1396 ;
  assign n1398 = ( ~n1365 & n1395 ) | ( ~n1365 & n1397 ) | ( n1395 & n1397 ) ;
  assign n1399 = ( x35 & ~x163 ) | ( x35 & n1398 ) | ( ~x163 & n1398 ) ;
  assign n1400 = ( n1392 & ~n1393 ) | ( n1392 & n1399 ) | ( ~n1393 & n1399 ) ;
  assign n1401 = x36 & ~x164 ;
  assign n1402 = ( x37 & ~x165 ) | ( x37 & n1401 ) | ( ~x165 & n1401 ) ;
  assign n1403 = ( ~x39 & x167 ) | ( ~x39 & n1357 ) | ( x167 & n1357 ) ;
  assign n1404 = x39 & ~x167 ;
  assign n1405 = ( n1402 & ~n1403 ) | ( n1402 & n1404 ) | ( ~n1403 & n1404 ) ;
  assign n1406 = ~n1354 & n1405 ;
  assign n1407 = ( ~n1354 & n1400 ) | ( ~n1354 & n1406 ) | ( n1400 & n1406 ) ;
  assign n1408 = ( n1354 & n1390 ) | ( n1354 & ~n1407 ) | ( n1390 & ~n1407 ) ;
  assign n1409 = x40 & ~x168 ;
  assign n1410 = ( x41 & ~x169 ) | ( x41 & n1409 ) | ( ~x169 & n1409 ) ;
  assign n1411 = x42 & ~x170 ;
  assign n1412 = ~n1348 & n1411 ;
  assign n1413 = ( ~n1348 & n1410 ) | ( ~n1348 & n1412 ) | ( n1410 & n1412 ) ;
  assign n1414 = ( x43 & ~x171 ) | ( x43 & n1413 ) | ( ~x171 & n1413 ) ;
  assign n1415 = ~n1346 & n1414 ;
  assign n1416 = x44 & ~x172 ;
  assign n1417 = ( x45 & ~x173 ) | ( x45 & n1416 ) | ( ~x173 & n1416 ) ;
  assign n1418 = ~n1342 & n1417 ;
  assign n1419 = x47 & ~x175 ;
  assign n1420 = x46 & ~x174 ;
  assign n1421 = ~n1340 & n1420 ;
  assign n1422 = n1419 | n1421 ;
  assign n1423 = n1418 | n1422 ;
  assign n1424 = n1415 | n1423 ;
  assign n1425 = ~n1339 & n1424 ;
  assign n1426 = ( n1339 & n1408 ) | ( n1339 & ~n1425 ) | ( n1408 & ~n1425 ) ;
  assign n1427 = ~x63 & x191 ;
  assign n1428 = ~x62 & x190 ;
  assign n1429 = n1427 | n1428 ;
  assign n1430 = ~x61 & x189 ;
  assign n1431 = ~x60 & x188 ;
  assign n1432 = n1430 | n1431 ;
  assign n1433 = n1429 | n1432 ;
  assign n1434 = ~x59 & x187 ;
  assign n1435 = ~x58 & x186 ;
  assign n1436 = n1434 | n1435 ;
  assign n1437 = ~x57 & x185 ;
  assign n1438 = ~x56 & x184 ;
  assign n1439 = n1437 | n1438 ;
  assign n1440 = n1436 | n1439 ;
  assign n1441 = n1433 | n1440 ;
  assign n1442 = x60 & ~x188 ;
  assign n1443 = ( x61 & ~x189 ) | ( x61 & n1442 ) | ( ~x189 & n1442 ) ;
  assign n1444 = ~n1429 & n1443 ;
  assign n1445 = x62 & ~x190 ;
  assign n1446 = ~n1427 & n1445 ;
  assign n1447 = n1444 | n1446 ;
  assign n1448 = n1441 & ~n1447 ;
  assign n1449 = x63 & ~x191 ;
  assign n1450 = x56 & ~x184 ;
  assign n1451 = ( x57 & ~x185 ) | ( x57 & n1450 ) | ( ~x185 & n1450 ) ;
  assign n1452 = x58 & ~x186 ;
  assign n1453 = ~n1435 & n1452 ;
  assign n1454 = ( ~n1435 & n1451 ) | ( ~n1435 & n1453 ) | ( n1451 & n1453 ) ;
  assign n1455 = ( x59 & ~x187 ) | ( x59 & n1454 ) | ( ~x187 & n1454 ) ;
  assign n1456 = n1433 & ~n1449 ;
  assign n1457 = ( n1449 & n1455 ) | ( n1449 & ~n1456 ) | ( n1455 & ~n1456 ) ;
  assign n1458 = n1448 & ~n1457 ;
  assign n1459 = ~x71 & x199 ;
  assign n1460 = x70 & ~x198 ;
  assign n1461 = ~n1459 & n1460 ;
  assign n1462 = ~x70 & x198 ;
  assign n1463 = n1459 | n1462 ;
  assign n1464 = ~x69 & x197 ;
  assign n1465 = ~x68 & x196 ;
  assign n1466 = n1464 | n1465 ;
  assign n1467 = n1463 | n1466 ;
  assign n1468 = ~x67 & x195 ;
  assign n1469 = ~x66 & x194 ;
  assign n1470 = n1468 | n1469 ;
  assign n1471 = ~x65 & x193 ;
  assign n1472 = ~x64 & x192 ;
  assign n1473 = n1471 | n1472 ;
  assign n1474 = n1470 | n1473 ;
  assign n1475 = n1467 | n1474 ;
  assign n1476 = x64 & ~x192 ;
  assign n1477 = ( x65 & ~x193 ) | ( x65 & n1476 ) | ( ~x193 & n1476 ) ;
  assign n1478 = x66 & ~x194 ;
  assign n1479 = ~n1469 & n1478 ;
  assign n1480 = ( ~n1469 & n1477 ) | ( ~n1469 & n1479 ) | ( n1477 & n1479 ) ;
  assign n1481 = ( x67 & ~x195 ) | ( x67 & n1480 ) | ( ~x195 & n1480 ) ;
  assign n1482 = ( n1467 & n1475 ) | ( n1467 & ~n1481 ) | ( n1475 & ~n1481 ) ;
  assign n1483 = ~n1461 & n1482 ;
  assign n1484 = ~x79 & x207 ;
  assign n1485 = ~x78 & x206 ;
  assign n1486 = n1484 | n1485 ;
  assign n1487 = ~x77 & x205 ;
  assign n1488 = ~x76 & x204 ;
  assign n1489 = n1487 | n1488 ;
  assign n1490 = n1486 | n1489 ;
  assign n1491 = ~x75 & x203 ;
  assign n1492 = ~x74 & x202 ;
  assign n1493 = n1491 | n1492 ;
  assign n1494 = ~x73 & x201 ;
  assign n1495 = ~x72 & x200 ;
  assign n1496 = n1494 | n1495 ;
  assign n1497 = n1493 | n1496 ;
  assign n1498 = x68 & ~x196 ;
  assign n1499 = ( x69 & ~x197 ) | ( x69 & n1498 ) | ( ~x197 & n1498 ) ;
  assign n1500 = ( ~x71 & x199 ) | ( ~x71 & n1462 ) | ( x199 & n1462 ) ;
  assign n1501 = x71 & ~x199 ;
  assign n1502 = ( n1499 & ~n1500 ) | ( n1499 & n1501 ) | ( ~n1500 & n1501 ) ;
  assign n1503 = ~n1497 & n1502 ;
  assign n1504 = x72 & ~x200 ;
  assign n1505 = ( x73 & ~x201 ) | ( x73 & n1504 ) | ( ~x201 & n1504 ) ;
  assign n1506 = x74 & ~x202 ;
  assign n1507 = ~n1492 & n1506 ;
  assign n1508 = ( ~n1492 & n1505 ) | ( ~n1492 & n1507 ) | ( n1505 & n1507 ) ;
  assign n1509 = ( x75 & ~x203 ) | ( x75 & n1508 ) | ( ~x203 & n1508 ) ;
  assign n1510 = ~n1490 & n1509 ;
  assign n1511 = ( ~n1490 & n1503 ) | ( ~n1490 & n1510 ) | ( n1503 & n1510 ) ;
  assign n1512 = n1490 | n1497 ;
  assign n1513 = ( n1490 & ~n1509 ) | ( n1490 & n1512 ) | ( ~n1509 & n1512 ) ;
  assign n1514 = ( n1483 & ~n1511 ) | ( n1483 & n1513 ) | ( ~n1511 & n1513 ) ;
  assign n1515 = ~n1461 & n1467 ;
  assign n1516 = ( n1461 & n1481 ) | ( n1461 & ~n1515 ) | ( n1481 & ~n1515 ) ;
  assign n1517 = ( n1511 & ~n1513 ) | ( n1511 & n1516 ) | ( ~n1513 & n1516 ) ;
  assign n1518 = ( n1458 & n1514 ) | ( n1458 & ~n1517 ) | ( n1514 & ~n1517 ) ;
  assign n1519 = ~x87 & x215 ;
  assign n1520 = ~x86 & x214 ;
  assign n1521 = n1519 | n1520 ;
  assign n1522 = ~x85 & x213 ;
  assign n1523 = ~x84 & x212 ;
  assign n1524 = n1522 | n1523 ;
  assign n1525 = n1521 | n1524 ;
  assign n1526 = ~x80 & x208 ;
  assign n1527 = ~x83 & x211 ;
  assign n1528 = ~x82 & x210 ;
  assign n1529 = n1527 | n1528 ;
  assign n1530 = ~x81 & x209 ;
  assign n1531 = x79 & ~x207 ;
  assign n1532 = ~n1530 & n1531 ;
  assign n1533 = ~n1529 & n1532 ;
  assign n1534 = ~n1526 & n1533 ;
  assign n1535 = n1526 | n1530 ;
  assign n1536 = n1529 | n1535 ;
  assign n1537 = x76 & ~x204 ;
  assign n1538 = ( ~x78 & x205 ) | ( ~x78 & x206 ) | ( x205 & x206 ) ;
  assign n1539 = ( x77 & x78 ) | ( x77 & ~x206 ) | ( x78 & ~x206 ) ;
  assign n1540 = ( n1537 & ~n1538 ) | ( n1537 & n1539 ) | ( ~n1538 & n1539 ) ;
  assign n1541 = ~n1484 & n1540 ;
  assign n1542 = ( n1534 & ~n1536 ) | ( n1534 & n1541 ) | ( ~n1536 & n1541 ) ;
  assign n1543 = x80 & ~x208 ;
  assign n1544 = ( x81 & ~x209 ) | ( x81 & n1543 ) | ( ~x209 & n1543 ) ;
  assign n1545 = x82 & ~x210 ;
  assign n1546 = ~n1528 & n1545 ;
  assign n1547 = ( ~n1528 & n1544 ) | ( ~n1528 & n1546 ) | ( n1544 & n1546 ) ;
  assign n1548 = ( x83 & ~x211 ) | ( x83 & n1547 ) | ( ~x211 & n1547 ) ;
  assign n1549 = ~n1525 & n1548 ;
  assign n1550 = ( ~n1525 & n1542 ) | ( ~n1525 & n1549 ) | ( n1542 & n1549 ) ;
  assign n1551 = x87 & ~x215 ;
  assign n1552 = x84 & ~x212 ;
  assign n1553 = ( ~x86 & x213 ) | ( ~x86 & x214 ) | ( x213 & x214 ) ;
  assign n1554 = ( x85 & x86 ) | ( x85 & ~x214 ) | ( x86 & ~x214 ) ;
  assign n1555 = ( n1552 & ~n1553 ) | ( n1552 & n1554 ) | ( ~n1553 & n1554 ) ;
  assign n1556 = n1519 & ~n1551 ;
  assign n1557 = ( n1551 & n1555 ) | ( n1551 & ~n1556 ) | ( n1555 & ~n1556 ) ;
  assign n1558 = n1550 | n1557 ;
  assign n1559 = ~x95 & x223 ;
  assign n1560 = x94 & ~x222 ;
  assign n1561 = ~n1559 & n1560 ;
  assign n1562 = ~x94 & x222 ;
  assign n1563 = n1559 | n1562 ;
  assign n1564 = ~x93 & x221 ;
  assign n1565 = ~x92 & x220 ;
  assign n1566 = n1564 | n1565 ;
  assign n1567 = n1563 | n1566 ;
  assign n1568 = ~x91 & x219 ;
  assign n1569 = ~x90 & x218 ;
  assign n1570 = n1568 | n1569 ;
  assign n1571 = ~x89 & x217 ;
  assign n1572 = ~x88 & x216 ;
  assign n1573 = n1571 | n1572 ;
  assign n1574 = n1570 | n1573 ;
  assign n1575 = n1567 | n1574 ;
  assign n1576 = x88 & ~x216 ;
  assign n1577 = ( x89 & ~x217 ) | ( x89 & n1576 ) | ( ~x217 & n1576 ) ;
  assign n1578 = x90 & ~x218 ;
  assign n1579 = ~n1569 & n1578 ;
  assign n1580 = ( ~n1569 & n1577 ) | ( ~n1569 & n1579 ) | ( n1577 & n1579 ) ;
  assign n1581 = ( x91 & ~x219 ) | ( x91 & n1580 ) | ( ~x219 & n1580 ) ;
  assign n1582 = ( n1567 & n1575 ) | ( n1567 & ~n1581 ) | ( n1575 & ~n1581 ) ;
  assign n1583 = ~n1561 & n1582 ;
  assign n1584 = ~x99 & x227 ;
  assign n1585 = ~x98 & x226 ;
  assign n1586 = n1584 | n1585 ;
  assign n1587 = ~x96 & x224 ;
  assign n1588 = ~x97 & x225 ;
  assign n1589 = n1587 | n1588 ;
  assign n1590 = n1586 | n1589 ;
  assign n1591 = x95 & ~x223 ;
  assign n1592 = n1563 & ~n1591 ;
  assign n1593 = x92 & ~x220 ;
  assign n1594 = ( x93 & ~x221 ) | ( x93 & n1593 ) | ( ~x221 & n1593 ) ;
  assign n1595 = ( n1591 & ~n1592 ) | ( n1591 & n1594 ) | ( ~n1592 & n1594 ) ;
  assign n1596 = ~n1590 & n1595 ;
  assign n1597 = ( n1583 & n1590 ) | ( n1583 & ~n1596 ) | ( n1590 & ~n1596 ) ;
  assign n1598 = ~n1561 & n1567 ;
  assign n1599 = ( n1561 & n1581 ) | ( n1561 & ~n1598 ) | ( n1581 & ~n1598 ) ;
  assign n1600 = ( ~n1590 & n1596 ) | ( ~n1590 & n1599 ) | ( n1596 & n1599 ) ;
  assign n1601 = ( n1558 & ~n1597 ) | ( n1558 & n1600 ) | ( ~n1597 & n1600 ) ;
  assign n1602 = ~n1519 & n1555 ;
  assign n1603 = n1525 | n1536 ;
  assign n1604 = ( n1525 & ~n1548 ) | ( n1525 & n1603 ) | ( ~n1548 & n1603 ) ;
  assign n1605 = ~n1602 & n1604 ;
  assign n1606 = n1551 & ~n1574 ;
  assign n1607 = n1581 | n1606 ;
  assign n1608 = ~n1567 & n1607 ;
  assign n1609 = ( n1582 & n1605 ) | ( n1582 & ~n1608 ) | ( n1605 & ~n1608 ) ;
  assign n1610 = ~n1561 & n1563 ;
  assign n1611 = ( n1561 & n1594 ) | ( n1561 & ~n1610 ) | ( n1594 & ~n1610 ) ;
  assign n1612 = n1586 | n1587 ;
  assign n1613 = ~n1588 & n1591 ;
  assign n1614 = ~n1612 & n1613 ;
  assign n1615 = ( ~n1590 & n1611 ) | ( ~n1590 & n1614 ) | ( n1611 & n1614 ) ;
  assign n1616 = ( n1590 & n1609 ) | ( n1590 & ~n1615 ) | ( n1609 & ~n1615 ) ;
  assign n1617 = ( n1518 & ~n1601 ) | ( n1518 & n1616 ) | ( ~n1601 & n1616 ) ;
  assign n1618 = x48 & ~x176 ;
  assign n1619 = ( x49 & ~x177 ) | ( x49 & n1618 ) | ( ~x177 & n1618 ) ;
  assign n1620 = x50 & ~x178 ;
  assign n1621 = ~n1335 & n1620 ;
  assign n1622 = ( ~n1335 & n1619 ) | ( ~n1335 & n1621 ) | ( n1619 & n1621 ) ;
  assign n1623 = ( x51 & ~x179 ) | ( x51 & n1622 ) | ( ~x179 & n1622 ) ;
  assign n1624 = ~n1332 & n1623 ;
  assign n1625 = x52 & ~x180 ;
  assign n1626 = ( x53 & ~x181 ) | ( x53 & n1625 ) | ( ~x181 & n1625 ) ;
  assign n1627 = x54 & ~x182 ;
  assign n1628 = ~n1327 & n1627 ;
  assign n1629 = ( ~n1327 & n1626 ) | ( ~n1327 & n1628 ) | ( n1626 & n1628 ) ;
  assign n1630 = ( x55 & ~x183 ) | ( x55 & n1629 ) | ( ~x183 & n1629 ) ;
  assign n1631 = ~n1441 & n1630 ;
  assign n1632 = ( ~n1441 & n1624 ) | ( ~n1441 & n1631 ) | ( n1624 & n1631 ) ;
  assign n1633 = ~n1433 & n1455 ;
  assign n1634 = n1447 | n1633 ;
  assign n1635 = n1632 | n1634 ;
  assign n1636 = n1449 & ~n1473 ;
  assign n1637 = ~n1470 & n1636 ;
  assign n1638 = n1481 | n1637 ;
  assign n1639 = ( n1461 & ~n1515 ) | ( n1461 & n1638 ) | ( ~n1515 & n1638 ) ;
  assign n1640 = ( n1511 & ~n1513 ) | ( n1511 & n1639 ) | ( ~n1513 & n1639 ) ;
  assign n1641 = ( ~n1514 & n1635 ) | ( ~n1514 & n1640 ) | ( n1635 & n1640 ) ;
  assign n1642 = ( n1601 & ~n1616 ) | ( n1601 & n1641 ) | ( ~n1616 & n1641 ) ;
  assign n1643 = ( n1426 & n1617 ) | ( n1426 & ~n1642 ) | ( n1617 & ~n1642 ) ;
  assign n1644 = ~x103 & x231 ;
  assign n1645 = x102 & ~x230 ;
  assign n1646 = ~n1644 & n1645 ;
  assign n1647 = ~x102 & x230 ;
  assign n1648 = n1644 | n1647 ;
  assign n1649 = ~x101 & x229 ;
  assign n1650 = ~x100 & x228 ;
  assign n1651 = n1649 | n1650 ;
  assign n1652 = n1648 | n1651 ;
  assign n1653 = ~n1646 & n1652 ;
  assign n1654 = x96 & ~x224 ;
  assign n1655 = ( x97 & ~x225 ) | ( x97 & n1654 ) | ( ~x225 & n1654 ) ;
  assign n1656 = x98 & ~x226 ;
  assign n1657 = ~n1585 & n1656 ;
  assign n1658 = ( ~n1585 & n1655 ) | ( ~n1585 & n1657 ) | ( n1655 & n1657 ) ;
  assign n1659 = ( x99 & ~x227 ) | ( x99 & n1658 ) | ( ~x227 & n1658 ) ;
  assign n1660 = ( n1646 & ~n1653 ) | ( n1646 & n1659 ) | ( ~n1653 & n1659 ) ;
  assign n1661 = x100 & ~x228 ;
  assign n1662 = ( x101 & ~x229 ) | ( x101 & n1661 ) | ( ~x229 & n1661 ) ;
  assign n1663 = ~n1648 & n1662 ;
  assign n1664 = x103 & ~x231 ;
  assign n1665 = n1663 | n1664 ;
  assign n1666 = n1660 | n1665 ;
  assign n1667 = ~x113 & x241 ;
  assign n1668 = ~x111 & x239 ;
  assign n1669 = ~x110 & x238 ;
  assign n1670 = n1668 | n1669 ;
  assign n1671 = x108 & ~x236 ;
  assign n1672 = ( x109 & ~x237 ) | ( x109 & n1671 ) | ( ~x237 & n1671 ) ;
  assign n1673 = ~n1670 & n1672 ;
  assign n1674 = x111 & ~x239 ;
  assign n1675 = x110 & ~x238 ;
  assign n1676 = ~n1668 & n1675 ;
  assign n1677 = n1674 | n1676 ;
  assign n1678 = n1673 | n1677 ;
  assign n1679 = ~n1667 & n1678 ;
  assign n1680 = ~x106 & x234 ;
  assign n1681 = x104 & ~x232 ;
  assign n1682 = ( x105 & ~x233 ) | ( x105 & n1681 ) | ( ~x233 & n1681 ) ;
  assign n1683 = x106 & ~x234 ;
  assign n1684 = ~n1680 & n1683 ;
  assign n1685 = ( ~n1680 & n1682 ) | ( ~n1680 & n1684 ) | ( n1682 & n1684 ) ;
  assign n1686 = ( x107 & ~x235 ) | ( x107 & n1685 ) | ( ~x235 & n1685 ) ;
  assign n1687 = ~x109 & x237 ;
  assign n1688 = ~x108 & x236 ;
  assign n1689 = n1687 | n1688 ;
  assign n1690 = n1670 | n1689 ;
  assign n1691 = ~x107 & x235 ;
  assign n1692 = n1680 | n1691 ;
  assign n1693 = ~x105 & x233 ;
  assign n1694 = ~x104 & x232 ;
  assign n1695 = n1693 | n1694 ;
  assign n1696 = n1692 | n1695 ;
  assign n1697 = n1690 | n1696 ;
  assign n1698 = ( ~n1686 & n1690 ) | ( ~n1686 & n1697 ) | ( n1690 & n1697 ) ;
  assign n1699 = ( n1667 & ~n1679 ) | ( n1667 & n1698 ) | ( ~n1679 & n1698 ) ;
  assign n1700 = n1686 & ~n1690 ;
  assign n1701 = ( ~n1667 & n1679 ) | ( ~n1667 & n1700 ) | ( n1679 & n1700 ) ;
  assign n1702 = ( n1666 & ~n1699 ) | ( n1666 & n1701 ) | ( ~n1699 & n1701 ) ;
  assign n1703 = ~x123 & x251 ;
  assign n1704 = ~x122 & x250 ;
  assign n1705 = n1703 | n1704 ;
  assign n1706 = ~x121 & x249 ;
  assign n1707 = ~x120 & x248 ;
  assign n1708 = n1706 | n1707 ;
  assign n1709 = n1705 | n1708 ;
  assign n1710 = x120 & ~x248 ;
  assign n1711 = ( x121 & ~x249 ) | ( x121 & n1710 ) | ( ~x249 & n1710 ) ;
  assign n1712 = x122 & ~x250 ;
  assign n1713 = ~n1704 & n1712 ;
  assign n1714 = ( ~n1704 & n1711 ) | ( ~n1704 & n1713 ) | ( n1711 & n1713 ) ;
  assign n1715 = ( x123 & ~x251 ) | ( x123 & n1714 ) | ( ~x251 & n1714 ) ;
  assign n1716 = n1709 & ~n1715 ;
  assign n1717 = ~x119 & x247 ;
  assign n1718 = ~x118 & x246 ;
  assign n1719 = n1717 | n1718 ;
  assign n1720 = ~x117 & x245 ;
  assign n1721 = ~x116 & x244 ;
  assign n1722 = n1720 | n1721 ;
  assign n1723 = n1719 | n1722 ;
  assign n1724 = ~x114 & x242 ;
  assign n1725 = x112 & ~x240 ;
  assign n1726 = ( x113 & ~x241 ) | ( x113 & n1725 ) | ( ~x241 & n1725 ) ;
  assign n1727 = x114 & ~x242 ;
  assign n1728 = ~n1724 & n1727 ;
  assign n1729 = ( ~n1724 & n1726 ) | ( ~n1724 & n1728 ) | ( n1726 & n1728 ) ;
  assign n1730 = ( x115 & ~x243 ) | ( x115 & n1729 ) | ( ~x243 & n1729 ) ;
  assign n1731 = ~x115 & x243 ;
  assign n1732 = n1724 | n1731 ;
  assign n1733 = ~x112 & x240 ;
  assign n1734 = n1732 | n1733 ;
  assign n1735 = n1723 | n1734 ;
  assign n1736 = ( n1723 & ~n1730 ) | ( n1723 & n1735 ) | ( ~n1730 & n1735 ) ;
  assign n1737 = x118 & ~x246 ;
  assign n1738 = ~n1717 & n1737 ;
  assign n1739 = x116 & ~x244 ;
  assign n1740 = ( x117 & ~x245 ) | ( x117 & n1739 ) | ( ~x245 & n1739 ) ;
  assign n1741 = ~n1719 & n1740 ;
  assign n1742 = n1738 | n1741 ;
  assign n1743 = n1736 & ~n1742 ;
  assign n1744 = x119 & ~x247 ;
  assign n1745 = ( n1715 & ~n1716 ) | ( n1715 & n1744 ) | ( ~n1716 & n1744 ) ;
  assign n1746 = ( n1716 & n1743 ) | ( n1716 & ~n1745 ) | ( n1743 & ~n1745 ) ;
  assign n1747 = n1723 & ~n1738 ;
  assign n1748 = ( n1730 & n1738 ) | ( n1730 & ~n1747 ) | ( n1738 & ~n1747 ) ;
  assign n1749 = n1741 | n1748 ;
  assign n1750 = ( ~n1716 & n1745 ) | ( ~n1716 & n1749 ) | ( n1745 & n1749 ) ;
  assign n1751 = ( n1702 & ~n1746 ) | ( n1702 & n1750 ) | ( ~n1746 & n1750 ) ;
  assign n1752 = x127 & ~x255 ;
  assign n1753 = x126 & ~x254 ;
  assign n1754 = ~n1752 & n1753 ;
  assign n1755 = ~x126 & x254 ;
  assign n1756 = x124 & ~x252 ;
  assign n1757 = ( x125 & ~x253 ) | ( x125 & n1756 ) | ( ~x253 & n1756 ) ;
  assign n1758 = ~n1755 & n1757 ;
  assign n1759 = ( ~n1752 & n1754 ) | ( ~n1752 & n1758 ) | ( n1754 & n1758 ) ;
  assign n1760 = ~x127 & x255 ;
  assign n1761 = ~x125 & x253 ;
  assign n1762 = n1755 | n1761 ;
  assign n1763 = ~x124 & x252 ;
  assign n1764 = n1752 | n1763 ;
  assign n1765 = n1762 | n1764 ;
  assign n1766 = ~n1760 & n1765 ;
  assign n1767 = ~n1759 & n1766 ;
  assign n1768 = x128 & n1767 ;
  assign n1769 = n1754 | n1760 ;
  assign n1770 = n1752 & ~n1760 ;
  assign n1771 = ( n1758 & n1769 ) | ( n1758 & ~n1770 ) | ( n1769 & ~n1770 ) ;
  assign n1772 = x128 & ~n1771 ;
  assign n1773 = ( ~n1751 & n1768 ) | ( ~n1751 & n1772 ) | ( n1768 & n1772 ) ;
  assign n1774 = ~n1686 & n1696 ;
  assign n1775 = ( n1664 & n1686 ) | ( n1664 & ~n1774 ) | ( n1686 & ~n1774 ) ;
  assign n1776 = ~n1676 & n1690 ;
  assign n1777 = ~n1673 & n1776 ;
  assign n1778 = n1673 | n1676 ;
  assign n1779 = ( n1774 & n1777 ) | ( n1774 & ~n1778 ) | ( n1777 & ~n1778 ) ;
  assign n1780 = n1653 & ~n1663 ;
  assign n1781 = ( n1777 & ~n1778 ) | ( n1777 & n1780 ) | ( ~n1778 & n1780 ) ;
  assign n1782 = ( ~n1775 & n1779 ) | ( ~n1775 & n1781 ) | ( n1779 & n1781 ) ;
  assign n1783 = ~n1674 & n1782 ;
  assign n1784 = n1741 | n1744 ;
  assign n1785 = ~n1709 & n1784 ;
  assign n1786 = n1715 | n1785 ;
  assign n1787 = ( ~n1716 & n1748 ) | ( ~n1716 & n1786 ) | ( n1748 & n1786 ) ;
  assign n1788 = ( n1768 & n1772 ) | ( n1768 & ~n1787 ) | ( n1772 & ~n1787 ) ;
  assign n1789 = n1667 | n1733 ;
  assign n1790 = n1732 | n1789 ;
  assign n1791 = n1723 | n1790 ;
  assign n1792 = ( n1723 & ~n1730 ) | ( n1723 & n1791 ) | ( ~n1730 & n1791 ) ;
  assign n1793 = ~n1738 & n1792 ;
  assign n1794 = ( n1716 & ~n1786 ) | ( n1716 & n1793 ) | ( ~n1786 & n1793 ) ;
  assign n1795 = ( n1768 & n1772 ) | ( n1768 & n1794 ) | ( n1772 & n1794 ) ;
  assign n1796 = ( n1783 & n1788 ) | ( n1783 & n1795 ) | ( n1788 & n1795 ) ;
  assign n1797 = ( n1643 & n1773 ) | ( n1643 & n1796 ) | ( n1773 & n1796 ) ;
  assign n1798 = n1400 | n1405 ;
  assign n1799 = n1385 | n1388 ;
  assign n1800 = x26 & ~x154 ;
  assign n1801 = ~x27 & x155 ;
  assign n1802 = n1800 & ~n1801 ;
  assign n1803 = x27 & ~x155 ;
  assign n1804 = ~n1375 & n1803 ;
  assign n1805 = ( ~n1375 & n1802 ) | ( ~n1375 & n1804 ) | ( n1802 & n1804 ) ;
  assign n1806 = n1372 | n1383 ;
  assign n1807 = n1370 & ~n1383 ;
  assign n1808 = ( n1805 & n1806 ) | ( n1805 & ~n1807 ) | ( n1806 & ~n1807 ) ;
  assign n1809 = n1378 & ~n1388 ;
  assign n1810 = ( n1381 & ~n1388 ) | ( n1381 & n1809 ) | ( ~n1388 & n1809 ) ;
  assign n1811 = ( n1799 & n1808 ) | ( n1799 & ~n1810 ) | ( n1808 & ~n1810 ) ;
  assign n1812 = ~n1369 & n1811 ;
  assign n1813 = n1798 | n1812 ;
  assign n1814 = n1418 | n1421 ;
  assign n1815 = n1415 | n1814 ;
  assign n1816 = ( ~n1339 & n1419 ) | ( ~n1339 & n1815 ) | ( n1419 & n1815 ) ;
  assign n1817 = n1354 & ~n1814 ;
  assign n1818 = ~n1415 & n1817 ;
  assign n1819 = ( n1339 & ~n1419 ) | ( n1339 & n1818 ) | ( ~n1419 & n1818 ) ;
  assign n1820 = ( n1813 & n1816 ) | ( n1813 & ~n1819 ) | ( n1816 & ~n1819 ) ;
  assign n1821 = ~n1339 & n1820 ;
  assign n1822 = ( ~n1617 & n1642 ) | ( ~n1617 & n1821 ) | ( n1642 & n1821 ) ;
  assign n1823 = ( n1773 & n1796 ) | ( n1773 & ~n1822 ) | ( n1796 & ~n1822 ) ;
  assign n1824 = ( ~n1324 & n1797 ) | ( ~n1324 & n1823 ) | ( n1797 & n1823 ) ;
  assign n1825 = x0 & ~n1767 ;
  assign n1826 = x0 & n1771 ;
  assign n1827 = ( n1751 & n1825 ) | ( n1751 & n1826 ) | ( n1825 & n1826 ) ;
  assign n1828 = ( n1787 & n1825 ) | ( n1787 & n1826 ) | ( n1825 & n1826 ) ;
  assign n1829 = ( ~n1794 & n1825 ) | ( ~n1794 & n1826 ) | ( n1825 & n1826 ) ;
  assign n1830 = ( ~n1783 & n1828 ) | ( ~n1783 & n1829 ) | ( n1828 & n1829 ) ;
  assign n1831 = ( ~n1643 & n1827 ) | ( ~n1643 & n1830 ) | ( n1827 & n1830 ) ;
  assign n1832 = ( n1822 & n1827 ) | ( n1822 & n1830 ) | ( n1827 & n1830 ) ;
  assign n1833 = ( n1324 & n1831 ) | ( n1324 & n1832 ) | ( n1831 & n1832 ) ;
  assign n1834 = n1824 | n1833 ;
  assign n1835 = ~n1170 & n1834 ;
  assign n1836 = n1193 & ~n1835 ;
  assign n1837 = x129 & n1767 ;
  assign n1838 = x129 & ~n1771 ;
  assign n1839 = ( ~n1751 & n1837 ) | ( ~n1751 & n1838 ) | ( n1837 & n1838 ) ;
  assign n1840 = ( ~n1787 & n1837 ) | ( ~n1787 & n1838 ) | ( n1837 & n1838 ) ;
  assign n1841 = ( n1794 & n1837 ) | ( n1794 & n1838 ) | ( n1837 & n1838 ) ;
  assign n1842 = ( n1783 & n1840 ) | ( n1783 & n1841 ) | ( n1840 & n1841 ) ;
  assign n1843 = ( n1643 & n1839 ) | ( n1643 & n1842 ) | ( n1839 & n1842 ) ;
  assign n1844 = ( ~n1822 & n1839 ) | ( ~n1822 & n1842 ) | ( n1839 & n1842 ) ;
  assign n1845 = ( ~n1324 & n1843 ) | ( ~n1324 & n1844 ) | ( n1843 & n1844 ) ;
  assign n1846 = x1 & ~n1767 ;
  assign n1847 = x1 & n1771 ;
  assign n1848 = ( n1751 & n1846 ) | ( n1751 & n1847 ) | ( n1846 & n1847 ) ;
  assign n1849 = ( n1787 & n1846 ) | ( n1787 & n1847 ) | ( n1846 & n1847 ) ;
  assign n1850 = ( ~n1794 & n1846 ) | ( ~n1794 & n1847 ) | ( n1846 & n1847 ) ;
  assign n1851 = ( ~n1783 & n1849 ) | ( ~n1783 & n1850 ) | ( n1849 & n1850 ) ;
  assign n1852 = ( ~n1643 & n1848 ) | ( ~n1643 & n1851 ) | ( n1848 & n1851 ) ;
  assign n1853 = ( n1822 & n1848 ) | ( n1822 & n1851 ) | ( n1848 & n1851 ) ;
  assign n1854 = ( n1324 & n1852 ) | ( n1324 & n1853 ) | ( n1852 & n1853 ) ;
  assign n1855 = n1845 | n1854 ;
  assign n1856 = n1193 & ~n1855 ;
  assign n1857 = ( n1835 & n1855 ) | ( n1835 & ~n1856 ) | ( n1855 & ~n1856 ) ;
  assign n1858 = ~n1836 & n1857 ;
  assign n1859 = x388 & n991 ;
  assign n1860 = x388 & ~n995 ;
  assign n1861 = ( ~n1104 & n1859 ) | ( ~n1104 & n1860 ) | ( n1859 & n1860 ) ;
  assign n1862 = ( ~n1119 & n1859 ) | ( ~n1119 & n1860 ) | ( n1859 & n1860 ) ;
  assign n1863 = ( n1126 & n1859 ) | ( n1126 & n1860 ) | ( n1859 & n1860 ) ;
  assign n1864 = ( n1115 & n1862 ) | ( n1115 & n1863 ) | ( n1862 & n1863 ) ;
  assign n1865 = ( n975 & n1861 ) | ( n975 & n1864 ) | ( n1861 & n1864 ) ;
  assign n1866 = ( ~n1154 & n1861 ) | ( ~n1154 & n1864 ) | ( n1861 & n1864 ) ;
  assign n1867 = ( x409 & n1865 ) | ( x409 & n1866 ) | ( n1865 & n1866 ) ;
  assign n1868 = ( ~x281 & n1865 ) | ( ~x281 & n1866 ) | ( n1865 & n1866 ) ;
  assign n1869 = ( ~n656 & n1867 ) | ( ~n656 & n1868 ) | ( n1867 & n1868 ) ;
  assign n1870 = x260 & ~n991 ;
  assign n1871 = x260 & n995 ;
  assign n1872 = ( n1104 & n1870 ) | ( n1104 & n1871 ) | ( n1870 & n1871 ) ;
  assign n1873 = ( n1119 & n1870 ) | ( n1119 & n1871 ) | ( n1870 & n1871 ) ;
  assign n1874 = ( ~n1126 & n1870 ) | ( ~n1126 & n1871 ) | ( n1870 & n1871 ) ;
  assign n1875 = ( ~n1115 & n1873 ) | ( ~n1115 & n1874 ) | ( n1873 & n1874 ) ;
  assign n1876 = ( ~n975 & n1872 ) | ( ~n975 & n1875 ) | ( n1872 & n1875 ) ;
  assign n1877 = ( n1154 & n1872 ) | ( n1154 & n1875 ) | ( n1872 & n1875 ) ;
  assign n1878 = ( ~x409 & n1876 ) | ( ~x409 & n1877 ) | ( n1876 & n1877 ) ;
  assign n1879 = ( x281 & n1876 ) | ( x281 & n1877 ) | ( n1876 & n1877 ) ;
  assign n1880 = ( n656 & n1878 ) | ( n656 & n1879 ) | ( n1878 & n1879 ) ;
  assign n1881 = n1869 | n1880 ;
  assign n1882 = x131 & n1767 ;
  assign n1883 = x131 & ~n1771 ;
  assign n1884 = ( ~n1751 & n1882 ) | ( ~n1751 & n1883 ) | ( n1882 & n1883 ) ;
  assign n1885 = ( ~n1787 & n1882 ) | ( ~n1787 & n1883 ) | ( n1882 & n1883 ) ;
  assign n1886 = ( n1794 & n1882 ) | ( n1794 & n1883 ) | ( n1882 & n1883 ) ;
  assign n1887 = ( n1783 & n1885 ) | ( n1783 & n1886 ) | ( n1885 & n1886 ) ;
  assign n1888 = ( n1643 & n1884 ) | ( n1643 & n1887 ) | ( n1884 & n1887 ) ;
  assign n1889 = ( ~n1822 & n1884 ) | ( ~n1822 & n1887 ) | ( n1884 & n1887 ) ;
  assign n1890 = ( ~n1324 & n1888 ) | ( ~n1324 & n1889 ) | ( n1888 & n1889 ) ;
  assign n1891 = x3 & ~n1767 ;
  assign n1892 = x3 & n1771 ;
  assign n1893 = ( n1751 & n1891 ) | ( n1751 & n1892 ) | ( n1891 & n1892 ) ;
  assign n1894 = ( n1787 & n1891 ) | ( n1787 & n1892 ) | ( n1891 & n1892 ) ;
  assign n1895 = ( ~n1794 & n1891 ) | ( ~n1794 & n1892 ) | ( n1891 & n1892 ) ;
  assign n1896 = ( ~n1783 & n1894 ) | ( ~n1783 & n1895 ) | ( n1894 & n1895 ) ;
  assign n1897 = ( ~n1643 & n1893 ) | ( ~n1643 & n1896 ) | ( n1893 & n1896 ) ;
  assign n1898 = ( n1822 & n1893 ) | ( n1822 & n1896 ) | ( n1893 & n1896 ) ;
  assign n1899 = ( n1324 & n1897 ) | ( n1324 & n1898 ) | ( n1897 & n1898 ) ;
  assign n1900 = n1890 | n1899 ;
  assign n1901 = x387 & n991 ;
  assign n1902 = x387 & ~n995 ;
  assign n1903 = ( ~n1104 & n1901 ) | ( ~n1104 & n1902 ) | ( n1901 & n1902 ) ;
  assign n1904 = ( ~n1119 & n1901 ) | ( ~n1119 & n1902 ) | ( n1901 & n1902 ) ;
  assign n1905 = ( n1126 & n1901 ) | ( n1126 & n1902 ) | ( n1901 & n1902 ) ;
  assign n1906 = ( n1115 & n1904 ) | ( n1115 & n1905 ) | ( n1904 & n1905 ) ;
  assign n1907 = ( n975 & n1903 ) | ( n975 & n1906 ) | ( n1903 & n1906 ) ;
  assign n1908 = ( ~n1154 & n1903 ) | ( ~n1154 & n1906 ) | ( n1903 & n1906 ) ;
  assign n1909 = ( x409 & n1907 ) | ( x409 & n1908 ) | ( n1907 & n1908 ) ;
  assign n1910 = ( ~x281 & n1907 ) | ( ~x281 & n1908 ) | ( n1907 & n1908 ) ;
  assign n1911 = ( ~n656 & n1909 ) | ( ~n656 & n1910 ) | ( n1909 & n1910 ) ;
  assign n1912 = x259 & ~n991 ;
  assign n1913 = x259 & n995 ;
  assign n1914 = ( n1104 & n1912 ) | ( n1104 & n1913 ) | ( n1912 & n1913 ) ;
  assign n1915 = ( n1119 & n1912 ) | ( n1119 & n1913 ) | ( n1912 & n1913 ) ;
  assign n1916 = ( ~n1126 & n1912 ) | ( ~n1126 & n1913 ) | ( n1912 & n1913 ) ;
  assign n1917 = ( ~n1115 & n1915 ) | ( ~n1115 & n1916 ) | ( n1915 & n1916 ) ;
  assign n1918 = ( ~n975 & n1914 ) | ( ~n975 & n1917 ) | ( n1914 & n1917 ) ;
  assign n1919 = ( n1154 & n1914 ) | ( n1154 & n1917 ) | ( n1914 & n1917 ) ;
  assign n1920 = ( ~x409 & n1918 ) | ( ~x409 & n1919 ) | ( n1918 & n1919 ) ;
  assign n1921 = ( x281 & n1918 ) | ( x281 & n1919 ) | ( n1918 & n1919 ) ;
  assign n1922 = ( n656 & n1920 ) | ( n656 & n1921 ) | ( n1920 & n1921 ) ;
  assign n1923 = n1911 | n1922 ;
  assign n1924 = ~n1900 & n1923 ;
  assign n1925 = x132 & n1767 ;
  assign n1926 = x132 & ~n1771 ;
  assign n1927 = ( ~n1751 & n1925 ) | ( ~n1751 & n1926 ) | ( n1925 & n1926 ) ;
  assign n1928 = ( ~n1787 & n1925 ) | ( ~n1787 & n1926 ) | ( n1925 & n1926 ) ;
  assign n1929 = ( n1794 & n1925 ) | ( n1794 & n1926 ) | ( n1925 & n1926 ) ;
  assign n1930 = ( n1783 & n1928 ) | ( n1783 & n1929 ) | ( n1928 & n1929 ) ;
  assign n1931 = ( n1643 & n1927 ) | ( n1643 & n1930 ) | ( n1927 & n1930 ) ;
  assign n1932 = ( ~n1822 & n1927 ) | ( ~n1822 & n1930 ) | ( n1927 & n1930 ) ;
  assign n1933 = ( ~n1324 & n1931 ) | ( ~n1324 & n1932 ) | ( n1931 & n1932 ) ;
  assign n1934 = x4 & ~n1767 ;
  assign n1935 = x4 & n1771 ;
  assign n1936 = ( n1751 & n1934 ) | ( n1751 & n1935 ) | ( n1934 & n1935 ) ;
  assign n1937 = ( n1787 & n1934 ) | ( n1787 & n1935 ) | ( n1934 & n1935 ) ;
  assign n1938 = ( ~n1794 & n1934 ) | ( ~n1794 & n1935 ) | ( n1934 & n1935 ) ;
  assign n1939 = ( ~n1783 & n1937 ) | ( ~n1783 & n1938 ) | ( n1937 & n1938 ) ;
  assign n1940 = ( ~n1643 & n1936 ) | ( ~n1643 & n1939 ) | ( n1936 & n1939 ) ;
  assign n1941 = ( n1822 & n1936 ) | ( n1822 & n1939 ) | ( n1936 & n1939 ) ;
  assign n1942 = ( n1324 & n1940 ) | ( n1324 & n1941 ) | ( n1940 & n1941 ) ;
  assign n1943 = n1933 | n1942 ;
  assign n1944 = ~n1881 & n1943 ;
  assign n1945 = ( n1881 & n1924 ) | ( n1881 & ~n1944 ) | ( n1924 & ~n1944 ) ;
  assign n1946 = n1900 & ~n1923 ;
  assign n1947 = ( ~n1881 & n1944 ) | ( ~n1881 & n1946 ) | ( n1944 & n1946 ) ;
  assign n1948 = x386 & n991 ;
  assign n1949 = x386 & ~n995 ;
  assign n1950 = ( ~n1104 & n1948 ) | ( ~n1104 & n1949 ) | ( n1948 & n1949 ) ;
  assign n1951 = ( ~n1119 & n1948 ) | ( ~n1119 & n1949 ) | ( n1948 & n1949 ) ;
  assign n1952 = ( n1126 & n1948 ) | ( n1126 & n1949 ) | ( n1948 & n1949 ) ;
  assign n1953 = ( n1115 & n1951 ) | ( n1115 & n1952 ) | ( n1951 & n1952 ) ;
  assign n1954 = ( n975 & n1950 ) | ( n975 & n1953 ) | ( n1950 & n1953 ) ;
  assign n1955 = ( ~n1154 & n1950 ) | ( ~n1154 & n1953 ) | ( n1950 & n1953 ) ;
  assign n1956 = ( x409 & n1954 ) | ( x409 & n1955 ) | ( n1954 & n1955 ) ;
  assign n1957 = ( ~x281 & n1954 ) | ( ~x281 & n1955 ) | ( n1954 & n1955 ) ;
  assign n1958 = ( ~n656 & n1956 ) | ( ~n656 & n1957 ) | ( n1956 & n1957 ) ;
  assign n1959 = x258 & ~n991 ;
  assign n1960 = x258 & n995 ;
  assign n1961 = ( n1104 & n1959 ) | ( n1104 & n1960 ) | ( n1959 & n1960 ) ;
  assign n1962 = ( n1119 & n1959 ) | ( n1119 & n1960 ) | ( n1959 & n1960 ) ;
  assign n1963 = ( ~n1126 & n1959 ) | ( ~n1126 & n1960 ) | ( n1959 & n1960 ) ;
  assign n1964 = ( ~n1115 & n1962 ) | ( ~n1115 & n1963 ) | ( n1962 & n1963 ) ;
  assign n1965 = ( ~n975 & n1961 ) | ( ~n975 & n1964 ) | ( n1961 & n1964 ) ;
  assign n1966 = ( n1154 & n1961 ) | ( n1154 & n1964 ) | ( n1961 & n1964 ) ;
  assign n1967 = ( ~x409 & n1965 ) | ( ~x409 & n1966 ) | ( n1965 & n1966 ) ;
  assign n1968 = ( x281 & n1965 ) | ( x281 & n1966 ) | ( n1965 & n1966 ) ;
  assign n1969 = ( n656 & n1967 ) | ( n656 & n1968 ) | ( n1967 & n1968 ) ;
  assign n1970 = n1958 | n1969 ;
  assign n1971 = ( n1945 & ~n1947 ) | ( n1945 & n1970 ) | ( ~n1947 & n1970 ) ;
  assign n1972 = x130 & n1767 ;
  assign n1973 = x130 & ~n1771 ;
  assign n1974 = ( ~n1751 & n1972 ) | ( ~n1751 & n1973 ) | ( n1972 & n1973 ) ;
  assign n1975 = ( ~n1787 & n1972 ) | ( ~n1787 & n1973 ) | ( n1972 & n1973 ) ;
  assign n1976 = ( n1794 & n1972 ) | ( n1794 & n1973 ) | ( n1972 & n1973 ) ;
  assign n1977 = ( n1783 & n1975 ) | ( n1783 & n1976 ) | ( n1975 & n1976 ) ;
  assign n1978 = ( n1643 & n1974 ) | ( n1643 & n1977 ) | ( n1974 & n1977 ) ;
  assign n1979 = ( ~n1822 & n1974 ) | ( ~n1822 & n1977 ) | ( n1974 & n1977 ) ;
  assign n1980 = ( ~n1324 & n1978 ) | ( ~n1324 & n1979 ) | ( n1978 & n1979 ) ;
  assign n1981 = x2 & ~n1767 ;
  assign n1982 = x2 & n1771 ;
  assign n1983 = ( n1751 & n1981 ) | ( n1751 & n1982 ) | ( n1981 & n1982 ) ;
  assign n1984 = ( n1787 & n1981 ) | ( n1787 & n1982 ) | ( n1981 & n1982 ) ;
  assign n1985 = ( ~n1794 & n1981 ) | ( ~n1794 & n1982 ) | ( n1981 & n1982 ) ;
  assign n1986 = ( ~n1783 & n1984 ) | ( ~n1783 & n1985 ) | ( n1984 & n1985 ) ;
  assign n1987 = ( ~n1643 & n1983 ) | ( ~n1643 & n1986 ) | ( n1983 & n1986 ) ;
  assign n1988 = ( n1822 & n1983 ) | ( n1822 & n1986 ) | ( n1983 & n1986 ) ;
  assign n1989 = ( n1324 & n1987 ) | ( n1324 & n1988 ) | ( n1987 & n1988 ) ;
  assign n1990 = n1980 | n1989 ;
  assign n1991 = ( ~n1945 & n1947 ) | ( ~n1945 & n1990 ) | ( n1947 & n1990 ) ;
  assign n1992 = ( n1858 & ~n1971 ) | ( n1858 & n1991 ) | ( ~n1971 & n1991 ) ;
  assign n1993 = ( ~n1924 & n1946 ) | ( ~n1924 & n1990 ) | ( n1946 & n1990 ) ;
  assign n1994 = n1943 & n1993 ;
  assign n1995 = ( n1924 & ~n1946 ) | ( n1924 & n1970 ) | ( ~n1946 & n1970 ) ;
  assign n1996 = n1943 & ~n1995 ;
  assign n1997 = ( n1858 & n1994 ) | ( n1858 & n1996 ) | ( n1994 & n1996 ) ;
  assign n1998 = n1992 | n1997 ;
  assign n1999 = x392 & n991 ;
  assign n2000 = x392 & ~n995 ;
  assign n2001 = ( ~n1104 & n1999 ) | ( ~n1104 & n2000 ) | ( n1999 & n2000 ) ;
  assign n2002 = ( ~n1119 & n1999 ) | ( ~n1119 & n2000 ) | ( n1999 & n2000 ) ;
  assign n2003 = ( n1126 & n1999 ) | ( n1126 & n2000 ) | ( n1999 & n2000 ) ;
  assign n2004 = ( n1115 & n2002 ) | ( n1115 & n2003 ) | ( n2002 & n2003 ) ;
  assign n2005 = ( n975 & n2001 ) | ( n975 & n2004 ) | ( n2001 & n2004 ) ;
  assign n2006 = ( ~n1154 & n2001 ) | ( ~n1154 & n2004 ) | ( n2001 & n2004 ) ;
  assign n2007 = ( x409 & n2005 ) | ( x409 & n2006 ) | ( n2005 & n2006 ) ;
  assign n2008 = ( ~x281 & n2005 ) | ( ~x281 & n2006 ) | ( n2005 & n2006 ) ;
  assign n2009 = ( ~n656 & n2007 ) | ( ~n656 & n2008 ) | ( n2007 & n2008 ) ;
  assign n2010 = x264 & ~n991 ;
  assign n2011 = x264 & n995 ;
  assign n2012 = ( n1104 & n2010 ) | ( n1104 & n2011 ) | ( n2010 & n2011 ) ;
  assign n2013 = ( n1119 & n2010 ) | ( n1119 & n2011 ) | ( n2010 & n2011 ) ;
  assign n2014 = ( ~n1126 & n2010 ) | ( ~n1126 & n2011 ) | ( n2010 & n2011 ) ;
  assign n2015 = ( ~n1115 & n2013 ) | ( ~n1115 & n2014 ) | ( n2013 & n2014 ) ;
  assign n2016 = ( ~n975 & n2012 ) | ( ~n975 & n2015 ) | ( n2012 & n2015 ) ;
  assign n2017 = ( n1154 & n2012 ) | ( n1154 & n2015 ) | ( n2012 & n2015 ) ;
  assign n2018 = ( ~x409 & n2016 ) | ( ~x409 & n2017 ) | ( n2016 & n2017 ) ;
  assign n2019 = ( x281 & n2016 ) | ( x281 & n2017 ) | ( n2016 & n2017 ) ;
  assign n2020 = ( n656 & n2018 ) | ( n656 & n2019 ) | ( n2018 & n2019 ) ;
  assign n2021 = n2009 | n2020 ;
  assign n2022 = x135 & n1767 ;
  assign n2023 = x135 & ~n1771 ;
  assign n2024 = ( ~n1751 & n2022 ) | ( ~n1751 & n2023 ) | ( n2022 & n2023 ) ;
  assign n2025 = ( ~n1787 & n2022 ) | ( ~n1787 & n2023 ) | ( n2022 & n2023 ) ;
  assign n2026 = ( n1794 & n2022 ) | ( n1794 & n2023 ) | ( n2022 & n2023 ) ;
  assign n2027 = ( n1783 & n2025 ) | ( n1783 & n2026 ) | ( n2025 & n2026 ) ;
  assign n2028 = ( n1643 & n2024 ) | ( n1643 & n2027 ) | ( n2024 & n2027 ) ;
  assign n2029 = ( ~n1822 & n2024 ) | ( ~n1822 & n2027 ) | ( n2024 & n2027 ) ;
  assign n2030 = ( ~n1324 & n2028 ) | ( ~n1324 & n2029 ) | ( n2028 & n2029 ) ;
  assign n2031 = x7 & ~n1767 ;
  assign n2032 = x7 & n1771 ;
  assign n2033 = ( n1751 & n2031 ) | ( n1751 & n2032 ) | ( n2031 & n2032 ) ;
  assign n2034 = ( n1787 & n2031 ) | ( n1787 & n2032 ) | ( n2031 & n2032 ) ;
  assign n2035 = ( ~n1794 & n2031 ) | ( ~n1794 & n2032 ) | ( n2031 & n2032 ) ;
  assign n2036 = ( ~n1783 & n2034 ) | ( ~n1783 & n2035 ) | ( n2034 & n2035 ) ;
  assign n2037 = ( ~n1643 & n2033 ) | ( ~n1643 & n2036 ) | ( n2033 & n2036 ) ;
  assign n2038 = ( n1822 & n2033 ) | ( n1822 & n2036 ) | ( n2033 & n2036 ) ;
  assign n2039 = ( n1324 & n2037 ) | ( n1324 & n2038 ) | ( n2037 & n2038 ) ;
  assign n2040 = n2030 | n2039 ;
  assign n2041 = x391 & n991 ;
  assign n2042 = x391 & ~n995 ;
  assign n2043 = ( ~n1104 & n2041 ) | ( ~n1104 & n2042 ) | ( n2041 & n2042 ) ;
  assign n2044 = ( ~n1119 & n2041 ) | ( ~n1119 & n2042 ) | ( n2041 & n2042 ) ;
  assign n2045 = ( n1126 & n2041 ) | ( n1126 & n2042 ) | ( n2041 & n2042 ) ;
  assign n2046 = ( n1115 & n2044 ) | ( n1115 & n2045 ) | ( n2044 & n2045 ) ;
  assign n2047 = ( n975 & n2043 ) | ( n975 & n2046 ) | ( n2043 & n2046 ) ;
  assign n2048 = ( ~n1154 & n2043 ) | ( ~n1154 & n2046 ) | ( n2043 & n2046 ) ;
  assign n2049 = ( x409 & n2047 ) | ( x409 & n2048 ) | ( n2047 & n2048 ) ;
  assign n2050 = ( ~x281 & n2047 ) | ( ~x281 & n2048 ) | ( n2047 & n2048 ) ;
  assign n2051 = ( ~n656 & n2049 ) | ( ~n656 & n2050 ) | ( n2049 & n2050 ) ;
  assign n2052 = x263 & ~n991 ;
  assign n2053 = x263 & n995 ;
  assign n2054 = ( n1104 & n2052 ) | ( n1104 & n2053 ) | ( n2052 & n2053 ) ;
  assign n2055 = ( n1119 & n2052 ) | ( n1119 & n2053 ) | ( n2052 & n2053 ) ;
  assign n2056 = ( ~n1126 & n2052 ) | ( ~n1126 & n2053 ) | ( n2052 & n2053 ) ;
  assign n2057 = ( ~n1115 & n2055 ) | ( ~n1115 & n2056 ) | ( n2055 & n2056 ) ;
  assign n2058 = ( ~n975 & n2054 ) | ( ~n975 & n2057 ) | ( n2054 & n2057 ) ;
  assign n2059 = ( n1154 & n2054 ) | ( n1154 & n2057 ) | ( n2054 & n2057 ) ;
  assign n2060 = ( ~x409 & n2058 ) | ( ~x409 & n2059 ) | ( n2058 & n2059 ) ;
  assign n2061 = ( x281 & n2058 ) | ( x281 & n2059 ) | ( n2058 & n2059 ) ;
  assign n2062 = ( n656 & n2060 ) | ( n656 & n2061 ) | ( n2060 & n2061 ) ;
  assign n2063 = n2051 | n2062 ;
  assign n2064 = ~n2040 & n2063 ;
  assign n2065 = x136 & n1767 ;
  assign n2066 = x136 & ~n1771 ;
  assign n2067 = ( ~n1751 & n2065 ) | ( ~n1751 & n2066 ) | ( n2065 & n2066 ) ;
  assign n2068 = ( ~n1787 & n2065 ) | ( ~n1787 & n2066 ) | ( n2065 & n2066 ) ;
  assign n2069 = ( n1794 & n2065 ) | ( n1794 & n2066 ) | ( n2065 & n2066 ) ;
  assign n2070 = ( n1783 & n2068 ) | ( n1783 & n2069 ) | ( n2068 & n2069 ) ;
  assign n2071 = ( n1643 & n2067 ) | ( n1643 & n2070 ) | ( n2067 & n2070 ) ;
  assign n2072 = ( ~n1822 & n2067 ) | ( ~n1822 & n2070 ) | ( n2067 & n2070 ) ;
  assign n2073 = ( ~n1324 & n2071 ) | ( ~n1324 & n2072 ) | ( n2071 & n2072 ) ;
  assign n2074 = x8 & ~n1767 ;
  assign n2075 = x8 & n1771 ;
  assign n2076 = ( n1751 & n2074 ) | ( n1751 & n2075 ) | ( n2074 & n2075 ) ;
  assign n2077 = ( n1787 & n2074 ) | ( n1787 & n2075 ) | ( n2074 & n2075 ) ;
  assign n2078 = ( ~n1794 & n2074 ) | ( ~n1794 & n2075 ) | ( n2074 & n2075 ) ;
  assign n2079 = ( ~n1783 & n2077 ) | ( ~n1783 & n2078 ) | ( n2077 & n2078 ) ;
  assign n2080 = ( ~n1643 & n2076 ) | ( ~n1643 & n2079 ) | ( n2076 & n2079 ) ;
  assign n2081 = ( n1822 & n2076 ) | ( n1822 & n2079 ) | ( n2076 & n2079 ) ;
  assign n2082 = ( n1324 & n2080 ) | ( n1324 & n2081 ) | ( n2080 & n2081 ) ;
  assign n2083 = n2073 | n2082 ;
  assign n2084 = ~n2021 & n2083 ;
  assign n2085 = ( n2021 & n2064 ) | ( n2021 & ~n2084 ) | ( n2064 & ~n2084 ) ;
  assign n2086 = n2040 & ~n2063 ;
  assign n2087 = ( ~n2021 & n2084 ) | ( ~n2021 & n2086 ) | ( n2084 & n2086 ) ;
  assign n2088 = x134 & n1767 ;
  assign n2089 = x134 & ~n1771 ;
  assign n2090 = ( ~n1751 & n2088 ) | ( ~n1751 & n2089 ) | ( n2088 & n2089 ) ;
  assign n2091 = ( ~n1787 & n2088 ) | ( ~n1787 & n2089 ) | ( n2088 & n2089 ) ;
  assign n2092 = ( n1794 & n2088 ) | ( n1794 & n2089 ) | ( n2088 & n2089 ) ;
  assign n2093 = ( n1783 & n2091 ) | ( n1783 & n2092 ) | ( n2091 & n2092 ) ;
  assign n2094 = ( n1643 & n2090 ) | ( n1643 & n2093 ) | ( n2090 & n2093 ) ;
  assign n2095 = ( ~n1822 & n2090 ) | ( ~n1822 & n2093 ) | ( n2090 & n2093 ) ;
  assign n2096 = ( ~n1324 & n2094 ) | ( ~n1324 & n2095 ) | ( n2094 & n2095 ) ;
  assign n2097 = x6 & ~n1767 ;
  assign n2098 = x6 & n1771 ;
  assign n2099 = ( n1751 & n2097 ) | ( n1751 & n2098 ) | ( n2097 & n2098 ) ;
  assign n2100 = ( n1787 & n2097 ) | ( n1787 & n2098 ) | ( n2097 & n2098 ) ;
  assign n2101 = ( ~n1794 & n2097 ) | ( ~n1794 & n2098 ) | ( n2097 & n2098 ) ;
  assign n2102 = ( ~n1783 & n2100 ) | ( ~n1783 & n2101 ) | ( n2100 & n2101 ) ;
  assign n2103 = ( ~n1643 & n2099 ) | ( ~n1643 & n2102 ) | ( n2099 & n2102 ) ;
  assign n2104 = ( n1822 & n2099 ) | ( n1822 & n2102 ) | ( n2099 & n2102 ) ;
  assign n2105 = ( n1324 & n2103 ) | ( n1324 & n2104 ) | ( n2103 & n2104 ) ;
  assign n2106 = n2096 | n2105 ;
  assign n2107 = x390 & n991 ;
  assign n2108 = x390 & ~n995 ;
  assign n2109 = ( ~n1104 & n2107 ) | ( ~n1104 & n2108 ) | ( n2107 & n2108 ) ;
  assign n2110 = ( ~n1119 & n2107 ) | ( ~n1119 & n2108 ) | ( n2107 & n2108 ) ;
  assign n2111 = ( n1126 & n2107 ) | ( n1126 & n2108 ) | ( n2107 & n2108 ) ;
  assign n2112 = ( n1115 & n2110 ) | ( n1115 & n2111 ) | ( n2110 & n2111 ) ;
  assign n2113 = ( n975 & n2109 ) | ( n975 & n2112 ) | ( n2109 & n2112 ) ;
  assign n2114 = ( ~n1154 & n2109 ) | ( ~n1154 & n2112 ) | ( n2109 & n2112 ) ;
  assign n2115 = ( x409 & n2113 ) | ( x409 & n2114 ) | ( n2113 & n2114 ) ;
  assign n2116 = ( ~x281 & n2113 ) | ( ~x281 & n2114 ) | ( n2113 & n2114 ) ;
  assign n2117 = ( ~n656 & n2115 ) | ( ~n656 & n2116 ) | ( n2115 & n2116 ) ;
  assign n2118 = x262 & ~n991 ;
  assign n2119 = x262 & n995 ;
  assign n2120 = ( n1104 & n2118 ) | ( n1104 & n2119 ) | ( n2118 & n2119 ) ;
  assign n2121 = ( n1119 & n2118 ) | ( n1119 & n2119 ) | ( n2118 & n2119 ) ;
  assign n2122 = ( ~n1126 & n2118 ) | ( ~n1126 & n2119 ) | ( n2118 & n2119 ) ;
  assign n2123 = ( ~n1115 & n2121 ) | ( ~n1115 & n2122 ) | ( n2121 & n2122 ) ;
  assign n2124 = ( ~n975 & n2120 ) | ( ~n975 & n2123 ) | ( n2120 & n2123 ) ;
  assign n2125 = ( n1154 & n2120 ) | ( n1154 & n2123 ) | ( n2120 & n2123 ) ;
  assign n2126 = ( ~x409 & n2124 ) | ( ~x409 & n2125 ) | ( n2124 & n2125 ) ;
  assign n2127 = ( x281 & n2124 ) | ( x281 & n2125 ) | ( n2124 & n2125 ) ;
  assign n2128 = ( n656 & n2126 ) | ( n656 & n2127 ) | ( n2126 & n2127 ) ;
  assign n2129 = n2117 | n2128 ;
  assign n2130 = x133 & n1767 ;
  assign n2131 = x133 & ~n1771 ;
  assign n2132 = ( ~n1751 & n2130 ) | ( ~n1751 & n2131 ) | ( n2130 & n2131 ) ;
  assign n2133 = ( ~n1787 & n2130 ) | ( ~n1787 & n2131 ) | ( n2130 & n2131 ) ;
  assign n2134 = ( n1794 & n2130 ) | ( n1794 & n2131 ) | ( n2130 & n2131 ) ;
  assign n2135 = ( n1783 & n2133 ) | ( n1783 & n2134 ) | ( n2133 & n2134 ) ;
  assign n2136 = ( n1643 & n2132 ) | ( n1643 & n2135 ) | ( n2132 & n2135 ) ;
  assign n2137 = ( ~n1822 & n2132 ) | ( ~n1822 & n2135 ) | ( n2132 & n2135 ) ;
  assign n2138 = ( ~n1324 & n2136 ) | ( ~n1324 & n2137 ) | ( n2136 & n2137 ) ;
  assign n2139 = x5 & ~n1767 ;
  assign n2140 = x5 & n1771 ;
  assign n2141 = ( n1751 & n2139 ) | ( n1751 & n2140 ) | ( n2139 & n2140 ) ;
  assign n2142 = ( n1787 & n2139 ) | ( n1787 & n2140 ) | ( n2139 & n2140 ) ;
  assign n2143 = ( ~n1794 & n2139 ) | ( ~n1794 & n2140 ) | ( n2139 & n2140 ) ;
  assign n2144 = ( ~n1783 & n2142 ) | ( ~n1783 & n2143 ) | ( n2142 & n2143 ) ;
  assign n2145 = ( ~n1643 & n2141 ) | ( ~n1643 & n2144 ) | ( n2141 & n2144 ) ;
  assign n2146 = ( n1822 & n2141 ) | ( n1822 & n2144 ) | ( n2141 & n2144 ) ;
  assign n2147 = ( n1324 & n2145 ) | ( n1324 & n2146 ) | ( n2145 & n2146 ) ;
  assign n2148 = n2138 | n2147 ;
  assign n2149 = ( n2106 & ~n2129 ) | ( n2106 & n2148 ) | ( ~n2129 & n2148 ) ;
  assign n2150 = ( ~n2085 & n2087 ) | ( ~n2085 & n2149 ) | ( n2087 & n2149 ) ;
  assign n2151 = x389 & n991 ;
  assign n2152 = x389 & ~n995 ;
  assign n2153 = ( ~n1104 & n2151 ) | ( ~n1104 & n2152 ) | ( n2151 & n2152 ) ;
  assign n2154 = ( ~n1119 & n2151 ) | ( ~n1119 & n2152 ) | ( n2151 & n2152 ) ;
  assign n2155 = ( n1126 & n2151 ) | ( n1126 & n2152 ) | ( n2151 & n2152 ) ;
  assign n2156 = ( n1115 & n2154 ) | ( n1115 & n2155 ) | ( n2154 & n2155 ) ;
  assign n2157 = ( n975 & n2153 ) | ( n975 & n2156 ) | ( n2153 & n2156 ) ;
  assign n2158 = ( ~n1154 & n2153 ) | ( ~n1154 & n2156 ) | ( n2153 & n2156 ) ;
  assign n2159 = ( x409 & n2157 ) | ( x409 & n2158 ) | ( n2157 & n2158 ) ;
  assign n2160 = ( ~x281 & n2157 ) | ( ~x281 & n2158 ) | ( n2157 & n2158 ) ;
  assign n2161 = ( ~n656 & n2159 ) | ( ~n656 & n2160 ) | ( n2159 & n2160 ) ;
  assign n2162 = x261 & ~n991 ;
  assign n2163 = x261 & n995 ;
  assign n2164 = ( n1104 & n2162 ) | ( n1104 & n2163 ) | ( n2162 & n2163 ) ;
  assign n2165 = ( n1119 & n2162 ) | ( n1119 & n2163 ) | ( n2162 & n2163 ) ;
  assign n2166 = ( ~n1126 & n2162 ) | ( ~n1126 & n2163 ) | ( n2162 & n2163 ) ;
  assign n2167 = ( ~n1115 & n2165 ) | ( ~n1115 & n2166 ) | ( n2165 & n2166 ) ;
  assign n2168 = ( ~n975 & n2164 ) | ( ~n975 & n2167 ) | ( n2164 & n2167 ) ;
  assign n2169 = ( n1154 & n2164 ) | ( n1154 & n2167 ) | ( n2164 & n2167 ) ;
  assign n2170 = ( ~x409 & n2168 ) | ( ~x409 & n2169 ) | ( n2168 & n2169 ) ;
  assign n2171 = ( x281 & n2168 ) | ( x281 & n2169 ) | ( n2168 & n2169 ) ;
  assign n2172 = ( n656 & n2170 ) | ( n656 & n2171 ) | ( n2170 & n2171 ) ;
  assign n2173 = n2161 | n2172 ;
  assign n2174 = ( ~n2106 & n2129 ) | ( ~n2106 & n2173 ) | ( n2129 & n2173 ) ;
  assign n2175 = ( n2085 & ~n2087 ) | ( n2085 & n2174 ) | ( ~n2087 & n2174 ) ;
  assign n2176 = ( n1998 & n2150 ) | ( n1998 & ~n2175 ) | ( n2150 & ~n2175 ) ;
  assign n2177 = ( n2064 & ~n2086 ) | ( n2064 & n2174 ) | ( ~n2086 & n2174 ) ;
  assign n2178 = n2083 & ~n2177 ;
  assign n2179 = ( ~n2064 & n2086 ) | ( ~n2064 & n2149 ) | ( n2086 & n2149 ) ;
  assign n2180 = n2083 & n2179 ;
  assign n2181 = ( n1998 & n2178 ) | ( n1998 & n2180 ) | ( n2178 & n2180 ) ;
  assign n2182 = n2176 | n2181 ;
  assign n2183 = x141 & n1767 ;
  assign n2184 = x141 & ~n1771 ;
  assign n2185 = ( ~n1751 & n2183 ) | ( ~n1751 & n2184 ) | ( n2183 & n2184 ) ;
  assign n2186 = ( ~n1787 & n2183 ) | ( ~n1787 & n2184 ) | ( n2183 & n2184 ) ;
  assign n2187 = ( n1794 & n2183 ) | ( n1794 & n2184 ) | ( n2183 & n2184 ) ;
  assign n2188 = ( n1783 & n2186 ) | ( n1783 & n2187 ) | ( n2186 & n2187 ) ;
  assign n2189 = ( n1643 & n2185 ) | ( n1643 & n2188 ) | ( n2185 & n2188 ) ;
  assign n2190 = ( ~n1822 & n2185 ) | ( ~n1822 & n2188 ) | ( n2185 & n2188 ) ;
  assign n2191 = ( ~n1324 & n2189 ) | ( ~n1324 & n2190 ) | ( n2189 & n2190 ) ;
  assign n2192 = x13 & ~n1767 ;
  assign n2193 = x13 & n1771 ;
  assign n2194 = ( n1751 & n2192 ) | ( n1751 & n2193 ) | ( n2192 & n2193 ) ;
  assign n2195 = ( n1787 & n2192 ) | ( n1787 & n2193 ) | ( n2192 & n2193 ) ;
  assign n2196 = ( ~n1794 & n2192 ) | ( ~n1794 & n2193 ) | ( n2192 & n2193 ) ;
  assign n2197 = ( ~n1783 & n2195 ) | ( ~n1783 & n2196 ) | ( n2195 & n2196 ) ;
  assign n2198 = ( ~n1643 & n2194 ) | ( ~n1643 & n2197 ) | ( n2194 & n2197 ) ;
  assign n2199 = ( n1822 & n2194 ) | ( n1822 & n2197 ) | ( n2194 & n2197 ) ;
  assign n2200 = ( n1324 & n2198 ) | ( n1324 & n2199 ) | ( n2198 & n2199 ) ;
  assign n2201 = n2191 | n2200 ;
  assign n2202 = x397 & n991 ;
  assign n2203 = x397 & ~n995 ;
  assign n2204 = ( ~n1104 & n2202 ) | ( ~n1104 & n2203 ) | ( n2202 & n2203 ) ;
  assign n2205 = ( ~n1119 & n2202 ) | ( ~n1119 & n2203 ) | ( n2202 & n2203 ) ;
  assign n2206 = ( n1126 & n2202 ) | ( n1126 & n2203 ) | ( n2202 & n2203 ) ;
  assign n2207 = ( n1115 & n2205 ) | ( n1115 & n2206 ) | ( n2205 & n2206 ) ;
  assign n2208 = ( n975 & n2204 ) | ( n975 & n2207 ) | ( n2204 & n2207 ) ;
  assign n2209 = ( ~n1154 & n2204 ) | ( ~n1154 & n2207 ) | ( n2204 & n2207 ) ;
  assign n2210 = ( x409 & n2208 ) | ( x409 & n2209 ) | ( n2208 & n2209 ) ;
  assign n2211 = ( ~x281 & n2208 ) | ( ~x281 & n2209 ) | ( n2208 & n2209 ) ;
  assign n2212 = ( ~n656 & n2210 ) | ( ~n656 & n2211 ) | ( n2210 & n2211 ) ;
  assign n2213 = x269 & ~n991 ;
  assign n2214 = x269 & n995 ;
  assign n2215 = ( n1104 & n2213 ) | ( n1104 & n2214 ) | ( n2213 & n2214 ) ;
  assign n2216 = ( n1119 & n2213 ) | ( n1119 & n2214 ) | ( n2213 & n2214 ) ;
  assign n2217 = ( ~n1126 & n2213 ) | ( ~n1126 & n2214 ) | ( n2213 & n2214 ) ;
  assign n2218 = ( ~n1115 & n2216 ) | ( ~n1115 & n2217 ) | ( n2216 & n2217 ) ;
  assign n2219 = ( ~n975 & n2215 ) | ( ~n975 & n2218 ) | ( n2215 & n2218 ) ;
  assign n2220 = ( n1154 & n2215 ) | ( n1154 & n2218 ) | ( n2215 & n2218 ) ;
  assign n2221 = ( ~x409 & n2219 ) | ( ~x409 & n2220 ) | ( n2219 & n2220 ) ;
  assign n2222 = ( x281 & n2219 ) | ( x281 & n2220 ) | ( n2219 & n2220 ) ;
  assign n2223 = ( n656 & n2221 ) | ( n656 & n2222 ) | ( n2221 & n2222 ) ;
  assign n2224 = n2212 | n2223 ;
  assign n2225 = ~n2201 & n2224 ;
  assign n2226 = x140 & n1767 ;
  assign n2227 = x140 & ~n1771 ;
  assign n2228 = ( ~n1751 & n2226 ) | ( ~n1751 & n2227 ) | ( n2226 & n2227 ) ;
  assign n2229 = ( ~n1787 & n2226 ) | ( ~n1787 & n2227 ) | ( n2226 & n2227 ) ;
  assign n2230 = ( n1794 & n2226 ) | ( n1794 & n2227 ) | ( n2226 & n2227 ) ;
  assign n2231 = ( n1783 & n2229 ) | ( n1783 & n2230 ) | ( n2229 & n2230 ) ;
  assign n2232 = ( n1643 & n2228 ) | ( n1643 & n2231 ) | ( n2228 & n2231 ) ;
  assign n2233 = ( ~n1822 & n2228 ) | ( ~n1822 & n2231 ) | ( n2228 & n2231 ) ;
  assign n2234 = ( ~n1324 & n2232 ) | ( ~n1324 & n2233 ) | ( n2232 & n2233 ) ;
  assign n2235 = x12 & ~n1767 ;
  assign n2236 = x12 & n1771 ;
  assign n2237 = ( n1751 & n2235 ) | ( n1751 & n2236 ) | ( n2235 & n2236 ) ;
  assign n2238 = ( n1787 & n2235 ) | ( n1787 & n2236 ) | ( n2235 & n2236 ) ;
  assign n2239 = ( ~n1794 & n2235 ) | ( ~n1794 & n2236 ) | ( n2235 & n2236 ) ;
  assign n2240 = ( ~n1783 & n2238 ) | ( ~n1783 & n2239 ) | ( n2238 & n2239 ) ;
  assign n2241 = ( ~n1643 & n2237 ) | ( ~n1643 & n2240 ) | ( n2237 & n2240 ) ;
  assign n2242 = ( n1822 & n2237 ) | ( n1822 & n2240 ) | ( n2237 & n2240 ) ;
  assign n2243 = ( n1324 & n2241 ) | ( n1324 & n2242 ) | ( n2241 & n2242 ) ;
  assign n2244 = n2234 | n2243 ;
  assign n2245 = x396 & n991 ;
  assign n2246 = x396 & ~n995 ;
  assign n2247 = ( ~n1104 & n2245 ) | ( ~n1104 & n2246 ) | ( n2245 & n2246 ) ;
  assign n2248 = ( ~n1119 & n2245 ) | ( ~n1119 & n2246 ) | ( n2245 & n2246 ) ;
  assign n2249 = ( n1126 & n2245 ) | ( n1126 & n2246 ) | ( n2245 & n2246 ) ;
  assign n2250 = ( n1115 & n2248 ) | ( n1115 & n2249 ) | ( n2248 & n2249 ) ;
  assign n2251 = ( n975 & n2247 ) | ( n975 & n2250 ) | ( n2247 & n2250 ) ;
  assign n2252 = ( ~n1154 & n2247 ) | ( ~n1154 & n2250 ) | ( n2247 & n2250 ) ;
  assign n2253 = ( x409 & n2251 ) | ( x409 & n2252 ) | ( n2251 & n2252 ) ;
  assign n2254 = ( ~x281 & n2251 ) | ( ~x281 & n2252 ) | ( n2251 & n2252 ) ;
  assign n2255 = ( ~n656 & n2253 ) | ( ~n656 & n2254 ) | ( n2253 & n2254 ) ;
  assign n2256 = x268 & ~n991 ;
  assign n2257 = x268 & n995 ;
  assign n2258 = ( n1104 & n2256 ) | ( n1104 & n2257 ) | ( n2256 & n2257 ) ;
  assign n2259 = ( n1119 & n2256 ) | ( n1119 & n2257 ) | ( n2256 & n2257 ) ;
  assign n2260 = ( ~n1126 & n2256 ) | ( ~n1126 & n2257 ) | ( n2256 & n2257 ) ;
  assign n2261 = ( ~n1115 & n2259 ) | ( ~n1115 & n2260 ) | ( n2259 & n2260 ) ;
  assign n2262 = ( ~n975 & n2258 ) | ( ~n975 & n2261 ) | ( n2258 & n2261 ) ;
  assign n2263 = ( n1154 & n2258 ) | ( n1154 & n2261 ) | ( n2258 & n2261 ) ;
  assign n2264 = ( ~x409 & n2262 ) | ( ~x409 & n2263 ) | ( n2262 & n2263 ) ;
  assign n2265 = ( x281 & n2262 ) | ( x281 & n2263 ) | ( n2262 & n2263 ) ;
  assign n2266 = ( n656 & n2264 ) | ( n656 & n2265 ) | ( n2264 & n2265 ) ;
  assign n2267 = n2255 | n2266 ;
  assign n2268 = n2244 & ~n2267 ;
  assign n2269 = ~n2225 & n2268 ;
  assign n2270 = x139 & n1767 ;
  assign n2271 = x139 & ~n1771 ;
  assign n2272 = ( ~n1751 & n2270 ) | ( ~n1751 & n2271 ) | ( n2270 & n2271 ) ;
  assign n2273 = ( ~n1787 & n2270 ) | ( ~n1787 & n2271 ) | ( n2270 & n2271 ) ;
  assign n2274 = ( n1794 & n2270 ) | ( n1794 & n2271 ) | ( n2270 & n2271 ) ;
  assign n2275 = ( n1783 & n2273 ) | ( n1783 & n2274 ) | ( n2273 & n2274 ) ;
  assign n2276 = ( n1643 & n2272 ) | ( n1643 & n2275 ) | ( n2272 & n2275 ) ;
  assign n2277 = ( ~n1822 & n2272 ) | ( ~n1822 & n2275 ) | ( n2272 & n2275 ) ;
  assign n2278 = ( ~n1324 & n2276 ) | ( ~n1324 & n2277 ) | ( n2276 & n2277 ) ;
  assign n2279 = x11 & ~n1767 ;
  assign n2280 = x11 & n1771 ;
  assign n2281 = ( n1751 & n2279 ) | ( n1751 & n2280 ) | ( n2279 & n2280 ) ;
  assign n2282 = ( n1787 & n2279 ) | ( n1787 & n2280 ) | ( n2279 & n2280 ) ;
  assign n2283 = ( ~n1794 & n2279 ) | ( ~n1794 & n2280 ) | ( n2279 & n2280 ) ;
  assign n2284 = ( ~n1783 & n2282 ) | ( ~n1783 & n2283 ) | ( n2282 & n2283 ) ;
  assign n2285 = ( ~n1643 & n2281 ) | ( ~n1643 & n2284 ) | ( n2281 & n2284 ) ;
  assign n2286 = ( n1822 & n2281 ) | ( n1822 & n2284 ) | ( n2281 & n2284 ) ;
  assign n2287 = ( n1324 & n2285 ) | ( n1324 & n2286 ) | ( n2285 & n2286 ) ;
  assign n2288 = n2278 | n2287 ;
  assign n2289 = x395 & n991 ;
  assign n2290 = x395 & ~n995 ;
  assign n2291 = ( ~n1104 & n2289 ) | ( ~n1104 & n2290 ) | ( n2289 & n2290 ) ;
  assign n2292 = ( ~n1119 & n2289 ) | ( ~n1119 & n2290 ) | ( n2289 & n2290 ) ;
  assign n2293 = ( n1126 & n2289 ) | ( n1126 & n2290 ) | ( n2289 & n2290 ) ;
  assign n2294 = ( n1115 & n2292 ) | ( n1115 & n2293 ) | ( n2292 & n2293 ) ;
  assign n2295 = ( n975 & n2291 ) | ( n975 & n2294 ) | ( n2291 & n2294 ) ;
  assign n2296 = ( ~n1154 & n2291 ) | ( ~n1154 & n2294 ) | ( n2291 & n2294 ) ;
  assign n2297 = ( x409 & n2295 ) | ( x409 & n2296 ) | ( n2295 & n2296 ) ;
  assign n2298 = ( ~x281 & n2295 ) | ( ~x281 & n2296 ) | ( n2295 & n2296 ) ;
  assign n2299 = ( ~n656 & n2297 ) | ( ~n656 & n2298 ) | ( n2297 & n2298 ) ;
  assign n2300 = x267 & ~n991 ;
  assign n2301 = x267 & n995 ;
  assign n2302 = ( n1104 & n2300 ) | ( n1104 & n2301 ) | ( n2300 & n2301 ) ;
  assign n2303 = ( n1119 & n2300 ) | ( n1119 & n2301 ) | ( n2300 & n2301 ) ;
  assign n2304 = ( ~n1126 & n2300 ) | ( ~n1126 & n2301 ) | ( n2300 & n2301 ) ;
  assign n2305 = ( ~n1115 & n2303 ) | ( ~n1115 & n2304 ) | ( n2303 & n2304 ) ;
  assign n2306 = ( ~n975 & n2302 ) | ( ~n975 & n2305 ) | ( n2302 & n2305 ) ;
  assign n2307 = ( n1154 & n2302 ) | ( n1154 & n2305 ) | ( n2302 & n2305 ) ;
  assign n2308 = ( ~x409 & n2306 ) | ( ~x409 & n2307 ) | ( n2306 & n2307 ) ;
  assign n2309 = ( x281 & n2306 ) | ( x281 & n2307 ) | ( n2306 & n2307 ) ;
  assign n2310 = ( n656 & n2308 ) | ( n656 & n2309 ) | ( n2308 & n2309 ) ;
  assign n2311 = n2299 | n2310 ;
  assign n2312 = x138 & n1767 ;
  assign n2313 = x138 & ~n1771 ;
  assign n2314 = ( ~n1751 & n2312 ) | ( ~n1751 & n2313 ) | ( n2312 & n2313 ) ;
  assign n2315 = ( ~n1787 & n2312 ) | ( ~n1787 & n2313 ) | ( n2312 & n2313 ) ;
  assign n2316 = ( n1794 & n2312 ) | ( n1794 & n2313 ) | ( n2312 & n2313 ) ;
  assign n2317 = ( n1783 & n2315 ) | ( n1783 & n2316 ) | ( n2315 & n2316 ) ;
  assign n2318 = ( n1643 & n2314 ) | ( n1643 & n2317 ) | ( n2314 & n2317 ) ;
  assign n2319 = ( ~n1822 & n2314 ) | ( ~n1822 & n2317 ) | ( n2314 & n2317 ) ;
  assign n2320 = ( ~n1324 & n2318 ) | ( ~n1324 & n2319 ) | ( n2318 & n2319 ) ;
  assign n2321 = x10 & ~n1767 ;
  assign n2322 = x10 & n1771 ;
  assign n2323 = ( n1751 & n2321 ) | ( n1751 & n2322 ) | ( n2321 & n2322 ) ;
  assign n2324 = ( n1787 & n2321 ) | ( n1787 & n2322 ) | ( n2321 & n2322 ) ;
  assign n2325 = ( ~n1794 & n2321 ) | ( ~n1794 & n2322 ) | ( n2321 & n2322 ) ;
  assign n2326 = ( ~n1783 & n2324 ) | ( ~n1783 & n2325 ) | ( n2324 & n2325 ) ;
  assign n2327 = ( ~n1643 & n2323 ) | ( ~n1643 & n2326 ) | ( n2323 & n2326 ) ;
  assign n2328 = ( n1822 & n2323 ) | ( n1822 & n2326 ) | ( n2323 & n2326 ) ;
  assign n2329 = ( n1324 & n2327 ) | ( n1324 & n2328 ) | ( n2327 & n2328 ) ;
  assign n2330 = n2320 | n2329 ;
  assign n2331 = x394 & n991 ;
  assign n2332 = x394 & ~n995 ;
  assign n2333 = ( ~n1104 & n2331 ) | ( ~n1104 & n2332 ) | ( n2331 & n2332 ) ;
  assign n2334 = ( ~n1119 & n2331 ) | ( ~n1119 & n2332 ) | ( n2331 & n2332 ) ;
  assign n2335 = ( n1126 & n2331 ) | ( n1126 & n2332 ) | ( n2331 & n2332 ) ;
  assign n2336 = ( n1115 & n2334 ) | ( n1115 & n2335 ) | ( n2334 & n2335 ) ;
  assign n2337 = ( n975 & n2333 ) | ( n975 & n2336 ) | ( n2333 & n2336 ) ;
  assign n2338 = ( ~n1154 & n2333 ) | ( ~n1154 & n2336 ) | ( n2333 & n2336 ) ;
  assign n2339 = ( x409 & n2337 ) | ( x409 & n2338 ) | ( n2337 & n2338 ) ;
  assign n2340 = ( ~x281 & n2337 ) | ( ~x281 & n2338 ) | ( n2337 & n2338 ) ;
  assign n2341 = ( ~n656 & n2339 ) | ( ~n656 & n2340 ) | ( n2339 & n2340 ) ;
  assign n2342 = x266 & ~n991 ;
  assign n2343 = x266 & n995 ;
  assign n2344 = ( n1104 & n2342 ) | ( n1104 & n2343 ) | ( n2342 & n2343 ) ;
  assign n2345 = ( n1119 & n2342 ) | ( n1119 & n2343 ) | ( n2342 & n2343 ) ;
  assign n2346 = ( ~n1126 & n2342 ) | ( ~n1126 & n2343 ) | ( n2342 & n2343 ) ;
  assign n2347 = ( ~n1115 & n2345 ) | ( ~n1115 & n2346 ) | ( n2345 & n2346 ) ;
  assign n2348 = ( ~n975 & n2344 ) | ( ~n975 & n2347 ) | ( n2344 & n2347 ) ;
  assign n2349 = ( n1154 & n2344 ) | ( n1154 & n2347 ) | ( n2344 & n2347 ) ;
  assign n2350 = ( ~x409 & n2348 ) | ( ~x409 & n2349 ) | ( n2348 & n2349 ) ;
  assign n2351 = ( x281 & n2348 ) | ( x281 & n2349 ) | ( n2348 & n2349 ) ;
  assign n2352 = ( n656 & n2350 ) | ( n656 & n2351 ) | ( n2350 & n2351 ) ;
  assign n2353 = n2341 | n2352 ;
  assign n2354 = ~n2330 & n2353 ;
  assign n2355 = ( ~n2288 & n2311 ) | ( ~n2288 & n2354 ) | ( n2311 & n2354 ) ;
  assign n2356 = ~n2244 & n2267 ;
  assign n2357 = n2225 | n2356 ;
  assign n2358 = ( ~n2269 & n2355 ) | ( ~n2269 & n2357 ) | ( n2355 & n2357 ) ;
  assign n2359 = x400 & n991 ;
  assign n2360 = x400 & ~n995 ;
  assign n2361 = ( ~n1104 & n2359 ) | ( ~n1104 & n2360 ) | ( n2359 & n2360 ) ;
  assign n2362 = ( ~n1119 & n2359 ) | ( ~n1119 & n2360 ) | ( n2359 & n2360 ) ;
  assign n2363 = ( n1126 & n2359 ) | ( n1126 & n2360 ) | ( n2359 & n2360 ) ;
  assign n2364 = ( n1115 & n2362 ) | ( n1115 & n2363 ) | ( n2362 & n2363 ) ;
  assign n2365 = ( n975 & n2361 ) | ( n975 & n2364 ) | ( n2361 & n2364 ) ;
  assign n2366 = ( ~n1154 & n2361 ) | ( ~n1154 & n2364 ) | ( n2361 & n2364 ) ;
  assign n2367 = ( x409 & n2365 ) | ( x409 & n2366 ) | ( n2365 & n2366 ) ;
  assign n2368 = ( ~x281 & n2365 ) | ( ~x281 & n2366 ) | ( n2365 & n2366 ) ;
  assign n2369 = ( ~n656 & n2367 ) | ( ~n656 & n2368 ) | ( n2367 & n2368 ) ;
  assign n2370 = x272 & ~n991 ;
  assign n2371 = x272 & n995 ;
  assign n2372 = ( n1104 & n2370 ) | ( n1104 & n2371 ) | ( n2370 & n2371 ) ;
  assign n2373 = ( n1119 & n2370 ) | ( n1119 & n2371 ) | ( n2370 & n2371 ) ;
  assign n2374 = ( ~n1126 & n2370 ) | ( ~n1126 & n2371 ) | ( n2370 & n2371 ) ;
  assign n2375 = ( ~n1115 & n2373 ) | ( ~n1115 & n2374 ) | ( n2373 & n2374 ) ;
  assign n2376 = ( ~n975 & n2372 ) | ( ~n975 & n2375 ) | ( n2372 & n2375 ) ;
  assign n2377 = ( n1154 & n2372 ) | ( n1154 & n2375 ) | ( n2372 & n2375 ) ;
  assign n2378 = ( ~x409 & n2376 ) | ( ~x409 & n2377 ) | ( n2376 & n2377 ) ;
  assign n2379 = ( x281 & n2376 ) | ( x281 & n2377 ) | ( n2376 & n2377 ) ;
  assign n2380 = ( n656 & n2378 ) | ( n656 & n2379 ) | ( n2378 & n2379 ) ;
  assign n2381 = n2369 | n2380 ;
  assign n2382 = x143 & n1767 ;
  assign n2383 = x143 & ~n1771 ;
  assign n2384 = ( ~n1751 & n2382 ) | ( ~n1751 & n2383 ) | ( n2382 & n2383 ) ;
  assign n2385 = ( ~n1787 & n2382 ) | ( ~n1787 & n2383 ) | ( n2382 & n2383 ) ;
  assign n2386 = ( n1794 & n2382 ) | ( n1794 & n2383 ) | ( n2382 & n2383 ) ;
  assign n2387 = ( n1783 & n2385 ) | ( n1783 & n2386 ) | ( n2385 & n2386 ) ;
  assign n2388 = ( n1643 & n2384 ) | ( n1643 & n2387 ) | ( n2384 & n2387 ) ;
  assign n2389 = ( ~n1822 & n2384 ) | ( ~n1822 & n2387 ) | ( n2384 & n2387 ) ;
  assign n2390 = ( ~n1324 & n2388 ) | ( ~n1324 & n2389 ) | ( n2388 & n2389 ) ;
  assign n2391 = x15 & ~n1767 ;
  assign n2392 = x15 & n1771 ;
  assign n2393 = ( n1751 & n2391 ) | ( n1751 & n2392 ) | ( n2391 & n2392 ) ;
  assign n2394 = ( n1787 & n2391 ) | ( n1787 & n2392 ) | ( n2391 & n2392 ) ;
  assign n2395 = ( ~n1794 & n2391 ) | ( ~n1794 & n2392 ) | ( n2391 & n2392 ) ;
  assign n2396 = ( ~n1783 & n2394 ) | ( ~n1783 & n2395 ) | ( n2394 & n2395 ) ;
  assign n2397 = ( ~n1643 & n2393 ) | ( ~n1643 & n2396 ) | ( n2393 & n2396 ) ;
  assign n2398 = ( n1822 & n2393 ) | ( n1822 & n2396 ) | ( n2393 & n2396 ) ;
  assign n2399 = ( n1324 & n2397 ) | ( n1324 & n2398 ) | ( n2397 & n2398 ) ;
  assign n2400 = n2390 | n2399 ;
  assign n2401 = x399 & n991 ;
  assign n2402 = x399 & ~n995 ;
  assign n2403 = ( ~n1104 & n2401 ) | ( ~n1104 & n2402 ) | ( n2401 & n2402 ) ;
  assign n2404 = ( ~n1119 & n2401 ) | ( ~n1119 & n2402 ) | ( n2401 & n2402 ) ;
  assign n2405 = ( n1126 & n2401 ) | ( n1126 & n2402 ) | ( n2401 & n2402 ) ;
  assign n2406 = ( n1115 & n2404 ) | ( n1115 & n2405 ) | ( n2404 & n2405 ) ;
  assign n2407 = ( n975 & n2403 ) | ( n975 & n2406 ) | ( n2403 & n2406 ) ;
  assign n2408 = ( ~n1154 & n2403 ) | ( ~n1154 & n2406 ) | ( n2403 & n2406 ) ;
  assign n2409 = ( x409 & n2407 ) | ( x409 & n2408 ) | ( n2407 & n2408 ) ;
  assign n2410 = ( ~x281 & n2407 ) | ( ~x281 & n2408 ) | ( n2407 & n2408 ) ;
  assign n2411 = ( ~n656 & n2409 ) | ( ~n656 & n2410 ) | ( n2409 & n2410 ) ;
  assign n2412 = x271 & ~n991 ;
  assign n2413 = x271 & n995 ;
  assign n2414 = ( n1104 & n2412 ) | ( n1104 & n2413 ) | ( n2412 & n2413 ) ;
  assign n2415 = ( n1119 & n2412 ) | ( n1119 & n2413 ) | ( n2412 & n2413 ) ;
  assign n2416 = ( ~n1126 & n2412 ) | ( ~n1126 & n2413 ) | ( n2412 & n2413 ) ;
  assign n2417 = ( ~n1115 & n2415 ) | ( ~n1115 & n2416 ) | ( n2415 & n2416 ) ;
  assign n2418 = ( ~n975 & n2414 ) | ( ~n975 & n2417 ) | ( n2414 & n2417 ) ;
  assign n2419 = ( n1154 & n2414 ) | ( n1154 & n2417 ) | ( n2414 & n2417 ) ;
  assign n2420 = ( ~x409 & n2418 ) | ( ~x409 & n2419 ) | ( n2418 & n2419 ) ;
  assign n2421 = ( x281 & n2418 ) | ( x281 & n2419 ) | ( n2418 & n2419 ) ;
  assign n2422 = ( n656 & n2420 ) | ( n656 & n2421 ) | ( n2420 & n2421 ) ;
  assign n2423 = n2411 | n2422 ;
  assign n2424 = ~n2400 & n2423 ;
  assign n2425 = x142 & n1767 ;
  assign n2426 = x142 & ~n1771 ;
  assign n2427 = ( ~n1751 & n2425 ) | ( ~n1751 & n2426 ) | ( n2425 & n2426 ) ;
  assign n2428 = ( ~n1787 & n2425 ) | ( ~n1787 & n2426 ) | ( n2425 & n2426 ) ;
  assign n2429 = ( n1794 & n2425 ) | ( n1794 & n2426 ) | ( n2425 & n2426 ) ;
  assign n2430 = ( n1783 & n2428 ) | ( n1783 & n2429 ) | ( n2428 & n2429 ) ;
  assign n2431 = ( n1643 & n2427 ) | ( n1643 & n2430 ) | ( n2427 & n2430 ) ;
  assign n2432 = ( ~n1822 & n2427 ) | ( ~n1822 & n2430 ) | ( n2427 & n2430 ) ;
  assign n2433 = ( ~n1324 & n2431 ) | ( ~n1324 & n2432 ) | ( n2431 & n2432 ) ;
  assign n2434 = x14 & ~n1767 ;
  assign n2435 = x14 & n1771 ;
  assign n2436 = ( n1751 & n2434 ) | ( n1751 & n2435 ) | ( n2434 & n2435 ) ;
  assign n2437 = ( n1787 & n2434 ) | ( n1787 & n2435 ) | ( n2434 & n2435 ) ;
  assign n2438 = ( ~n1794 & n2434 ) | ( ~n1794 & n2435 ) | ( n2434 & n2435 ) ;
  assign n2439 = ( ~n1783 & n2437 ) | ( ~n1783 & n2438 ) | ( n2437 & n2438 ) ;
  assign n2440 = ( ~n1643 & n2436 ) | ( ~n1643 & n2439 ) | ( n2436 & n2439 ) ;
  assign n2441 = ( n1822 & n2436 ) | ( n1822 & n2439 ) | ( n2436 & n2439 ) ;
  assign n2442 = ( n1324 & n2440 ) | ( n1324 & n2441 ) | ( n2440 & n2441 ) ;
  assign n2443 = n2433 | n2442 ;
  assign n2444 = x398 & n991 ;
  assign n2445 = x398 & ~n995 ;
  assign n2446 = ( ~n1104 & n2444 ) | ( ~n1104 & n2445 ) | ( n2444 & n2445 ) ;
  assign n2447 = ( ~n1119 & n2444 ) | ( ~n1119 & n2445 ) | ( n2444 & n2445 ) ;
  assign n2448 = ( n1126 & n2444 ) | ( n1126 & n2445 ) | ( n2444 & n2445 ) ;
  assign n2449 = ( n1115 & n2447 ) | ( n1115 & n2448 ) | ( n2447 & n2448 ) ;
  assign n2450 = ( n975 & n2446 ) | ( n975 & n2449 ) | ( n2446 & n2449 ) ;
  assign n2451 = ( ~n1154 & n2446 ) | ( ~n1154 & n2449 ) | ( n2446 & n2449 ) ;
  assign n2452 = ( x409 & n2450 ) | ( x409 & n2451 ) | ( n2450 & n2451 ) ;
  assign n2453 = ( ~x281 & n2450 ) | ( ~x281 & n2451 ) | ( n2450 & n2451 ) ;
  assign n2454 = ( ~n656 & n2452 ) | ( ~n656 & n2453 ) | ( n2452 & n2453 ) ;
  assign n2455 = x270 & ~n991 ;
  assign n2456 = x270 & n995 ;
  assign n2457 = ( n1104 & n2455 ) | ( n1104 & n2456 ) | ( n2455 & n2456 ) ;
  assign n2458 = ( n1119 & n2455 ) | ( n1119 & n2456 ) | ( n2455 & n2456 ) ;
  assign n2459 = ( ~n1126 & n2455 ) | ( ~n1126 & n2456 ) | ( n2455 & n2456 ) ;
  assign n2460 = ( ~n1115 & n2458 ) | ( ~n1115 & n2459 ) | ( n2458 & n2459 ) ;
  assign n2461 = ( ~n975 & n2457 ) | ( ~n975 & n2460 ) | ( n2457 & n2460 ) ;
  assign n2462 = ( n1154 & n2457 ) | ( n1154 & n2460 ) | ( n2457 & n2460 ) ;
  assign n2463 = ( ~x409 & n2461 ) | ( ~x409 & n2462 ) | ( n2461 & n2462 ) ;
  assign n2464 = ( x281 & n2461 ) | ( x281 & n2462 ) | ( n2461 & n2462 ) ;
  assign n2465 = ( n656 & n2463 ) | ( n656 & n2464 ) | ( n2463 & n2464 ) ;
  assign n2466 = n2454 | n2465 ;
  assign n2467 = ~n2443 & n2466 ;
  assign n2468 = n2201 & ~n2224 ;
  assign n2469 = ~n2467 & n2468 ;
  assign n2470 = n2443 & ~n2466 ;
  assign n2471 = ~n2424 & n2470 ;
  assign n2472 = ( ~n2424 & n2469 ) | ( ~n2424 & n2471 ) | ( n2469 & n2471 ) ;
  assign n2473 = n2400 & ~n2423 ;
  assign n2474 = x144 & n1767 ;
  assign n2475 = x144 & ~n1771 ;
  assign n2476 = ( ~n1751 & n2474 ) | ( ~n1751 & n2475 ) | ( n2474 & n2475 ) ;
  assign n2477 = ( ~n1787 & n2474 ) | ( ~n1787 & n2475 ) | ( n2474 & n2475 ) ;
  assign n2478 = ( n1794 & n2474 ) | ( n1794 & n2475 ) | ( n2474 & n2475 ) ;
  assign n2479 = ( n1783 & n2477 ) | ( n1783 & n2478 ) | ( n2477 & n2478 ) ;
  assign n2480 = ( n1643 & n2476 ) | ( n1643 & n2479 ) | ( n2476 & n2479 ) ;
  assign n2481 = ( ~n1822 & n2476 ) | ( ~n1822 & n2479 ) | ( n2476 & n2479 ) ;
  assign n2482 = ( ~n1324 & n2480 ) | ( ~n1324 & n2481 ) | ( n2480 & n2481 ) ;
  assign n2483 = x16 & ~n1767 ;
  assign n2484 = x16 & n1771 ;
  assign n2485 = ( n1751 & n2483 ) | ( n1751 & n2484 ) | ( n2483 & n2484 ) ;
  assign n2486 = ( n1787 & n2483 ) | ( n1787 & n2484 ) | ( n2483 & n2484 ) ;
  assign n2487 = ( ~n1794 & n2483 ) | ( ~n1794 & n2484 ) | ( n2483 & n2484 ) ;
  assign n2488 = ( ~n1783 & n2486 ) | ( ~n1783 & n2487 ) | ( n2486 & n2487 ) ;
  assign n2489 = ( ~n1643 & n2485 ) | ( ~n1643 & n2488 ) | ( n2485 & n2488 ) ;
  assign n2490 = ( n1822 & n2485 ) | ( n1822 & n2488 ) | ( n2485 & n2488 ) ;
  assign n2491 = ( n1324 & n2489 ) | ( n1324 & n2490 ) | ( n2489 & n2490 ) ;
  assign n2492 = n2482 | n2491 ;
  assign n2493 = ~n2381 & n2492 ;
  assign n2494 = ( ~n2381 & n2473 ) | ( ~n2381 & n2493 ) | ( n2473 & n2493 ) ;
  assign n2495 = ( ~n2381 & n2472 ) | ( ~n2381 & n2494 ) | ( n2472 & n2494 ) ;
  assign n2496 = n2467 & ~n2470 ;
  assign n2497 = n2424 | n2496 ;
  assign n2498 = ( n2381 & ~n2494 ) | ( n2381 & n2497 ) | ( ~n2494 & n2497 ) ;
  assign n2499 = ( n2358 & ~n2495 ) | ( n2358 & n2498 ) | ( ~n2495 & n2498 ) ;
  assign n2500 = n2424 & ~n2473 ;
  assign n2501 = ( ~n2473 & n2496 ) | ( ~n2473 & n2500 ) | ( n2496 & n2500 ) ;
  assign n2502 = ( n2381 & ~n2493 ) | ( n2381 & n2501 ) | ( ~n2493 & n2501 ) ;
  assign n2503 = n2381 & ~n2493 ;
  assign n2504 = ( n2471 & n2494 ) | ( n2471 & ~n2503 ) | ( n2494 & ~n2503 ) ;
  assign n2505 = n2330 & ~n2353 ;
  assign n2506 = ~n2288 & n2311 ;
  assign n2507 = n2505 & ~n2506 ;
  assign n2508 = n2288 & ~n2311 ;
  assign n2509 = ~n2356 & n2508 ;
  assign n2510 = ( ~n2356 & n2507 ) | ( ~n2356 & n2509 ) | ( n2507 & n2509 ) ;
  assign n2511 = n2269 | n2468 ;
  assign n2512 = n2225 & ~n2468 ;
  assign n2513 = ( n2510 & n2511 ) | ( n2510 & ~n2512 ) | ( n2511 & ~n2512 ) ;
  assign n2514 = ( ~n2502 & n2504 ) | ( ~n2502 & n2513 ) | ( n2504 & n2513 ) ;
  assign n2515 = x393 & n991 ;
  assign n2516 = x393 & ~n995 ;
  assign n2517 = ( ~n1104 & n2515 ) | ( ~n1104 & n2516 ) | ( n2515 & n2516 ) ;
  assign n2518 = ( ~n1119 & n2515 ) | ( ~n1119 & n2516 ) | ( n2515 & n2516 ) ;
  assign n2519 = ( n1126 & n2515 ) | ( n1126 & n2516 ) | ( n2515 & n2516 ) ;
  assign n2520 = ( n1115 & n2518 ) | ( n1115 & n2519 ) | ( n2518 & n2519 ) ;
  assign n2521 = ( n975 & n2517 ) | ( n975 & n2520 ) | ( n2517 & n2520 ) ;
  assign n2522 = ( ~n1154 & n2517 ) | ( ~n1154 & n2520 ) | ( n2517 & n2520 ) ;
  assign n2523 = ( x409 & n2521 ) | ( x409 & n2522 ) | ( n2521 & n2522 ) ;
  assign n2524 = ( ~x281 & n2521 ) | ( ~x281 & n2522 ) | ( n2521 & n2522 ) ;
  assign n2525 = ( ~n656 & n2523 ) | ( ~n656 & n2524 ) | ( n2523 & n2524 ) ;
  assign n2526 = x265 & ~n991 ;
  assign n2527 = x265 & n995 ;
  assign n2528 = ( n1104 & n2526 ) | ( n1104 & n2527 ) | ( n2526 & n2527 ) ;
  assign n2529 = ( n1119 & n2526 ) | ( n1119 & n2527 ) | ( n2526 & n2527 ) ;
  assign n2530 = ( ~n1126 & n2526 ) | ( ~n1126 & n2527 ) | ( n2526 & n2527 ) ;
  assign n2531 = ( ~n1115 & n2529 ) | ( ~n1115 & n2530 ) | ( n2529 & n2530 ) ;
  assign n2532 = ( ~n975 & n2528 ) | ( ~n975 & n2531 ) | ( n2528 & n2531 ) ;
  assign n2533 = ( n1154 & n2528 ) | ( n1154 & n2531 ) | ( n2528 & n2531 ) ;
  assign n2534 = ( ~x409 & n2532 ) | ( ~x409 & n2533 ) | ( n2532 & n2533 ) ;
  assign n2535 = ( x281 & n2532 ) | ( x281 & n2533 ) | ( n2532 & n2533 ) ;
  assign n2536 = ( n656 & n2534 ) | ( n656 & n2535 ) | ( n2534 & n2535 ) ;
  assign n2537 = n2525 | n2536 ;
  assign n2538 = ( n2499 & ~n2514 ) | ( n2499 & n2537 ) | ( ~n2514 & n2537 ) ;
  assign n2539 = x137 & n1767 ;
  assign n2540 = x137 & ~n1771 ;
  assign n2541 = ( ~n1751 & n2539 ) | ( ~n1751 & n2540 ) | ( n2539 & n2540 ) ;
  assign n2542 = ( ~n1787 & n2539 ) | ( ~n1787 & n2540 ) | ( n2539 & n2540 ) ;
  assign n2543 = ( n1794 & n2539 ) | ( n1794 & n2540 ) | ( n2539 & n2540 ) ;
  assign n2544 = ( n1783 & n2542 ) | ( n1783 & n2543 ) | ( n2542 & n2543 ) ;
  assign n2545 = ( n1643 & n2541 ) | ( n1643 & n2544 ) | ( n2541 & n2544 ) ;
  assign n2546 = ( ~n1822 & n2541 ) | ( ~n1822 & n2544 ) | ( n2541 & n2544 ) ;
  assign n2547 = ( ~n1324 & n2545 ) | ( ~n1324 & n2546 ) | ( n2545 & n2546 ) ;
  assign n2548 = x9 & ~n1767 ;
  assign n2549 = x9 & n1771 ;
  assign n2550 = ( n1751 & n2548 ) | ( n1751 & n2549 ) | ( n2548 & n2549 ) ;
  assign n2551 = ( n1787 & n2548 ) | ( n1787 & n2549 ) | ( n2548 & n2549 ) ;
  assign n2552 = ( ~n1794 & n2548 ) | ( ~n1794 & n2549 ) | ( n2548 & n2549 ) ;
  assign n2553 = ( ~n1783 & n2551 ) | ( ~n1783 & n2552 ) | ( n2551 & n2552 ) ;
  assign n2554 = ( ~n1643 & n2550 ) | ( ~n1643 & n2553 ) | ( n2550 & n2553 ) ;
  assign n2555 = ( n1822 & n2550 ) | ( n1822 & n2553 ) | ( n2550 & n2553 ) ;
  assign n2556 = ( n1324 & n2554 ) | ( n1324 & n2555 ) | ( n2554 & n2555 ) ;
  assign n2557 = n2547 | n2556 ;
  assign n2558 = ( ~n2499 & n2514 ) | ( ~n2499 & n2557 ) | ( n2514 & n2557 ) ;
  assign n2559 = ( n2182 & ~n2538 ) | ( n2182 & n2558 ) | ( ~n2538 & n2558 ) ;
  assign n2560 = n2492 & ~n2501 ;
  assign n2561 = n2400 & n2492 ;
  assign n2562 = ~n2423 & n2561 ;
  assign n2563 = ( n2471 & n2492 ) | ( n2471 & n2562 ) | ( n2492 & n2562 ) ;
  assign n2564 = ( n2513 & n2560 ) | ( n2513 & n2563 ) | ( n2560 & n2563 ) ;
  assign n2565 = ( n2472 & n2492 ) | ( n2472 & n2562 ) | ( n2492 & n2562 ) ;
  assign n2566 = ( ~n2424 & n2492 ) | ( ~n2424 & n2562 ) | ( n2492 & n2562 ) ;
  assign n2567 = n2492 & n2562 ;
  assign n2568 = ( ~n2496 & n2566 ) | ( ~n2496 & n2567 ) | ( n2566 & n2567 ) ;
  assign n2569 = ( ~n2358 & n2565 ) | ( ~n2358 & n2568 ) | ( n2565 & n2568 ) ;
  assign n2570 = ( ~n2537 & n2564 ) | ( ~n2537 & n2569 ) | ( n2564 & n2569 ) ;
  assign n2571 = ( n2557 & n2564 ) | ( n2557 & n2569 ) | ( n2564 & n2569 ) ;
  assign n2572 = ( n2182 & n2570 ) | ( n2182 & n2571 ) | ( n2570 & n2571 ) ;
  assign n2573 = n2559 | n2572 ;
  assign n2574 = x149 & n1767 ;
  assign n2575 = x149 & ~n1771 ;
  assign n2576 = ( ~n1751 & n2574 ) | ( ~n1751 & n2575 ) | ( n2574 & n2575 ) ;
  assign n2577 = ( ~n1787 & n2574 ) | ( ~n1787 & n2575 ) | ( n2574 & n2575 ) ;
  assign n2578 = ( n1794 & n2574 ) | ( n1794 & n2575 ) | ( n2574 & n2575 ) ;
  assign n2579 = ( n1783 & n2577 ) | ( n1783 & n2578 ) | ( n2577 & n2578 ) ;
  assign n2580 = ( n1643 & n2576 ) | ( n1643 & n2579 ) | ( n2576 & n2579 ) ;
  assign n2581 = ( ~n1822 & n2576 ) | ( ~n1822 & n2579 ) | ( n2576 & n2579 ) ;
  assign n2582 = ( ~n1324 & n2580 ) | ( ~n1324 & n2581 ) | ( n2580 & n2581 ) ;
  assign n2583 = x21 & ~n1767 ;
  assign n2584 = x21 & n1771 ;
  assign n2585 = ( n1751 & n2583 ) | ( n1751 & n2584 ) | ( n2583 & n2584 ) ;
  assign n2586 = ( n1787 & n2583 ) | ( n1787 & n2584 ) | ( n2583 & n2584 ) ;
  assign n2587 = ( ~n1794 & n2583 ) | ( ~n1794 & n2584 ) | ( n2583 & n2584 ) ;
  assign n2588 = ( ~n1783 & n2586 ) | ( ~n1783 & n2587 ) | ( n2586 & n2587 ) ;
  assign n2589 = ( ~n1643 & n2585 ) | ( ~n1643 & n2588 ) | ( n2585 & n2588 ) ;
  assign n2590 = ( n1822 & n2585 ) | ( n1822 & n2588 ) | ( n2585 & n2588 ) ;
  assign n2591 = ( n1324 & n2589 ) | ( n1324 & n2590 ) | ( n2589 & n2590 ) ;
  assign n2592 = n2582 | n2591 ;
  assign n2593 = x405 & n991 ;
  assign n2594 = x405 & ~n995 ;
  assign n2595 = ( ~n1104 & n2593 ) | ( ~n1104 & n2594 ) | ( n2593 & n2594 ) ;
  assign n2596 = ( ~n1119 & n2593 ) | ( ~n1119 & n2594 ) | ( n2593 & n2594 ) ;
  assign n2597 = ( n1126 & n2593 ) | ( n1126 & n2594 ) | ( n2593 & n2594 ) ;
  assign n2598 = ( n1115 & n2596 ) | ( n1115 & n2597 ) | ( n2596 & n2597 ) ;
  assign n2599 = ( n975 & n2595 ) | ( n975 & n2598 ) | ( n2595 & n2598 ) ;
  assign n2600 = ( ~n1154 & n2595 ) | ( ~n1154 & n2598 ) | ( n2595 & n2598 ) ;
  assign n2601 = ( x409 & n2599 ) | ( x409 & n2600 ) | ( n2599 & n2600 ) ;
  assign n2602 = ( ~x281 & n2599 ) | ( ~x281 & n2600 ) | ( n2599 & n2600 ) ;
  assign n2603 = ( ~n656 & n2601 ) | ( ~n656 & n2602 ) | ( n2601 & n2602 ) ;
  assign n2604 = x277 & ~n991 ;
  assign n2605 = x277 & n995 ;
  assign n2606 = ( n1104 & n2604 ) | ( n1104 & n2605 ) | ( n2604 & n2605 ) ;
  assign n2607 = ( n1119 & n2604 ) | ( n1119 & n2605 ) | ( n2604 & n2605 ) ;
  assign n2608 = ( ~n1126 & n2604 ) | ( ~n1126 & n2605 ) | ( n2604 & n2605 ) ;
  assign n2609 = ( ~n1115 & n2607 ) | ( ~n1115 & n2608 ) | ( n2607 & n2608 ) ;
  assign n2610 = ( ~n975 & n2606 ) | ( ~n975 & n2609 ) | ( n2606 & n2609 ) ;
  assign n2611 = ( n1154 & n2606 ) | ( n1154 & n2609 ) | ( n2606 & n2609 ) ;
  assign n2612 = ( ~x409 & n2610 ) | ( ~x409 & n2611 ) | ( n2610 & n2611 ) ;
  assign n2613 = ( x281 & n2610 ) | ( x281 & n2611 ) | ( n2610 & n2611 ) ;
  assign n2614 = ( n656 & n2612 ) | ( n656 & n2613 ) | ( n2612 & n2613 ) ;
  assign n2615 = n2603 | n2614 ;
  assign n2616 = ~n2592 & n2615 ;
  assign n2617 = x148 & n1767 ;
  assign n2618 = x148 & ~n1771 ;
  assign n2619 = ( ~n1751 & n2617 ) | ( ~n1751 & n2618 ) | ( n2617 & n2618 ) ;
  assign n2620 = ( ~n1787 & n2617 ) | ( ~n1787 & n2618 ) | ( n2617 & n2618 ) ;
  assign n2621 = ( n1794 & n2617 ) | ( n1794 & n2618 ) | ( n2617 & n2618 ) ;
  assign n2622 = ( n1783 & n2620 ) | ( n1783 & n2621 ) | ( n2620 & n2621 ) ;
  assign n2623 = ( n1643 & n2619 ) | ( n1643 & n2622 ) | ( n2619 & n2622 ) ;
  assign n2624 = ( ~n1822 & n2619 ) | ( ~n1822 & n2622 ) | ( n2619 & n2622 ) ;
  assign n2625 = ( ~n1324 & n2623 ) | ( ~n1324 & n2624 ) | ( n2623 & n2624 ) ;
  assign n2626 = x20 & ~n1767 ;
  assign n2627 = x20 & n1771 ;
  assign n2628 = ( n1751 & n2626 ) | ( n1751 & n2627 ) | ( n2626 & n2627 ) ;
  assign n2629 = ( n1787 & n2626 ) | ( n1787 & n2627 ) | ( n2626 & n2627 ) ;
  assign n2630 = ( ~n1794 & n2626 ) | ( ~n1794 & n2627 ) | ( n2626 & n2627 ) ;
  assign n2631 = ( ~n1783 & n2629 ) | ( ~n1783 & n2630 ) | ( n2629 & n2630 ) ;
  assign n2632 = ( ~n1643 & n2628 ) | ( ~n1643 & n2631 ) | ( n2628 & n2631 ) ;
  assign n2633 = ( n1822 & n2628 ) | ( n1822 & n2631 ) | ( n2628 & n2631 ) ;
  assign n2634 = ( n1324 & n2632 ) | ( n1324 & n2633 ) | ( n2632 & n2633 ) ;
  assign n2635 = n2625 | n2634 ;
  assign n2636 = x404 & n991 ;
  assign n2637 = x404 & ~n995 ;
  assign n2638 = ( ~n1104 & n2636 ) | ( ~n1104 & n2637 ) | ( n2636 & n2637 ) ;
  assign n2639 = ( ~n1119 & n2636 ) | ( ~n1119 & n2637 ) | ( n2636 & n2637 ) ;
  assign n2640 = ( n1126 & n2636 ) | ( n1126 & n2637 ) | ( n2636 & n2637 ) ;
  assign n2641 = ( n1115 & n2639 ) | ( n1115 & n2640 ) | ( n2639 & n2640 ) ;
  assign n2642 = ( n975 & n2638 ) | ( n975 & n2641 ) | ( n2638 & n2641 ) ;
  assign n2643 = ( ~n1154 & n2638 ) | ( ~n1154 & n2641 ) | ( n2638 & n2641 ) ;
  assign n2644 = ( x409 & n2642 ) | ( x409 & n2643 ) | ( n2642 & n2643 ) ;
  assign n2645 = ( ~x281 & n2642 ) | ( ~x281 & n2643 ) | ( n2642 & n2643 ) ;
  assign n2646 = ( ~n656 & n2644 ) | ( ~n656 & n2645 ) | ( n2644 & n2645 ) ;
  assign n2647 = x276 & ~n991 ;
  assign n2648 = x276 & n995 ;
  assign n2649 = ( n1104 & n2647 ) | ( n1104 & n2648 ) | ( n2647 & n2648 ) ;
  assign n2650 = ( n1119 & n2647 ) | ( n1119 & n2648 ) | ( n2647 & n2648 ) ;
  assign n2651 = ( ~n1126 & n2647 ) | ( ~n1126 & n2648 ) | ( n2647 & n2648 ) ;
  assign n2652 = ( ~n1115 & n2650 ) | ( ~n1115 & n2651 ) | ( n2650 & n2651 ) ;
  assign n2653 = ( ~n975 & n2649 ) | ( ~n975 & n2652 ) | ( n2649 & n2652 ) ;
  assign n2654 = ( n1154 & n2649 ) | ( n1154 & n2652 ) | ( n2649 & n2652 ) ;
  assign n2655 = ( ~x409 & n2653 ) | ( ~x409 & n2654 ) | ( n2653 & n2654 ) ;
  assign n2656 = ( x281 & n2653 ) | ( x281 & n2654 ) | ( n2653 & n2654 ) ;
  assign n2657 = ( n656 & n2655 ) | ( n656 & n2656 ) | ( n2655 & n2656 ) ;
  assign n2658 = n2646 | n2657 ;
  assign n2659 = n2635 & ~n2658 ;
  assign n2660 = ~n2616 & n2659 ;
  assign n2661 = x147 & n1767 ;
  assign n2662 = x147 & ~n1771 ;
  assign n2663 = ( ~n1751 & n2661 ) | ( ~n1751 & n2662 ) | ( n2661 & n2662 ) ;
  assign n2664 = ( ~n1787 & n2661 ) | ( ~n1787 & n2662 ) | ( n2661 & n2662 ) ;
  assign n2665 = ( n1794 & n2661 ) | ( n1794 & n2662 ) | ( n2661 & n2662 ) ;
  assign n2666 = ( n1783 & n2664 ) | ( n1783 & n2665 ) | ( n2664 & n2665 ) ;
  assign n2667 = ( n1643 & n2663 ) | ( n1643 & n2666 ) | ( n2663 & n2666 ) ;
  assign n2668 = ( ~n1822 & n2663 ) | ( ~n1822 & n2666 ) | ( n2663 & n2666 ) ;
  assign n2669 = ( ~n1324 & n2667 ) | ( ~n1324 & n2668 ) | ( n2667 & n2668 ) ;
  assign n2670 = x19 & ~n1767 ;
  assign n2671 = x19 & n1771 ;
  assign n2672 = ( n1751 & n2670 ) | ( n1751 & n2671 ) | ( n2670 & n2671 ) ;
  assign n2673 = ( n1787 & n2670 ) | ( n1787 & n2671 ) | ( n2670 & n2671 ) ;
  assign n2674 = ( ~n1794 & n2670 ) | ( ~n1794 & n2671 ) | ( n2670 & n2671 ) ;
  assign n2675 = ( ~n1783 & n2673 ) | ( ~n1783 & n2674 ) | ( n2673 & n2674 ) ;
  assign n2676 = ( ~n1643 & n2672 ) | ( ~n1643 & n2675 ) | ( n2672 & n2675 ) ;
  assign n2677 = ( n1822 & n2672 ) | ( n1822 & n2675 ) | ( n2672 & n2675 ) ;
  assign n2678 = ( n1324 & n2676 ) | ( n1324 & n2677 ) | ( n2676 & n2677 ) ;
  assign n2679 = n2669 | n2678 ;
  assign n2680 = x403 & n991 ;
  assign n2681 = x403 & ~n995 ;
  assign n2682 = ( ~n1104 & n2680 ) | ( ~n1104 & n2681 ) | ( n2680 & n2681 ) ;
  assign n2683 = ( ~n1119 & n2680 ) | ( ~n1119 & n2681 ) | ( n2680 & n2681 ) ;
  assign n2684 = ( n1126 & n2680 ) | ( n1126 & n2681 ) | ( n2680 & n2681 ) ;
  assign n2685 = ( n1115 & n2683 ) | ( n1115 & n2684 ) | ( n2683 & n2684 ) ;
  assign n2686 = ( n975 & n2682 ) | ( n975 & n2685 ) | ( n2682 & n2685 ) ;
  assign n2687 = ( ~n1154 & n2682 ) | ( ~n1154 & n2685 ) | ( n2682 & n2685 ) ;
  assign n2688 = ( x409 & n2686 ) | ( x409 & n2687 ) | ( n2686 & n2687 ) ;
  assign n2689 = ( ~x281 & n2686 ) | ( ~x281 & n2687 ) | ( n2686 & n2687 ) ;
  assign n2690 = ( ~n656 & n2688 ) | ( ~n656 & n2689 ) | ( n2688 & n2689 ) ;
  assign n2691 = x275 & ~n991 ;
  assign n2692 = x275 & n995 ;
  assign n2693 = ( n1104 & n2691 ) | ( n1104 & n2692 ) | ( n2691 & n2692 ) ;
  assign n2694 = ( n1119 & n2691 ) | ( n1119 & n2692 ) | ( n2691 & n2692 ) ;
  assign n2695 = ( ~n1126 & n2691 ) | ( ~n1126 & n2692 ) | ( n2691 & n2692 ) ;
  assign n2696 = ( ~n1115 & n2694 ) | ( ~n1115 & n2695 ) | ( n2694 & n2695 ) ;
  assign n2697 = ( ~n975 & n2693 ) | ( ~n975 & n2696 ) | ( n2693 & n2696 ) ;
  assign n2698 = ( n1154 & n2693 ) | ( n1154 & n2696 ) | ( n2693 & n2696 ) ;
  assign n2699 = ( ~x409 & n2697 ) | ( ~x409 & n2698 ) | ( n2697 & n2698 ) ;
  assign n2700 = ( x281 & n2697 ) | ( x281 & n2698 ) | ( n2697 & n2698 ) ;
  assign n2701 = ( n656 & n2699 ) | ( n656 & n2700 ) | ( n2699 & n2700 ) ;
  assign n2702 = n2690 | n2701 ;
  assign n2703 = x146 & n1767 ;
  assign n2704 = x146 & ~n1771 ;
  assign n2705 = ( ~n1751 & n2703 ) | ( ~n1751 & n2704 ) | ( n2703 & n2704 ) ;
  assign n2706 = ( ~n1787 & n2703 ) | ( ~n1787 & n2704 ) | ( n2703 & n2704 ) ;
  assign n2707 = ( n1794 & n2703 ) | ( n1794 & n2704 ) | ( n2703 & n2704 ) ;
  assign n2708 = ( n1783 & n2706 ) | ( n1783 & n2707 ) | ( n2706 & n2707 ) ;
  assign n2709 = ( n1643 & n2705 ) | ( n1643 & n2708 ) | ( n2705 & n2708 ) ;
  assign n2710 = ( ~n1822 & n2705 ) | ( ~n1822 & n2708 ) | ( n2705 & n2708 ) ;
  assign n2711 = ( ~n1324 & n2709 ) | ( ~n1324 & n2710 ) | ( n2709 & n2710 ) ;
  assign n2712 = x18 & ~n1767 ;
  assign n2713 = x18 & n1771 ;
  assign n2714 = ( n1751 & n2712 ) | ( n1751 & n2713 ) | ( n2712 & n2713 ) ;
  assign n2715 = ( n1787 & n2712 ) | ( n1787 & n2713 ) | ( n2712 & n2713 ) ;
  assign n2716 = ( ~n1794 & n2712 ) | ( ~n1794 & n2713 ) | ( n2712 & n2713 ) ;
  assign n2717 = ( ~n1783 & n2715 ) | ( ~n1783 & n2716 ) | ( n2715 & n2716 ) ;
  assign n2718 = ( ~n1643 & n2714 ) | ( ~n1643 & n2717 ) | ( n2714 & n2717 ) ;
  assign n2719 = ( n1822 & n2714 ) | ( n1822 & n2717 ) | ( n2714 & n2717 ) ;
  assign n2720 = ( n1324 & n2718 ) | ( n1324 & n2719 ) | ( n2718 & n2719 ) ;
  assign n2721 = n2711 | n2720 ;
  assign n2722 = x402 & n991 ;
  assign n2723 = x402 & ~n995 ;
  assign n2724 = ( ~n1104 & n2722 ) | ( ~n1104 & n2723 ) | ( n2722 & n2723 ) ;
  assign n2725 = ( ~n1119 & n2722 ) | ( ~n1119 & n2723 ) | ( n2722 & n2723 ) ;
  assign n2726 = ( n1126 & n2722 ) | ( n1126 & n2723 ) | ( n2722 & n2723 ) ;
  assign n2727 = ( n1115 & n2725 ) | ( n1115 & n2726 ) | ( n2725 & n2726 ) ;
  assign n2728 = ( n975 & n2724 ) | ( n975 & n2727 ) | ( n2724 & n2727 ) ;
  assign n2729 = ( ~n1154 & n2724 ) | ( ~n1154 & n2727 ) | ( n2724 & n2727 ) ;
  assign n2730 = ( x409 & n2728 ) | ( x409 & n2729 ) | ( n2728 & n2729 ) ;
  assign n2731 = ( ~x281 & n2728 ) | ( ~x281 & n2729 ) | ( n2728 & n2729 ) ;
  assign n2732 = ( ~n656 & n2730 ) | ( ~n656 & n2731 ) | ( n2730 & n2731 ) ;
  assign n2733 = x274 & ~n991 ;
  assign n2734 = x274 & n995 ;
  assign n2735 = ( n1104 & n2733 ) | ( n1104 & n2734 ) | ( n2733 & n2734 ) ;
  assign n2736 = ( n1119 & n2733 ) | ( n1119 & n2734 ) | ( n2733 & n2734 ) ;
  assign n2737 = ( ~n1126 & n2733 ) | ( ~n1126 & n2734 ) | ( n2733 & n2734 ) ;
  assign n2738 = ( ~n1115 & n2736 ) | ( ~n1115 & n2737 ) | ( n2736 & n2737 ) ;
  assign n2739 = ( ~n975 & n2735 ) | ( ~n975 & n2738 ) | ( n2735 & n2738 ) ;
  assign n2740 = ( n1154 & n2735 ) | ( n1154 & n2738 ) | ( n2735 & n2738 ) ;
  assign n2741 = ( ~x409 & n2739 ) | ( ~x409 & n2740 ) | ( n2739 & n2740 ) ;
  assign n2742 = ( x281 & n2739 ) | ( x281 & n2740 ) | ( n2739 & n2740 ) ;
  assign n2743 = ( n656 & n2741 ) | ( n656 & n2742 ) | ( n2741 & n2742 ) ;
  assign n2744 = n2732 | n2743 ;
  assign n2745 = ~n2721 & n2744 ;
  assign n2746 = ( ~n2679 & n2702 ) | ( ~n2679 & n2745 ) | ( n2702 & n2745 ) ;
  assign n2747 = ~n2635 & n2658 ;
  assign n2748 = n2616 | n2747 ;
  assign n2749 = ( ~n2660 & n2746 ) | ( ~n2660 & n2748 ) | ( n2746 & n2748 ) ;
  assign n2750 = x408 & n991 ;
  assign n2751 = x408 & ~n995 ;
  assign n2752 = ( ~n1104 & n2750 ) | ( ~n1104 & n2751 ) | ( n2750 & n2751 ) ;
  assign n2753 = ( ~n1119 & n2750 ) | ( ~n1119 & n2751 ) | ( n2750 & n2751 ) ;
  assign n2754 = ( n1126 & n2750 ) | ( n1126 & n2751 ) | ( n2750 & n2751 ) ;
  assign n2755 = ( n1115 & n2753 ) | ( n1115 & n2754 ) | ( n2753 & n2754 ) ;
  assign n2756 = ( n975 & n2752 ) | ( n975 & n2755 ) | ( n2752 & n2755 ) ;
  assign n2757 = ( ~n1154 & n2752 ) | ( ~n1154 & n2755 ) | ( n2752 & n2755 ) ;
  assign n2758 = ( x409 & n2756 ) | ( x409 & n2757 ) | ( n2756 & n2757 ) ;
  assign n2759 = ( ~x281 & n2756 ) | ( ~x281 & n2757 ) | ( n2756 & n2757 ) ;
  assign n2760 = ( ~n656 & n2758 ) | ( ~n656 & n2759 ) | ( n2758 & n2759 ) ;
  assign n2761 = x280 & ~n991 ;
  assign n2762 = x280 & n995 ;
  assign n2763 = ( n1104 & n2761 ) | ( n1104 & n2762 ) | ( n2761 & n2762 ) ;
  assign n2764 = ( n1119 & n2761 ) | ( n1119 & n2762 ) | ( n2761 & n2762 ) ;
  assign n2765 = ( ~n1126 & n2761 ) | ( ~n1126 & n2762 ) | ( n2761 & n2762 ) ;
  assign n2766 = ( ~n1115 & n2764 ) | ( ~n1115 & n2765 ) | ( n2764 & n2765 ) ;
  assign n2767 = ( ~n975 & n2763 ) | ( ~n975 & n2766 ) | ( n2763 & n2766 ) ;
  assign n2768 = ( n1154 & n2763 ) | ( n1154 & n2766 ) | ( n2763 & n2766 ) ;
  assign n2769 = ( ~x409 & n2767 ) | ( ~x409 & n2768 ) | ( n2767 & n2768 ) ;
  assign n2770 = ( x281 & n2767 ) | ( x281 & n2768 ) | ( n2767 & n2768 ) ;
  assign n2771 = ( n656 & n2769 ) | ( n656 & n2770 ) | ( n2769 & n2770 ) ;
  assign n2772 = n2760 | n2771 ;
  assign n2773 = x151 & n1767 ;
  assign n2774 = x151 & ~n1771 ;
  assign n2775 = ( ~n1751 & n2773 ) | ( ~n1751 & n2774 ) | ( n2773 & n2774 ) ;
  assign n2776 = ( ~n1787 & n2773 ) | ( ~n1787 & n2774 ) | ( n2773 & n2774 ) ;
  assign n2777 = ( n1794 & n2773 ) | ( n1794 & n2774 ) | ( n2773 & n2774 ) ;
  assign n2778 = ( n1783 & n2776 ) | ( n1783 & n2777 ) | ( n2776 & n2777 ) ;
  assign n2779 = ( n1643 & n2775 ) | ( n1643 & n2778 ) | ( n2775 & n2778 ) ;
  assign n2780 = ( ~n1822 & n2775 ) | ( ~n1822 & n2778 ) | ( n2775 & n2778 ) ;
  assign n2781 = ( ~n1324 & n2779 ) | ( ~n1324 & n2780 ) | ( n2779 & n2780 ) ;
  assign n2782 = x23 & ~n1767 ;
  assign n2783 = x23 & n1771 ;
  assign n2784 = ( n1751 & n2782 ) | ( n1751 & n2783 ) | ( n2782 & n2783 ) ;
  assign n2785 = ( n1787 & n2782 ) | ( n1787 & n2783 ) | ( n2782 & n2783 ) ;
  assign n2786 = ( ~n1794 & n2782 ) | ( ~n1794 & n2783 ) | ( n2782 & n2783 ) ;
  assign n2787 = ( ~n1783 & n2785 ) | ( ~n1783 & n2786 ) | ( n2785 & n2786 ) ;
  assign n2788 = ( ~n1643 & n2784 ) | ( ~n1643 & n2787 ) | ( n2784 & n2787 ) ;
  assign n2789 = ( n1822 & n2784 ) | ( n1822 & n2787 ) | ( n2784 & n2787 ) ;
  assign n2790 = ( n1324 & n2788 ) | ( n1324 & n2789 ) | ( n2788 & n2789 ) ;
  assign n2791 = n2781 | n2790 ;
  assign n2792 = x407 & n991 ;
  assign n2793 = x407 & ~n995 ;
  assign n2794 = ( ~n1104 & n2792 ) | ( ~n1104 & n2793 ) | ( n2792 & n2793 ) ;
  assign n2795 = ( ~n1119 & n2792 ) | ( ~n1119 & n2793 ) | ( n2792 & n2793 ) ;
  assign n2796 = ( n1126 & n2792 ) | ( n1126 & n2793 ) | ( n2792 & n2793 ) ;
  assign n2797 = ( n1115 & n2795 ) | ( n1115 & n2796 ) | ( n2795 & n2796 ) ;
  assign n2798 = ( n975 & n2794 ) | ( n975 & n2797 ) | ( n2794 & n2797 ) ;
  assign n2799 = ( ~n1154 & n2794 ) | ( ~n1154 & n2797 ) | ( n2794 & n2797 ) ;
  assign n2800 = ( x409 & n2798 ) | ( x409 & n2799 ) | ( n2798 & n2799 ) ;
  assign n2801 = ( ~x281 & n2798 ) | ( ~x281 & n2799 ) | ( n2798 & n2799 ) ;
  assign n2802 = ( ~n656 & n2800 ) | ( ~n656 & n2801 ) | ( n2800 & n2801 ) ;
  assign n2803 = x279 & ~n991 ;
  assign n2804 = x279 & n995 ;
  assign n2805 = ( n1104 & n2803 ) | ( n1104 & n2804 ) | ( n2803 & n2804 ) ;
  assign n2806 = ( n1119 & n2803 ) | ( n1119 & n2804 ) | ( n2803 & n2804 ) ;
  assign n2807 = ( ~n1126 & n2803 ) | ( ~n1126 & n2804 ) | ( n2803 & n2804 ) ;
  assign n2808 = ( ~n1115 & n2806 ) | ( ~n1115 & n2807 ) | ( n2806 & n2807 ) ;
  assign n2809 = ( ~n975 & n2805 ) | ( ~n975 & n2808 ) | ( n2805 & n2808 ) ;
  assign n2810 = ( n1154 & n2805 ) | ( n1154 & n2808 ) | ( n2805 & n2808 ) ;
  assign n2811 = ( ~x409 & n2809 ) | ( ~x409 & n2810 ) | ( n2809 & n2810 ) ;
  assign n2812 = ( x281 & n2809 ) | ( x281 & n2810 ) | ( n2809 & n2810 ) ;
  assign n2813 = ( n656 & n2811 ) | ( n656 & n2812 ) | ( n2811 & n2812 ) ;
  assign n2814 = n2802 | n2813 ;
  assign n2815 = ~n2791 & n2814 ;
  assign n2816 = x150 & n1767 ;
  assign n2817 = x150 & ~n1771 ;
  assign n2818 = ( ~n1751 & n2816 ) | ( ~n1751 & n2817 ) | ( n2816 & n2817 ) ;
  assign n2819 = ( ~n1787 & n2816 ) | ( ~n1787 & n2817 ) | ( n2816 & n2817 ) ;
  assign n2820 = ( n1794 & n2816 ) | ( n1794 & n2817 ) | ( n2816 & n2817 ) ;
  assign n2821 = ( n1783 & n2819 ) | ( n1783 & n2820 ) | ( n2819 & n2820 ) ;
  assign n2822 = ( n1643 & n2818 ) | ( n1643 & n2821 ) | ( n2818 & n2821 ) ;
  assign n2823 = ( ~n1822 & n2818 ) | ( ~n1822 & n2821 ) | ( n2818 & n2821 ) ;
  assign n2824 = ( ~n1324 & n2822 ) | ( ~n1324 & n2823 ) | ( n2822 & n2823 ) ;
  assign n2825 = x22 & ~n1767 ;
  assign n2826 = x22 & n1771 ;
  assign n2827 = ( n1751 & n2825 ) | ( n1751 & n2826 ) | ( n2825 & n2826 ) ;
  assign n2828 = ( n1787 & n2825 ) | ( n1787 & n2826 ) | ( n2825 & n2826 ) ;
  assign n2829 = ( ~n1794 & n2825 ) | ( ~n1794 & n2826 ) | ( n2825 & n2826 ) ;
  assign n2830 = ( ~n1783 & n2828 ) | ( ~n1783 & n2829 ) | ( n2828 & n2829 ) ;
  assign n2831 = ( ~n1643 & n2827 ) | ( ~n1643 & n2830 ) | ( n2827 & n2830 ) ;
  assign n2832 = ( n1822 & n2827 ) | ( n1822 & n2830 ) | ( n2827 & n2830 ) ;
  assign n2833 = ( n1324 & n2831 ) | ( n1324 & n2832 ) | ( n2831 & n2832 ) ;
  assign n2834 = n2824 | n2833 ;
  assign n2835 = x406 & n991 ;
  assign n2836 = x406 & ~n995 ;
  assign n2837 = ( ~n1104 & n2835 ) | ( ~n1104 & n2836 ) | ( n2835 & n2836 ) ;
  assign n2838 = ( ~n1119 & n2835 ) | ( ~n1119 & n2836 ) | ( n2835 & n2836 ) ;
  assign n2839 = ( n1126 & n2835 ) | ( n1126 & n2836 ) | ( n2835 & n2836 ) ;
  assign n2840 = ( n1115 & n2838 ) | ( n1115 & n2839 ) | ( n2838 & n2839 ) ;
  assign n2841 = ( n975 & n2837 ) | ( n975 & n2840 ) | ( n2837 & n2840 ) ;
  assign n2842 = ( ~n1154 & n2837 ) | ( ~n1154 & n2840 ) | ( n2837 & n2840 ) ;
  assign n2843 = ( x409 & n2841 ) | ( x409 & n2842 ) | ( n2841 & n2842 ) ;
  assign n2844 = ( ~x281 & n2841 ) | ( ~x281 & n2842 ) | ( n2841 & n2842 ) ;
  assign n2845 = ( ~n656 & n2843 ) | ( ~n656 & n2844 ) | ( n2843 & n2844 ) ;
  assign n2846 = x278 & ~n991 ;
  assign n2847 = x278 & n995 ;
  assign n2848 = ( n1104 & n2846 ) | ( n1104 & n2847 ) | ( n2846 & n2847 ) ;
  assign n2849 = ( n1119 & n2846 ) | ( n1119 & n2847 ) | ( n2846 & n2847 ) ;
  assign n2850 = ( ~n1126 & n2846 ) | ( ~n1126 & n2847 ) | ( n2846 & n2847 ) ;
  assign n2851 = ( ~n1115 & n2849 ) | ( ~n1115 & n2850 ) | ( n2849 & n2850 ) ;
  assign n2852 = ( ~n975 & n2848 ) | ( ~n975 & n2851 ) | ( n2848 & n2851 ) ;
  assign n2853 = ( n1154 & n2848 ) | ( n1154 & n2851 ) | ( n2848 & n2851 ) ;
  assign n2854 = ( ~x409 & n2852 ) | ( ~x409 & n2853 ) | ( n2852 & n2853 ) ;
  assign n2855 = ( x281 & n2852 ) | ( x281 & n2853 ) | ( n2852 & n2853 ) ;
  assign n2856 = ( n656 & n2854 ) | ( n656 & n2855 ) | ( n2854 & n2855 ) ;
  assign n2857 = n2845 | n2856 ;
  assign n2858 = ~n2834 & n2857 ;
  assign n2859 = n2592 & ~n2615 ;
  assign n2860 = ~n2858 & n2859 ;
  assign n2861 = n2834 & ~n2857 ;
  assign n2862 = ~n2815 & n2861 ;
  assign n2863 = ( ~n2815 & n2860 ) | ( ~n2815 & n2862 ) | ( n2860 & n2862 ) ;
  assign n2864 = n2791 & ~n2814 ;
  assign n2865 = x152 & n1767 ;
  assign n2866 = x152 & ~n1771 ;
  assign n2867 = ( ~n1751 & n2865 ) | ( ~n1751 & n2866 ) | ( n2865 & n2866 ) ;
  assign n2868 = ( ~n1787 & n2865 ) | ( ~n1787 & n2866 ) | ( n2865 & n2866 ) ;
  assign n2869 = ( n1794 & n2865 ) | ( n1794 & n2866 ) | ( n2865 & n2866 ) ;
  assign n2870 = ( n1783 & n2868 ) | ( n1783 & n2869 ) | ( n2868 & n2869 ) ;
  assign n2871 = ( n1643 & n2867 ) | ( n1643 & n2870 ) | ( n2867 & n2870 ) ;
  assign n2872 = ( ~n1822 & n2867 ) | ( ~n1822 & n2870 ) | ( n2867 & n2870 ) ;
  assign n2873 = ( ~n1324 & n2871 ) | ( ~n1324 & n2872 ) | ( n2871 & n2872 ) ;
  assign n2874 = x24 & ~n1767 ;
  assign n2875 = x24 & n1771 ;
  assign n2876 = ( n1751 & n2874 ) | ( n1751 & n2875 ) | ( n2874 & n2875 ) ;
  assign n2877 = ( n1787 & n2874 ) | ( n1787 & n2875 ) | ( n2874 & n2875 ) ;
  assign n2878 = ( ~n1794 & n2874 ) | ( ~n1794 & n2875 ) | ( n2874 & n2875 ) ;
  assign n2879 = ( ~n1783 & n2877 ) | ( ~n1783 & n2878 ) | ( n2877 & n2878 ) ;
  assign n2880 = ( ~n1643 & n2876 ) | ( ~n1643 & n2879 ) | ( n2876 & n2879 ) ;
  assign n2881 = ( n1822 & n2876 ) | ( n1822 & n2879 ) | ( n2876 & n2879 ) ;
  assign n2882 = ( n1324 & n2880 ) | ( n1324 & n2881 ) | ( n2880 & n2881 ) ;
  assign n2883 = n2873 | n2882 ;
  assign n2884 = ~n2772 & n2883 ;
  assign n2885 = ( ~n2772 & n2864 ) | ( ~n2772 & n2884 ) | ( n2864 & n2884 ) ;
  assign n2886 = ( ~n2772 & n2863 ) | ( ~n2772 & n2885 ) | ( n2863 & n2885 ) ;
  assign n2887 = n2858 & ~n2861 ;
  assign n2888 = n2815 | n2887 ;
  assign n2889 = ( n2772 & ~n2885 ) | ( n2772 & n2888 ) | ( ~n2885 & n2888 ) ;
  assign n2890 = ( n2749 & ~n2886 ) | ( n2749 & n2889 ) | ( ~n2886 & n2889 ) ;
  assign n2891 = n2815 & ~n2864 ;
  assign n2892 = ( ~n2864 & n2887 ) | ( ~n2864 & n2891 ) | ( n2887 & n2891 ) ;
  assign n2893 = ( n2772 & ~n2884 ) | ( n2772 & n2892 ) | ( ~n2884 & n2892 ) ;
  assign n2894 = n2772 & ~n2884 ;
  assign n2895 = ( n2862 & n2885 ) | ( n2862 & ~n2894 ) | ( n2885 & ~n2894 ) ;
  assign n2896 = n2721 & ~n2744 ;
  assign n2897 = ~n2679 & n2702 ;
  assign n2898 = n2896 & ~n2897 ;
  assign n2899 = n2679 & ~n2702 ;
  assign n2900 = ~n2747 & n2899 ;
  assign n2901 = ( ~n2747 & n2898 ) | ( ~n2747 & n2900 ) | ( n2898 & n2900 ) ;
  assign n2902 = n2660 | n2859 ;
  assign n2903 = n2616 & ~n2859 ;
  assign n2904 = ( n2901 & n2902 ) | ( n2901 & ~n2903 ) | ( n2902 & ~n2903 ) ;
  assign n2905 = ( ~n2893 & n2895 ) | ( ~n2893 & n2904 ) | ( n2895 & n2904 ) ;
  assign n2906 = x401 & n991 ;
  assign n2907 = x401 & ~n995 ;
  assign n2908 = ( ~n1104 & n2906 ) | ( ~n1104 & n2907 ) | ( n2906 & n2907 ) ;
  assign n2909 = ( ~n1119 & n2906 ) | ( ~n1119 & n2907 ) | ( n2906 & n2907 ) ;
  assign n2910 = ( n1126 & n2906 ) | ( n1126 & n2907 ) | ( n2906 & n2907 ) ;
  assign n2911 = ( n1115 & n2909 ) | ( n1115 & n2910 ) | ( n2909 & n2910 ) ;
  assign n2912 = ( n975 & n2908 ) | ( n975 & n2911 ) | ( n2908 & n2911 ) ;
  assign n2913 = ( ~n1154 & n2908 ) | ( ~n1154 & n2911 ) | ( n2908 & n2911 ) ;
  assign n2914 = ( x409 & n2912 ) | ( x409 & n2913 ) | ( n2912 & n2913 ) ;
  assign n2915 = ( ~x281 & n2912 ) | ( ~x281 & n2913 ) | ( n2912 & n2913 ) ;
  assign n2916 = ( ~n656 & n2914 ) | ( ~n656 & n2915 ) | ( n2914 & n2915 ) ;
  assign n2917 = x273 & ~n991 ;
  assign n2918 = x273 & n995 ;
  assign n2919 = ( n1104 & n2917 ) | ( n1104 & n2918 ) | ( n2917 & n2918 ) ;
  assign n2920 = ( n1119 & n2917 ) | ( n1119 & n2918 ) | ( n2917 & n2918 ) ;
  assign n2921 = ( ~n1126 & n2917 ) | ( ~n1126 & n2918 ) | ( n2917 & n2918 ) ;
  assign n2922 = ( ~n1115 & n2920 ) | ( ~n1115 & n2921 ) | ( n2920 & n2921 ) ;
  assign n2923 = ( ~n975 & n2919 ) | ( ~n975 & n2922 ) | ( n2919 & n2922 ) ;
  assign n2924 = ( n1154 & n2919 ) | ( n1154 & n2922 ) | ( n2919 & n2922 ) ;
  assign n2925 = ( ~x409 & n2923 ) | ( ~x409 & n2924 ) | ( n2923 & n2924 ) ;
  assign n2926 = ( x281 & n2923 ) | ( x281 & n2924 ) | ( n2923 & n2924 ) ;
  assign n2927 = ( n656 & n2925 ) | ( n656 & n2926 ) | ( n2925 & n2926 ) ;
  assign n2928 = n2916 | n2927 ;
  assign n2929 = ( n2890 & ~n2905 ) | ( n2890 & n2928 ) | ( ~n2905 & n2928 ) ;
  assign n2930 = x145 & n1767 ;
  assign n2931 = x145 & ~n1771 ;
  assign n2932 = ( ~n1751 & n2930 ) | ( ~n1751 & n2931 ) | ( n2930 & n2931 ) ;
  assign n2933 = ( ~n1787 & n2930 ) | ( ~n1787 & n2931 ) | ( n2930 & n2931 ) ;
  assign n2934 = ( n1794 & n2930 ) | ( n1794 & n2931 ) | ( n2930 & n2931 ) ;
  assign n2935 = ( n1783 & n2933 ) | ( n1783 & n2934 ) | ( n2933 & n2934 ) ;
  assign n2936 = ( n1643 & n2932 ) | ( n1643 & n2935 ) | ( n2932 & n2935 ) ;
  assign n2937 = ( ~n1822 & n2932 ) | ( ~n1822 & n2935 ) | ( n2932 & n2935 ) ;
  assign n2938 = ( ~n1324 & n2936 ) | ( ~n1324 & n2937 ) | ( n2936 & n2937 ) ;
  assign n2939 = x17 & ~n1767 ;
  assign n2940 = x17 & n1771 ;
  assign n2941 = ( n1751 & n2939 ) | ( n1751 & n2940 ) | ( n2939 & n2940 ) ;
  assign n2942 = ( n1787 & n2939 ) | ( n1787 & n2940 ) | ( n2939 & n2940 ) ;
  assign n2943 = ( ~n1794 & n2939 ) | ( ~n1794 & n2940 ) | ( n2939 & n2940 ) ;
  assign n2944 = ( ~n1783 & n2942 ) | ( ~n1783 & n2943 ) | ( n2942 & n2943 ) ;
  assign n2945 = ( ~n1643 & n2941 ) | ( ~n1643 & n2944 ) | ( n2941 & n2944 ) ;
  assign n2946 = ( n1822 & n2941 ) | ( n1822 & n2944 ) | ( n2941 & n2944 ) ;
  assign n2947 = ( n1324 & n2945 ) | ( n1324 & n2946 ) | ( n2945 & n2946 ) ;
  assign n2948 = n2938 | n2947 ;
  assign n2949 = ( ~n2890 & n2905 ) | ( ~n2890 & n2948 ) | ( n2905 & n2948 ) ;
  assign n2950 = ( n2573 & ~n2929 ) | ( n2573 & n2949 ) | ( ~n2929 & n2949 ) ;
  assign n2951 = n2883 & ~n2892 ;
  assign n2952 = n2791 & n2883 ;
  assign n2953 = ~n2814 & n2952 ;
  assign n2954 = ( n2862 & n2883 ) | ( n2862 & n2953 ) | ( n2883 & n2953 ) ;
  assign n2955 = ( n2904 & n2951 ) | ( n2904 & n2954 ) | ( n2951 & n2954 ) ;
  assign n2956 = ( n2863 & n2883 ) | ( n2863 & n2953 ) | ( n2883 & n2953 ) ;
  assign n2957 = ( ~n2815 & n2883 ) | ( ~n2815 & n2953 ) | ( n2883 & n2953 ) ;
  assign n2958 = n2883 & n2953 ;
  assign n2959 = ( ~n2887 & n2957 ) | ( ~n2887 & n2958 ) | ( n2957 & n2958 ) ;
  assign n2960 = ( ~n2749 & n2956 ) | ( ~n2749 & n2959 ) | ( n2956 & n2959 ) ;
  assign n2961 = ( ~n2928 & n2955 ) | ( ~n2928 & n2960 ) | ( n2955 & n2960 ) ;
  assign n2962 = ( n2948 & n2955 ) | ( n2948 & n2960 ) | ( n2955 & n2960 ) ;
  assign n2963 = ( n2573 & n2961 ) | ( n2573 & n2962 ) | ( n2961 & n2962 ) ;
  assign n2964 = n2950 | n2963 ;
  assign n2965 = x153 & n1767 ;
  assign n2966 = x153 & ~n1771 ;
  assign n2967 = ( ~n1751 & n2965 ) | ( ~n1751 & n2966 ) | ( n2965 & n2966 ) ;
  assign n2968 = ( ~n1787 & n2965 ) | ( ~n1787 & n2966 ) | ( n2965 & n2966 ) ;
  assign n2969 = ( n1794 & n2965 ) | ( n1794 & n2966 ) | ( n2965 & n2966 ) ;
  assign n2970 = ( n1783 & n2968 ) | ( n1783 & n2969 ) | ( n2968 & n2969 ) ;
  assign n2971 = ( n1643 & n2967 ) | ( n1643 & n2970 ) | ( n2967 & n2970 ) ;
  assign n2972 = ( ~n1822 & n2967 ) | ( ~n1822 & n2970 ) | ( n2967 & n2970 ) ;
  assign n2973 = ( ~n1324 & n2971 ) | ( ~n1324 & n2972 ) | ( n2971 & n2972 ) ;
  assign n2974 = x25 & ~n1767 ;
  assign n2975 = x25 & n1771 ;
  assign n2976 = ( n1751 & n2974 ) | ( n1751 & n2975 ) | ( n2974 & n2975 ) ;
  assign n2977 = ( n1787 & n2974 ) | ( n1787 & n2975 ) | ( n2974 & n2975 ) ;
  assign n2978 = ( ~n1794 & n2974 ) | ( ~n1794 & n2975 ) | ( n2974 & n2975 ) ;
  assign n2979 = ( ~n1783 & n2977 ) | ( ~n1783 & n2978 ) | ( n2977 & n2978 ) ;
  assign n2980 = ( ~n1643 & n2976 ) | ( ~n1643 & n2979 ) | ( n2976 & n2979 ) ;
  assign n2981 = ( n1822 & n2976 ) | ( n1822 & n2979 ) | ( n2976 & n2979 ) ;
  assign n2982 = ( n1324 & n2980 ) | ( n1324 & n2981 ) | ( n2980 & n2981 ) ;
  assign n2983 = n2973 | n2982 ;
  assign n2984 = x409 & n991 ;
  assign n2985 = x409 & ~n995 ;
  assign n2986 = ( ~n1104 & n2984 ) | ( ~n1104 & n2985 ) | ( n2984 & n2985 ) ;
  assign n2987 = ( ~n1119 & n2984 ) | ( ~n1119 & n2985 ) | ( n2984 & n2985 ) ;
  assign n2988 = ( n1126 & n2984 ) | ( n1126 & n2985 ) | ( n2984 & n2985 ) ;
  assign n2989 = ( n1115 & n2987 ) | ( n1115 & n2988 ) | ( n2987 & n2988 ) ;
  assign n2990 = ( n975 & n2986 ) | ( n975 & n2989 ) | ( n2986 & n2989 ) ;
  assign n2991 = ( ~n1154 & n2986 ) | ( ~n1154 & n2989 ) | ( n2986 & n2989 ) ;
  assign n2992 = ( x409 & n2990 ) | ( x409 & n2991 ) | ( n2990 & n2991 ) ;
  assign n2993 = ( ~x281 & n2990 ) | ( ~x281 & n2991 ) | ( n2990 & n2991 ) ;
  assign n2994 = ( ~n656 & n2992 ) | ( ~n656 & n2993 ) | ( n2992 & n2993 ) ;
  assign n2995 = x281 & ~n991 ;
  assign n2996 = x281 & n995 ;
  assign n2997 = ( n1104 & n2995 ) | ( n1104 & n2996 ) | ( n2995 & n2996 ) ;
  assign n2998 = ( n1119 & n2995 ) | ( n1119 & n2996 ) | ( n2995 & n2996 ) ;
  assign n2999 = ( ~n1126 & n2995 ) | ( ~n1126 & n2996 ) | ( n2995 & n2996 ) ;
  assign n3000 = ( ~n1115 & n2998 ) | ( ~n1115 & n2999 ) | ( n2998 & n2999 ) ;
  assign n3001 = ( ~n975 & n2997 ) | ( ~n975 & n3000 ) | ( n2997 & n3000 ) ;
  assign n3002 = ( n1154 & n2997 ) | ( n1154 & n3000 ) | ( n2997 & n3000 ) ;
  assign n3003 = ( ~x409 & n3001 ) | ( ~x409 & n3002 ) | ( n3001 & n3002 ) ;
  assign n3004 = ( x281 & n3001 ) | ( x281 & n3002 ) | ( n3001 & n3002 ) ;
  assign n3005 = ( n656 & n3003 ) | ( n656 & n3004 ) | ( n3003 & n3004 ) ;
  assign n3006 = n2994 | n3005 ;
  assign n3007 = ( n2964 & n2983 ) | ( n2964 & ~n3006 ) | ( n2983 & ~n3006 ) ;
  assign n3008 = x239 & n1767 ;
  assign n3009 = x239 & ~n1771 ;
  assign n3010 = ( ~n1751 & n3008 ) | ( ~n1751 & n3009 ) | ( n3008 & n3009 ) ;
  assign n3011 = ( ~n1787 & n3008 ) | ( ~n1787 & n3009 ) | ( n3008 & n3009 ) ;
  assign n3012 = ( n1794 & n3008 ) | ( n1794 & n3009 ) | ( n3008 & n3009 ) ;
  assign n3013 = ( n1783 & n3011 ) | ( n1783 & n3012 ) | ( n3011 & n3012 ) ;
  assign n3014 = ( n1643 & n3010 ) | ( n1643 & n3013 ) | ( n3010 & n3013 ) ;
  assign n3015 = ( ~n1822 & n3010 ) | ( ~n1822 & n3013 ) | ( n3010 & n3013 ) ;
  assign n3016 = ( ~n1324 & n3014 ) | ( ~n1324 & n3015 ) | ( n3014 & n3015 ) ;
  assign n3017 = x111 & ~n1767 ;
  assign n3018 = x111 & n1771 ;
  assign n3019 = ( n1751 & n3017 ) | ( n1751 & n3018 ) | ( n3017 & n3018 ) ;
  assign n3020 = ( n1787 & n3017 ) | ( n1787 & n3018 ) | ( n3017 & n3018 ) ;
  assign n3021 = ( ~n1794 & n3017 ) | ( ~n1794 & n3018 ) | ( n3017 & n3018 ) ;
  assign n3022 = ( ~n1783 & n3020 ) | ( ~n1783 & n3021 ) | ( n3020 & n3021 ) ;
  assign n3023 = ( ~n1643 & n3019 ) | ( ~n1643 & n3022 ) | ( n3019 & n3022 ) ;
  assign n3024 = ( n1822 & n3019 ) | ( n1822 & n3022 ) | ( n3019 & n3022 ) ;
  assign n3025 = ( n1324 & n3023 ) | ( n1324 & n3024 ) | ( n3023 & n3024 ) ;
  assign n3026 = n3016 | n3025 ;
  assign n3027 = x495 & n991 ;
  assign n3028 = x495 & ~n995 ;
  assign n3029 = ( ~n1104 & n3027 ) | ( ~n1104 & n3028 ) | ( n3027 & n3028 ) ;
  assign n3030 = ( ~n1119 & n3027 ) | ( ~n1119 & n3028 ) | ( n3027 & n3028 ) ;
  assign n3031 = ( n1126 & n3027 ) | ( n1126 & n3028 ) | ( n3027 & n3028 ) ;
  assign n3032 = ( n1115 & n3030 ) | ( n1115 & n3031 ) | ( n3030 & n3031 ) ;
  assign n3033 = ( n975 & n3029 ) | ( n975 & n3032 ) | ( n3029 & n3032 ) ;
  assign n3034 = ( ~n1154 & n3029 ) | ( ~n1154 & n3032 ) | ( n3029 & n3032 ) ;
  assign n3035 = ( x409 & n3033 ) | ( x409 & n3034 ) | ( n3033 & n3034 ) ;
  assign n3036 = ( ~x281 & n3033 ) | ( ~x281 & n3034 ) | ( n3033 & n3034 ) ;
  assign n3037 = ( ~n656 & n3035 ) | ( ~n656 & n3036 ) | ( n3035 & n3036 ) ;
  assign n3038 = x367 & ~n991 ;
  assign n3039 = x367 & n995 ;
  assign n3040 = ( n1104 & n3038 ) | ( n1104 & n3039 ) | ( n3038 & n3039 ) ;
  assign n3041 = ( n1119 & n3038 ) | ( n1119 & n3039 ) | ( n3038 & n3039 ) ;
  assign n3042 = ( ~n1126 & n3038 ) | ( ~n1126 & n3039 ) | ( n3038 & n3039 ) ;
  assign n3043 = ( ~n1115 & n3041 ) | ( ~n1115 & n3042 ) | ( n3041 & n3042 ) ;
  assign n3044 = ( ~n975 & n3040 ) | ( ~n975 & n3043 ) | ( n3040 & n3043 ) ;
  assign n3045 = ( n1154 & n3040 ) | ( n1154 & n3043 ) | ( n3040 & n3043 ) ;
  assign n3046 = ( ~x409 & n3044 ) | ( ~x409 & n3045 ) | ( n3044 & n3045 ) ;
  assign n3047 = ( x281 & n3044 ) | ( x281 & n3045 ) | ( n3044 & n3045 ) ;
  assign n3048 = ( n656 & n3046 ) | ( n656 & n3047 ) | ( n3046 & n3047 ) ;
  assign n3049 = n3037 | n3048 ;
  assign n3050 = ~n3026 & n3049 ;
  assign n3051 = x494 & n991 ;
  assign n3052 = x494 & ~n995 ;
  assign n3053 = ( ~n1104 & n3051 ) | ( ~n1104 & n3052 ) | ( n3051 & n3052 ) ;
  assign n3054 = ( ~n1119 & n3051 ) | ( ~n1119 & n3052 ) | ( n3051 & n3052 ) ;
  assign n3055 = ( n1126 & n3051 ) | ( n1126 & n3052 ) | ( n3051 & n3052 ) ;
  assign n3056 = ( n1115 & n3054 ) | ( n1115 & n3055 ) | ( n3054 & n3055 ) ;
  assign n3057 = ( n975 & n3053 ) | ( n975 & n3056 ) | ( n3053 & n3056 ) ;
  assign n3058 = ( ~n1154 & n3053 ) | ( ~n1154 & n3056 ) | ( n3053 & n3056 ) ;
  assign n3059 = ( x409 & n3057 ) | ( x409 & n3058 ) | ( n3057 & n3058 ) ;
  assign n3060 = ( ~x281 & n3057 ) | ( ~x281 & n3058 ) | ( n3057 & n3058 ) ;
  assign n3061 = ( ~n656 & n3059 ) | ( ~n656 & n3060 ) | ( n3059 & n3060 ) ;
  assign n3062 = x366 & ~n991 ;
  assign n3063 = x366 & n995 ;
  assign n3064 = ( n1104 & n3062 ) | ( n1104 & n3063 ) | ( n3062 & n3063 ) ;
  assign n3065 = ( n1119 & n3062 ) | ( n1119 & n3063 ) | ( n3062 & n3063 ) ;
  assign n3066 = ( ~n1126 & n3062 ) | ( ~n1126 & n3063 ) | ( n3062 & n3063 ) ;
  assign n3067 = ( ~n1115 & n3065 ) | ( ~n1115 & n3066 ) | ( n3065 & n3066 ) ;
  assign n3068 = ( ~n975 & n3064 ) | ( ~n975 & n3067 ) | ( n3064 & n3067 ) ;
  assign n3069 = ( n1154 & n3064 ) | ( n1154 & n3067 ) | ( n3064 & n3067 ) ;
  assign n3070 = ( ~x409 & n3068 ) | ( ~x409 & n3069 ) | ( n3068 & n3069 ) ;
  assign n3071 = ( x281 & n3068 ) | ( x281 & n3069 ) | ( n3068 & n3069 ) ;
  assign n3072 = ( n656 & n3070 ) | ( n656 & n3071 ) | ( n3070 & n3071 ) ;
  assign n3073 = n3061 | n3072 ;
  assign n3074 = x238 & n1767 ;
  assign n3075 = x238 & ~n1771 ;
  assign n3076 = ( ~n1751 & n3074 ) | ( ~n1751 & n3075 ) | ( n3074 & n3075 ) ;
  assign n3077 = ( ~n1787 & n3074 ) | ( ~n1787 & n3075 ) | ( n3074 & n3075 ) ;
  assign n3078 = ( n1794 & n3074 ) | ( n1794 & n3075 ) | ( n3074 & n3075 ) ;
  assign n3079 = ( n1783 & n3077 ) | ( n1783 & n3078 ) | ( n3077 & n3078 ) ;
  assign n3080 = ( n1643 & n3076 ) | ( n1643 & n3079 ) | ( n3076 & n3079 ) ;
  assign n3081 = ( ~n1822 & n3076 ) | ( ~n1822 & n3079 ) | ( n3076 & n3079 ) ;
  assign n3082 = ( ~n1324 & n3080 ) | ( ~n1324 & n3081 ) | ( n3080 & n3081 ) ;
  assign n3083 = x110 & ~n1767 ;
  assign n3084 = x110 & n1771 ;
  assign n3085 = ( n1751 & n3083 ) | ( n1751 & n3084 ) | ( n3083 & n3084 ) ;
  assign n3086 = ( n1787 & n3083 ) | ( n1787 & n3084 ) | ( n3083 & n3084 ) ;
  assign n3087 = ( ~n1794 & n3083 ) | ( ~n1794 & n3084 ) | ( n3083 & n3084 ) ;
  assign n3088 = ( ~n1783 & n3086 ) | ( ~n1783 & n3087 ) | ( n3086 & n3087 ) ;
  assign n3089 = ( ~n1643 & n3085 ) | ( ~n1643 & n3088 ) | ( n3085 & n3088 ) ;
  assign n3090 = ( n1822 & n3085 ) | ( n1822 & n3088 ) | ( n3085 & n3088 ) ;
  assign n3091 = ( n1324 & n3089 ) | ( n1324 & n3090 ) | ( n3089 & n3090 ) ;
  assign n3092 = n3082 | n3091 ;
  assign n3093 = ~n3073 & n3092 ;
  assign n3094 = ~n3050 & n3093 ;
  assign n3095 = n3073 & ~n3092 ;
  assign n3096 = n3050 | n3095 ;
  assign n3097 = x237 & n1767 ;
  assign n3098 = x237 & ~n1771 ;
  assign n3099 = ( ~n1751 & n3097 ) | ( ~n1751 & n3098 ) | ( n3097 & n3098 ) ;
  assign n3100 = ( ~n1787 & n3097 ) | ( ~n1787 & n3098 ) | ( n3097 & n3098 ) ;
  assign n3101 = ( n1794 & n3097 ) | ( n1794 & n3098 ) | ( n3097 & n3098 ) ;
  assign n3102 = ( n1783 & n3100 ) | ( n1783 & n3101 ) | ( n3100 & n3101 ) ;
  assign n3103 = ( n1643 & n3099 ) | ( n1643 & n3102 ) | ( n3099 & n3102 ) ;
  assign n3104 = ( ~n1822 & n3099 ) | ( ~n1822 & n3102 ) | ( n3099 & n3102 ) ;
  assign n3105 = ( ~n1324 & n3103 ) | ( ~n1324 & n3104 ) | ( n3103 & n3104 ) ;
  assign n3106 = x109 & ~n1767 ;
  assign n3107 = x109 & n1771 ;
  assign n3108 = ( n1751 & n3106 ) | ( n1751 & n3107 ) | ( n3106 & n3107 ) ;
  assign n3109 = ( n1787 & n3106 ) | ( n1787 & n3107 ) | ( n3106 & n3107 ) ;
  assign n3110 = ( ~n1794 & n3106 ) | ( ~n1794 & n3107 ) | ( n3106 & n3107 ) ;
  assign n3111 = ( ~n1783 & n3109 ) | ( ~n1783 & n3110 ) | ( n3109 & n3110 ) ;
  assign n3112 = ( ~n1643 & n3108 ) | ( ~n1643 & n3111 ) | ( n3108 & n3111 ) ;
  assign n3113 = ( n1822 & n3108 ) | ( n1822 & n3111 ) | ( n3108 & n3111 ) ;
  assign n3114 = ( n1324 & n3112 ) | ( n1324 & n3113 ) | ( n3112 & n3113 ) ;
  assign n3115 = n3105 | n3114 ;
  assign n3116 = x493 & n991 ;
  assign n3117 = x493 & ~n995 ;
  assign n3118 = ( ~n1104 & n3116 ) | ( ~n1104 & n3117 ) | ( n3116 & n3117 ) ;
  assign n3119 = ( ~n1119 & n3116 ) | ( ~n1119 & n3117 ) | ( n3116 & n3117 ) ;
  assign n3120 = ( n1126 & n3116 ) | ( n1126 & n3117 ) | ( n3116 & n3117 ) ;
  assign n3121 = ( n1115 & n3119 ) | ( n1115 & n3120 ) | ( n3119 & n3120 ) ;
  assign n3122 = ( n975 & n3118 ) | ( n975 & n3121 ) | ( n3118 & n3121 ) ;
  assign n3123 = ( ~n1154 & n3118 ) | ( ~n1154 & n3121 ) | ( n3118 & n3121 ) ;
  assign n3124 = ( x409 & n3122 ) | ( x409 & n3123 ) | ( n3122 & n3123 ) ;
  assign n3125 = ( ~x281 & n3122 ) | ( ~x281 & n3123 ) | ( n3122 & n3123 ) ;
  assign n3126 = ( ~n656 & n3124 ) | ( ~n656 & n3125 ) | ( n3124 & n3125 ) ;
  assign n3127 = x365 & ~n991 ;
  assign n3128 = x365 & n995 ;
  assign n3129 = ( n1104 & n3127 ) | ( n1104 & n3128 ) | ( n3127 & n3128 ) ;
  assign n3130 = ( n1119 & n3127 ) | ( n1119 & n3128 ) | ( n3127 & n3128 ) ;
  assign n3131 = ( ~n1126 & n3127 ) | ( ~n1126 & n3128 ) | ( n3127 & n3128 ) ;
  assign n3132 = ( ~n1115 & n3130 ) | ( ~n1115 & n3131 ) | ( n3130 & n3131 ) ;
  assign n3133 = ( ~n975 & n3129 ) | ( ~n975 & n3132 ) | ( n3129 & n3132 ) ;
  assign n3134 = ( n1154 & n3129 ) | ( n1154 & n3132 ) | ( n3129 & n3132 ) ;
  assign n3135 = ( ~x409 & n3133 ) | ( ~x409 & n3134 ) | ( n3133 & n3134 ) ;
  assign n3136 = ( x281 & n3133 ) | ( x281 & n3134 ) | ( n3133 & n3134 ) ;
  assign n3137 = ( n656 & n3135 ) | ( n656 & n3136 ) | ( n3135 & n3136 ) ;
  assign n3138 = n3126 | n3137 ;
  assign n3139 = ~n3115 & n3138 ;
  assign n3140 = x236 & n1767 ;
  assign n3141 = x236 & ~n1771 ;
  assign n3142 = ( ~n1751 & n3140 ) | ( ~n1751 & n3141 ) | ( n3140 & n3141 ) ;
  assign n3143 = ( ~n1787 & n3140 ) | ( ~n1787 & n3141 ) | ( n3140 & n3141 ) ;
  assign n3144 = ( n1794 & n3140 ) | ( n1794 & n3141 ) | ( n3140 & n3141 ) ;
  assign n3145 = ( n1783 & n3143 ) | ( n1783 & n3144 ) | ( n3143 & n3144 ) ;
  assign n3146 = ( n1643 & n3142 ) | ( n1643 & n3145 ) | ( n3142 & n3145 ) ;
  assign n3147 = ( ~n1822 & n3142 ) | ( ~n1822 & n3145 ) | ( n3142 & n3145 ) ;
  assign n3148 = ( ~n1324 & n3146 ) | ( ~n1324 & n3147 ) | ( n3146 & n3147 ) ;
  assign n3149 = x108 & ~n1767 ;
  assign n3150 = x108 & n1771 ;
  assign n3151 = ( n1751 & n3149 ) | ( n1751 & n3150 ) | ( n3149 & n3150 ) ;
  assign n3152 = ( n1787 & n3149 ) | ( n1787 & n3150 ) | ( n3149 & n3150 ) ;
  assign n3153 = ( ~n1794 & n3149 ) | ( ~n1794 & n3150 ) | ( n3149 & n3150 ) ;
  assign n3154 = ( ~n1783 & n3152 ) | ( ~n1783 & n3153 ) | ( n3152 & n3153 ) ;
  assign n3155 = ( ~n1643 & n3151 ) | ( ~n1643 & n3154 ) | ( n3151 & n3154 ) ;
  assign n3156 = ( n1822 & n3151 ) | ( n1822 & n3154 ) | ( n3151 & n3154 ) ;
  assign n3157 = ( n1324 & n3155 ) | ( n1324 & n3156 ) | ( n3155 & n3156 ) ;
  assign n3158 = n3148 | n3157 ;
  assign n3159 = x492 & n991 ;
  assign n3160 = x492 & ~n995 ;
  assign n3161 = ( ~n1104 & n3159 ) | ( ~n1104 & n3160 ) | ( n3159 & n3160 ) ;
  assign n3162 = ( ~n1119 & n3159 ) | ( ~n1119 & n3160 ) | ( n3159 & n3160 ) ;
  assign n3163 = ( n1126 & n3159 ) | ( n1126 & n3160 ) | ( n3159 & n3160 ) ;
  assign n3164 = ( n1115 & n3162 ) | ( n1115 & n3163 ) | ( n3162 & n3163 ) ;
  assign n3165 = ( n975 & n3161 ) | ( n975 & n3164 ) | ( n3161 & n3164 ) ;
  assign n3166 = ( ~n1154 & n3161 ) | ( ~n1154 & n3164 ) | ( n3161 & n3164 ) ;
  assign n3167 = ( x409 & n3165 ) | ( x409 & n3166 ) | ( n3165 & n3166 ) ;
  assign n3168 = ( ~x281 & n3165 ) | ( ~x281 & n3166 ) | ( n3165 & n3166 ) ;
  assign n3169 = ( ~n656 & n3167 ) | ( ~n656 & n3168 ) | ( n3167 & n3168 ) ;
  assign n3170 = x364 & ~n991 ;
  assign n3171 = x364 & n995 ;
  assign n3172 = ( n1104 & n3170 ) | ( n1104 & n3171 ) | ( n3170 & n3171 ) ;
  assign n3173 = ( n1119 & n3170 ) | ( n1119 & n3171 ) | ( n3170 & n3171 ) ;
  assign n3174 = ( ~n1126 & n3170 ) | ( ~n1126 & n3171 ) | ( n3170 & n3171 ) ;
  assign n3175 = ( ~n1115 & n3173 ) | ( ~n1115 & n3174 ) | ( n3173 & n3174 ) ;
  assign n3176 = ( ~n975 & n3172 ) | ( ~n975 & n3175 ) | ( n3172 & n3175 ) ;
  assign n3177 = ( n1154 & n3172 ) | ( n1154 & n3175 ) | ( n3172 & n3175 ) ;
  assign n3178 = ( ~x409 & n3176 ) | ( ~x409 & n3177 ) | ( n3176 & n3177 ) ;
  assign n3179 = ( x281 & n3176 ) | ( x281 & n3177 ) | ( n3176 & n3177 ) ;
  assign n3180 = ( n656 & n3178 ) | ( n656 & n3179 ) | ( n3178 & n3179 ) ;
  assign n3181 = n3169 | n3180 ;
  assign n3182 = ~n3158 & n3181 ;
  assign n3183 = n3139 | n3182 ;
  assign n3184 = n3096 | n3183 ;
  assign n3185 = ~n3094 & n3184 ;
  assign n3186 = x235 & n1767 ;
  assign n3187 = x235 & ~n1771 ;
  assign n3188 = ( ~n1751 & n3186 ) | ( ~n1751 & n3187 ) | ( n3186 & n3187 ) ;
  assign n3189 = ( ~n1787 & n3186 ) | ( ~n1787 & n3187 ) | ( n3186 & n3187 ) ;
  assign n3190 = ( n1794 & n3186 ) | ( n1794 & n3187 ) | ( n3186 & n3187 ) ;
  assign n3191 = ( n1783 & n3189 ) | ( n1783 & n3190 ) | ( n3189 & n3190 ) ;
  assign n3192 = ( n1643 & n3188 ) | ( n1643 & n3191 ) | ( n3188 & n3191 ) ;
  assign n3193 = ( ~n1822 & n3188 ) | ( ~n1822 & n3191 ) | ( n3188 & n3191 ) ;
  assign n3194 = ( ~n1324 & n3192 ) | ( ~n1324 & n3193 ) | ( n3192 & n3193 ) ;
  assign n3195 = x107 & ~n1767 ;
  assign n3196 = x107 & n1771 ;
  assign n3197 = ( n1751 & n3195 ) | ( n1751 & n3196 ) | ( n3195 & n3196 ) ;
  assign n3198 = ( n1787 & n3195 ) | ( n1787 & n3196 ) | ( n3195 & n3196 ) ;
  assign n3199 = ( ~n1794 & n3195 ) | ( ~n1794 & n3196 ) | ( n3195 & n3196 ) ;
  assign n3200 = ( ~n1783 & n3198 ) | ( ~n1783 & n3199 ) | ( n3198 & n3199 ) ;
  assign n3201 = ( ~n1643 & n3197 ) | ( ~n1643 & n3200 ) | ( n3197 & n3200 ) ;
  assign n3202 = ( n1822 & n3197 ) | ( n1822 & n3200 ) | ( n3197 & n3200 ) ;
  assign n3203 = ( n1324 & n3201 ) | ( n1324 & n3202 ) | ( n3201 & n3202 ) ;
  assign n3204 = n3194 | n3203 ;
  assign n3205 = x491 & n991 ;
  assign n3206 = x491 & ~n995 ;
  assign n3207 = ( ~n1104 & n3205 ) | ( ~n1104 & n3206 ) | ( n3205 & n3206 ) ;
  assign n3208 = ( ~n1119 & n3205 ) | ( ~n1119 & n3206 ) | ( n3205 & n3206 ) ;
  assign n3209 = ( n1126 & n3205 ) | ( n1126 & n3206 ) | ( n3205 & n3206 ) ;
  assign n3210 = ( n1115 & n3208 ) | ( n1115 & n3209 ) | ( n3208 & n3209 ) ;
  assign n3211 = ( n975 & n3207 ) | ( n975 & n3210 ) | ( n3207 & n3210 ) ;
  assign n3212 = ( ~n1154 & n3207 ) | ( ~n1154 & n3210 ) | ( n3207 & n3210 ) ;
  assign n3213 = ( x409 & n3211 ) | ( x409 & n3212 ) | ( n3211 & n3212 ) ;
  assign n3214 = ( ~x281 & n3211 ) | ( ~x281 & n3212 ) | ( n3211 & n3212 ) ;
  assign n3215 = ( ~n656 & n3213 ) | ( ~n656 & n3214 ) | ( n3213 & n3214 ) ;
  assign n3216 = x363 & ~n991 ;
  assign n3217 = x363 & n995 ;
  assign n3218 = ( n1104 & n3216 ) | ( n1104 & n3217 ) | ( n3216 & n3217 ) ;
  assign n3219 = ( n1119 & n3216 ) | ( n1119 & n3217 ) | ( n3216 & n3217 ) ;
  assign n3220 = ( ~n1126 & n3216 ) | ( ~n1126 & n3217 ) | ( n3216 & n3217 ) ;
  assign n3221 = ( ~n1115 & n3219 ) | ( ~n1115 & n3220 ) | ( n3219 & n3220 ) ;
  assign n3222 = ( ~n975 & n3218 ) | ( ~n975 & n3221 ) | ( n3218 & n3221 ) ;
  assign n3223 = ( n1154 & n3218 ) | ( n1154 & n3221 ) | ( n3218 & n3221 ) ;
  assign n3224 = ( ~x409 & n3222 ) | ( ~x409 & n3223 ) | ( n3222 & n3223 ) ;
  assign n3225 = ( x281 & n3222 ) | ( x281 & n3223 ) | ( n3222 & n3223 ) ;
  assign n3226 = ( n656 & n3224 ) | ( n656 & n3225 ) | ( n3224 & n3225 ) ;
  assign n3227 = n3215 | n3226 ;
  assign n3228 = x490 & n991 ;
  assign n3229 = x490 & ~n995 ;
  assign n3230 = ( ~n1104 & n3228 ) | ( ~n1104 & n3229 ) | ( n3228 & n3229 ) ;
  assign n3231 = ( ~n1119 & n3228 ) | ( ~n1119 & n3229 ) | ( n3228 & n3229 ) ;
  assign n3232 = ( n1126 & n3228 ) | ( n1126 & n3229 ) | ( n3228 & n3229 ) ;
  assign n3233 = ( n1115 & n3231 ) | ( n1115 & n3232 ) | ( n3231 & n3232 ) ;
  assign n3234 = ( n975 & n3230 ) | ( n975 & n3233 ) | ( n3230 & n3233 ) ;
  assign n3235 = ( ~n1154 & n3230 ) | ( ~n1154 & n3233 ) | ( n3230 & n3233 ) ;
  assign n3236 = ( x409 & n3234 ) | ( x409 & n3235 ) | ( n3234 & n3235 ) ;
  assign n3237 = ( ~x281 & n3234 ) | ( ~x281 & n3235 ) | ( n3234 & n3235 ) ;
  assign n3238 = ( ~n656 & n3236 ) | ( ~n656 & n3237 ) | ( n3236 & n3237 ) ;
  assign n3239 = x362 & ~n991 ;
  assign n3240 = x362 & n995 ;
  assign n3241 = ( n1104 & n3239 ) | ( n1104 & n3240 ) | ( n3239 & n3240 ) ;
  assign n3242 = ( n1119 & n3239 ) | ( n1119 & n3240 ) | ( n3239 & n3240 ) ;
  assign n3243 = ( ~n1126 & n3239 ) | ( ~n1126 & n3240 ) | ( n3239 & n3240 ) ;
  assign n3244 = ( ~n1115 & n3242 ) | ( ~n1115 & n3243 ) | ( n3242 & n3243 ) ;
  assign n3245 = ( ~n975 & n3241 ) | ( ~n975 & n3244 ) | ( n3241 & n3244 ) ;
  assign n3246 = ( n1154 & n3241 ) | ( n1154 & n3244 ) | ( n3241 & n3244 ) ;
  assign n3247 = ( ~x409 & n3245 ) | ( ~x409 & n3246 ) | ( n3245 & n3246 ) ;
  assign n3248 = ( x281 & n3245 ) | ( x281 & n3246 ) | ( n3245 & n3246 ) ;
  assign n3249 = ( n656 & n3247 ) | ( n656 & n3248 ) | ( n3247 & n3248 ) ;
  assign n3250 = n3238 | n3249 ;
  assign n3251 = x234 & n1767 ;
  assign n3252 = x234 & ~n1771 ;
  assign n3253 = ( ~n1751 & n3251 ) | ( ~n1751 & n3252 ) | ( n3251 & n3252 ) ;
  assign n3254 = ( ~n1787 & n3251 ) | ( ~n1787 & n3252 ) | ( n3251 & n3252 ) ;
  assign n3255 = ( n1794 & n3251 ) | ( n1794 & n3252 ) | ( n3251 & n3252 ) ;
  assign n3256 = ( n1783 & n3254 ) | ( n1783 & n3255 ) | ( n3254 & n3255 ) ;
  assign n3257 = ( n1643 & n3253 ) | ( n1643 & n3256 ) | ( n3253 & n3256 ) ;
  assign n3258 = ( ~n1822 & n3253 ) | ( ~n1822 & n3256 ) | ( n3253 & n3256 ) ;
  assign n3259 = ( ~n1324 & n3257 ) | ( ~n1324 & n3258 ) | ( n3257 & n3258 ) ;
  assign n3260 = x106 & ~n1767 ;
  assign n3261 = x106 & n1771 ;
  assign n3262 = ( n1751 & n3260 ) | ( n1751 & n3261 ) | ( n3260 & n3261 ) ;
  assign n3263 = ( n1787 & n3260 ) | ( n1787 & n3261 ) | ( n3260 & n3261 ) ;
  assign n3264 = ( ~n1794 & n3260 ) | ( ~n1794 & n3261 ) | ( n3260 & n3261 ) ;
  assign n3265 = ( ~n1783 & n3263 ) | ( ~n1783 & n3264 ) | ( n3263 & n3264 ) ;
  assign n3266 = ( ~n1643 & n3262 ) | ( ~n1643 & n3265 ) | ( n3262 & n3265 ) ;
  assign n3267 = ( n1822 & n3262 ) | ( n1822 & n3265 ) | ( n3262 & n3265 ) ;
  assign n3268 = ( n1324 & n3266 ) | ( n1324 & n3267 ) | ( n3266 & n3267 ) ;
  assign n3269 = n3259 | n3268 ;
  assign n3270 = n3250 & ~n3269 ;
  assign n3271 = x233 & n1767 ;
  assign n3272 = x233 & ~n1771 ;
  assign n3273 = ( ~n1751 & n3271 ) | ( ~n1751 & n3272 ) | ( n3271 & n3272 ) ;
  assign n3274 = ( ~n1787 & n3271 ) | ( ~n1787 & n3272 ) | ( n3271 & n3272 ) ;
  assign n3275 = ( n1794 & n3271 ) | ( n1794 & n3272 ) | ( n3271 & n3272 ) ;
  assign n3276 = ( n1783 & n3274 ) | ( n1783 & n3275 ) | ( n3274 & n3275 ) ;
  assign n3277 = ( n1643 & n3273 ) | ( n1643 & n3276 ) | ( n3273 & n3276 ) ;
  assign n3278 = ( ~n1822 & n3273 ) | ( ~n1822 & n3276 ) | ( n3273 & n3276 ) ;
  assign n3279 = ( ~n1324 & n3277 ) | ( ~n1324 & n3278 ) | ( n3277 & n3278 ) ;
  assign n3280 = x105 & ~n1767 ;
  assign n3281 = x105 & n1771 ;
  assign n3282 = ( n1751 & n3280 ) | ( n1751 & n3281 ) | ( n3280 & n3281 ) ;
  assign n3283 = ( n1787 & n3280 ) | ( n1787 & n3281 ) | ( n3280 & n3281 ) ;
  assign n3284 = ( ~n1794 & n3280 ) | ( ~n1794 & n3281 ) | ( n3280 & n3281 ) ;
  assign n3285 = ( ~n1783 & n3283 ) | ( ~n1783 & n3284 ) | ( n3283 & n3284 ) ;
  assign n3286 = ( ~n1643 & n3282 ) | ( ~n1643 & n3285 ) | ( n3282 & n3285 ) ;
  assign n3287 = ( n1822 & n3282 ) | ( n1822 & n3285 ) | ( n3282 & n3285 ) ;
  assign n3288 = ( n1324 & n3286 ) | ( n1324 & n3287 ) | ( n3286 & n3287 ) ;
  assign n3289 = n3279 | n3288 ;
  assign n3290 = x489 & n991 ;
  assign n3291 = x489 & ~n995 ;
  assign n3292 = ( ~n1104 & n3290 ) | ( ~n1104 & n3291 ) | ( n3290 & n3291 ) ;
  assign n3293 = ( ~n1119 & n3290 ) | ( ~n1119 & n3291 ) | ( n3290 & n3291 ) ;
  assign n3294 = ( n1126 & n3290 ) | ( n1126 & n3291 ) | ( n3290 & n3291 ) ;
  assign n3295 = ( n1115 & n3293 ) | ( n1115 & n3294 ) | ( n3293 & n3294 ) ;
  assign n3296 = ( n975 & n3292 ) | ( n975 & n3295 ) | ( n3292 & n3295 ) ;
  assign n3297 = ( ~n1154 & n3292 ) | ( ~n1154 & n3295 ) | ( n3292 & n3295 ) ;
  assign n3298 = ( x409 & n3296 ) | ( x409 & n3297 ) | ( n3296 & n3297 ) ;
  assign n3299 = ( ~x281 & n3296 ) | ( ~x281 & n3297 ) | ( n3296 & n3297 ) ;
  assign n3300 = ( ~n656 & n3298 ) | ( ~n656 & n3299 ) | ( n3298 & n3299 ) ;
  assign n3301 = x361 & ~n991 ;
  assign n3302 = x361 & n995 ;
  assign n3303 = ( n1104 & n3301 ) | ( n1104 & n3302 ) | ( n3301 & n3302 ) ;
  assign n3304 = ( n1119 & n3301 ) | ( n1119 & n3302 ) | ( n3301 & n3302 ) ;
  assign n3305 = ( ~n1126 & n3301 ) | ( ~n1126 & n3302 ) | ( n3301 & n3302 ) ;
  assign n3306 = ( ~n1115 & n3304 ) | ( ~n1115 & n3305 ) | ( n3304 & n3305 ) ;
  assign n3307 = ( ~n975 & n3303 ) | ( ~n975 & n3306 ) | ( n3303 & n3306 ) ;
  assign n3308 = ( n1154 & n3303 ) | ( n1154 & n3306 ) | ( n3303 & n3306 ) ;
  assign n3309 = ( ~x409 & n3307 ) | ( ~x409 & n3308 ) | ( n3307 & n3308 ) ;
  assign n3310 = ( x281 & n3307 ) | ( x281 & n3308 ) | ( n3307 & n3308 ) ;
  assign n3311 = ( n656 & n3309 ) | ( n656 & n3310 ) | ( n3309 & n3310 ) ;
  assign n3312 = n3300 | n3311 ;
  assign n3313 = x488 & n991 ;
  assign n3314 = x488 & ~n995 ;
  assign n3315 = ( ~n1104 & n3313 ) | ( ~n1104 & n3314 ) | ( n3313 & n3314 ) ;
  assign n3316 = ( ~n1119 & n3313 ) | ( ~n1119 & n3314 ) | ( n3313 & n3314 ) ;
  assign n3317 = ( n1126 & n3313 ) | ( n1126 & n3314 ) | ( n3313 & n3314 ) ;
  assign n3318 = ( n1115 & n3316 ) | ( n1115 & n3317 ) | ( n3316 & n3317 ) ;
  assign n3319 = ( n975 & n3315 ) | ( n975 & n3318 ) | ( n3315 & n3318 ) ;
  assign n3320 = ( ~n1154 & n3315 ) | ( ~n1154 & n3318 ) | ( n3315 & n3318 ) ;
  assign n3321 = ( x409 & n3319 ) | ( x409 & n3320 ) | ( n3319 & n3320 ) ;
  assign n3322 = ( ~x281 & n3319 ) | ( ~x281 & n3320 ) | ( n3319 & n3320 ) ;
  assign n3323 = ( ~n656 & n3321 ) | ( ~n656 & n3322 ) | ( n3321 & n3322 ) ;
  assign n3324 = x360 & ~n991 ;
  assign n3325 = x360 & n995 ;
  assign n3326 = ( n1104 & n3324 ) | ( n1104 & n3325 ) | ( n3324 & n3325 ) ;
  assign n3327 = ( n1119 & n3324 ) | ( n1119 & n3325 ) | ( n3324 & n3325 ) ;
  assign n3328 = ( ~n1126 & n3324 ) | ( ~n1126 & n3325 ) | ( n3324 & n3325 ) ;
  assign n3329 = ( ~n1115 & n3327 ) | ( ~n1115 & n3328 ) | ( n3327 & n3328 ) ;
  assign n3330 = ( ~n975 & n3326 ) | ( ~n975 & n3329 ) | ( n3326 & n3329 ) ;
  assign n3331 = ( n1154 & n3326 ) | ( n1154 & n3329 ) | ( n3326 & n3329 ) ;
  assign n3332 = ( ~x409 & n3330 ) | ( ~x409 & n3331 ) | ( n3330 & n3331 ) ;
  assign n3333 = ( x281 & n3330 ) | ( x281 & n3331 ) | ( n3330 & n3331 ) ;
  assign n3334 = ( n656 & n3332 ) | ( n656 & n3333 ) | ( n3332 & n3333 ) ;
  assign n3335 = n3323 | n3334 ;
  assign n3336 = x232 & n1767 ;
  assign n3337 = x232 & ~n1771 ;
  assign n3338 = ( ~n1751 & n3336 ) | ( ~n1751 & n3337 ) | ( n3336 & n3337 ) ;
  assign n3339 = ( ~n1787 & n3336 ) | ( ~n1787 & n3337 ) | ( n3336 & n3337 ) ;
  assign n3340 = ( n1794 & n3336 ) | ( n1794 & n3337 ) | ( n3336 & n3337 ) ;
  assign n3341 = ( n1783 & n3339 ) | ( n1783 & n3340 ) | ( n3339 & n3340 ) ;
  assign n3342 = ( n1643 & n3338 ) | ( n1643 & n3341 ) | ( n3338 & n3341 ) ;
  assign n3343 = ( ~n1822 & n3338 ) | ( ~n1822 & n3341 ) | ( n3338 & n3341 ) ;
  assign n3344 = ( ~n1324 & n3342 ) | ( ~n1324 & n3343 ) | ( n3342 & n3343 ) ;
  assign n3345 = x104 & ~n1767 ;
  assign n3346 = x104 & n1771 ;
  assign n3347 = ( n1751 & n3345 ) | ( n1751 & n3346 ) | ( n3345 & n3346 ) ;
  assign n3348 = ( n1787 & n3345 ) | ( n1787 & n3346 ) | ( n3345 & n3346 ) ;
  assign n3349 = ( ~n1794 & n3345 ) | ( ~n1794 & n3346 ) | ( n3345 & n3346 ) ;
  assign n3350 = ( ~n1783 & n3348 ) | ( ~n1783 & n3349 ) | ( n3348 & n3349 ) ;
  assign n3351 = ( ~n1643 & n3347 ) | ( ~n1643 & n3350 ) | ( n3347 & n3350 ) ;
  assign n3352 = ( n1822 & n3347 ) | ( n1822 & n3350 ) | ( n3347 & n3350 ) ;
  assign n3353 = ( n1324 & n3351 ) | ( n1324 & n3352 ) | ( n3351 & n3352 ) ;
  assign n3354 = n3344 | n3353 ;
  assign n3355 = ~n3335 & n3354 ;
  assign n3356 = ( n3289 & ~n3312 ) | ( n3289 & n3355 ) | ( ~n3312 & n3355 ) ;
  assign n3357 = ~n3250 & n3269 ;
  assign n3358 = ~n3270 & n3357 ;
  assign n3359 = ( ~n3270 & n3356 ) | ( ~n3270 & n3358 ) | ( n3356 & n3358 ) ;
  assign n3360 = ( n3204 & ~n3227 ) | ( n3204 & n3359 ) | ( ~n3227 & n3359 ) ;
  assign n3361 = ( n3094 & ~n3185 ) | ( n3094 & n3360 ) | ( ~n3185 & n3360 ) ;
  assign n3362 = n3026 & ~n3049 ;
  assign n3363 = n3158 & ~n3181 ;
  assign n3364 = ( n3115 & ~n3138 ) | ( n3115 & n3363 ) | ( ~n3138 & n3363 ) ;
  assign n3365 = ~n3096 & n3364 ;
  assign n3366 = n3362 | n3365 ;
  assign n3367 = n3361 | n3366 ;
  assign n3368 = x251 & n1767 ;
  assign n3369 = x251 & ~n1771 ;
  assign n3370 = ( ~n1751 & n3368 ) | ( ~n1751 & n3369 ) | ( n3368 & n3369 ) ;
  assign n3371 = ( ~n1787 & n3368 ) | ( ~n1787 & n3369 ) | ( n3368 & n3369 ) ;
  assign n3372 = ( n1794 & n3368 ) | ( n1794 & n3369 ) | ( n3368 & n3369 ) ;
  assign n3373 = ( n1783 & n3371 ) | ( n1783 & n3372 ) | ( n3371 & n3372 ) ;
  assign n3374 = ( n1643 & n3370 ) | ( n1643 & n3373 ) | ( n3370 & n3373 ) ;
  assign n3375 = ( ~n1822 & n3370 ) | ( ~n1822 & n3373 ) | ( n3370 & n3373 ) ;
  assign n3376 = ( ~n1324 & n3374 ) | ( ~n1324 & n3375 ) | ( n3374 & n3375 ) ;
  assign n3377 = x123 & ~n1767 ;
  assign n3378 = x123 & n1771 ;
  assign n3379 = ( n1751 & n3377 ) | ( n1751 & n3378 ) | ( n3377 & n3378 ) ;
  assign n3380 = ( n1787 & n3377 ) | ( n1787 & n3378 ) | ( n3377 & n3378 ) ;
  assign n3381 = ( ~n1794 & n3377 ) | ( ~n1794 & n3378 ) | ( n3377 & n3378 ) ;
  assign n3382 = ( ~n1783 & n3380 ) | ( ~n1783 & n3381 ) | ( n3380 & n3381 ) ;
  assign n3383 = ( ~n1643 & n3379 ) | ( ~n1643 & n3382 ) | ( n3379 & n3382 ) ;
  assign n3384 = ( n1822 & n3379 ) | ( n1822 & n3382 ) | ( n3379 & n3382 ) ;
  assign n3385 = ( n1324 & n3383 ) | ( n1324 & n3384 ) | ( n3383 & n3384 ) ;
  assign n3386 = n3376 | n3385 ;
  assign n3387 = x507 & n991 ;
  assign n3388 = x507 & ~n995 ;
  assign n3389 = ( ~n1104 & n3387 ) | ( ~n1104 & n3388 ) | ( n3387 & n3388 ) ;
  assign n3390 = ( ~n1119 & n3387 ) | ( ~n1119 & n3388 ) | ( n3387 & n3388 ) ;
  assign n3391 = ( n1126 & n3387 ) | ( n1126 & n3388 ) | ( n3387 & n3388 ) ;
  assign n3392 = ( n1115 & n3390 ) | ( n1115 & n3391 ) | ( n3390 & n3391 ) ;
  assign n3393 = ( n975 & n3389 ) | ( n975 & n3392 ) | ( n3389 & n3392 ) ;
  assign n3394 = ( ~n1154 & n3389 ) | ( ~n1154 & n3392 ) | ( n3389 & n3392 ) ;
  assign n3395 = ( x409 & n3393 ) | ( x409 & n3394 ) | ( n3393 & n3394 ) ;
  assign n3396 = ( ~x281 & n3393 ) | ( ~x281 & n3394 ) | ( n3393 & n3394 ) ;
  assign n3397 = ( ~n656 & n3395 ) | ( ~n656 & n3396 ) | ( n3395 & n3396 ) ;
  assign n3398 = x379 & ~n991 ;
  assign n3399 = x379 & n995 ;
  assign n3400 = ( n1104 & n3398 ) | ( n1104 & n3399 ) | ( n3398 & n3399 ) ;
  assign n3401 = ( n1119 & n3398 ) | ( n1119 & n3399 ) | ( n3398 & n3399 ) ;
  assign n3402 = ( ~n1126 & n3398 ) | ( ~n1126 & n3399 ) | ( n3398 & n3399 ) ;
  assign n3403 = ( ~n1115 & n3401 ) | ( ~n1115 & n3402 ) | ( n3401 & n3402 ) ;
  assign n3404 = ( ~n975 & n3400 ) | ( ~n975 & n3403 ) | ( n3400 & n3403 ) ;
  assign n3405 = ( n1154 & n3400 ) | ( n1154 & n3403 ) | ( n3400 & n3403 ) ;
  assign n3406 = ( ~x409 & n3404 ) | ( ~x409 & n3405 ) | ( n3404 & n3405 ) ;
  assign n3407 = ( x281 & n3404 ) | ( x281 & n3405 ) | ( n3404 & n3405 ) ;
  assign n3408 = ( n656 & n3406 ) | ( n656 & n3407 ) | ( n3406 & n3407 ) ;
  assign n3409 = n3397 | n3408 ;
  assign n3410 = ~n3386 & n3409 ;
  assign n3411 = x506 & n991 ;
  assign n3412 = x506 & ~n995 ;
  assign n3413 = ( ~n1104 & n3411 ) | ( ~n1104 & n3412 ) | ( n3411 & n3412 ) ;
  assign n3414 = ( ~n1119 & n3411 ) | ( ~n1119 & n3412 ) | ( n3411 & n3412 ) ;
  assign n3415 = ( n1126 & n3411 ) | ( n1126 & n3412 ) | ( n3411 & n3412 ) ;
  assign n3416 = ( n1115 & n3414 ) | ( n1115 & n3415 ) | ( n3414 & n3415 ) ;
  assign n3417 = ( n975 & n3413 ) | ( n975 & n3416 ) | ( n3413 & n3416 ) ;
  assign n3418 = ( ~n1154 & n3413 ) | ( ~n1154 & n3416 ) | ( n3413 & n3416 ) ;
  assign n3419 = ( x409 & n3417 ) | ( x409 & n3418 ) | ( n3417 & n3418 ) ;
  assign n3420 = ( ~x281 & n3417 ) | ( ~x281 & n3418 ) | ( n3417 & n3418 ) ;
  assign n3421 = ( ~n656 & n3419 ) | ( ~n656 & n3420 ) | ( n3419 & n3420 ) ;
  assign n3422 = x378 & ~n991 ;
  assign n3423 = x378 & n995 ;
  assign n3424 = ( n1104 & n3422 ) | ( n1104 & n3423 ) | ( n3422 & n3423 ) ;
  assign n3425 = ( n1119 & n3422 ) | ( n1119 & n3423 ) | ( n3422 & n3423 ) ;
  assign n3426 = ( ~n1126 & n3422 ) | ( ~n1126 & n3423 ) | ( n3422 & n3423 ) ;
  assign n3427 = ( ~n1115 & n3425 ) | ( ~n1115 & n3426 ) | ( n3425 & n3426 ) ;
  assign n3428 = ( ~n975 & n3424 ) | ( ~n975 & n3427 ) | ( n3424 & n3427 ) ;
  assign n3429 = ( n1154 & n3424 ) | ( n1154 & n3427 ) | ( n3424 & n3427 ) ;
  assign n3430 = ( ~x409 & n3428 ) | ( ~x409 & n3429 ) | ( n3428 & n3429 ) ;
  assign n3431 = ( x281 & n3428 ) | ( x281 & n3429 ) | ( n3428 & n3429 ) ;
  assign n3432 = ( n656 & n3430 ) | ( n656 & n3431 ) | ( n3430 & n3431 ) ;
  assign n3433 = n3421 | n3432 ;
  assign n3434 = x250 & n1767 ;
  assign n3435 = x250 & ~n1771 ;
  assign n3436 = ( ~n1751 & n3434 ) | ( ~n1751 & n3435 ) | ( n3434 & n3435 ) ;
  assign n3437 = ( ~n1787 & n3434 ) | ( ~n1787 & n3435 ) | ( n3434 & n3435 ) ;
  assign n3438 = ( n1794 & n3434 ) | ( n1794 & n3435 ) | ( n3434 & n3435 ) ;
  assign n3439 = ( n1783 & n3437 ) | ( n1783 & n3438 ) | ( n3437 & n3438 ) ;
  assign n3440 = ( n1643 & n3436 ) | ( n1643 & n3439 ) | ( n3436 & n3439 ) ;
  assign n3441 = ( ~n1822 & n3436 ) | ( ~n1822 & n3439 ) | ( n3436 & n3439 ) ;
  assign n3442 = ( ~n1324 & n3440 ) | ( ~n1324 & n3441 ) | ( n3440 & n3441 ) ;
  assign n3443 = x122 & ~n1767 ;
  assign n3444 = x122 & n1771 ;
  assign n3445 = ( n1751 & n3443 ) | ( n1751 & n3444 ) | ( n3443 & n3444 ) ;
  assign n3446 = ( n1787 & n3443 ) | ( n1787 & n3444 ) | ( n3443 & n3444 ) ;
  assign n3447 = ( ~n1794 & n3443 ) | ( ~n1794 & n3444 ) | ( n3443 & n3444 ) ;
  assign n3448 = ( ~n1783 & n3446 ) | ( ~n1783 & n3447 ) | ( n3446 & n3447 ) ;
  assign n3449 = ( ~n1643 & n3445 ) | ( ~n1643 & n3448 ) | ( n3445 & n3448 ) ;
  assign n3450 = ( n1822 & n3445 ) | ( n1822 & n3448 ) | ( n3445 & n3448 ) ;
  assign n3451 = ( n1324 & n3449 ) | ( n1324 & n3450 ) | ( n3449 & n3450 ) ;
  assign n3452 = n3442 | n3451 ;
  assign n3453 = n3433 & ~n3452 ;
  assign n3454 = n3410 | n3453 ;
  assign n3455 = x249 & n1767 ;
  assign n3456 = x249 & ~n1771 ;
  assign n3457 = ( ~n1751 & n3455 ) | ( ~n1751 & n3456 ) | ( n3455 & n3456 ) ;
  assign n3458 = ( ~n1787 & n3455 ) | ( ~n1787 & n3456 ) | ( n3455 & n3456 ) ;
  assign n3459 = ( n1794 & n3455 ) | ( n1794 & n3456 ) | ( n3455 & n3456 ) ;
  assign n3460 = ( n1783 & n3458 ) | ( n1783 & n3459 ) | ( n3458 & n3459 ) ;
  assign n3461 = ( n1643 & n3457 ) | ( n1643 & n3460 ) | ( n3457 & n3460 ) ;
  assign n3462 = ( ~n1822 & n3457 ) | ( ~n1822 & n3460 ) | ( n3457 & n3460 ) ;
  assign n3463 = ( ~n1324 & n3461 ) | ( ~n1324 & n3462 ) | ( n3461 & n3462 ) ;
  assign n3464 = x121 & ~n1767 ;
  assign n3465 = x121 & n1771 ;
  assign n3466 = ( n1751 & n3464 ) | ( n1751 & n3465 ) | ( n3464 & n3465 ) ;
  assign n3467 = ( n1787 & n3464 ) | ( n1787 & n3465 ) | ( n3464 & n3465 ) ;
  assign n3468 = ( ~n1794 & n3464 ) | ( ~n1794 & n3465 ) | ( n3464 & n3465 ) ;
  assign n3469 = ( ~n1783 & n3467 ) | ( ~n1783 & n3468 ) | ( n3467 & n3468 ) ;
  assign n3470 = ( ~n1643 & n3466 ) | ( ~n1643 & n3469 ) | ( n3466 & n3469 ) ;
  assign n3471 = ( n1822 & n3466 ) | ( n1822 & n3469 ) | ( n3466 & n3469 ) ;
  assign n3472 = ( n1324 & n3470 ) | ( n1324 & n3471 ) | ( n3470 & n3471 ) ;
  assign n3473 = n3463 | n3472 ;
  assign n3474 = x505 & n991 ;
  assign n3475 = x505 & ~n995 ;
  assign n3476 = ( ~n1104 & n3474 ) | ( ~n1104 & n3475 ) | ( n3474 & n3475 ) ;
  assign n3477 = ( ~n1119 & n3474 ) | ( ~n1119 & n3475 ) | ( n3474 & n3475 ) ;
  assign n3478 = ( n1126 & n3474 ) | ( n1126 & n3475 ) | ( n3474 & n3475 ) ;
  assign n3479 = ( n1115 & n3477 ) | ( n1115 & n3478 ) | ( n3477 & n3478 ) ;
  assign n3480 = ( n975 & n3476 ) | ( n975 & n3479 ) | ( n3476 & n3479 ) ;
  assign n3481 = ( ~n1154 & n3476 ) | ( ~n1154 & n3479 ) | ( n3476 & n3479 ) ;
  assign n3482 = ( x409 & n3480 ) | ( x409 & n3481 ) | ( n3480 & n3481 ) ;
  assign n3483 = ( ~x281 & n3480 ) | ( ~x281 & n3481 ) | ( n3480 & n3481 ) ;
  assign n3484 = ( ~n656 & n3482 ) | ( ~n656 & n3483 ) | ( n3482 & n3483 ) ;
  assign n3485 = x377 & ~n991 ;
  assign n3486 = x377 & n995 ;
  assign n3487 = ( n1104 & n3485 ) | ( n1104 & n3486 ) | ( n3485 & n3486 ) ;
  assign n3488 = ( n1119 & n3485 ) | ( n1119 & n3486 ) | ( n3485 & n3486 ) ;
  assign n3489 = ( ~n1126 & n3485 ) | ( ~n1126 & n3486 ) | ( n3485 & n3486 ) ;
  assign n3490 = ( ~n1115 & n3488 ) | ( ~n1115 & n3489 ) | ( n3488 & n3489 ) ;
  assign n3491 = ( ~n975 & n3487 ) | ( ~n975 & n3490 ) | ( n3487 & n3490 ) ;
  assign n3492 = ( n1154 & n3487 ) | ( n1154 & n3490 ) | ( n3487 & n3490 ) ;
  assign n3493 = ( ~x409 & n3491 ) | ( ~x409 & n3492 ) | ( n3491 & n3492 ) ;
  assign n3494 = ( x281 & n3491 ) | ( x281 & n3492 ) | ( n3491 & n3492 ) ;
  assign n3495 = ( n656 & n3493 ) | ( n656 & n3494 ) | ( n3493 & n3494 ) ;
  assign n3496 = n3484 | n3495 ;
  assign n3497 = ~n3473 & n3496 ;
  assign n3498 = x504 & n991 ;
  assign n3499 = x504 & ~n995 ;
  assign n3500 = ( ~n1104 & n3498 ) | ( ~n1104 & n3499 ) | ( n3498 & n3499 ) ;
  assign n3501 = ( ~n1119 & n3498 ) | ( ~n1119 & n3499 ) | ( n3498 & n3499 ) ;
  assign n3502 = ( n1126 & n3498 ) | ( n1126 & n3499 ) | ( n3498 & n3499 ) ;
  assign n3503 = ( n1115 & n3501 ) | ( n1115 & n3502 ) | ( n3501 & n3502 ) ;
  assign n3504 = ( n975 & n3500 ) | ( n975 & n3503 ) | ( n3500 & n3503 ) ;
  assign n3505 = ( ~n1154 & n3500 ) | ( ~n1154 & n3503 ) | ( n3500 & n3503 ) ;
  assign n3506 = ( x409 & n3504 ) | ( x409 & n3505 ) | ( n3504 & n3505 ) ;
  assign n3507 = ( ~x281 & n3504 ) | ( ~x281 & n3505 ) | ( n3504 & n3505 ) ;
  assign n3508 = ( ~n656 & n3506 ) | ( ~n656 & n3507 ) | ( n3506 & n3507 ) ;
  assign n3509 = x376 & ~n991 ;
  assign n3510 = x376 & n995 ;
  assign n3511 = ( n1104 & n3509 ) | ( n1104 & n3510 ) | ( n3509 & n3510 ) ;
  assign n3512 = ( n1119 & n3509 ) | ( n1119 & n3510 ) | ( n3509 & n3510 ) ;
  assign n3513 = ( ~n1126 & n3509 ) | ( ~n1126 & n3510 ) | ( n3509 & n3510 ) ;
  assign n3514 = ( ~n1115 & n3512 ) | ( ~n1115 & n3513 ) | ( n3512 & n3513 ) ;
  assign n3515 = ( ~n975 & n3511 ) | ( ~n975 & n3514 ) | ( n3511 & n3514 ) ;
  assign n3516 = ( n1154 & n3511 ) | ( n1154 & n3514 ) | ( n3511 & n3514 ) ;
  assign n3517 = ( ~x409 & n3515 ) | ( ~x409 & n3516 ) | ( n3515 & n3516 ) ;
  assign n3518 = ( x281 & n3515 ) | ( x281 & n3516 ) | ( n3515 & n3516 ) ;
  assign n3519 = ( n656 & n3517 ) | ( n656 & n3518 ) | ( n3517 & n3518 ) ;
  assign n3520 = n3508 | n3519 ;
  assign n3521 = x248 & n1767 ;
  assign n3522 = x248 & ~n1771 ;
  assign n3523 = ( ~n1751 & n3521 ) | ( ~n1751 & n3522 ) | ( n3521 & n3522 ) ;
  assign n3524 = ( ~n1787 & n3521 ) | ( ~n1787 & n3522 ) | ( n3521 & n3522 ) ;
  assign n3525 = ( n1794 & n3521 ) | ( n1794 & n3522 ) | ( n3521 & n3522 ) ;
  assign n3526 = ( n1783 & n3524 ) | ( n1783 & n3525 ) | ( n3524 & n3525 ) ;
  assign n3527 = ( n1643 & n3523 ) | ( n1643 & n3526 ) | ( n3523 & n3526 ) ;
  assign n3528 = ( ~n1822 & n3523 ) | ( ~n1822 & n3526 ) | ( n3523 & n3526 ) ;
  assign n3529 = ( ~n1324 & n3527 ) | ( ~n1324 & n3528 ) | ( n3527 & n3528 ) ;
  assign n3530 = x120 & ~n1767 ;
  assign n3531 = x120 & n1771 ;
  assign n3532 = ( n1751 & n3530 ) | ( n1751 & n3531 ) | ( n3530 & n3531 ) ;
  assign n3533 = ( n1787 & n3530 ) | ( n1787 & n3531 ) | ( n3530 & n3531 ) ;
  assign n3534 = ( ~n1794 & n3530 ) | ( ~n1794 & n3531 ) | ( n3530 & n3531 ) ;
  assign n3535 = ( ~n1783 & n3533 ) | ( ~n1783 & n3534 ) | ( n3533 & n3534 ) ;
  assign n3536 = ( ~n1643 & n3532 ) | ( ~n1643 & n3535 ) | ( n3532 & n3535 ) ;
  assign n3537 = ( n1822 & n3532 ) | ( n1822 & n3535 ) | ( n3532 & n3535 ) ;
  assign n3538 = ( n1324 & n3536 ) | ( n1324 & n3537 ) | ( n3536 & n3537 ) ;
  assign n3539 = n3529 | n3538 ;
  assign n3540 = n3520 & ~n3539 ;
  assign n3541 = n3497 | n3540 ;
  assign n3542 = n3454 | n3541 ;
  assign n3543 = x247 & n1767 ;
  assign n3544 = x247 & ~n1771 ;
  assign n3545 = ( ~n1751 & n3543 ) | ( ~n1751 & n3544 ) | ( n3543 & n3544 ) ;
  assign n3546 = ( ~n1787 & n3543 ) | ( ~n1787 & n3544 ) | ( n3543 & n3544 ) ;
  assign n3547 = ( n1794 & n3543 ) | ( n1794 & n3544 ) | ( n3543 & n3544 ) ;
  assign n3548 = ( n1783 & n3546 ) | ( n1783 & n3547 ) | ( n3546 & n3547 ) ;
  assign n3549 = ( n1643 & n3545 ) | ( n1643 & n3548 ) | ( n3545 & n3548 ) ;
  assign n3550 = ( ~n1822 & n3545 ) | ( ~n1822 & n3548 ) | ( n3545 & n3548 ) ;
  assign n3551 = ( ~n1324 & n3549 ) | ( ~n1324 & n3550 ) | ( n3549 & n3550 ) ;
  assign n3552 = x119 & ~n1767 ;
  assign n3553 = x119 & n1771 ;
  assign n3554 = ( n1751 & n3552 ) | ( n1751 & n3553 ) | ( n3552 & n3553 ) ;
  assign n3555 = ( n1787 & n3552 ) | ( n1787 & n3553 ) | ( n3552 & n3553 ) ;
  assign n3556 = ( ~n1794 & n3552 ) | ( ~n1794 & n3553 ) | ( n3552 & n3553 ) ;
  assign n3557 = ( ~n1783 & n3555 ) | ( ~n1783 & n3556 ) | ( n3555 & n3556 ) ;
  assign n3558 = ( ~n1643 & n3554 ) | ( ~n1643 & n3557 ) | ( n3554 & n3557 ) ;
  assign n3559 = ( n1822 & n3554 ) | ( n1822 & n3557 ) | ( n3554 & n3557 ) ;
  assign n3560 = ( n1324 & n3558 ) | ( n1324 & n3559 ) | ( n3558 & n3559 ) ;
  assign n3561 = n3551 | n3560 ;
  assign n3562 = x503 & n991 ;
  assign n3563 = x503 & ~n995 ;
  assign n3564 = ( ~n1104 & n3562 ) | ( ~n1104 & n3563 ) | ( n3562 & n3563 ) ;
  assign n3565 = ( ~n1119 & n3562 ) | ( ~n1119 & n3563 ) | ( n3562 & n3563 ) ;
  assign n3566 = ( n1126 & n3562 ) | ( n1126 & n3563 ) | ( n3562 & n3563 ) ;
  assign n3567 = ( n1115 & n3565 ) | ( n1115 & n3566 ) | ( n3565 & n3566 ) ;
  assign n3568 = ( n975 & n3564 ) | ( n975 & n3567 ) | ( n3564 & n3567 ) ;
  assign n3569 = ( ~n1154 & n3564 ) | ( ~n1154 & n3567 ) | ( n3564 & n3567 ) ;
  assign n3570 = ( x409 & n3568 ) | ( x409 & n3569 ) | ( n3568 & n3569 ) ;
  assign n3571 = ( ~x281 & n3568 ) | ( ~x281 & n3569 ) | ( n3568 & n3569 ) ;
  assign n3572 = ( ~n656 & n3570 ) | ( ~n656 & n3571 ) | ( n3570 & n3571 ) ;
  assign n3573 = x375 & ~n991 ;
  assign n3574 = x375 & n995 ;
  assign n3575 = ( n1104 & n3573 ) | ( n1104 & n3574 ) | ( n3573 & n3574 ) ;
  assign n3576 = ( n1119 & n3573 ) | ( n1119 & n3574 ) | ( n3573 & n3574 ) ;
  assign n3577 = ( ~n1126 & n3573 ) | ( ~n1126 & n3574 ) | ( n3573 & n3574 ) ;
  assign n3578 = ( ~n1115 & n3576 ) | ( ~n1115 & n3577 ) | ( n3576 & n3577 ) ;
  assign n3579 = ( ~n975 & n3575 ) | ( ~n975 & n3578 ) | ( n3575 & n3578 ) ;
  assign n3580 = ( n1154 & n3575 ) | ( n1154 & n3578 ) | ( n3575 & n3578 ) ;
  assign n3581 = ( ~x409 & n3579 ) | ( ~x409 & n3580 ) | ( n3579 & n3580 ) ;
  assign n3582 = ( x281 & n3579 ) | ( x281 & n3580 ) | ( n3579 & n3580 ) ;
  assign n3583 = ( n656 & n3581 ) | ( n656 & n3582 ) | ( n3581 & n3582 ) ;
  assign n3584 = n3572 | n3583 ;
  assign n3585 = ~n3561 & n3584 ;
  assign n3586 = x502 & n991 ;
  assign n3587 = x502 & ~n995 ;
  assign n3588 = ( ~n1104 & n3586 ) | ( ~n1104 & n3587 ) | ( n3586 & n3587 ) ;
  assign n3589 = ( ~n1119 & n3586 ) | ( ~n1119 & n3587 ) | ( n3586 & n3587 ) ;
  assign n3590 = ( n1126 & n3586 ) | ( n1126 & n3587 ) | ( n3586 & n3587 ) ;
  assign n3591 = ( n1115 & n3589 ) | ( n1115 & n3590 ) | ( n3589 & n3590 ) ;
  assign n3592 = ( n975 & n3588 ) | ( n975 & n3591 ) | ( n3588 & n3591 ) ;
  assign n3593 = ( ~n1154 & n3588 ) | ( ~n1154 & n3591 ) | ( n3588 & n3591 ) ;
  assign n3594 = ( x409 & n3592 ) | ( x409 & n3593 ) | ( n3592 & n3593 ) ;
  assign n3595 = ( ~x281 & n3592 ) | ( ~x281 & n3593 ) | ( n3592 & n3593 ) ;
  assign n3596 = ( ~n656 & n3594 ) | ( ~n656 & n3595 ) | ( n3594 & n3595 ) ;
  assign n3597 = x374 & ~n991 ;
  assign n3598 = x374 & n995 ;
  assign n3599 = ( n1104 & n3597 ) | ( n1104 & n3598 ) | ( n3597 & n3598 ) ;
  assign n3600 = ( n1119 & n3597 ) | ( n1119 & n3598 ) | ( n3597 & n3598 ) ;
  assign n3601 = ( ~n1126 & n3597 ) | ( ~n1126 & n3598 ) | ( n3597 & n3598 ) ;
  assign n3602 = ( ~n1115 & n3600 ) | ( ~n1115 & n3601 ) | ( n3600 & n3601 ) ;
  assign n3603 = ( ~n975 & n3599 ) | ( ~n975 & n3602 ) | ( n3599 & n3602 ) ;
  assign n3604 = ( n1154 & n3599 ) | ( n1154 & n3602 ) | ( n3599 & n3602 ) ;
  assign n3605 = ( ~x409 & n3603 ) | ( ~x409 & n3604 ) | ( n3603 & n3604 ) ;
  assign n3606 = ( x281 & n3603 ) | ( x281 & n3604 ) | ( n3603 & n3604 ) ;
  assign n3607 = ( n656 & n3605 ) | ( n656 & n3606 ) | ( n3605 & n3606 ) ;
  assign n3608 = n3596 | n3607 ;
  assign n3609 = x246 & n1767 ;
  assign n3610 = x246 & ~n1771 ;
  assign n3611 = ( ~n1751 & n3609 ) | ( ~n1751 & n3610 ) | ( n3609 & n3610 ) ;
  assign n3612 = ( ~n1787 & n3609 ) | ( ~n1787 & n3610 ) | ( n3609 & n3610 ) ;
  assign n3613 = ( n1794 & n3609 ) | ( n1794 & n3610 ) | ( n3609 & n3610 ) ;
  assign n3614 = ( n1783 & n3612 ) | ( n1783 & n3613 ) | ( n3612 & n3613 ) ;
  assign n3615 = ( n1643 & n3611 ) | ( n1643 & n3614 ) | ( n3611 & n3614 ) ;
  assign n3616 = ( ~n1822 & n3611 ) | ( ~n1822 & n3614 ) | ( n3611 & n3614 ) ;
  assign n3617 = ( ~n1324 & n3615 ) | ( ~n1324 & n3616 ) | ( n3615 & n3616 ) ;
  assign n3618 = x118 & ~n1767 ;
  assign n3619 = x118 & n1771 ;
  assign n3620 = ( n1751 & n3618 ) | ( n1751 & n3619 ) | ( n3618 & n3619 ) ;
  assign n3621 = ( n1787 & n3618 ) | ( n1787 & n3619 ) | ( n3618 & n3619 ) ;
  assign n3622 = ( ~n1794 & n3618 ) | ( ~n1794 & n3619 ) | ( n3618 & n3619 ) ;
  assign n3623 = ( ~n1783 & n3621 ) | ( ~n1783 & n3622 ) | ( n3621 & n3622 ) ;
  assign n3624 = ( ~n1643 & n3620 ) | ( ~n1643 & n3623 ) | ( n3620 & n3623 ) ;
  assign n3625 = ( n1822 & n3620 ) | ( n1822 & n3623 ) | ( n3620 & n3623 ) ;
  assign n3626 = ( n1324 & n3624 ) | ( n1324 & n3625 ) | ( n3624 & n3625 ) ;
  assign n3627 = n3617 | n3626 ;
  assign n3628 = n3608 & ~n3627 ;
  assign n3629 = n3585 | n3628 ;
  assign n3630 = x245 & n1767 ;
  assign n3631 = x245 & ~n1771 ;
  assign n3632 = ( ~n1751 & n3630 ) | ( ~n1751 & n3631 ) | ( n3630 & n3631 ) ;
  assign n3633 = ( ~n1787 & n3630 ) | ( ~n1787 & n3631 ) | ( n3630 & n3631 ) ;
  assign n3634 = ( n1794 & n3630 ) | ( n1794 & n3631 ) | ( n3630 & n3631 ) ;
  assign n3635 = ( n1783 & n3633 ) | ( n1783 & n3634 ) | ( n3633 & n3634 ) ;
  assign n3636 = ( n1643 & n3632 ) | ( n1643 & n3635 ) | ( n3632 & n3635 ) ;
  assign n3637 = ( ~n1822 & n3632 ) | ( ~n1822 & n3635 ) | ( n3632 & n3635 ) ;
  assign n3638 = ( ~n1324 & n3636 ) | ( ~n1324 & n3637 ) | ( n3636 & n3637 ) ;
  assign n3639 = x117 & ~n1767 ;
  assign n3640 = x117 & n1771 ;
  assign n3641 = ( n1751 & n3639 ) | ( n1751 & n3640 ) | ( n3639 & n3640 ) ;
  assign n3642 = ( n1787 & n3639 ) | ( n1787 & n3640 ) | ( n3639 & n3640 ) ;
  assign n3643 = ( ~n1794 & n3639 ) | ( ~n1794 & n3640 ) | ( n3639 & n3640 ) ;
  assign n3644 = ( ~n1783 & n3642 ) | ( ~n1783 & n3643 ) | ( n3642 & n3643 ) ;
  assign n3645 = ( ~n1643 & n3641 ) | ( ~n1643 & n3644 ) | ( n3641 & n3644 ) ;
  assign n3646 = ( n1822 & n3641 ) | ( n1822 & n3644 ) | ( n3641 & n3644 ) ;
  assign n3647 = ( n1324 & n3645 ) | ( n1324 & n3646 ) | ( n3645 & n3646 ) ;
  assign n3648 = n3638 | n3647 ;
  assign n3649 = x501 & n991 ;
  assign n3650 = x501 & ~n995 ;
  assign n3651 = ( ~n1104 & n3649 ) | ( ~n1104 & n3650 ) | ( n3649 & n3650 ) ;
  assign n3652 = ( ~n1119 & n3649 ) | ( ~n1119 & n3650 ) | ( n3649 & n3650 ) ;
  assign n3653 = ( n1126 & n3649 ) | ( n1126 & n3650 ) | ( n3649 & n3650 ) ;
  assign n3654 = ( n1115 & n3652 ) | ( n1115 & n3653 ) | ( n3652 & n3653 ) ;
  assign n3655 = ( n975 & n3651 ) | ( n975 & n3654 ) | ( n3651 & n3654 ) ;
  assign n3656 = ( ~n1154 & n3651 ) | ( ~n1154 & n3654 ) | ( n3651 & n3654 ) ;
  assign n3657 = ( x409 & n3655 ) | ( x409 & n3656 ) | ( n3655 & n3656 ) ;
  assign n3658 = ( ~x281 & n3655 ) | ( ~x281 & n3656 ) | ( n3655 & n3656 ) ;
  assign n3659 = ( ~n656 & n3657 ) | ( ~n656 & n3658 ) | ( n3657 & n3658 ) ;
  assign n3660 = x373 & ~n991 ;
  assign n3661 = x373 & n995 ;
  assign n3662 = ( n1104 & n3660 ) | ( n1104 & n3661 ) | ( n3660 & n3661 ) ;
  assign n3663 = ( n1119 & n3660 ) | ( n1119 & n3661 ) | ( n3660 & n3661 ) ;
  assign n3664 = ( ~n1126 & n3660 ) | ( ~n1126 & n3661 ) | ( n3660 & n3661 ) ;
  assign n3665 = ( ~n1115 & n3663 ) | ( ~n1115 & n3664 ) | ( n3663 & n3664 ) ;
  assign n3666 = ( ~n975 & n3662 ) | ( ~n975 & n3665 ) | ( n3662 & n3665 ) ;
  assign n3667 = ( n1154 & n3662 ) | ( n1154 & n3665 ) | ( n3662 & n3665 ) ;
  assign n3668 = ( ~x409 & n3666 ) | ( ~x409 & n3667 ) | ( n3666 & n3667 ) ;
  assign n3669 = ( x281 & n3666 ) | ( x281 & n3667 ) | ( n3666 & n3667 ) ;
  assign n3670 = ( n656 & n3668 ) | ( n656 & n3669 ) | ( n3668 & n3669 ) ;
  assign n3671 = n3659 | n3670 ;
  assign n3672 = x244 & n1767 ;
  assign n3673 = x244 & ~n1771 ;
  assign n3674 = ( ~n1751 & n3672 ) | ( ~n1751 & n3673 ) | ( n3672 & n3673 ) ;
  assign n3675 = ( ~n1787 & n3672 ) | ( ~n1787 & n3673 ) | ( n3672 & n3673 ) ;
  assign n3676 = ( n1794 & n3672 ) | ( n1794 & n3673 ) | ( n3672 & n3673 ) ;
  assign n3677 = ( n1783 & n3675 ) | ( n1783 & n3676 ) | ( n3675 & n3676 ) ;
  assign n3678 = ( n1643 & n3674 ) | ( n1643 & n3677 ) | ( n3674 & n3677 ) ;
  assign n3679 = ( ~n1822 & n3674 ) | ( ~n1822 & n3677 ) | ( n3674 & n3677 ) ;
  assign n3680 = ( ~n1324 & n3678 ) | ( ~n1324 & n3679 ) | ( n3678 & n3679 ) ;
  assign n3681 = x116 & ~n1767 ;
  assign n3682 = x116 & n1771 ;
  assign n3683 = ( n1751 & n3681 ) | ( n1751 & n3682 ) | ( n3681 & n3682 ) ;
  assign n3684 = ( n1787 & n3681 ) | ( n1787 & n3682 ) | ( n3681 & n3682 ) ;
  assign n3685 = ( ~n1794 & n3681 ) | ( ~n1794 & n3682 ) | ( n3681 & n3682 ) ;
  assign n3686 = ( ~n1783 & n3684 ) | ( ~n1783 & n3685 ) | ( n3684 & n3685 ) ;
  assign n3687 = ( ~n1643 & n3683 ) | ( ~n1643 & n3686 ) | ( n3683 & n3686 ) ;
  assign n3688 = ( n1822 & n3683 ) | ( n1822 & n3686 ) | ( n3683 & n3686 ) ;
  assign n3689 = ( n1324 & n3687 ) | ( n1324 & n3688 ) | ( n3687 & n3688 ) ;
  assign n3690 = n3680 | n3689 ;
  assign n3691 = x500 & n991 ;
  assign n3692 = x500 & ~n995 ;
  assign n3693 = ( ~n1104 & n3691 ) | ( ~n1104 & n3692 ) | ( n3691 & n3692 ) ;
  assign n3694 = ( ~n1119 & n3691 ) | ( ~n1119 & n3692 ) | ( n3691 & n3692 ) ;
  assign n3695 = ( n1126 & n3691 ) | ( n1126 & n3692 ) | ( n3691 & n3692 ) ;
  assign n3696 = ( n1115 & n3694 ) | ( n1115 & n3695 ) | ( n3694 & n3695 ) ;
  assign n3697 = ( n975 & n3693 ) | ( n975 & n3696 ) | ( n3693 & n3696 ) ;
  assign n3698 = ( ~n1154 & n3693 ) | ( ~n1154 & n3696 ) | ( n3693 & n3696 ) ;
  assign n3699 = ( x409 & n3697 ) | ( x409 & n3698 ) | ( n3697 & n3698 ) ;
  assign n3700 = ( ~x281 & n3697 ) | ( ~x281 & n3698 ) | ( n3697 & n3698 ) ;
  assign n3701 = ( ~n656 & n3699 ) | ( ~n656 & n3700 ) | ( n3699 & n3700 ) ;
  assign n3702 = x372 & ~n991 ;
  assign n3703 = x372 & n995 ;
  assign n3704 = ( n1104 & n3702 ) | ( n1104 & n3703 ) | ( n3702 & n3703 ) ;
  assign n3705 = ( n1119 & n3702 ) | ( n1119 & n3703 ) | ( n3702 & n3703 ) ;
  assign n3706 = ( ~n1126 & n3702 ) | ( ~n1126 & n3703 ) | ( n3702 & n3703 ) ;
  assign n3707 = ( ~n1115 & n3705 ) | ( ~n1115 & n3706 ) | ( n3705 & n3706 ) ;
  assign n3708 = ( ~n975 & n3704 ) | ( ~n975 & n3707 ) | ( n3704 & n3707 ) ;
  assign n3709 = ( n1154 & n3704 ) | ( n1154 & n3707 ) | ( n3704 & n3707 ) ;
  assign n3710 = ( ~x409 & n3708 ) | ( ~x409 & n3709 ) | ( n3708 & n3709 ) ;
  assign n3711 = ( x281 & n3708 ) | ( x281 & n3709 ) | ( n3708 & n3709 ) ;
  assign n3712 = ( n656 & n3710 ) | ( n656 & n3711 ) | ( n3710 & n3711 ) ;
  assign n3713 = n3701 | n3712 ;
  assign n3714 = n3690 & ~n3713 ;
  assign n3715 = ( n3648 & ~n3671 ) | ( n3648 & n3714 ) | ( ~n3671 & n3714 ) ;
  assign n3716 = ~n3629 & n3715 ;
  assign n3717 = n3561 & ~n3584 ;
  assign n3718 = ~n3608 & n3627 ;
  assign n3719 = ~n3585 & n3718 ;
  assign n3720 = n3717 | n3719 ;
  assign n3721 = n3716 | n3720 ;
  assign n3722 = ~n3542 & n3721 ;
  assign n3723 = ~n3648 & n3671 ;
  assign n3724 = ~n3690 & n3713 ;
  assign n3725 = n3723 | n3724 ;
  assign n3726 = n3629 | n3725 ;
  assign n3727 = x243 & n1767 ;
  assign n3728 = x243 & ~n1771 ;
  assign n3729 = ( ~n1751 & n3727 ) | ( ~n1751 & n3728 ) | ( n3727 & n3728 ) ;
  assign n3730 = ( ~n1787 & n3727 ) | ( ~n1787 & n3728 ) | ( n3727 & n3728 ) ;
  assign n3731 = ( n1794 & n3727 ) | ( n1794 & n3728 ) | ( n3727 & n3728 ) ;
  assign n3732 = ( n1783 & n3730 ) | ( n1783 & n3731 ) | ( n3730 & n3731 ) ;
  assign n3733 = ( n1643 & n3729 ) | ( n1643 & n3732 ) | ( n3729 & n3732 ) ;
  assign n3734 = ( ~n1822 & n3729 ) | ( ~n1822 & n3732 ) | ( n3729 & n3732 ) ;
  assign n3735 = ( ~n1324 & n3733 ) | ( ~n1324 & n3734 ) | ( n3733 & n3734 ) ;
  assign n3736 = x115 & ~n1767 ;
  assign n3737 = x115 & n1771 ;
  assign n3738 = ( n1751 & n3736 ) | ( n1751 & n3737 ) | ( n3736 & n3737 ) ;
  assign n3739 = ( n1787 & n3736 ) | ( n1787 & n3737 ) | ( n3736 & n3737 ) ;
  assign n3740 = ( ~n1794 & n3736 ) | ( ~n1794 & n3737 ) | ( n3736 & n3737 ) ;
  assign n3741 = ( ~n1783 & n3739 ) | ( ~n1783 & n3740 ) | ( n3739 & n3740 ) ;
  assign n3742 = ( ~n1643 & n3738 ) | ( ~n1643 & n3741 ) | ( n3738 & n3741 ) ;
  assign n3743 = ( n1822 & n3738 ) | ( n1822 & n3741 ) | ( n3738 & n3741 ) ;
  assign n3744 = ( n1324 & n3742 ) | ( n1324 & n3743 ) | ( n3742 & n3743 ) ;
  assign n3745 = n3735 | n3744 ;
  assign n3746 = x499 & n991 ;
  assign n3747 = x499 & ~n995 ;
  assign n3748 = ( ~n1104 & n3746 ) | ( ~n1104 & n3747 ) | ( n3746 & n3747 ) ;
  assign n3749 = ( ~n1119 & n3746 ) | ( ~n1119 & n3747 ) | ( n3746 & n3747 ) ;
  assign n3750 = ( n1126 & n3746 ) | ( n1126 & n3747 ) | ( n3746 & n3747 ) ;
  assign n3751 = ( n1115 & n3749 ) | ( n1115 & n3750 ) | ( n3749 & n3750 ) ;
  assign n3752 = ( n975 & n3748 ) | ( n975 & n3751 ) | ( n3748 & n3751 ) ;
  assign n3753 = ( ~n1154 & n3748 ) | ( ~n1154 & n3751 ) | ( n3748 & n3751 ) ;
  assign n3754 = ( x409 & n3752 ) | ( x409 & n3753 ) | ( n3752 & n3753 ) ;
  assign n3755 = ( ~x281 & n3752 ) | ( ~x281 & n3753 ) | ( n3752 & n3753 ) ;
  assign n3756 = ( ~n656 & n3754 ) | ( ~n656 & n3755 ) | ( n3754 & n3755 ) ;
  assign n3757 = x371 & ~n991 ;
  assign n3758 = x371 & n995 ;
  assign n3759 = ( n1104 & n3757 ) | ( n1104 & n3758 ) | ( n3757 & n3758 ) ;
  assign n3760 = ( n1119 & n3757 ) | ( n1119 & n3758 ) | ( n3757 & n3758 ) ;
  assign n3761 = ( ~n1126 & n3757 ) | ( ~n1126 & n3758 ) | ( n3757 & n3758 ) ;
  assign n3762 = ( ~n1115 & n3760 ) | ( ~n1115 & n3761 ) | ( n3760 & n3761 ) ;
  assign n3763 = ( ~n975 & n3759 ) | ( ~n975 & n3762 ) | ( n3759 & n3762 ) ;
  assign n3764 = ( n1154 & n3759 ) | ( n1154 & n3762 ) | ( n3759 & n3762 ) ;
  assign n3765 = ( ~x409 & n3763 ) | ( ~x409 & n3764 ) | ( n3763 & n3764 ) ;
  assign n3766 = ( x281 & n3763 ) | ( x281 & n3764 ) | ( n3763 & n3764 ) ;
  assign n3767 = ( n656 & n3765 ) | ( n656 & n3766 ) | ( n3765 & n3766 ) ;
  assign n3768 = n3756 | n3767 ;
  assign n3769 = x498 & n991 ;
  assign n3770 = x498 & ~n995 ;
  assign n3771 = ( ~n1104 & n3769 ) | ( ~n1104 & n3770 ) | ( n3769 & n3770 ) ;
  assign n3772 = ( ~n1119 & n3769 ) | ( ~n1119 & n3770 ) | ( n3769 & n3770 ) ;
  assign n3773 = ( n1126 & n3769 ) | ( n1126 & n3770 ) | ( n3769 & n3770 ) ;
  assign n3774 = ( n1115 & n3772 ) | ( n1115 & n3773 ) | ( n3772 & n3773 ) ;
  assign n3775 = ( n975 & n3771 ) | ( n975 & n3774 ) | ( n3771 & n3774 ) ;
  assign n3776 = ( ~n1154 & n3771 ) | ( ~n1154 & n3774 ) | ( n3771 & n3774 ) ;
  assign n3777 = ( x409 & n3775 ) | ( x409 & n3776 ) | ( n3775 & n3776 ) ;
  assign n3778 = ( ~x281 & n3775 ) | ( ~x281 & n3776 ) | ( n3775 & n3776 ) ;
  assign n3779 = ( ~n656 & n3777 ) | ( ~n656 & n3778 ) | ( n3777 & n3778 ) ;
  assign n3780 = x370 & ~n991 ;
  assign n3781 = x370 & n995 ;
  assign n3782 = ( n1104 & n3780 ) | ( n1104 & n3781 ) | ( n3780 & n3781 ) ;
  assign n3783 = ( n1119 & n3780 ) | ( n1119 & n3781 ) | ( n3780 & n3781 ) ;
  assign n3784 = ( ~n1126 & n3780 ) | ( ~n1126 & n3781 ) | ( n3780 & n3781 ) ;
  assign n3785 = ( ~n1115 & n3783 ) | ( ~n1115 & n3784 ) | ( n3783 & n3784 ) ;
  assign n3786 = ( ~n975 & n3782 ) | ( ~n975 & n3785 ) | ( n3782 & n3785 ) ;
  assign n3787 = ( n1154 & n3782 ) | ( n1154 & n3785 ) | ( n3782 & n3785 ) ;
  assign n3788 = ( ~x409 & n3786 ) | ( ~x409 & n3787 ) | ( n3786 & n3787 ) ;
  assign n3789 = ( x281 & n3786 ) | ( x281 & n3787 ) | ( n3786 & n3787 ) ;
  assign n3790 = ( n656 & n3788 ) | ( n656 & n3789 ) | ( n3788 & n3789 ) ;
  assign n3791 = n3779 | n3790 ;
  assign n3792 = x242 & n1767 ;
  assign n3793 = x242 & ~n1771 ;
  assign n3794 = ( ~n1751 & n3792 ) | ( ~n1751 & n3793 ) | ( n3792 & n3793 ) ;
  assign n3795 = ( ~n1787 & n3792 ) | ( ~n1787 & n3793 ) | ( n3792 & n3793 ) ;
  assign n3796 = ( n1794 & n3792 ) | ( n1794 & n3793 ) | ( n3792 & n3793 ) ;
  assign n3797 = ( n1783 & n3795 ) | ( n1783 & n3796 ) | ( n3795 & n3796 ) ;
  assign n3798 = ( n1643 & n3794 ) | ( n1643 & n3797 ) | ( n3794 & n3797 ) ;
  assign n3799 = ( ~n1822 & n3794 ) | ( ~n1822 & n3797 ) | ( n3794 & n3797 ) ;
  assign n3800 = ( ~n1324 & n3798 ) | ( ~n1324 & n3799 ) | ( n3798 & n3799 ) ;
  assign n3801 = x114 & ~n1767 ;
  assign n3802 = x114 & n1771 ;
  assign n3803 = ( n1751 & n3801 ) | ( n1751 & n3802 ) | ( n3801 & n3802 ) ;
  assign n3804 = ( n1787 & n3801 ) | ( n1787 & n3802 ) | ( n3801 & n3802 ) ;
  assign n3805 = ( ~n1794 & n3801 ) | ( ~n1794 & n3802 ) | ( n3801 & n3802 ) ;
  assign n3806 = ( ~n1783 & n3804 ) | ( ~n1783 & n3805 ) | ( n3804 & n3805 ) ;
  assign n3807 = ( ~n1643 & n3803 ) | ( ~n1643 & n3806 ) | ( n3803 & n3806 ) ;
  assign n3808 = ( n1822 & n3803 ) | ( n1822 & n3806 ) | ( n3803 & n3806 ) ;
  assign n3809 = ( n1324 & n3807 ) | ( n1324 & n3808 ) | ( n3807 & n3808 ) ;
  assign n3810 = n3800 | n3809 ;
  assign n3811 = n3791 & ~n3810 ;
  assign n3812 = x241 & n1767 ;
  assign n3813 = x241 & ~n1771 ;
  assign n3814 = ( ~n1751 & n3812 ) | ( ~n1751 & n3813 ) | ( n3812 & n3813 ) ;
  assign n3815 = ( ~n1787 & n3812 ) | ( ~n1787 & n3813 ) | ( n3812 & n3813 ) ;
  assign n3816 = ( n1794 & n3812 ) | ( n1794 & n3813 ) | ( n3812 & n3813 ) ;
  assign n3817 = ( n1783 & n3815 ) | ( n1783 & n3816 ) | ( n3815 & n3816 ) ;
  assign n3818 = ( n1643 & n3814 ) | ( n1643 & n3817 ) | ( n3814 & n3817 ) ;
  assign n3819 = ( ~n1822 & n3814 ) | ( ~n1822 & n3817 ) | ( n3814 & n3817 ) ;
  assign n3820 = ( ~n1324 & n3818 ) | ( ~n1324 & n3819 ) | ( n3818 & n3819 ) ;
  assign n3821 = x113 & ~n1767 ;
  assign n3822 = x113 & n1771 ;
  assign n3823 = ( n1751 & n3821 ) | ( n1751 & n3822 ) | ( n3821 & n3822 ) ;
  assign n3824 = ( n1787 & n3821 ) | ( n1787 & n3822 ) | ( n3821 & n3822 ) ;
  assign n3825 = ( ~n1794 & n3821 ) | ( ~n1794 & n3822 ) | ( n3821 & n3822 ) ;
  assign n3826 = ( ~n1783 & n3824 ) | ( ~n1783 & n3825 ) | ( n3824 & n3825 ) ;
  assign n3827 = ( ~n1643 & n3823 ) | ( ~n1643 & n3826 ) | ( n3823 & n3826 ) ;
  assign n3828 = ( n1822 & n3823 ) | ( n1822 & n3826 ) | ( n3823 & n3826 ) ;
  assign n3829 = ( n1324 & n3827 ) | ( n1324 & n3828 ) | ( n3827 & n3828 ) ;
  assign n3830 = n3820 | n3829 ;
  assign n3831 = x497 & n991 ;
  assign n3832 = x497 & ~n995 ;
  assign n3833 = ( ~n1104 & n3831 ) | ( ~n1104 & n3832 ) | ( n3831 & n3832 ) ;
  assign n3834 = ( ~n1119 & n3831 ) | ( ~n1119 & n3832 ) | ( n3831 & n3832 ) ;
  assign n3835 = ( n1126 & n3831 ) | ( n1126 & n3832 ) | ( n3831 & n3832 ) ;
  assign n3836 = ( n1115 & n3834 ) | ( n1115 & n3835 ) | ( n3834 & n3835 ) ;
  assign n3837 = ( n975 & n3833 ) | ( n975 & n3836 ) | ( n3833 & n3836 ) ;
  assign n3838 = ( ~n1154 & n3833 ) | ( ~n1154 & n3836 ) | ( n3833 & n3836 ) ;
  assign n3839 = ( x409 & n3837 ) | ( x409 & n3838 ) | ( n3837 & n3838 ) ;
  assign n3840 = ( ~x281 & n3837 ) | ( ~x281 & n3838 ) | ( n3837 & n3838 ) ;
  assign n3841 = ( ~n656 & n3839 ) | ( ~n656 & n3840 ) | ( n3839 & n3840 ) ;
  assign n3842 = x369 & ~n991 ;
  assign n3843 = x369 & n995 ;
  assign n3844 = ( n1104 & n3842 ) | ( n1104 & n3843 ) | ( n3842 & n3843 ) ;
  assign n3845 = ( n1119 & n3842 ) | ( n1119 & n3843 ) | ( n3842 & n3843 ) ;
  assign n3846 = ( ~n1126 & n3842 ) | ( ~n1126 & n3843 ) | ( n3842 & n3843 ) ;
  assign n3847 = ( ~n1115 & n3845 ) | ( ~n1115 & n3846 ) | ( n3845 & n3846 ) ;
  assign n3848 = ( ~n975 & n3844 ) | ( ~n975 & n3847 ) | ( n3844 & n3847 ) ;
  assign n3849 = ( n1154 & n3844 ) | ( n1154 & n3847 ) | ( n3844 & n3847 ) ;
  assign n3850 = ( ~x409 & n3848 ) | ( ~x409 & n3849 ) | ( n3848 & n3849 ) ;
  assign n3851 = ( x281 & n3848 ) | ( x281 & n3849 ) | ( n3848 & n3849 ) ;
  assign n3852 = ( n656 & n3850 ) | ( n656 & n3851 ) | ( n3850 & n3851 ) ;
  assign n3853 = n3841 | n3852 ;
  assign n3854 = x496 & n991 ;
  assign n3855 = x496 & ~n995 ;
  assign n3856 = ( ~n1104 & n3854 ) | ( ~n1104 & n3855 ) | ( n3854 & n3855 ) ;
  assign n3857 = ( ~n1119 & n3854 ) | ( ~n1119 & n3855 ) | ( n3854 & n3855 ) ;
  assign n3858 = ( n1126 & n3854 ) | ( n1126 & n3855 ) | ( n3854 & n3855 ) ;
  assign n3859 = ( n1115 & n3857 ) | ( n1115 & n3858 ) | ( n3857 & n3858 ) ;
  assign n3860 = ( n975 & n3856 ) | ( n975 & n3859 ) | ( n3856 & n3859 ) ;
  assign n3861 = ( ~n1154 & n3856 ) | ( ~n1154 & n3859 ) | ( n3856 & n3859 ) ;
  assign n3862 = ( x409 & n3860 ) | ( x409 & n3861 ) | ( n3860 & n3861 ) ;
  assign n3863 = ( ~x281 & n3860 ) | ( ~x281 & n3861 ) | ( n3860 & n3861 ) ;
  assign n3864 = ( ~n656 & n3862 ) | ( ~n656 & n3863 ) | ( n3862 & n3863 ) ;
  assign n3865 = x368 & ~n991 ;
  assign n3866 = x368 & n995 ;
  assign n3867 = ( n1104 & n3865 ) | ( n1104 & n3866 ) | ( n3865 & n3866 ) ;
  assign n3868 = ( n1119 & n3865 ) | ( n1119 & n3866 ) | ( n3865 & n3866 ) ;
  assign n3869 = ( ~n1126 & n3865 ) | ( ~n1126 & n3866 ) | ( n3865 & n3866 ) ;
  assign n3870 = ( ~n1115 & n3868 ) | ( ~n1115 & n3869 ) | ( n3868 & n3869 ) ;
  assign n3871 = ( ~n975 & n3867 ) | ( ~n975 & n3870 ) | ( n3867 & n3870 ) ;
  assign n3872 = ( n1154 & n3867 ) | ( n1154 & n3870 ) | ( n3867 & n3870 ) ;
  assign n3873 = ( ~x409 & n3871 ) | ( ~x409 & n3872 ) | ( n3871 & n3872 ) ;
  assign n3874 = ( x281 & n3871 ) | ( x281 & n3872 ) | ( n3871 & n3872 ) ;
  assign n3875 = ( n656 & n3873 ) | ( n656 & n3874 ) | ( n3873 & n3874 ) ;
  assign n3876 = n3864 | n3875 ;
  assign n3877 = x240 & n1767 ;
  assign n3878 = x240 & ~n1771 ;
  assign n3879 = ( ~n1751 & n3877 ) | ( ~n1751 & n3878 ) | ( n3877 & n3878 ) ;
  assign n3880 = ( ~n1787 & n3877 ) | ( ~n1787 & n3878 ) | ( n3877 & n3878 ) ;
  assign n3881 = ( n1794 & n3877 ) | ( n1794 & n3878 ) | ( n3877 & n3878 ) ;
  assign n3882 = ( n1783 & n3880 ) | ( n1783 & n3881 ) | ( n3880 & n3881 ) ;
  assign n3883 = ( n1643 & n3879 ) | ( n1643 & n3882 ) | ( n3879 & n3882 ) ;
  assign n3884 = ( ~n1822 & n3879 ) | ( ~n1822 & n3882 ) | ( n3879 & n3882 ) ;
  assign n3885 = ( ~n1324 & n3883 ) | ( ~n1324 & n3884 ) | ( n3883 & n3884 ) ;
  assign n3886 = x112 & ~n1767 ;
  assign n3887 = x112 & n1771 ;
  assign n3888 = ( n1751 & n3886 ) | ( n1751 & n3887 ) | ( n3886 & n3887 ) ;
  assign n3889 = ( n1787 & n3886 ) | ( n1787 & n3887 ) | ( n3886 & n3887 ) ;
  assign n3890 = ( ~n1794 & n3886 ) | ( ~n1794 & n3887 ) | ( n3886 & n3887 ) ;
  assign n3891 = ( ~n1783 & n3889 ) | ( ~n1783 & n3890 ) | ( n3889 & n3890 ) ;
  assign n3892 = ( ~n1643 & n3888 ) | ( ~n1643 & n3891 ) | ( n3888 & n3891 ) ;
  assign n3893 = ( n1822 & n3888 ) | ( n1822 & n3891 ) | ( n3888 & n3891 ) ;
  assign n3894 = ( n1324 & n3892 ) | ( n1324 & n3893 ) | ( n3892 & n3893 ) ;
  assign n3895 = n3885 | n3894 ;
  assign n3896 = ~n3876 & n3895 ;
  assign n3897 = ( n3830 & ~n3853 ) | ( n3830 & n3896 ) | ( ~n3853 & n3896 ) ;
  assign n3898 = ~n3791 & n3810 ;
  assign n3899 = ~n3811 & n3898 ;
  assign n3900 = ( ~n3811 & n3897 ) | ( ~n3811 & n3899 ) | ( n3897 & n3899 ) ;
  assign n3901 = ( n3745 & ~n3768 ) | ( n3745 & n3900 ) | ( ~n3768 & n3900 ) ;
  assign n3902 = ~n3745 & n3768 ;
  assign n3903 = n3811 | n3902 ;
  assign n3904 = ~n3830 & n3853 ;
  assign n3905 = n3876 & ~n3895 ;
  assign n3906 = n3904 | n3905 ;
  assign n3907 = n3903 | n3906 ;
  assign n3908 = n3726 | n3907 ;
  assign n3909 = ( n3726 & ~n3901 ) | ( n3726 & n3908 ) | ( ~n3901 & n3908 ) ;
  assign n3910 = ( n3542 & ~n3722 ) | ( n3542 & n3909 ) | ( ~n3722 & n3909 ) ;
  assign n3911 = ~n3726 & n3901 ;
  assign n3912 = ( ~n3542 & n3722 ) | ( ~n3542 & n3911 ) | ( n3722 & n3911 ) ;
  assign n3913 = ( n3367 & ~n3910 ) | ( n3367 & n3912 ) | ( ~n3910 & n3912 ) ;
  assign n3914 = x254 & n1767 ;
  assign n3915 = x254 & ~n1771 ;
  assign n3916 = ( ~n1751 & n3914 ) | ( ~n1751 & n3915 ) | ( n3914 & n3915 ) ;
  assign n3917 = ( ~n1787 & n3914 ) | ( ~n1787 & n3915 ) | ( n3914 & n3915 ) ;
  assign n3918 = ( n1794 & n3914 ) | ( n1794 & n3915 ) | ( n3914 & n3915 ) ;
  assign n3919 = ( n1783 & n3917 ) | ( n1783 & n3918 ) | ( n3917 & n3918 ) ;
  assign n3920 = ( n1643 & n3916 ) | ( n1643 & n3919 ) | ( n3916 & n3919 ) ;
  assign n3921 = ( ~n1822 & n3916 ) | ( ~n1822 & n3919 ) | ( n3916 & n3919 ) ;
  assign n3922 = ( ~n1324 & n3920 ) | ( ~n1324 & n3921 ) | ( n3920 & n3921 ) ;
  assign n3923 = x126 & ~n1767 ;
  assign n3924 = x126 & n1771 ;
  assign n3925 = ( n1751 & n3923 ) | ( n1751 & n3924 ) | ( n3923 & n3924 ) ;
  assign n3926 = ( n1787 & n3923 ) | ( n1787 & n3924 ) | ( n3923 & n3924 ) ;
  assign n3927 = ( ~n1794 & n3923 ) | ( ~n1794 & n3924 ) | ( n3923 & n3924 ) ;
  assign n3928 = ( ~n1783 & n3926 ) | ( ~n1783 & n3927 ) | ( n3926 & n3927 ) ;
  assign n3929 = ( ~n1643 & n3925 ) | ( ~n1643 & n3928 ) | ( n3925 & n3928 ) ;
  assign n3930 = ( n1822 & n3925 ) | ( n1822 & n3928 ) | ( n3925 & n3928 ) ;
  assign n3931 = ( n1324 & n3929 ) | ( n1324 & n3930 ) | ( n3929 & n3930 ) ;
  assign n3932 = n3922 | n3931 ;
  assign n3933 = x510 & n991 ;
  assign n3934 = x510 & ~n995 ;
  assign n3935 = ( ~n1104 & n3933 ) | ( ~n1104 & n3934 ) | ( n3933 & n3934 ) ;
  assign n3936 = ( ~n1119 & n3933 ) | ( ~n1119 & n3934 ) | ( n3933 & n3934 ) ;
  assign n3937 = ( n1126 & n3933 ) | ( n1126 & n3934 ) | ( n3933 & n3934 ) ;
  assign n3938 = ( n1115 & n3936 ) | ( n1115 & n3937 ) | ( n3936 & n3937 ) ;
  assign n3939 = ( n975 & n3935 ) | ( n975 & n3938 ) | ( n3935 & n3938 ) ;
  assign n3940 = ( ~n1154 & n3935 ) | ( ~n1154 & n3938 ) | ( n3935 & n3938 ) ;
  assign n3941 = ( x409 & n3939 ) | ( x409 & n3940 ) | ( n3939 & n3940 ) ;
  assign n3942 = ( ~x281 & n3939 ) | ( ~x281 & n3940 ) | ( n3939 & n3940 ) ;
  assign n3943 = ( ~n656 & n3941 ) | ( ~n656 & n3942 ) | ( n3941 & n3942 ) ;
  assign n3944 = x382 & ~n991 ;
  assign n3945 = x382 & n995 ;
  assign n3946 = ( n1104 & n3944 ) | ( n1104 & n3945 ) | ( n3944 & n3945 ) ;
  assign n3947 = ( n1119 & n3944 ) | ( n1119 & n3945 ) | ( n3944 & n3945 ) ;
  assign n3948 = ( ~n1126 & n3944 ) | ( ~n1126 & n3945 ) | ( n3944 & n3945 ) ;
  assign n3949 = ( ~n1115 & n3947 ) | ( ~n1115 & n3948 ) | ( n3947 & n3948 ) ;
  assign n3950 = ( ~n975 & n3946 ) | ( ~n975 & n3949 ) | ( n3946 & n3949 ) ;
  assign n3951 = ( n1154 & n3946 ) | ( n1154 & n3949 ) | ( n3946 & n3949 ) ;
  assign n3952 = ( ~x409 & n3950 ) | ( ~x409 & n3951 ) | ( n3950 & n3951 ) ;
  assign n3953 = ( x281 & n3950 ) | ( x281 & n3951 ) | ( n3950 & n3951 ) ;
  assign n3954 = ( n656 & n3952 ) | ( n656 & n3953 ) | ( n3952 & n3953 ) ;
  assign n3955 = n3943 | n3954 ;
  assign n3956 = ~n3932 & n3955 ;
  assign n3957 = x253 & n1767 ;
  assign n3958 = x253 & ~n1771 ;
  assign n3959 = ( ~n1751 & n3957 ) | ( ~n1751 & n3958 ) | ( n3957 & n3958 ) ;
  assign n3960 = ( ~n1787 & n3957 ) | ( ~n1787 & n3958 ) | ( n3957 & n3958 ) ;
  assign n3961 = ( n1794 & n3957 ) | ( n1794 & n3958 ) | ( n3957 & n3958 ) ;
  assign n3962 = ( n1783 & n3960 ) | ( n1783 & n3961 ) | ( n3960 & n3961 ) ;
  assign n3963 = ( n1643 & n3959 ) | ( n1643 & n3962 ) | ( n3959 & n3962 ) ;
  assign n3964 = ( ~n1822 & n3959 ) | ( ~n1822 & n3962 ) | ( n3959 & n3962 ) ;
  assign n3965 = ( ~n1324 & n3963 ) | ( ~n1324 & n3964 ) | ( n3963 & n3964 ) ;
  assign n3966 = x125 & ~n1767 ;
  assign n3967 = x125 & n1771 ;
  assign n3968 = ( n1751 & n3966 ) | ( n1751 & n3967 ) | ( n3966 & n3967 ) ;
  assign n3969 = ( n1787 & n3966 ) | ( n1787 & n3967 ) | ( n3966 & n3967 ) ;
  assign n3970 = ( ~n1794 & n3966 ) | ( ~n1794 & n3967 ) | ( n3966 & n3967 ) ;
  assign n3971 = ( ~n1783 & n3969 ) | ( ~n1783 & n3970 ) | ( n3969 & n3970 ) ;
  assign n3972 = ( ~n1643 & n3968 ) | ( ~n1643 & n3971 ) | ( n3968 & n3971 ) ;
  assign n3973 = ( n1822 & n3968 ) | ( n1822 & n3971 ) | ( n3968 & n3971 ) ;
  assign n3974 = ( n1324 & n3972 ) | ( n1324 & n3973 ) | ( n3972 & n3973 ) ;
  assign n3975 = n3965 | n3974 ;
  assign n3976 = x509 & n991 ;
  assign n3977 = x509 & ~n995 ;
  assign n3978 = ( ~n1104 & n3976 ) | ( ~n1104 & n3977 ) | ( n3976 & n3977 ) ;
  assign n3979 = ( ~n1119 & n3976 ) | ( ~n1119 & n3977 ) | ( n3976 & n3977 ) ;
  assign n3980 = ( n1126 & n3976 ) | ( n1126 & n3977 ) | ( n3976 & n3977 ) ;
  assign n3981 = ( n1115 & n3979 ) | ( n1115 & n3980 ) | ( n3979 & n3980 ) ;
  assign n3982 = ( n975 & n3978 ) | ( n975 & n3981 ) | ( n3978 & n3981 ) ;
  assign n3983 = ( ~n1154 & n3978 ) | ( ~n1154 & n3981 ) | ( n3978 & n3981 ) ;
  assign n3984 = ( x409 & n3982 ) | ( x409 & n3983 ) | ( n3982 & n3983 ) ;
  assign n3985 = ( ~x281 & n3982 ) | ( ~x281 & n3983 ) | ( n3982 & n3983 ) ;
  assign n3986 = ( ~n656 & n3984 ) | ( ~n656 & n3985 ) | ( n3984 & n3985 ) ;
  assign n3987 = x381 & ~n991 ;
  assign n3988 = x381 & n995 ;
  assign n3989 = ( n1104 & n3987 ) | ( n1104 & n3988 ) | ( n3987 & n3988 ) ;
  assign n3990 = ( n1119 & n3987 ) | ( n1119 & n3988 ) | ( n3987 & n3988 ) ;
  assign n3991 = ( ~n1126 & n3987 ) | ( ~n1126 & n3988 ) | ( n3987 & n3988 ) ;
  assign n3992 = ( ~n1115 & n3990 ) | ( ~n1115 & n3991 ) | ( n3990 & n3991 ) ;
  assign n3993 = ( ~n975 & n3989 ) | ( ~n975 & n3992 ) | ( n3989 & n3992 ) ;
  assign n3994 = ( n1154 & n3989 ) | ( n1154 & n3992 ) | ( n3989 & n3992 ) ;
  assign n3995 = ( ~x409 & n3993 ) | ( ~x409 & n3994 ) | ( n3993 & n3994 ) ;
  assign n3996 = ( x281 & n3993 ) | ( x281 & n3994 ) | ( n3993 & n3994 ) ;
  assign n3997 = ( n656 & n3995 ) | ( n656 & n3996 ) | ( n3995 & n3996 ) ;
  assign n3998 = n3986 | n3997 ;
  assign n3999 = ~n3975 & n3998 ;
  assign n4000 = n3956 | n3999 ;
  assign n4001 = x252 & n1767 ;
  assign n4002 = x252 & ~n1771 ;
  assign n4003 = ( ~n1751 & n4001 ) | ( ~n1751 & n4002 ) | ( n4001 & n4002 ) ;
  assign n4004 = ( ~n1787 & n4001 ) | ( ~n1787 & n4002 ) | ( n4001 & n4002 ) ;
  assign n4005 = ( n1794 & n4001 ) | ( n1794 & n4002 ) | ( n4001 & n4002 ) ;
  assign n4006 = ( n1783 & n4004 ) | ( n1783 & n4005 ) | ( n4004 & n4005 ) ;
  assign n4007 = ( n1643 & n4003 ) | ( n1643 & n4006 ) | ( n4003 & n4006 ) ;
  assign n4008 = ( ~n1822 & n4003 ) | ( ~n1822 & n4006 ) | ( n4003 & n4006 ) ;
  assign n4009 = ( ~n1324 & n4007 ) | ( ~n1324 & n4008 ) | ( n4007 & n4008 ) ;
  assign n4010 = x124 & ~n1767 ;
  assign n4011 = x124 & n1771 ;
  assign n4012 = ( n1751 & n4010 ) | ( n1751 & n4011 ) | ( n4010 & n4011 ) ;
  assign n4013 = ( n1787 & n4010 ) | ( n1787 & n4011 ) | ( n4010 & n4011 ) ;
  assign n4014 = ( ~n1794 & n4010 ) | ( ~n1794 & n4011 ) | ( n4010 & n4011 ) ;
  assign n4015 = ( ~n1783 & n4013 ) | ( ~n1783 & n4014 ) | ( n4013 & n4014 ) ;
  assign n4016 = ( ~n1643 & n4012 ) | ( ~n1643 & n4015 ) | ( n4012 & n4015 ) ;
  assign n4017 = ( n1822 & n4012 ) | ( n1822 & n4015 ) | ( n4012 & n4015 ) ;
  assign n4018 = ( n1324 & n4016 ) | ( n1324 & n4017 ) | ( n4016 & n4017 ) ;
  assign n4019 = n4009 | n4018 ;
  assign n4020 = x508 & n991 ;
  assign n4021 = x508 & ~n995 ;
  assign n4022 = ( ~n1104 & n4020 ) | ( ~n1104 & n4021 ) | ( n4020 & n4021 ) ;
  assign n4023 = ( ~n1119 & n4020 ) | ( ~n1119 & n4021 ) | ( n4020 & n4021 ) ;
  assign n4024 = ( n1126 & n4020 ) | ( n1126 & n4021 ) | ( n4020 & n4021 ) ;
  assign n4025 = ( n1115 & n4023 ) | ( n1115 & n4024 ) | ( n4023 & n4024 ) ;
  assign n4026 = ( n975 & n4022 ) | ( n975 & n4025 ) | ( n4022 & n4025 ) ;
  assign n4027 = ( ~n1154 & n4022 ) | ( ~n1154 & n4025 ) | ( n4022 & n4025 ) ;
  assign n4028 = ( x409 & n4026 ) | ( x409 & n4027 ) | ( n4026 & n4027 ) ;
  assign n4029 = ( ~x281 & n4026 ) | ( ~x281 & n4027 ) | ( n4026 & n4027 ) ;
  assign n4030 = ( ~n656 & n4028 ) | ( ~n656 & n4029 ) | ( n4028 & n4029 ) ;
  assign n4031 = x380 & ~n991 ;
  assign n4032 = x380 & n995 ;
  assign n4033 = ( n1104 & n4031 ) | ( n1104 & n4032 ) | ( n4031 & n4032 ) ;
  assign n4034 = ( n1119 & n4031 ) | ( n1119 & n4032 ) | ( n4031 & n4032 ) ;
  assign n4035 = ( ~n1126 & n4031 ) | ( ~n1126 & n4032 ) | ( n4031 & n4032 ) ;
  assign n4036 = ( ~n1115 & n4034 ) | ( ~n1115 & n4035 ) | ( n4034 & n4035 ) ;
  assign n4037 = ( ~n975 & n4033 ) | ( ~n975 & n4036 ) | ( n4033 & n4036 ) ;
  assign n4038 = ( n1154 & n4033 ) | ( n1154 & n4036 ) | ( n4033 & n4036 ) ;
  assign n4039 = ( ~x409 & n4037 ) | ( ~x409 & n4038 ) | ( n4037 & n4038 ) ;
  assign n4040 = ( x281 & n4037 ) | ( x281 & n4038 ) | ( n4037 & n4038 ) ;
  assign n4041 = ( n656 & n4039 ) | ( n656 & n4040 ) | ( n4039 & n4040 ) ;
  assign n4042 = n4030 | n4041 ;
  assign n4043 = ~n4019 & n4042 ;
  assign n4044 = ~x255 & n1765 ;
  assign n4045 = ~n1759 & n4044 ;
  assign n4046 = x127 & ~n4045 ;
  assign n4047 = x255 | n1754 ;
  assign n4048 = ~x255 & n1752 ;
  assign n4049 = ( n1758 & n4047 ) | ( n1758 & ~n4048 ) | ( n4047 & ~n4048 ) ;
  assign n4050 = x127 & n4049 ;
  assign n4051 = ( n1751 & n4046 ) | ( n1751 & n4050 ) | ( n4046 & n4050 ) ;
  assign n4052 = ( n1787 & n4046 ) | ( n1787 & n4050 ) | ( n4046 & n4050 ) ;
  assign n4053 = ( ~n1794 & n4046 ) | ( ~n1794 & n4050 ) | ( n4046 & n4050 ) ;
  assign n4054 = ( ~n1783 & n4052 ) | ( ~n1783 & n4053 ) | ( n4052 & n4053 ) ;
  assign n4055 = ( ~n1643 & n4051 ) | ( ~n1643 & n4054 ) | ( n4051 & n4054 ) ;
  assign n4056 = ( n1822 & n4051 ) | ( n1822 & n4054 ) | ( n4051 & n4054 ) ;
  assign n4057 = ( n1324 & n4055 ) | ( n1324 & n4056 ) | ( n4055 & n4056 ) ;
  assign n4058 = ~x511 & n989 ;
  assign n4059 = ~n983 & n4058 ;
  assign n4060 = x383 & ~n4059 ;
  assign n4061 = x511 | n978 ;
  assign n4062 = ~x511 & n976 ;
  assign n4063 = ( n982 & n4061 ) | ( n982 & ~n4062 ) | ( n4061 & ~n4062 ) ;
  assign n4064 = x383 & n4063 ;
  assign n4065 = ( n1104 & n4060 ) | ( n1104 & n4064 ) | ( n4060 & n4064 ) ;
  assign n4066 = ( n1119 & n4060 ) | ( n1119 & n4064 ) | ( n4060 & n4064 ) ;
  assign n4067 = ( ~n1126 & n4060 ) | ( ~n1126 & n4064 ) | ( n4060 & n4064 ) ;
  assign n4068 = ( ~n1115 & n4066 ) | ( ~n1115 & n4067 ) | ( n4066 & n4067 ) ;
  assign n4069 = ( ~n975 & n4065 ) | ( ~n975 & n4068 ) | ( n4065 & n4068 ) ;
  assign n4070 = ( n1154 & n4065 ) | ( n1154 & n4068 ) | ( n4065 & n4068 ) ;
  assign n4071 = ( ~x409 & n4069 ) | ( ~x409 & n4070 ) | ( n4069 & n4070 ) ;
  assign n4072 = ( x281 & n4069 ) | ( x281 & n4070 ) | ( n4069 & n4070 ) ;
  assign n4073 = ( n656 & n4071 ) | ( n656 & n4072 ) | ( n4071 & n4072 ) ;
  assign n4074 = n4057 & ~n4073 ;
  assign n4075 = n4043 | n4074 ;
  assign n4076 = n4000 | n4075 ;
  assign n4077 = ~n3520 & n3539 ;
  assign n4078 = ( n3473 & ~n3496 ) | ( n3473 & n4077 ) | ( ~n3496 & n4077 ) ;
  assign n4079 = ~n3433 & n3452 ;
  assign n4080 = ~n3453 & n4079 ;
  assign n4081 = ( ~n3453 & n4078 ) | ( ~n3453 & n4080 ) | ( n4078 & n4080 ) ;
  assign n4082 = ( n3386 & ~n3409 ) | ( n3386 & n4081 ) | ( ~n3409 & n4081 ) ;
  assign n4083 = ~n4076 & n4082 ;
  assign n4084 = n4019 & ~n4042 ;
  assign n4085 = ( n3975 & ~n3998 ) | ( n3975 & n4084 ) | ( ~n3998 & n4084 ) ;
  assign n4086 = ~n3956 & n4085 ;
  assign n4087 = ~n4057 & n4073 ;
  assign n4088 = n4074 & ~n4087 ;
  assign n4089 = n3932 & ~n3955 ;
  assign n4090 = ( n4087 & ~n4088 ) | ( n4087 & n4089 ) | ( ~n4088 & n4089 ) ;
  assign n4091 = ( n4086 & ~n4088 ) | ( n4086 & n4090 ) | ( ~n4088 & n4090 ) ;
  assign n4092 = n4083 | n4091 ;
  assign n4093 = n4076 & ~n4091 ;
  assign n4094 = ( n3913 & n4092 ) | ( n3913 & ~n4093 ) | ( n4092 & ~n4093 ) ;
  assign n4095 = n3542 | n4076 ;
  assign n4096 = ( n4076 & ~n4082 ) | ( n4076 & n4095 ) | ( ~n4082 & n4095 ) ;
  assign n4097 = ~n4091 & n4096 ;
  assign n4098 = n3185 & ~n3365 ;
  assign n4099 = n3362 & ~n3904 ;
  assign n4100 = ~n3903 & n4099 ;
  assign n4101 = ~n3905 & n4100 ;
  assign n4102 = n3901 | n4101 ;
  assign n4103 = ~n3901 & n3907 ;
  assign n4104 = ( n4098 & ~n4102 ) | ( n4098 & n4103 ) | ( ~n4102 & n4103 ) ;
  assign n4105 = ~n3719 & n3726 ;
  assign n4106 = n3716 | n3717 ;
  assign n4107 = n4105 & ~n4106 ;
  assign n4108 = ( ~n3721 & n4104 ) | ( ~n3721 & n4107 ) | ( n4104 & n4107 ) ;
  assign n4109 = ( ~n4092 & n4097 ) | ( ~n4092 & n4108 ) | ( n4097 & n4108 ) ;
  assign n4110 = ~n3204 & n3227 ;
  assign n4111 = n3270 | n4110 ;
  assign n4112 = ~n3289 & n3312 ;
  assign n4113 = n3335 & ~n3354 ;
  assign n4114 = n4112 | n4113 ;
  assign n4115 = n4111 | n4114 ;
  assign n4116 = x231 & n1767 ;
  assign n4117 = x231 & ~n1771 ;
  assign n4118 = ( ~n1751 & n4116 ) | ( ~n1751 & n4117 ) | ( n4116 & n4117 ) ;
  assign n4119 = ( ~n1787 & n4116 ) | ( ~n1787 & n4117 ) | ( n4116 & n4117 ) ;
  assign n4120 = ( n1794 & n4116 ) | ( n1794 & n4117 ) | ( n4116 & n4117 ) ;
  assign n4121 = ( n1783 & n4119 ) | ( n1783 & n4120 ) | ( n4119 & n4120 ) ;
  assign n4122 = ( n1643 & n4118 ) | ( n1643 & n4121 ) | ( n4118 & n4121 ) ;
  assign n4123 = ( ~n1822 & n4118 ) | ( ~n1822 & n4121 ) | ( n4118 & n4121 ) ;
  assign n4124 = ( ~n1324 & n4122 ) | ( ~n1324 & n4123 ) | ( n4122 & n4123 ) ;
  assign n4125 = x103 & ~n1767 ;
  assign n4126 = x103 & n1771 ;
  assign n4127 = ( n1751 & n4125 ) | ( n1751 & n4126 ) | ( n4125 & n4126 ) ;
  assign n4128 = ( n1787 & n4125 ) | ( n1787 & n4126 ) | ( n4125 & n4126 ) ;
  assign n4129 = ( ~n1794 & n4125 ) | ( ~n1794 & n4126 ) | ( n4125 & n4126 ) ;
  assign n4130 = ( ~n1783 & n4128 ) | ( ~n1783 & n4129 ) | ( n4128 & n4129 ) ;
  assign n4131 = ( ~n1643 & n4127 ) | ( ~n1643 & n4130 ) | ( n4127 & n4130 ) ;
  assign n4132 = ( n1822 & n4127 ) | ( n1822 & n4130 ) | ( n4127 & n4130 ) ;
  assign n4133 = ( n1324 & n4131 ) | ( n1324 & n4132 ) | ( n4131 & n4132 ) ;
  assign n4134 = n4124 | n4133 ;
  assign n4135 = x487 & n991 ;
  assign n4136 = x487 & ~n995 ;
  assign n4137 = ( ~n1104 & n4135 ) | ( ~n1104 & n4136 ) | ( n4135 & n4136 ) ;
  assign n4138 = ( ~n1119 & n4135 ) | ( ~n1119 & n4136 ) | ( n4135 & n4136 ) ;
  assign n4139 = ( n1126 & n4135 ) | ( n1126 & n4136 ) | ( n4135 & n4136 ) ;
  assign n4140 = ( n1115 & n4138 ) | ( n1115 & n4139 ) | ( n4138 & n4139 ) ;
  assign n4141 = ( n975 & n4137 ) | ( n975 & n4140 ) | ( n4137 & n4140 ) ;
  assign n4142 = ( ~n1154 & n4137 ) | ( ~n1154 & n4140 ) | ( n4137 & n4140 ) ;
  assign n4143 = ( x409 & n4141 ) | ( x409 & n4142 ) | ( n4141 & n4142 ) ;
  assign n4144 = ( ~x281 & n4141 ) | ( ~x281 & n4142 ) | ( n4141 & n4142 ) ;
  assign n4145 = ( ~n656 & n4143 ) | ( ~n656 & n4144 ) | ( n4143 & n4144 ) ;
  assign n4146 = x359 & ~n991 ;
  assign n4147 = x359 & n995 ;
  assign n4148 = ( n1104 & n4146 ) | ( n1104 & n4147 ) | ( n4146 & n4147 ) ;
  assign n4149 = ( n1119 & n4146 ) | ( n1119 & n4147 ) | ( n4146 & n4147 ) ;
  assign n4150 = ( ~n1126 & n4146 ) | ( ~n1126 & n4147 ) | ( n4146 & n4147 ) ;
  assign n4151 = ( ~n1115 & n4149 ) | ( ~n1115 & n4150 ) | ( n4149 & n4150 ) ;
  assign n4152 = ( ~n975 & n4148 ) | ( ~n975 & n4151 ) | ( n4148 & n4151 ) ;
  assign n4153 = ( n1154 & n4148 ) | ( n1154 & n4151 ) | ( n4148 & n4151 ) ;
  assign n4154 = ( ~x409 & n4152 ) | ( ~x409 & n4153 ) | ( n4152 & n4153 ) ;
  assign n4155 = ( x281 & n4152 ) | ( x281 & n4153 ) | ( n4152 & n4153 ) ;
  assign n4156 = ( n656 & n4154 ) | ( n656 & n4155 ) | ( n4154 & n4155 ) ;
  assign n4157 = n4145 | n4156 ;
  assign n4158 = n4134 & ~n4157 ;
  assign n4159 = ~n4115 & n4158 ;
  assign n4160 = x215 & n1767 ;
  assign n4161 = x215 & ~n1771 ;
  assign n4162 = ( ~n1751 & n4160 ) | ( ~n1751 & n4161 ) | ( n4160 & n4161 ) ;
  assign n4163 = ( ~n1787 & n4160 ) | ( ~n1787 & n4161 ) | ( n4160 & n4161 ) ;
  assign n4164 = ( n1794 & n4160 ) | ( n1794 & n4161 ) | ( n4160 & n4161 ) ;
  assign n4165 = ( n1783 & n4163 ) | ( n1783 & n4164 ) | ( n4163 & n4164 ) ;
  assign n4166 = ( n1643 & n4162 ) | ( n1643 & n4165 ) | ( n4162 & n4165 ) ;
  assign n4167 = ( ~n1822 & n4162 ) | ( ~n1822 & n4165 ) | ( n4162 & n4165 ) ;
  assign n4168 = ( ~n1324 & n4166 ) | ( ~n1324 & n4167 ) | ( n4166 & n4167 ) ;
  assign n4169 = x87 & ~n1767 ;
  assign n4170 = x87 & n1771 ;
  assign n4171 = ( n1751 & n4169 ) | ( n1751 & n4170 ) | ( n4169 & n4170 ) ;
  assign n4172 = ( n1787 & n4169 ) | ( n1787 & n4170 ) | ( n4169 & n4170 ) ;
  assign n4173 = ( ~n1794 & n4169 ) | ( ~n1794 & n4170 ) | ( n4169 & n4170 ) ;
  assign n4174 = ( ~n1783 & n4172 ) | ( ~n1783 & n4173 ) | ( n4172 & n4173 ) ;
  assign n4175 = ( ~n1643 & n4171 ) | ( ~n1643 & n4174 ) | ( n4171 & n4174 ) ;
  assign n4176 = ( n1822 & n4171 ) | ( n1822 & n4174 ) | ( n4171 & n4174 ) ;
  assign n4177 = ( n1324 & n4175 ) | ( n1324 & n4176 ) | ( n4175 & n4176 ) ;
  assign n4178 = n4168 | n4177 ;
  assign n4179 = x471 & n991 ;
  assign n4180 = x471 & ~n995 ;
  assign n4181 = ( ~n1104 & n4179 ) | ( ~n1104 & n4180 ) | ( n4179 & n4180 ) ;
  assign n4182 = ( ~n1119 & n4179 ) | ( ~n1119 & n4180 ) | ( n4179 & n4180 ) ;
  assign n4183 = ( n1126 & n4179 ) | ( n1126 & n4180 ) | ( n4179 & n4180 ) ;
  assign n4184 = ( n1115 & n4182 ) | ( n1115 & n4183 ) | ( n4182 & n4183 ) ;
  assign n4185 = ( n975 & n4181 ) | ( n975 & n4184 ) | ( n4181 & n4184 ) ;
  assign n4186 = ( ~n1154 & n4181 ) | ( ~n1154 & n4184 ) | ( n4181 & n4184 ) ;
  assign n4187 = ( x409 & n4185 ) | ( x409 & n4186 ) | ( n4185 & n4186 ) ;
  assign n4188 = ( ~x281 & n4185 ) | ( ~x281 & n4186 ) | ( n4185 & n4186 ) ;
  assign n4189 = ( ~n656 & n4187 ) | ( ~n656 & n4188 ) | ( n4187 & n4188 ) ;
  assign n4190 = x343 & ~n991 ;
  assign n4191 = x343 & n995 ;
  assign n4192 = ( n1104 & n4190 ) | ( n1104 & n4191 ) | ( n4190 & n4191 ) ;
  assign n4193 = ( n1119 & n4190 ) | ( n1119 & n4191 ) | ( n4190 & n4191 ) ;
  assign n4194 = ( ~n1126 & n4190 ) | ( ~n1126 & n4191 ) | ( n4190 & n4191 ) ;
  assign n4195 = ( ~n1115 & n4193 ) | ( ~n1115 & n4194 ) | ( n4193 & n4194 ) ;
  assign n4196 = ( ~n975 & n4192 ) | ( ~n975 & n4195 ) | ( n4192 & n4195 ) ;
  assign n4197 = ( n1154 & n4192 ) | ( n1154 & n4195 ) | ( n4192 & n4195 ) ;
  assign n4198 = ( ~x409 & n4196 ) | ( ~x409 & n4197 ) | ( n4196 & n4197 ) ;
  assign n4199 = ( x281 & n4196 ) | ( x281 & n4197 ) | ( n4196 & n4197 ) ;
  assign n4200 = ( n656 & n4198 ) | ( n656 & n4199 ) | ( n4198 & n4199 ) ;
  assign n4201 = n4189 | n4200 ;
  assign n4202 = ~n4178 & n4201 ;
  assign n4203 = x470 & n991 ;
  assign n4204 = x470 & ~n995 ;
  assign n4205 = ( ~n1104 & n4203 ) | ( ~n1104 & n4204 ) | ( n4203 & n4204 ) ;
  assign n4206 = ( ~n1119 & n4203 ) | ( ~n1119 & n4204 ) | ( n4203 & n4204 ) ;
  assign n4207 = ( n1126 & n4203 ) | ( n1126 & n4204 ) | ( n4203 & n4204 ) ;
  assign n4208 = ( n1115 & n4206 ) | ( n1115 & n4207 ) | ( n4206 & n4207 ) ;
  assign n4209 = ( n975 & n4205 ) | ( n975 & n4208 ) | ( n4205 & n4208 ) ;
  assign n4210 = ( ~n1154 & n4205 ) | ( ~n1154 & n4208 ) | ( n4205 & n4208 ) ;
  assign n4211 = ( x409 & n4209 ) | ( x409 & n4210 ) | ( n4209 & n4210 ) ;
  assign n4212 = ( ~x281 & n4209 ) | ( ~x281 & n4210 ) | ( n4209 & n4210 ) ;
  assign n4213 = ( ~n656 & n4211 ) | ( ~n656 & n4212 ) | ( n4211 & n4212 ) ;
  assign n4214 = x342 & ~n991 ;
  assign n4215 = x342 & n995 ;
  assign n4216 = ( n1104 & n4214 ) | ( n1104 & n4215 ) | ( n4214 & n4215 ) ;
  assign n4217 = ( n1119 & n4214 ) | ( n1119 & n4215 ) | ( n4214 & n4215 ) ;
  assign n4218 = ( ~n1126 & n4214 ) | ( ~n1126 & n4215 ) | ( n4214 & n4215 ) ;
  assign n4219 = ( ~n1115 & n4217 ) | ( ~n1115 & n4218 ) | ( n4217 & n4218 ) ;
  assign n4220 = ( ~n975 & n4216 ) | ( ~n975 & n4219 ) | ( n4216 & n4219 ) ;
  assign n4221 = ( n1154 & n4216 ) | ( n1154 & n4219 ) | ( n4216 & n4219 ) ;
  assign n4222 = ( ~x409 & n4220 ) | ( ~x409 & n4221 ) | ( n4220 & n4221 ) ;
  assign n4223 = ( x281 & n4220 ) | ( x281 & n4221 ) | ( n4220 & n4221 ) ;
  assign n4224 = ( n656 & n4222 ) | ( n656 & n4223 ) | ( n4222 & n4223 ) ;
  assign n4225 = n4213 | n4224 ;
  assign n4226 = x214 & n1767 ;
  assign n4227 = x214 & ~n1771 ;
  assign n4228 = ( ~n1751 & n4226 ) | ( ~n1751 & n4227 ) | ( n4226 & n4227 ) ;
  assign n4229 = ( ~n1787 & n4226 ) | ( ~n1787 & n4227 ) | ( n4226 & n4227 ) ;
  assign n4230 = ( n1794 & n4226 ) | ( n1794 & n4227 ) | ( n4226 & n4227 ) ;
  assign n4231 = ( n1783 & n4229 ) | ( n1783 & n4230 ) | ( n4229 & n4230 ) ;
  assign n4232 = ( n1643 & n4228 ) | ( n1643 & n4231 ) | ( n4228 & n4231 ) ;
  assign n4233 = ( ~n1822 & n4228 ) | ( ~n1822 & n4231 ) | ( n4228 & n4231 ) ;
  assign n4234 = ( ~n1324 & n4232 ) | ( ~n1324 & n4233 ) | ( n4232 & n4233 ) ;
  assign n4235 = x86 & ~n1767 ;
  assign n4236 = x86 & n1771 ;
  assign n4237 = ( n1751 & n4235 ) | ( n1751 & n4236 ) | ( n4235 & n4236 ) ;
  assign n4238 = ( n1787 & n4235 ) | ( n1787 & n4236 ) | ( n4235 & n4236 ) ;
  assign n4239 = ( ~n1794 & n4235 ) | ( ~n1794 & n4236 ) | ( n4235 & n4236 ) ;
  assign n4240 = ( ~n1783 & n4238 ) | ( ~n1783 & n4239 ) | ( n4238 & n4239 ) ;
  assign n4241 = ( ~n1643 & n4237 ) | ( ~n1643 & n4240 ) | ( n4237 & n4240 ) ;
  assign n4242 = ( n1822 & n4237 ) | ( n1822 & n4240 ) | ( n4237 & n4240 ) ;
  assign n4243 = ( n1324 & n4241 ) | ( n1324 & n4242 ) | ( n4241 & n4242 ) ;
  assign n4244 = n4234 | n4243 ;
  assign n4245 = n4225 & ~n4244 ;
  assign n4246 = n4202 | n4245 ;
  assign n4247 = x213 & n1767 ;
  assign n4248 = x213 & ~n1771 ;
  assign n4249 = ( ~n1751 & n4247 ) | ( ~n1751 & n4248 ) | ( n4247 & n4248 ) ;
  assign n4250 = ( ~n1787 & n4247 ) | ( ~n1787 & n4248 ) | ( n4247 & n4248 ) ;
  assign n4251 = ( n1794 & n4247 ) | ( n1794 & n4248 ) | ( n4247 & n4248 ) ;
  assign n4252 = ( n1783 & n4250 ) | ( n1783 & n4251 ) | ( n4250 & n4251 ) ;
  assign n4253 = ( n1643 & n4249 ) | ( n1643 & n4252 ) | ( n4249 & n4252 ) ;
  assign n4254 = ( ~n1822 & n4249 ) | ( ~n1822 & n4252 ) | ( n4249 & n4252 ) ;
  assign n4255 = ( ~n1324 & n4253 ) | ( ~n1324 & n4254 ) | ( n4253 & n4254 ) ;
  assign n4256 = x85 & ~n1767 ;
  assign n4257 = x85 & n1771 ;
  assign n4258 = ( n1751 & n4256 ) | ( n1751 & n4257 ) | ( n4256 & n4257 ) ;
  assign n4259 = ( n1787 & n4256 ) | ( n1787 & n4257 ) | ( n4256 & n4257 ) ;
  assign n4260 = ( ~n1794 & n4256 ) | ( ~n1794 & n4257 ) | ( n4256 & n4257 ) ;
  assign n4261 = ( ~n1783 & n4259 ) | ( ~n1783 & n4260 ) | ( n4259 & n4260 ) ;
  assign n4262 = ( ~n1643 & n4258 ) | ( ~n1643 & n4261 ) | ( n4258 & n4261 ) ;
  assign n4263 = ( n1822 & n4258 ) | ( n1822 & n4261 ) | ( n4258 & n4261 ) ;
  assign n4264 = ( n1324 & n4262 ) | ( n1324 & n4263 ) | ( n4262 & n4263 ) ;
  assign n4265 = n4255 | n4264 ;
  assign n4266 = x469 & n991 ;
  assign n4267 = x469 & ~n995 ;
  assign n4268 = ( ~n1104 & n4266 ) | ( ~n1104 & n4267 ) | ( n4266 & n4267 ) ;
  assign n4269 = ( ~n1119 & n4266 ) | ( ~n1119 & n4267 ) | ( n4266 & n4267 ) ;
  assign n4270 = ( n1126 & n4266 ) | ( n1126 & n4267 ) | ( n4266 & n4267 ) ;
  assign n4271 = ( n1115 & n4269 ) | ( n1115 & n4270 ) | ( n4269 & n4270 ) ;
  assign n4272 = ( n975 & n4268 ) | ( n975 & n4271 ) | ( n4268 & n4271 ) ;
  assign n4273 = ( ~n1154 & n4268 ) | ( ~n1154 & n4271 ) | ( n4268 & n4271 ) ;
  assign n4274 = ( x409 & n4272 ) | ( x409 & n4273 ) | ( n4272 & n4273 ) ;
  assign n4275 = ( ~x281 & n4272 ) | ( ~x281 & n4273 ) | ( n4272 & n4273 ) ;
  assign n4276 = ( ~n656 & n4274 ) | ( ~n656 & n4275 ) | ( n4274 & n4275 ) ;
  assign n4277 = x341 & ~n991 ;
  assign n4278 = x341 & n995 ;
  assign n4279 = ( n1104 & n4277 ) | ( n1104 & n4278 ) | ( n4277 & n4278 ) ;
  assign n4280 = ( n1119 & n4277 ) | ( n1119 & n4278 ) | ( n4277 & n4278 ) ;
  assign n4281 = ( ~n1126 & n4277 ) | ( ~n1126 & n4278 ) | ( n4277 & n4278 ) ;
  assign n4282 = ( ~n1115 & n4280 ) | ( ~n1115 & n4281 ) | ( n4280 & n4281 ) ;
  assign n4283 = ( ~n975 & n4279 ) | ( ~n975 & n4282 ) | ( n4279 & n4282 ) ;
  assign n4284 = ( n1154 & n4279 ) | ( n1154 & n4282 ) | ( n4279 & n4282 ) ;
  assign n4285 = ( ~x409 & n4283 ) | ( ~x409 & n4284 ) | ( n4283 & n4284 ) ;
  assign n4286 = ( x281 & n4283 ) | ( x281 & n4284 ) | ( n4283 & n4284 ) ;
  assign n4287 = ( n656 & n4285 ) | ( n656 & n4286 ) | ( n4285 & n4286 ) ;
  assign n4288 = n4276 | n4287 ;
  assign n4289 = ~n4265 & n4288 ;
  assign n4290 = x212 & n1767 ;
  assign n4291 = x212 & ~n1771 ;
  assign n4292 = ( ~n1751 & n4290 ) | ( ~n1751 & n4291 ) | ( n4290 & n4291 ) ;
  assign n4293 = ( ~n1787 & n4290 ) | ( ~n1787 & n4291 ) | ( n4290 & n4291 ) ;
  assign n4294 = ( n1794 & n4290 ) | ( n1794 & n4291 ) | ( n4290 & n4291 ) ;
  assign n4295 = ( n1783 & n4293 ) | ( n1783 & n4294 ) | ( n4293 & n4294 ) ;
  assign n4296 = ( n1643 & n4292 ) | ( n1643 & n4295 ) | ( n4292 & n4295 ) ;
  assign n4297 = ( ~n1822 & n4292 ) | ( ~n1822 & n4295 ) | ( n4292 & n4295 ) ;
  assign n4298 = ( ~n1324 & n4296 ) | ( ~n1324 & n4297 ) | ( n4296 & n4297 ) ;
  assign n4299 = x84 & ~n1767 ;
  assign n4300 = x84 & n1771 ;
  assign n4301 = ( n1751 & n4299 ) | ( n1751 & n4300 ) | ( n4299 & n4300 ) ;
  assign n4302 = ( n1787 & n4299 ) | ( n1787 & n4300 ) | ( n4299 & n4300 ) ;
  assign n4303 = ( ~n1794 & n4299 ) | ( ~n1794 & n4300 ) | ( n4299 & n4300 ) ;
  assign n4304 = ( ~n1783 & n4302 ) | ( ~n1783 & n4303 ) | ( n4302 & n4303 ) ;
  assign n4305 = ( ~n1643 & n4301 ) | ( ~n1643 & n4304 ) | ( n4301 & n4304 ) ;
  assign n4306 = ( n1822 & n4301 ) | ( n1822 & n4304 ) | ( n4301 & n4304 ) ;
  assign n4307 = ( n1324 & n4305 ) | ( n1324 & n4306 ) | ( n4305 & n4306 ) ;
  assign n4308 = n4298 | n4307 ;
  assign n4309 = x468 & n991 ;
  assign n4310 = x468 & ~n995 ;
  assign n4311 = ( ~n1104 & n4309 ) | ( ~n1104 & n4310 ) | ( n4309 & n4310 ) ;
  assign n4312 = ( ~n1119 & n4309 ) | ( ~n1119 & n4310 ) | ( n4309 & n4310 ) ;
  assign n4313 = ( n1126 & n4309 ) | ( n1126 & n4310 ) | ( n4309 & n4310 ) ;
  assign n4314 = ( n1115 & n4312 ) | ( n1115 & n4313 ) | ( n4312 & n4313 ) ;
  assign n4315 = ( n975 & n4311 ) | ( n975 & n4314 ) | ( n4311 & n4314 ) ;
  assign n4316 = ( ~n1154 & n4311 ) | ( ~n1154 & n4314 ) | ( n4311 & n4314 ) ;
  assign n4317 = ( x409 & n4315 ) | ( x409 & n4316 ) | ( n4315 & n4316 ) ;
  assign n4318 = ( ~x281 & n4315 ) | ( ~x281 & n4316 ) | ( n4315 & n4316 ) ;
  assign n4319 = ( ~n656 & n4317 ) | ( ~n656 & n4318 ) | ( n4317 & n4318 ) ;
  assign n4320 = x340 & ~n991 ;
  assign n4321 = x340 & n995 ;
  assign n4322 = ( n1104 & n4320 ) | ( n1104 & n4321 ) | ( n4320 & n4321 ) ;
  assign n4323 = ( n1119 & n4320 ) | ( n1119 & n4321 ) | ( n4320 & n4321 ) ;
  assign n4324 = ( ~n1126 & n4320 ) | ( ~n1126 & n4321 ) | ( n4320 & n4321 ) ;
  assign n4325 = ( ~n1115 & n4323 ) | ( ~n1115 & n4324 ) | ( n4323 & n4324 ) ;
  assign n4326 = ( ~n975 & n4322 ) | ( ~n975 & n4325 ) | ( n4322 & n4325 ) ;
  assign n4327 = ( n1154 & n4322 ) | ( n1154 & n4325 ) | ( n4322 & n4325 ) ;
  assign n4328 = ( ~x409 & n4326 ) | ( ~x409 & n4327 ) | ( n4326 & n4327 ) ;
  assign n4329 = ( x281 & n4326 ) | ( x281 & n4327 ) | ( n4326 & n4327 ) ;
  assign n4330 = ( n656 & n4328 ) | ( n656 & n4329 ) | ( n4328 & n4329 ) ;
  assign n4331 = n4319 | n4330 ;
  assign n4332 = ~n4308 & n4331 ;
  assign n4333 = n4289 | n4332 ;
  assign n4334 = n4246 | n4333 ;
  assign n4335 = x211 & n1767 ;
  assign n4336 = x211 & ~n1771 ;
  assign n4337 = ( ~n1751 & n4335 ) | ( ~n1751 & n4336 ) | ( n4335 & n4336 ) ;
  assign n4338 = ( ~n1787 & n4335 ) | ( ~n1787 & n4336 ) | ( n4335 & n4336 ) ;
  assign n4339 = ( n1794 & n4335 ) | ( n1794 & n4336 ) | ( n4335 & n4336 ) ;
  assign n4340 = ( n1783 & n4338 ) | ( n1783 & n4339 ) | ( n4338 & n4339 ) ;
  assign n4341 = ( n1643 & n4337 ) | ( n1643 & n4340 ) | ( n4337 & n4340 ) ;
  assign n4342 = ( ~n1822 & n4337 ) | ( ~n1822 & n4340 ) | ( n4337 & n4340 ) ;
  assign n4343 = ( ~n1324 & n4341 ) | ( ~n1324 & n4342 ) | ( n4341 & n4342 ) ;
  assign n4344 = x83 & ~n1767 ;
  assign n4345 = x83 & n1771 ;
  assign n4346 = ( n1751 & n4344 ) | ( n1751 & n4345 ) | ( n4344 & n4345 ) ;
  assign n4347 = ( n1787 & n4344 ) | ( n1787 & n4345 ) | ( n4344 & n4345 ) ;
  assign n4348 = ( ~n1794 & n4344 ) | ( ~n1794 & n4345 ) | ( n4344 & n4345 ) ;
  assign n4349 = ( ~n1783 & n4347 ) | ( ~n1783 & n4348 ) | ( n4347 & n4348 ) ;
  assign n4350 = ( ~n1643 & n4346 ) | ( ~n1643 & n4349 ) | ( n4346 & n4349 ) ;
  assign n4351 = ( n1822 & n4346 ) | ( n1822 & n4349 ) | ( n4346 & n4349 ) ;
  assign n4352 = ( n1324 & n4350 ) | ( n1324 & n4351 ) | ( n4350 & n4351 ) ;
  assign n4353 = n4343 | n4352 ;
  assign n4354 = x467 & n991 ;
  assign n4355 = x467 & ~n995 ;
  assign n4356 = ( ~n1104 & n4354 ) | ( ~n1104 & n4355 ) | ( n4354 & n4355 ) ;
  assign n4357 = ( ~n1119 & n4354 ) | ( ~n1119 & n4355 ) | ( n4354 & n4355 ) ;
  assign n4358 = ( n1126 & n4354 ) | ( n1126 & n4355 ) | ( n4354 & n4355 ) ;
  assign n4359 = ( n1115 & n4357 ) | ( n1115 & n4358 ) | ( n4357 & n4358 ) ;
  assign n4360 = ( n975 & n4356 ) | ( n975 & n4359 ) | ( n4356 & n4359 ) ;
  assign n4361 = ( ~n1154 & n4356 ) | ( ~n1154 & n4359 ) | ( n4356 & n4359 ) ;
  assign n4362 = ( x409 & n4360 ) | ( x409 & n4361 ) | ( n4360 & n4361 ) ;
  assign n4363 = ( ~x281 & n4360 ) | ( ~x281 & n4361 ) | ( n4360 & n4361 ) ;
  assign n4364 = ( ~n656 & n4362 ) | ( ~n656 & n4363 ) | ( n4362 & n4363 ) ;
  assign n4365 = x339 & ~n991 ;
  assign n4366 = x339 & n995 ;
  assign n4367 = ( n1104 & n4365 ) | ( n1104 & n4366 ) | ( n4365 & n4366 ) ;
  assign n4368 = ( n1119 & n4365 ) | ( n1119 & n4366 ) | ( n4365 & n4366 ) ;
  assign n4369 = ( ~n1126 & n4365 ) | ( ~n1126 & n4366 ) | ( n4365 & n4366 ) ;
  assign n4370 = ( ~n1115 & n4368 ) | ( ~n1115 & n4369 ) | ( n4368 & n4369 ) ;
  assign n4371 = ( ~n975 & n4367 ) | ( ~n975 & n4370 ) | ( n4367 & n4370 ) ;
  assign n4372 = ( n1154 & n4367 ) | ( n1154 & n4370 ) | ( n4367 & n4370 ) ;
  assign n4373 = ( ~x409 & n4371 ) | ( ~x409 & n4372 ) | ( n4371 & n4372 ) ;
  assign n4374 = ( x281 & n4371 ) | ( x281 & n4372 ) | ( n4371 & n4372 ) ;
  assign n4375 = ( n656 & n4373 ) | ( n656 & n4374 ) | ( n4373 & n4374 ) ;
  assign n4376 = n4364 | n4375 ;
  assign n4377 = ~n4353 & n4376 ;
  assign n4378 = x466 & n991 ;
  assign n4379 = x466 & ~n995 ;
  assign n4380 = ( ~n1104 & n4378 ) | ( ~n1104 & n4379 ) | ( n4378 & n4379 ) ;
  assign n4381 = ( ~n1119 & n4378 ) | ( ~n1119 & n4379 ) | ( n4378 & n4379 ) ;
  assign n4382 = ( n1126 & n4378 ) | ( n1126 & n4379 ) | ( n4378 & n4379 ) ;
  assign n4383 = ( n1115 & n4381 ) | ( n1115 & n4382 ) | ( n4381 & n4382 ) ;
  assign n4384 = ( n975 & n4380 ) | ( n975 & n4383 ) | ( n4380 & n4383 ) ;
  assign n4385 = ( ~n1154 & n4380 ) | ( ~n1154 & n4383 ) | ( n4380 & n4383 ) ;
  assign n4386 = ( x409 & n4384 ) | ( x409 & n4385 ) | ( n4384 & n4385 ) ;
  assign n4387 = ( ~x281 & n4384 ) | ( ~x281 & n4385 ) | ( n4384 & n4385 ) ;
  assign n4388 = ( ~n656 & n4386 ) | ( ~n656 & n4387 ) | ( n4386 & n4387 ) ;
  assign n4389 = x338 & ~n991 ;
  assign n4390 = x338 & n995 ;
  assign n4391 = ( n1104 & n4389 ) | ( n1104 & n4390 ) | ( n4389 & n4390 ) ;
  assign n4392 = ( n1119 & n4389 ) | ( n1119 & n4390 ) | ( n4389 & n4390 ) ;
  assign n4393 = ( ~n1126 & n4389 ) | ( ~n1126 & n4390 ) | ( n4389 & n4390 ) ;
  assign n4394 = ( ~n1115 & n4392 ) | ( ~n1115 & n4393 ) | ( n4392 & n4393 ) ;
  assign n4395 = ( ~n975 & n4391 ) | ( ~n975 & n4394 ) | ( n4391 & n4394 ) ;
  assign n4396 = ( n1154 & n4391 ) | ( n1154 & n4394 ) | ( n4391 & n4394 ) ;
  assign n4397 = ( ~x409 & n4395 ) | ( ~x409 & n4396 ) | ( n4395 & n4396 ) ;
  assign n4398 = ( x281 & n4395 ) | ( x281 & n4396 ) | ( n4395 & n4396 ) ;
  assign n4399 = ( n656 & n4397 ) | ( n656 & n4398 ) | ( n4397 & n4398 ) ;
  assign n4400 = n4388 | n4399 ;
  assign n4401 = x210 & n1767 ;
  assign n4402 = x210 & ~n1771 ;
  assign n4403 = ( ~n1751 & n4401 ) | ( ~n1751 & n4402 ) | ( n4401 & n4402 ) ;
  assign n4404 = ( ~n1787 & n4401 ) | ( ~n1787 & n4402 ) | ( n4401 & n4402 ) ;
  assign n4405 = ( n1794 & n4401 ) | ( n1794 & n4402 ) | ( n4401 & n4402 ) ;
  assign n4406 = ( n1783 & n4404 ) | ( n1783 & n4405 ) | ( n4404 & n4405 ) ;
  assign n4407 = ( n1643 & n4403 ) | ( n1643 & n4406 ) | ( n4403 & n4406 ) ;
  assign n4408 = ( ~n1822 & n4403 ) | ( ~n1822 & n4406 ) | ( n4403 & n4406 ) ;
  assign n4409 = ( ~n1324 & n4407 ) | ( ~n1324 & n4408 ) | ( n4407 & n4408 ) ;
  assign n4410 = x82 & ~n1767 ;
  assign n4411 = x82 & n1771 ;
  assign n4412 = ( n1751 & n4410 ) | ( n1751 & n4411 ) | ( n4410 & n4411 ) ;
  assign n4413 = ( n1787 & n4410 ) | ( n1787 & n4411 ) | ( n4410 & n4411 ) ;
  assign n4414 = ( ~n1794 & n4410 ) | ( ~n1794 & n4411 ) | ( n4410 & n4411 ) ;
  assign n4415 = ( ~n1783 & n4413 ) | ( ~n1783 & n4414 ) | ( n4413 & n4414 ) ;
  assign n4416 = ( ~n1643 & n4412 ) | ( ~n1643 & n4415 ) | ( n4412 & n4415 ) ;
  assign n4417 = ( n1822 & n4412 ) | ( n1822 & n4415 ) | ( n4412 & n4415 ) ;
  assign n4418 = ( n1324 & n4416 ) | ( n1324 & n4417 ) | ( n4416 & n4417 ) ;
  assign n4419 = n4409 | n4418 ;
  assign n4420 = n4400 & ~n4419 ;
  assign n4421 = n4377 | n4420 ;
  assign n4422 = x464 & n991 ;
  assign n4423 = x464 & ~n995 ;
  assign n4424 = ( ~n1104 & n4422 ) | ( ~n1104 & n4423 ) | ( n4422 & n4423 ) ;
  assign n4425 = ( ~n1119 & n4422 ) | ( ~n1119 & n4423 ) | ( n4422 & n4423 ) ;
  assign n4426 = ( n1126 & n4422 ) | ( n1126 & n4423 ) | ( n4422 & n4423 ) ;
  assign n4427 = ( n1115 & n4425 ) | ( n1115 & n4426 ) | ( n4425 & n4426 ) ;
  assign n4428 = ( n975 & n4424 ) | ( n975 & n4427 ) | ( n4424 & n4427 ) ;
  assign n4429 = ( ~n1154 & n4424 ) | ( ~n1154 & n4427 ) | ( n4424 & n4427 ) ;
  assign n4430 = ( x409 & n4428 ) | ( x409 & n4429 ) | ( n4428 & n4429 ) ;
  assign n4431 = ( ~x281 & n4428 ) | ( ~x281 & n4429 ) | ( n4428 & n4429 ) ;
  assign n4432 = ( ~n656 & n4430 ) | ( ~n656 & n4431 ) | ( n4430 & n4431 ) ;
  assign n4433 = x336 & ~n991 ;
  assign n4434 = x336 & n995 ;
  assign n4435 = ( n1104 & n4433 ) | ( n1104 & n4434 ) | ( n4433 & n4434 ) ;
  assign n4436 = ( n1119 & n4433 ) | ( n1119 & n4434 ) | ( n4433 & n4434 ) ;
  assign n4437 = ( ~n1126 & n4433 ) | ( ~n1126 & n4434 ) | ( n4433 & n4434 ) ;
  assign n4438 = ( ~n1115 & n4436 ) | ( ~n1115 & n4437 ) | ( n4436 & n4437 ) ;
  assign n4439 = ( ~n975 & n4435 ) | ( ~n975 & n4438 ) | ( n4435 & n4438 ) ;
  assign n4440 = ( n1154 & n4435 ) | ( n1154 & n4438 ) | ( n4435 & n4438 ) ;
  assign n4441 = ( ~x409 & n4439 ) | ( ~x409 & n4440 ) | ( n4439 & n4440 ) ;
  assign n4442 = ( x281 & n4439 ) | ( x281 & n4440 ) | ( n4439 & n4440 ) ;
  assign n4443 = ( n656 & n4441 ) | ( n656 & n4442 ) | ( n4441 & n4442 ) ;
  assign n4444 = n4432 | n4443 ;
  assign n4445 = x208 & n1767 ;
  assign n4446 = x208 & ~n1771 ;
  assign n4447 = ( ~n1751 & n4445 ) | ( ~n1751 & n4446 ) | ( n4445 & n4446 ) ;
  assign n4448 = ( ~n1787 & n4445 ) | ( ~n1787 & n4446 ) | ( n4445 & n4446 ) ;
  assign n4449 = ( n1794 & n4445 ) | ( n1794 & n4446 ) | ( n4445 & n4446 ) ;
  assign n4450 = ( n1783 & n4448 ) | ( n1783 & n4449 ) | ( n4448 & n4449 ) ;
  assign n4451 = ( n1643 & n4447 ) | ( n1643 & n4450 ) | ( n4447 & n4450 ) ;
  assign n4452 = ( ~n1822 & n4447 ) | ( ~n1822 & n4450 ) | ( n4447 & n4450 ) ;
  assign n4453 = ( ~n1324 & n4451 ) | ( ~n1324 & n4452 ) | ( n4451 & n4452 ) ;
  assign n4454 = x80 & ~n1767 ;
  assign n4455 = x80 & n1771 ;
  assign n4456 = ( n1751 & n4454 ) | ( n1751 & n4455 ) | ( n4454 & n4455 ) ;
  assign n4457 = ( n1787 & n4454 ) | ( n1787 & n4455 ) | ( n4454 & n4455 ) ;
  assign n4458 = ( ~n1794 & n4454 ) | ( ~n1794 & n4455 ) | ( n4454 & n4455 ) ;
  assign n4459 = ( ~n1783 & n4457 ) | ( ~n1783 & n4458 ) | ( n4457 & n4458 ) ;
  assign n4460 = ( ~n1643 & n4456 ) | ( ~n1643 & n4459 ) | ( n4456 & n4459 ) ;
  assign n4461 = ( n1822 & n4456 ) | ( n1822 & n4459 ) | ( n4456 & n4459 ) ;
  assign n4462 = ( n1324 & n4460 ) | ( n1324 & n4461 ) | ( n4460 & n4461 ) ;
  assign n4463 = n4453 | n4462 ;
  assign n4464 = n4444 & ~n4463 ;
  assign n4465 = n4421 | n4464 ;
  assign n4466 = n4334 | n4465 ;
  assign n4467 = x209 & n1767 ;
  assign n4468 = x209 & ~n1771 ;
  assign n4469 = ( ~n1751 & n4467 ) | ( ~n1751 & n4468 ) | ( n4467 & n4468 ) ;
  assign n4470 = ( ~n1787 & n4467 ) | ( ~n1787 & n4468 ) | ( n4467 & n4468 ) ;
  assign n4471 = ( n1794 & n4467 ) | ( n1794 & n4468 ) | ( n4467 & n4468 ) ;
  assign n4472 = ( n1783 & n4470 ) | ( n1783 & n4471 ) | ( n4470 & n4471 ) ;
  assign n4473 = ( n1643 & n4469 ) | ( n1643 & n4472 ) | ( n4469 & n4472 ) ;
  assign n4474 = ( ~n1822 & n4469 ) | ( ~n1822 & n4472 ) | ( n4469 & n4472 ) ;
  assign n4475 = ( ~n1324 & n4473 ) | ( ~n1324 & n4474 ) | ( n4473 & n4474 ) ;
  assign n4476 = x81 & ~n1767 ;
  assign n4477 = x81 & n1771 ;
  assign n4478 = ( n1751 & n4476 ) | ( n1751 & n4477 ) | ( n4476 & n4477 ) ;
  assign n4479 = ( n1787 & n4476 ) | ( n1787 & n4477 ) | ( n4476 & n4477 ) ;
  assign n4480 = ( ~n1794 & n4476 ) | ( ~n1794 & n4477 ) | ( n4476 & n4477 ) ;
  assign n4481 = ( ~n1783 & n4479 ) | ( ~n1783 & n4480 ) | ( n4479 & n4480 ) ;
  assign n4482 = ( ~n1643 & n4478 ) | ( ~n1643 & n4481 ) | ( n4478 & n4481 ) ;
  assign n4483 = ( n1822 & n4478 ) | ( n1822 & n4481 ) | ( n4478 & n4481 ) ;
  assign n4484 = ( n1324 & n4482 ) | ( n1324 & n4483 ) | ( n4482 & n4483 ) ;
  assign n4485 = n4475 | n4484 ;
  assign n4486 = x465 & n991 ;
  assign n4487 = x465 & ~n995 ;
  assign n4488 = ( ~n1104 & n4486 ) | ( ~n1104 & n4487 ) | ( n4486 & n4487 ) ;
  assign n4489 = ( ~n1119 & n4486 ) | ( ~n1119 & n4487 ) | ( n4486 & n4487 ) ;
  assign n4490 = ( n1126 & n4486 ) | ( n1126 & n4487 ) | ( n4486 & n4487 ) ;
  assign n4491 = ( n1115 & n4489 ) | ( n1115 & n4490 ) | ( n4489 & n4490 ) ;
  assign n4492 = ( n975 & n4488 ) | ( n975 & n4491 ) | ( n4488 & n4491 ) ;
  assign n4493 = ( ~n1154 & n4488 ) | ( ~n1154 & n4491 ) | ( n4488 & n4491 ) ;
  assign n4494 = ( x409 & n4492 ) | ( x409 & n4493 ) | ( n4492 & n4493 ) ;
  assign n4495 = ( ~x281 & n4492 ) | ( ~x281 & n4493 ) | ( n4492 & n4493 ) ;
  assign n4496 = ( ~n656 & n4494 ) | ( ~n656 & n4495 ) | ( n4494 & n4495 ) ;
  assign n4497 = x337 & ~n991 ;
  assign n4498 = x337 & n995 ;
  assign n4499 = ( n1104 & n4497 ) | ( n1104 & n4498 ) | ( n4497 & n4498 ) ;
  assign n4500 = ( n1119 & n4497 ) | ( n1119 & n4498 ) | ( n4497 & n4498 ) ;
  assign n4501 = ( ~n1126 & n4497 ) | ( ~n1126 & n4498 ) | ( n4497 & n4498 ) ;
  assign n4502 = ( ~n1115 & n4500 ) | ( ~n1115 & n4501 ) | ( n4500 & n4501 ) ;
  assign n4503 = ( ~n975 & n4499 ) | ( ~n975 & n4502 ) | ( n4499 & n4502 ) ;
  assign n4504 = ( n1154 & n4499 ) | ( n1154 & n4502 ) | ( n4499 & n4502 ) ;
  assign n4505 = ( ~x409 & n4503 ) | ( ~x409 & n4504 ) | ( n4503 & n4504 ) ;
  assign n4506 = ( x281 & n4503 ) | ( x281 & n4504 ) | ( n4503 & n4504 ) ;
  assign n4507 = ( n656 & n4505 ) | ( n656 & n4506 ) | ( n4505 & n4506 ) ;
  assign n4508 = n4496 | n4507 ;
  assign n4509 = ~n4444 & n4463 ;
  assign n4510 = ( n4485 & ~n4508 ) | ( n4485 & n4509 ) | ( ~n4508 & n4509 ) ;
  assign n4511 = ~n4400 & n4419 ;
  assign n4512 = ~n4420 & n4511 ;
  assign n4513 = ( ~n4420 & n4510 ) | ( ~n4420 & n4512 ) | ( n4510 & n4512 ) ;
  assign n4514 = ( n4353 & ~n4376 ) | ( n4353 & n4513 ) | ( ~n4376 & n4513 ) ;
  assign n4515 = ( n4334 & n4466 ) | ( n4334 & ~n4514 ) | ( n4466 & ~n4514 ) ;
  assign n4516 = ~n4225 & n4244 ;
  assign n4517 = ~n4202 & n4516 ;
  assign n4518 = n4246 & ~n4517 ;
  assign n4519 = n4308 & ~n4331 ;
  assign n4520 = ( n4265 & ~n4288 ) | ( n4265 & n4519 ) | ( ~n4288 & n4519 ) ;
  assign n4521 = ( n4517 & ~n4518 ) | ( n4517 & n4520 ) | ( ~n4518 & n4520 ) ;
  assign n4522 = n4515 & ~n4521 ;
  assign n4523 = x223 & n1767 ;
  assign n4524 = x223 & ~n1771 ;
  assign n4525 = ( ~n1751 & n4523 ) | ( ~n1751 & n4524 ) | ( n4523 & n4524 ) ;
  assign n4526 = ( ~n1787 & n4523 ) | ( ~n1787 & n4524 ) | ( n4523 & n4524 ) ;
  assign n4527 = ( n1794 & n4523 ) | ( n1794 & n4524 ) | ( n4523 & n4524 ) ;
  assign n4528 = ( n1783 & n4526 ) | ( n1783 & n4527 ) | ( n4526 & n4527 ) ;
  assign n4529 = ( n1643 & n4525 ) | ( n1643 & n4528 ) | ( n4525 & n4528 ) ;
  assign n4530 = ( ~n1822 & n4525 ) | ( ~n1822 & n4528 ) | ( n4525 & n4528 ) ;
  assign n4531 = ( ~n1324 & n4529 ) | ( ~n1324 & n4530 ) | ( n4529 & n4530 ) ;
  assign n4532 = x95 & ~n1767 ;
  assign n4533 = x95 & n1771 ;
  assign n4534 = ( n1751 & n4532 ) | ( n1751 & n4533 ) | ( n4532 & n4533 ) ;
  assign n4535 = ( n1787 & n4532 ) | ( n1787 & n4533 ) | ( n4532 & n4533 ) ;
  assign n4536 = ( ~n1794 & n4532 ) | ( ~n1794 & n4533 ) | ( n4532 & n4533 ) ;
  assign n4537 = ( ~n1783 & n4535 ) | ( ~n1783 & n4536 ) | ( n4535 & n4536 ) ;
  assign n4538 = ( ~n1643 & n4534 ) | ( ~n1643 & n4537 ) | ( n4534 & n4537 ) ;
  assign n4539 = ( n1822 & n4534 ) | ( n1822 & n4537 ) | ( n4534 & n4537 ) ;
  assign n4540 = ( n1324 & n4538 ) | ( n1324 & n4539 ) | ( n4538 & n4539 ) ;
  assign n4541 = n4531 | n4540 ;
  assign n4542 = x479 & n991 ;
  assign n4543 = x479 & ~n995 ;
  assign n4544 = ( ~n1104 & n4542 ) | ( ~n1104 & n4543 ) | ( n4542 & n4543 ) ;
  assign n4545 = ( ~n1119 & n4542 ) | ( ~n1119 & n4543 ) | ( n4542 & n4543 ) ;
  assign n4546 = ( n1126 & n4542 ) | ( n1126 & n4543 ) | ( n4542 & n4543 ) ;
  assign n4547 = ( n1115 & n4545 ) | ( n1115 & n4546 ) | ( n4545 & n4546 ) ;
  assign n4548 = ( n975 & n4544 ) | ( n975 & n4547 ) | ( n4544 & n4547 ) ;
  assign n4549 = ( ~n1154 & n4544 ) | ( ~n1154 & n4547 ) | ( n4544 & n4547 ) ;
  assign n4550 = ( x409 & n4548 ) | ( x409 & n4549 ) | ( n4548 & n4549 ) ;
  assign n4551 = ( ~x281 & n4548 ) | ( ~x281 & n4549 ) | ( n4548 & n4549 ) ;
  assign n4552 = ( ~n656 & n4550 ) | ( ~n656 & n4551 ) | ( n4550 & n4551 ) ;
  assign n4553 = x351 & ~n991 ;
  assign n4554 = x351 & n995 ;
  assign n4555 = ( n1104 & n4553 ) | ( n1104 & n4554 ) | ( n4553 & n4554 ) ;
  assign n4556 = ( n1119 & n4553 ) | ( n1119 & n4554 ) | ( n4553 & n4554 ) ;
  assign n4557 = ( ~n1126 & n4553 ) | ( ~n1126 & n4554 ) | ( n4553 & n4554 ) ;
  assign n4558 = ( ~n1115 & n4556 ) | ( ~n1115 & n4557 ) | ( n4556 & n4557 ) ;
  assign n4559 = ( ~n975 & n4555 ) | ( ~n975 & n4558 ) | ( n4555 & n4558 ) ;
  assign n4560 = ( n1154 & n4555 ) | ( n1154 & n4558 ) | ( n4555 & n4558 ) ;
  assign n4561 = ( ~x409 & n4559 ) | ( ~x409 & n4560 ) | ( n4559 & n4560 ) ;
  assign n4562 = ( x281 & n4559 ) | ( x281 & n4560 ) | ( n4559 & n4560 ) ;
  assign n4563 = ( n656 & n4561 ) | ( n656 & n4562 ) | ( n4561 & n4562 ) ;
  assign n4564 = n4552 | n4563 ;
  assign n4565 = ~n4541 & n4564 ;
  assign n4566 = x478 & n991 ;
  assign n4567 = x478 & ~n995 ;
  assign n4568 = ( ~n1104 & n4566 ) | ( ~n1104 & n4567 ) | ( n4566 & n4567 ) ;
  assign n4569 = ( ~n1119 & n4566 ) | ( ~n1119 & n4567 ) | ( n4566 & n4567 ) ;
  assign n4570 = ( n1126 & n4566 ) | ( n1126 & n4567 ) | ( n4566 & n4567 ) ;
  assign n4571 = ( n1115 & n4569 ) | ( n1115 & n4570 ) | ( n4569 & n4570 ) ;
  assign n4572 = ( n975 & n4568 ) | ( n975 & n4571 ) | ( n4568 & n4571 ) ;
  assign n4573 = ( ~n1154 & n4568 ) | ( ~n1154 & n4571 ) | ( n4568 & n4571 ) ;
  assign n4574 = ( x409 & n4572 ) | ( x409 & n4573 ) | ( n4572 & n4573 ) ;
  assign n4575 = ( ~x281 & n4572 ) | ( ~x281 & n4573 ) | ( n4572 & n4573 ) ;
  assign n4576 = ( ~n656 & n4574 ) | ( ~n656 & n4575 ) | ( n4574 & n4575 ) ;
  assign n4577 = x350 & ~n991 ;
  assign n4578 = x350 & n995 ;
  assign n4579 = ( n1104 & n4577 ) | ( n1104 & n4578 ) | ( n4577 & n4578 ) ;
  assign n4580 = ( n1119 & n4577 ) | ( n1119 & n4578 ) | ( n4577 & n4578 ) ;
  assign n4581 = ( ~n1126 & n4577 ) | ( ~n1126 & n4578 ) | ( n4577 & n4578 ) ;
  assign n4582 = ( ~n1115 & n4580 ) | ( ~n1115 & n4581 ) | ( n4580 & n4581 ) ;
  assign n4583 = ( ~n975 & n4579 ) | ( ~n975 & n4582 ) | ( n4579 & n4582 ) ;
  assign n4584 = ( n1154 & n4579 ) | ( n1154 & n4582 ) | ( n4579 & n4582 ) ;
  assign n4585 = ( ~x409 & n4583 ) | ( ~x409 & n4584 ) | ( n4583 & n4584 ) ;
  assign n4586 = ( x281 & n4583 ) | ( x281 & n4584 ) | ( n4583 & n4584 ) ;
  assign n4587 = ( n656 & n4585 ) | ( n656 & n4586 ) | ( n4585 & n4586 ) ;
  assign n4588 = n4576 | n4587 ;
  assign n4589 = x222 & n1767 ;
  assign n4590 = x222 & ~n1771 ;
  assign n4591 = ( ~n1751 & n4589 ) | ( ~n1751 & n4590 ) | ( n4589 & n4590 ) ;
  assign n4592 = ( ~n1787 & n4589 ) | ( ~n1787 & n4590 ) | ( n4589 & n4590 ) ;
  assign n4593 = ( n1794 & n4589 ) | ( n1794 & n4590 ) | ( n4589 & n4590 ) ;
  assign n4594 = ( n1783 & n4592 ) | ( n1783 & n4593 ) | ( n4592 & n4593 ) ;
  assign n4595 = ( n1643 & n4591 ) | ( n1643 & n4594 ) | ( n4591 & n4594 ) ;
  assign n4596 = ( ~n1822 & n4591 ) | ( ~n1822 & n4594 ) | ( n4591 & n4594 ) ;
  assign n4597 = ( ~n1324 & n4595 ) | ( ~n1324 & n4596 ) | ( n4595 & n4596 ) ;
  assign n4598 = x94 & ~n1767 ;
  assign n4599 = x94 & n1771 ;
  assign n4600 = ( n1751 & n4598 ) | ( n1751 & n4599 ) | ( n4598 & n4599 ) ;
  assign n4601 = ( n1787 & n4598 ) | ( n1787 & n4599 ) | ( n4598 & n4599 ) ;
  assign n4602 = ( ~n1794 & n4598 ) | ( ~n1794 & n4599 ) | ( n4598 & n4599 ) ;
  assign n4603 = ( ~n1783 & n4601 ) | ( ~n1783 & n4602 ) | ( n4601 & n4602 ) ;
  assign n4604 = ( ~n1643 & n4600 ) | ( ~n1643 & n4603 ) | ( n4600 & n4603 ) ;
  assign n4605 = ( n1822 & n4600 ) | ( n1822 & n4603 ) | ( n4600 & n4603 ) ;
  assign n4606 = ( n1324 & n4604 ) | ( n1324 & n4605 ) | ( n4604 & n4605 ) ;
  assign n4607 = n4597 | n4606 ;
  assign n4608 = n4588 & ~n4607 ;
  assign n4609 = n4565 | n4608 ;
  assign n4610 = x221 & n1767 ;
  assign n4611 = x221 & ~n1771 ;
  assign n4612 = ( ~n1751 & n4610 ) | ( ~n1751 & n4611 ) | ( n4610 & n4611 ) ;
  assign n4613 = ( ~n1787 & n4610 ) | ( ~n1787 & n4611 ) | ( n4610 & n4611 ) ;
  assign n4614 = ( n1794 & n4610 ) | ( n1794 & n4611 ) | ( n4610 & n4611 ) ;
  assign n4615 = ( n1783 & n4613 ) | ( n1783 & n4614 ) | ( n4613 & n4614 ) ;
  assign n4616 = ( n1643 & n4612 ) | ( n1643 & n4615 ) | ( n4612 & n4615 ) ;
  assign n4617 = ( ~n1822 & n4612 ) | ( ~n1822 & n4615 ) | ( n4612 & n4615 ) ;
  assign n4618 = ( ~n1324 & n4616 ) | ( ~n1324 & n4617 ) | ( n4616 & n4617 ) ;
  assign n4619 = x93 & ~n1767 ;
  assign n4620 = x93 & n1771 ;
  assign n4621 = ( n1751 & n4619 ) | ( n1751 & n4620 ) | ( n4619 & n4620 ) ;
  assign n4622 = ( n1787 & n4619 ) | ( n1787 & n4620 ) | ( n4619 & n4620 ) ;
  assign n4623 = ( ~n1794 & n4619 ) | ( ~n1794 & n4620 ) | ( n4619 & n4620 ) ;
  assign n4624 = ( ~n1783 & n4622 ) | ( ~n1783 & n4623 ) | ( n4622 & n4623 ) ;
  assign n4625 = ( ~n1643 & n4621 ) | ( ~n1643 & n4624 ) | ( n4621 & n4624 ) ;
  assign n4626 = ( n1822 & n4621 ) | ( n1822 & n4624 ) | ( n4621 & n4624 ) ;
  assign n4627 = ( n1324 & n4625 ) | ( n1324 & n4626 ) | ( n4625 & n4626 ) ;
  assign n4628 = n4618 | n4627 ;
  assign n4629 = x477 & n991 ;
  assign n4630 = x477 & ~n995 ;
  assign n4631 = ( ~n1104 & n4629 ) | ( ~n1104 & n4630 ) | ( n4629 & n4630 ) ;
  assign n4632 = ( ~n1119 & n4629 ) | ( ~n1119 & n4630 ) | ( n4629 & n4630 ) ;
  assign n4633 = ( n1126 & n4629 ) | ( n1126 & n4630 ) | ( n4629 & n4630 ) ;
  assign n4634 = ( n1115 & n4632 ) | ( n1115 & n4633 ) | ( n4632 & n4633 ) ;
  assign n4635 = ( n975 & n4631 ) | ( n975 & n4634 ) | ( n4631 & n4634 ) ;
  assign n4636 = ( ~n1154 & n4631 ) | ( ~n1154 & n4634 ) | ( n4631 & n4634 ) ;
  assign n4637 = ( x409 & n4635 ) | ( x409 & n4636 ) | ( n4635 & n4636 ) ;
  assign n4638 = ( ~x281 & n4635 ) | ( ~x281 & n4636 ) | ( n4635 & n4636 ) ;
  assign n4639 = ( ~n656 & n4637 ) | ( ~n656 & n4638 ) | ( n4637 & n4638 ) ;
  assign n4640 = x349 & ~n991 ;
  assign n4641 = x349 & n995 ;
  assign n4642 = ( n1104 & n4640 ) | ( n1104 & n4641 ) | ( n4640 & n4641 ) ;
  assign n4643 = ( n1119 & n4640 ) | ( n1119 & n4641 ) | ( n4640 & n4641 ) ;
  assign n4644 = ( ~n1126 & n4640 ) | ( ~n1126 & n4641 ) | ( n4640 & n4641 ) ;
  assign n4645 = ( ~n1115 & n4643 ) | ( ~n1115 & n4644 ) | ( n4643 & n4644 ) ;
  assign n4646 = ( ~n975 & n4642 ) | ( ~n975 & n4645 ) | ( n4642 & n4645 ) ;
  assign n4647 = ( n1154 & n4642 ) | ( n1154 & n4645 ) | ( n4642 & n4645 ) ;
  assign n4648 = ( ~x409 & n4646 ) | ( ~x409 & n4647 ) | ( n4646 & n4647 ) ;
  assign n4649 = ( x281 & n4646 ) | ( x281 & n4647 ) | ( n4646 & n4647 ) ;
  assign n4650 = ( n656 & n4648 ) | ( n656 & n4649 ) | ( n4648 & n4649 ) ;
  assign n4651 = n4639 | n4650 ;
  assign n4652 = ~n4628 & n4651 ;
  assign n4653 = x220 & n1767 ;
  assign n4654 = x220 & ~n1771 ;
  assign n4655 = ( ~n1751 & n4653 ) | ( ~n1751 & n4654 ) | ( n4653 & n4654 ) ;
  assign n4656 = ( ~n1787 & n4653 ) | ( ~n1787 & n4654 ) | ( n4653 & n4654 ) ;
  assign n4657 = ( n1794 & n4653 ) | ( n1794 & n4654 ) | ( n4653 & n4654 ) ;
  assign n4658 = ( n1783 & n4656 ) | ( n1783 & n4657 ) | ( n4656 & n4657 ) ;
  assign n4659 = ( n1643 & n4655 ) | ( n1643 & n4658 ) | ( n4655 & n4658 ) ;
  assign n4660 = ( ~n1822 & n4655 ) | ( ~n1822 & n4658 ) | ( n4655 & n4658 ) ;
  assign n4661 = ( ~n1324 & n4659 ) | ( ~n1324 & n4660 ) | ( n4659 & n4660 ) ;
  assign n4662 = x92 & ~n1767 ;
  assign n4663 = x92 & n1771 ;
  assign n4664 = ( n1751 & n4662 ) | ( n1751 & n4663 ) | ( n4662 & n4663 ) ;
  assign n4665 = ( n1787 & n4662 ) | ( n1787 & n4663 ) | ( n4662 & n4663 ) ;
  assign n4666 = ( ~n1794 & n4662 ) | ( ~n1794 & n4663 ) | ( n4662 & n4663 ) ;
  assign n4667 = ( ~n1783 & n4665 ) | ( ~n1783 & n4666 ) | ( n4665 & n4666 ) ;
  assign n4668 = ( ~n1643 & n4664 ) | ( ~n1643 & n4667 ) | ( n4664 & n4667 ) ;
  assign n4669 = ( n1822 & n4664 ) | ( n1822 & n4667 ) | ( n4664 & n4667 ) ;
  assign n4670 = ( n1324 & n4668 ) | ( n1324 & n4669 ) | ( n4668 & n4669 ) ;
  assign n4671 = n4661 | n4670 ;
  assign n4672 = x476 & n991 ;
  assign n4673 = x476 & ~n995 ;
  assign n4674 = ( ~n1104 & n4672 ) | ( ~n1104 & n4673 ) | ( n4672 & n4673 ) ;
  assign n4675 = ( ~n1119 & n4672 ) | ( ~n1119 & n4673 ) | ( n4672 & n4673 ) ;
  assign n4676 = ( n1126 & n4672 ) | ( n1126 & n4673 ) | ( n4672 & n4673 ) ;
  assign n4677 = ( n1115 & n4675 ) | ( n1115 & n4676 ) | ( n4675 & n4676 ) ;
  assign n4678 = ( n975 & n4674 ) | ( n975 & n4677 ) | ( n4674 & n4677 ) ;
  assign n4679 = ( ~n1154 & n4674 ) | ( ~n1154 & n4677 ) | ( n4674 & n4677 ) ;
  assign n4680 = ( x409 & n4678 ) | ( x409 & n4679 ) | ( n4678 & n4679 ) ;
  assign n4681 = ( ~x281 & n4678 ) | ( ~x281 & n4679 ) | ( n4678 & n4679 ) ;
  assign n4682 = ( ~n656 & n4680 ) | ( ~n656 & n4681 ) | ( n4680 & n4681 ) ;
  assign n4683 = x348 & ~n991 ;
  assign n4684 = x348 & n995 ;
  assign n4685 = ( n1104 & n4683 ) | ( n1104 & n4684 ) | ( n4683 & n4684 ) ;
  assign n4686 = ( n1119 & n4683 ) | ( n1119 & n4684 ) | ( n4683 & n4684 ) ;
  assign n4687 = ( ~n1126 & n4683 ) | ( ~n1126 & n4684 ) | ( n4683 & n4684 ) ;
  assign n4688 = ( ~n1115 & n4686 ) | ( ~n1115 & n4687 ) | ( n4686 & n4687 ) ;
  assign n4689 = ( ~n975 & n4685 ) | ( ~n975 & n4688 ) | ( n4685 & n4688 ) ;
  assign n4690 = ( n1154 & n4685 ) | ( n1154 & n4688 ) | ( n4685 & n4688 ) ;
  assign n4691 = ( ~x409 & n4689 ) | ( ~x409 & n4690 ) | ( n4689 & n4690 ) ;
  assign n4692 = ( x281 & n4689 ) | ( x281 & n4690 ) | ( n4689 & n4690 ) ;
  assign n4693 = ( n656 & n4691 ) | ( n656 & n4692 ) | ( n4691 & n4692 ) ;
  assign n4694 = n4682 | n4693 ;
  assign n4695 = ~n4671 & n4694 ;
  assign n4696 = n4652 | n4695 ;
  assign n4697 = n4609 | n4696 ;
  assign n4698 = n4178 & ~n4201 ;
  assign n4699 = x219 & n1767 ;
  assign n4700 = x219 & ~n1771 ;
  assign n4701 = ( ~n1751 & n4699 ) | ( ~n1751 & n4700 ) | ( n4699 & n4700 ) ;
  assign n4702 = ( ~n1787 & n4699 ) | ( ~n1787 & n4700 ) | ( n4699 & n4700 ) ;
  assign n4703 = ( n1794 & n4699 ) | ( n1794 & n4700 ) | ( n4699 & n4700 ) ;
  assign n4704 = ( n1783 & n4702 ) | ( n1783 & n4703 ) | ( n4702 & n4703 ) ;
  assign n4705 = ( n1643 & n4701 ) | ( n1643 & n4704 ) | ( n4701 & n4704 ) ;
  assign n4706 = ( ~n1822 & n4701 ) | ( ~n1822 & n4704 ) | ( n4701 & n4704 ) ;
  assign n4707 = ( ~n1324 & n4705 ) | ( ~n1324 & n4706 ) | ( n4705 & n4706 ) ;
  assign n4708 = x91 & ~n1767 ;
  assign n4709 = x91 & n1771 ;
  assign n4710 = ( n1751 & n4708 ) | ( n1751 & n4709 ) | ( n4708 & n4709 ) ;
  assign n4711 = ( n1787 & n4708 ) | ( n1787 & n4709 ) | ( n4708 & n4709 ) ;
  assign n4712 = ( ~n1794 & n4708 ) | ( ~n1794 & n4709 ) | ( n4708 & n4709 ) ;
  assign n4713 = ( ~n1783 & n4711 ) | ( ~n1783 & n4712 ) | ( n4711 & n4712 ) ;
  assign n4714 = ( ~n1643 & n4710 ) | ( ~n1643 & n4713 ) | ( n4710 & n4713 ) ;
  assign n4715 = ( n1822 & n4710 ) | ( n1822 & n4713 ) | ( n4710 & n4713 ) ;
  assign n4716 = ( n1324 & n4714 ) | ( n1324 & n4715 ) | ( n4714 & n4715 ) ;
  assign n4717 = n4707 | n4716 ;
  assign n4718 = x475 & n991 ;
  assign n4719 = x475 & ~n995 ;
  assign n4720 = ( ~n1104 & n4718 ) | ( ~n1104 & n4719 ) | ( n4718 & n4719 ) ;
  assign n4721 = ( ~n1119 & n4718 ) | ( ~n1119 & n4719 ) | ( n4718 & n4719 ) ;
  assign n4722 = ( n1126 & n4718 ) | ( n1126 & n4719 ) | ( n4718 & n4719 ) ;
  assign n4723 = ( n1115 & n4721 ) | ( n1115 & n4722 ) | ( n4721 & n4722 ) ;
  assign n4724 = ( n975 & n4720 ) | ( n975 & n4723 ) | ( n4720 & n4723 ) ;
  assign n4725 = ( ~n1154 & n4720 ) | ( ~n1154 & n4723 ) | ( n4720 & n4723 ) ;
  assign n4726 = ( x409 & n4724 ) | ( x409 & n4725 ) | ( n4724 & n4725 ) ;
  assign n4727 = ( ~x281 & n4724 ) | ( ~x281 & n4725 ) | ( n4724 & n4725 ) ;
  assign n4728 = ( ~n656 & n4726 ) | ( ~n656 & n4727 ) | ( n4726 & n4727 ) ;
  assign n4729 = x347 & ~n991 ;
  assign n4730 = x347 & n995 ;
  assign n4731 = ( n1104 & n4729 ) | ( n1104 & n4730 ) | ( n4729 & n4730 ) ;
  assign n4732 = ( n1119 & n4729 ) | ( n1119 & n4730 ) | ( n4729 & n4730 ) ;
  assign n4733 = ( ~n1126 & n4729 ) | ( ~n1126 & n4730 ) | ( n4729 & n4730 ) ;
  assign n4734 = ( ~n1115 & n4732 ) | ( ~n1115 & n4733 ) | ( n4732 & n4733 ) ;
  assign n4735 = ( ~n975 & n4731 ) | ( ~n975 & n4734 ) | ( n4731 & n4734 ) ;
  assign n4736 = ( n1154 & n4731 ) | ( n1154 & n4734 ) | ( n4731 & n4734 ) ;
  assign n4737 = ( ~x409 & n4735 ) | ( ~x409 & n4736 ) | ( n4735 & n4736 ) ;
  assign n4738 = ( x281 & n4735 ) | ( x281 & n4736 ) | ( n4735 & n4736 ) ;
  assign n4739 = ( n656 & n4737 ) | ( n656 & n4738 ) | ( n4737 & n4738 ) ;
  assign n4740 = n4728 | n4739 ;
  assign n4741 = ~n4717 & n4740 ;
  assign n4742 = x474 & n991 ;
  assign n4743 = x474 & ~n995 ;
  assign n4744 = ( ~n1104 & n4742 ) | ( ~n1104 & n4743 ) | ( n4742 & n4743 ) ;
  assign n4745 = ( ~n1119 & n4742 ) | ( ~n1119 & n4743 ) | ( n4742 & n4743 ) ;
  assign n4746 = ( n1126 & n4742 ) | ( n1126 & n4743 ) | ( n4742 & n4743 ) ;
  assign n4747 = ( n1115 & n4745 ) | ( n1115 & n4746 ) | ( n4745 & n4746 ) ;
  assign n4748 = ( n975 & n4744 ) | ( n975 & n4747 ) | ( n4744 & n4747 ) ;
  assign n4749 = ( ~n1154 & n4744 ) | ( ~n1154 & n4747 ) | ( n4744 & n4747 ) ;
  assign n4750 = ( x409 & n4748 ) | ( x409 & n4749 ) | ( n4748 & n4749 ) ;
  assign n4751 = ( ~x281 & n4748 ) | ( ~x281 & n4749 ) | ( n4748 & n4749 ) ;
  assign n4752 = ( ~n656 & n4750 ) | ( ~n656 & n4751 ) | ( n4750 & n4751 ) ;
  assign n4753 = x346 & ~n991 ;
  assign n4754 = x346 & n995 ;
  assign n4755 = ( n1104 & n4753 ) | ( n1104 & n4754 ) | ( n4753 & n4754 ) ;
  assign n4756 = ( n1119 & n4753 ) | ( n1119 & n4754 ) | ( n4753 & n4754 ) ;
  assign n4757 = ( ~n1126 & n4753 ) | ( ~n1126 & n4754 ) | ( n4753 & n4754 ) ;
  assign n4758 = ( ~n1115 & n4756 ) | ( ~n1115 & n4757 ) | ( n4756 & n4757 ) ;
  assign n4759 = ( ~n975 & n4755 ) | ( ~n975 & n4758 ) | ( n4755 & n4758 ) ;
  assign n4760 = ( n1154 & n4755 ) | ( n1154 & n4758 ) | ( n4755 & n4758 ) ;
  assign n4761 = ( ~x409 & n4759 ) | ( ~x409 & n4760 ) | ( n4759 & n4760 ) ;
  assign n4762 = ( x281 & n4759 ) | ( x281 & n4760 ) | ( n4759 & n4760 ) ;
  assign n4763 = ( n656 & n4761 ) | ( n656 & n4762 ) | ( n4761 & n4762 ) ;
  assign n4764 = n4752 | n4763 ;
  assign n4765 = x218 & n1767 ;
  assign n4766 = x218 & ~n1771 ;
  assign n4767 = ( ~n1751 & n4765 ) | ( ~n1751 & n4766 ) | ( n4765 & n4766 ) ;
  assign n4768 = ( ~n1787 & n4765 ) | ( ~n1787 & n4766 ) | ( n4765 & n4766 ) ;
  assign n4769 = ( n1794 & n4765 ) | ( n1794 & n4766 ) | ( n4765 & n4766 ) ;
  assign n4770 = ( n1783 & n4768 ) | ( n1783 & n4769 ) | ( n4768 & n4769 ) ;
  assign n4771 = ( n1643 & n4767 ) | ( n1643 & n4770 ) | ( n4767 & n4770 ) ;
  assign n4772 = ( ~n1822 & n4767 ) | ( ~n1822 & n4770 ) | ( n4767 & n4770 ) ;
  assign n4773 = ( ~n1324 & n4771 ) | ( ~n1324 & n4772 ) | ( n4771 & n4772 ) ;
  assign n4774 = x90 & ~n1767 ;
  assign n4775 = x90 & n1771 ;
  assign n4776 = ( n1751 & n4774 ) | ( n1751 & n4775 ) | ( n4774 & n4775 ) ;
  assign n4777 = ( n1787 & n4774 ) | ( n1787 & n4775 ) | ( n4774 & n4775 ) ;
  assign n4778 = ( ~n1794 & n4774 ) | ( ~n1794 & n4775 ) | ( n4774 & n4775 ) ;
  assign n4779 = ( ~n1783 & n4777 ) | ( ~n1783 & n4778 ) | ( n4777 & n4778 ) ;
  assign n4780 = ( ~n1643 & n4776 ) | ( ~n1643 & n4779 ) | ( n4776 & n4779 ) ;
  assign n4781 = ( n1822 & n4776 ) | ( n1822 & n4779 ) | ( n4776 & n4779 ) ;
  assign n4782 = ( n1324 & n4780 ) | ( n1324 & n4781 ) | ( n4780 & n4781 ) ;
  assign n4783 = n4773 | n4782 ;
  assign n4784 = n4764 & ~n4783 ;
  assign n4785 = n4741 | n4784 ;
  assign n4786 = x217 & n1767 ;
  assign n4787 = x217 & ~n1771 ;
  assign n4788 = ( ~n1751 & n4786 ) | ( ~n1751 & n4787 ) | ( n4786 & n4787 ) ;
  assign n4789 = ( ~n1787 & n4786 ) | ( ~n1787 & n4787 ) | ( n4786 & n4787 ) ;
  assign n4790 = ( n1794 & n4786 ) | ( n1794 & n4787 ) | ( n4786 & n4787 ) ;
  assign n4791 = ( n1783 & n4789 ) | ( n1783 & n4790 ) | ( n4789 & n4790 ) ;
  assign n4792 = ( n1643 & n4788 ) | ( n1643 & n4791 ) | ( n4788 & n4791 ) ;
  assign n4793 = ( ~n1822 & n4788 ) | ( ~n1822 & n4791 ) | ( n4788 & n4791 ) ;
  assign n4794 = ( ~n1324 & n4792 ) | ( ~n1324 & n4793 ) | ( n4792 & n4793 ) ;
  assign n4795 = x89 & ~n1767 ;
  assign n4796 = x89 & n1771 ;
  assign n4797 = ( n1751 & n4795 ) | ( n1751 & n4796 ) | ( n4795 & n4796 ) ;
  assign n4798 = ( n1787 & n4795 ) | ( n1787 & n4796 ) | ( n4795 & n4796 ) ;
  assign n4799 = ( ~n1794 & n4795 ) | ( ~n1794 & n4796 ) | ( n4795 & n4796 ) ;
  assign n4800 = ( ~n1783 & n4798 ) | ( ~n1783 & n4799 ) | ( n4798 & n4799 ) ;
  assign n4801 = ( ~n1643 & n4797 ) | ( ~n1643 & n4800 ) | ( n4797 & n4800 ) ;
  assign n4802 = ( n1822 & n4797 ) | ( n1822 & n4800 ) | ( n4797 & n4800 ) ;
  assign n4803 = ( n1324 & n4801 ) | ( n1324 & n4802 ) | ( n4801 & n4802 ) ;
  assign n4804 = n4794 | n4803 ;
  assign n4805 = x473 & n991 ;
  assign n4806 = x473 & ~n995 ;
  assign n4807 = ( ~n1104 & n4805 ) | ( ~n1104 & n4806 ) | ( n4805 & n4806 ) ;
  assign n4808 = ( ~n1119 & n4805 ) | ( ~n1119 & n4806 ) | ( n4805 & n4806 ) ;
  assign n4809 = ( n1126 & n4805 ) | ( n1126 & n4806 ) | ( n4805 & n4806 ) ;
  assign n4810 = ( n1115 & n4808 ) | ( n1115 & n4809 ) | ( n4808 & n4809 ) ;
  assign n4811 = ( n975 & n4807 ) | ( n975 & n4810 ) | ( n4807 & n4810 ) ;
  assign n4812 = ( ~n1154 & n4807 ) | ( ~n1154 & n4810 ) | ( n4807 & n4810 ) ;
  assign n4813 = ( x409 & n4811 ) | ( x409 & n4812 ) | ( n4811 & n4812 ) ;
  assign n4814 = ( ~x281 & n4811 ) | ( ~x281 & n4812 ) | ( n4811 & n4812 ) ;
  assign n4815 = ( ~n656 & n4813 ) | ( ~n656 & n4814 ) | ( n4813 & n4814 ) ;
  assign n4816 = x345 & ~n991 ;
  assign n4817 = x345 & n995 ;
  assign n4818 = ( n1104 & n4816 ) | ( n1104 & n4817 ) | ( n4816 & n4817 ) ;
  assign n4819 = ( n1119 & n4816 ) | ( n1119 & n4817 ) | ( n4816 & n4817 ) ;
  assign n4820 = ( ~n1126 & n4816 ) | ( ~n1126 & n4817 ) | ( n4816 & n4817 ) ;
  assign n4821 = ( ~n1115 & n4819 ) | ( ~n1115 & n4820 ) | ( n4819 & n4820 ) ;
  assign n4822 = ( ~n975 & n4818 ) | ( ~n975 & n4821 ) | ( n4818 & n4821 ) ;
  assign n4823 = ( n1154 & n4818 ) | ( n1154 & n4821 ) | ( n4818 & n4821 ) ;
  assign n4824 = ( ~x409 & n4822 ) | ( ~x409 & n4823 ) | ( n4822 & n4823 ) ;
  assign n4825 = ( x281 & n4822 ) | ( x281 & n4823 ) | ( n4822 & n4823 ) ;
  assign n4826 = ( n656 & n4824 ) | ( n656 & n4825 ) | ( n4824 & n4825 ) ;
  assign n4827 = n4815 | n4826 ;
  assign n4828 = ~n4804 & n4827 ;
  assign n4829 = x472 & n991 ;
  assign n4830 = x472 & ~n995 ;
  assign n4831 = ( ~n1104 & n4829 ) | ( ~n1104 & n4830 ) | ( n4829 & n4830 ) ;
  assign n4832 = ( ~n1119 & n4829 ) | ( ~n1119 & n4830 ) | ( n4829 & n4830 ) ;
  assign n4833 = ( n1126 & n4829 ) | ( n1126 & n4830 ) | ( n4829 & n4830 ) ;
  assign n4834 = ( n1115 & n4832 ) | ( n1115 & n4833 ) | ( n4832 & n4833 ) ;
  assign n4835 = ( n975 & n4831 ) | ( n975 & n4834 ) | ( n4831 & n4834 ) ;
  assign n4836 = ( ~n1154 & n4831 ) | ( ~n1154 & n4834 ) | ( n4831 & n4834 ) ;
  assign n4837 = ( x409 & n4835 ) | ( x409 & n4836 ) | ( n4835 & n4836 ) ;
  assign n4838 = ( ~x281 & n4835 ) | ( ~x281 & n4836 ) | ( n4835 & n4836 ) ;
  assign n4839 = ( ~n656 & n4837 ) | ( ~n656 & n4838 ) | ( n4837 & n4838 ) ;
  assign n4840 = x344 & ~n991 ;
  assign n4841 = x344 & n995 ;
  assign n4842 = ( n1104 & n4840 ) | ( n1104 & n4841 ) | ( n4840 & n4841 ) ;
  assign n4843 = ( n1119 & n4840 ) | ( n1119 & n4841 ) | ( n4840 & n4841 ) ;
  assign n4844 = ( ~n1126 & n4840 ) | ( ~n1126 & n4841 ) | ( n4840 & n4841 ) ;
  assign n4845 = ( ~n1115 & n4843 ) | ( ~n1115 & n4844 ) | ( n4843 & n4844 ) ;
  assign n4846 = ( ~n975 & n4842 ) | ( ~n975 & n4845 ) | ( n4842 & n4845 ) ;
  assign n4847 = ( n1154 & n4842 ) | ( n1154 & n4845 ) | ( n4842 & n4845 ) ;
  assign n4848 = ( ~x409 & n4846 ) | ( ~x409 & n4847 ) | ( n4846 & n4847 ) ;
  assign n4849 = ( x281 & n4846 ) | ( x281 & n4847 ) | ( n4846 & n4847 ) ;
  assign n4850 = ( n656 & n4848 ) | ( n656 & n4849 ) | ( n4848 & n4849 ) ;
  assign n4851 = n4839 | n4850 ;
  assign n4852 = x216 & n1767 ;
  assign n4853 = x216 & ~n1771 ;
  assign n4854 = ( ~n1751 & n4852 ) | ( ~n1751 & n4853 ) | ( n4852 & n4853 ) ;
  assign n4855 = ( ~n1787 & n4852 ) | ( ~n1787 & n4853 ) | ( n4852 & n4853 ) ;
  assign n4856 = ( n1794 & n4852 ) | ( n1794 & n4853 ) | ( n4852 & n4853 ) ;
  assign n4857 = ( n1783 & n4855 ) | ( n1783 & n4856 ) | ( n4855 & n4856 ) ;
  assign n4858 = ( n1643 & n4854 ) | ( n1643 & n4857 ) | ( n4854 & n4857 ) ;
  assign n4859 = ( ~n1822 & n4854 ) | ( ~n1822 & n4857 ) | ( n4854 & n4857 ) ;
  assign n4860 = ( ~n1324 & n4858 ) | ( ~n1324 & n4859 ) | ( n4858 & n4859 ) ;
  assign n4861 = x88 & ~n1767 ;
  assign n4862 = x88 & n1771 ;
  assign n4863 = ( n1751 & n4861 ) | ( n1751 & n4862 ) | ( n4861 & n4862 ) ;
  assign n4864 = ( n1787 & n4861 ) | ( n1787 & n4862 ) | ( n4861 & n4862 ) ;
  assign n4865 = ( ~n1794 & n4861 ) | ( ~n1794 & n4862 ) | ( n4861 & n4862 ) ;
  assign n4866 = ( ~n1783 & n4864 ) | ( ~n1783 & n4865 ) | ( n4864 & n4865 ) ;
  assign n4867 = ( ~n1643 & n4863 ) | ( ~n1643 & n4866 ) | ( n4863 & n4866 ) ;
  assign n4868 = ( n1822 & n4863 ) | ( n1822 & n4866 ) | ( n4863 & n4866 ) ;
  assign n4869 = ( n1324 & n4867 ) | ( n1324 & n4868 ) | ( n4867 & n4868 ) ;
  assign n4870 = n4860 | n4869 ;
  assign n4871 = n4851 & ~n4870 ;
  assign n4872 = n4828 | n4871 ;
  assign n4873 = n4785 | n4872 ;
  assign n4874 = n4698 & ~n4873 ;
  assign n4875 = ~n4851 & n4870 ;
  assign n4876 = ( n4804 & ~n4827 ) | ( n4804 & n4875 ) | ( ~n4827 & n4875 ) ;
  assign n4877 = ~n4764 & n4783 ;
  assign n4878 = ~n4784 & n4877 ;
  assign n4879 = ( ~n4784 & n4876 ) | ( ~n4784 & n4878 ) | ( n4876 & n4878 ) ;
  assign n4880 = ( n4717 & ~n4740 ) | ( n4717 & n4879 ) | ( ~n4740 & n4879 ) ;
  assign n4881 = n4874 | n4880 ;
  assign n4882 = ~n4697 & n4881 ;
  assign n4883 = n4697 | n4873 ;
  assign n4884 = ( n4697 & ~n4880 ) | ( n4697 & n4883 ) | ( ~n4880 & n4883 ) ;
  assign n4885 = ( n4522 & ~n4882 ) | ( n4522 & n4884 ) | ( ~n4882 & n4884 ) ;
  assign n4886 = ~n4134 & n4157 ;
  assign n4887 = x486 & n991 ;
  assign n4888 = x486 & ~n995 ;
  assign n4889 = ( ~n1104 & n4887 ) | ( ~n1104 & n4888 ) | ( n4887 & n4888 ) ;
  assign n4890 = ( ~n1119 & n4887 ) | ( ~n1119 & n4888 ) | ( n4887 & n4888 ) ;
  assign n4891 = ( n1126 & n4887 ) | ( n1126 & n4888 ) | ( n4887 & n4888 ) ;
  assign n4892 = ( n1115 & n4890 ) | ( n1115 & n4891 ) | ( n4890 & n4891 ) ;
  assign n4893 = ( n975 & n4889 ) | ( n975 & n4892 ) | ( n4889 & n4892 ) ;
  assign n4894 = ( ~n1154 & n4889 ) | ( ~n1154 & n4892 ) | ( n4889 & n4892 ) ;
  assign n4895 = ( x409 & n4893 ) | ( x409 & n4894 ) | ( n4893 & n4894 ) ;
  assign n4896 = ( ~x281 & n4893 ) | ( ~x281 & n4894 ) | ( n4893 & n4894 ) ;
  assign n4897 = ( ~n656 & n4895 ) | ( ~n656 & n4896 ) | ( n4895 & n4896 ) ;
  assign n4898 = x358 & ~n991 ;
  assign n4899 = x358 & n995 ;
  assign n4900 = ( n1104 & n4898 ) | ( n1104 & n4899 ) | ( n4898 & n4899 ) ;
  assign n4901 = ( n1119 & n4898 ) | ( n1119 & n4899 ) | ( n4898 & n4899 ) ;
  assign n4902 = ( ~n1126 & n4898 ) | ( ~n1126 & n4899 ) | ( n4898 & n4899 ) ;
  assign n4903 = ( ~n1115 & n4901 ) | ( ~n1115 & n4902 ) | ( n4901 & n4902 ) ;
  assign n4904 = ( ~n975 & n4900 ) | ( ~n975 & n4903 ) | ( n4900 & n4903 ) ;
  assign n4905 = ( n1154 & n4900 ) | ( n1154 & n4903 ) | ( n4900 & n4903 ) ;
  assign n4906 = ( ~x409 & n4904 ) | ( ~x409 & n4905 ) | ( n4904 & n4905 ) ;
  assign n4907 = ( x281 & n4904 ) | ( x281 & n4905 ) | ( n4904 & n4905 ) ;
  assign n4908 = ( n656 & n4906 ) | ( n656 & n4907 ) | ( n4906 & n4907 ) ;
  assign n4909 = n4897 | n4908 ;
  assign n4910 = x230 & n1767 ;
  assign n4911 = x230 & ~n1771 ;
  assign n4912 = ( ~n1751 & n4910 ) | ( ~n1751 & n4911 ) | ( n4910 & n4911 ) ;
  assign n4913 = ( ~n1787 & n4910 ) | ( ~n1787 & n4911 ) | ( n4910 & n4911 ) ;
  assign n4914 = ( n1794 & n4910 ) | ( n1794 & n4911 ) | ( n4910 & n4911 ) ;
  assign n4915 = ( n1783 & n4913 ) | ( n1783 & n4914 ) | ( n4913 & n4914 ) ;
  assign n4916 = ( n1643 & n4912 ) | ( n1643 & n4915 ) | ( n4912 & n4915 ) ;
  assign n4917 = ( ~n1822 & n4912 ) | ( ~n1822 & n4915 ) | ( n4912 & n4915 ) ;
  assign n4918 = ( ~n1324 & n4916 ) | ( ~n1324 & n4917 ) | ( n4916 & n4917 ) ;
  assign n4919 = x102 & ~n1767 ;
  assign n4920 = x102 & n1771 ;
  assign n4921 = ( n1751 & n4919 ) | ( n1751 & n4920 ) | ( n4919 & n4920 ) ;
  assign n4922 = ( n1787 & n4919 ) | ( n1787 & n4920 ) | ( n4919 & n4920 ) ;
  assign n4923 = ( ~n1794 & n4919 ) | ( ~n1794 & n4920 ) | ( n4919 & n4920 ) ;
  assign n4924 = ( ~n1783 & n4922 ) | ( ~n1783 & n4923 ) | ( n4922 & n4923 ) ;
  assign n4925 = ( ~n1643 & n4921 ) | ( ~n1643 & n4924 ) | ( n4921 & n4924 ) ;
  assign n4926 = ( n1822 & n4921 ) | ( n1822 & n4924 ) | ( n4921 & n4924 ) ;
  assign n4927 = ( n1324 & n4925 ) | ( n1324 & n4926 ) | ( n4925 & n4926 ) ;
  assign n4928 = n4918 | n4927 ;
  assign n4929 = n4909 & ~n4928 ;
  assign n4930 = n4886 | n4929 ;
  assign n4931 = x229 & n1767 ;
  assign n4932 = x229 & ~n1771 ;
  assign n4933 = ( ~n1751 & n4931 ) | ( ~n1751 & n4932 ) | ( n4931 & n4932 ) ;
  assign n4934 = ( ~n1787 & n4931 ) | ( ~n1787 & n4932 ) | ( n4931 & n4932 ) ;
  assign n4935 = ( n1794 & n4931 ) | ( n1794 & n4932 ) | ( n4931 & n4932 ) ;
  assign n4936 = ( n1783 & n4934 ) | ( n1783 & n4935 ) | ( n4934 & n4935 ) ;
  assign n4937 = ( n1643 & n4933 ) | ( n1643 & n4936 ) | ( n4933 & n4936 ) ;
  assign n4938 = ( ~n1822 & n4933 ) | ( ~n1822 & n4936 ) | ( n4933 & n4936 ) ;
  assign n4939 = ( ~n1324 & n4937 ) | ( ~n1324 & n4938 ) | ( n4937 & n4938 ) ;
  assign n4940 = x101 & ~n1767 ;
  assign n4941 = x101 & n1771 ;
  assign n4942 = ( n1751 & n4940 ) | ( n1751 & n4941 ) | ( n4940 & n4941 ) ;
  assign n4943 = ( n1787 & n4940 ) | ( n1787 & n4941 ) | ( n4940 & n4941 ) ;
  assign n4944 = ( ~n1794 & n4940 ) | ( ~n1794 & n4941 ) | ( n4940 & n4941 ) ;
  assign n4945 = ( ~n1783 & n4943 ) | ( ~n1783 & n4944 ) | ( n4943 & n4944 ) ;
  assign n4946 = ( ~n1643 & n4942 ) | ( ~n1643 & n4945 ) | ( n4942 & n4945 ) ;
  assign n4947 = ( n1822 & n4942 ) | ( n1822 & n4945 ) | ( n4942 & n4945 ) ;
  assign n4948 = ( n1324 & n4946 ) | ( n1324 & n4947 ) | ( n4946 & n4947 ) ;
  assign n4949 = n4939 | n4948 ;
  assign n4950 = x485 & n991 ;
  assign n4951 = x485 & ~n995 ;
  assign n4952 = ( ~n1104 & n4950 ) | ( ~n1104 & n4951 ) | ( n4950 & n4951 ) ;
  assign n4953 = ( ~n1119 & n4950 ) | ( ~n1119 & n4951 ) | ( n4950 & n4951 ) ;
  assign n4954 = ( n1126 & n4950 ) | ( n1126 & n4951 ) | ( n4950 & n4951 ) ;
  assign n4955 = ( n1115 & n4953 ) | ( n1115 & n4954 ) | ( n4953 & n4954 ) ;
  assign n4956 = ( n975 & n4952 ) | ( n975 & n4955 ) | ( n4952 & n4955 ) ;
  assign n4957 = ( ~n1154 & n4952 ) | ( ~n1154 & n4955 ) | ( n4952 & n4955 ) ;
  assign n4958 = ( x409 & n4956 ) | ( x409 & n4957 ) | ( n4956 & n4957 ) ;
  assign n4959 = ( ~x281 & n4956 ) | ( ~x281 & n4957 ) | ( n4956 & n4957 ) ;
  assign n4960 = ( ~n656 & n4958 ) | ( ~n656 & n4959 ) | ( n4958 & n4959 ) ;
  assign n4961 = x357 & ~n991 ;
  assign n4962 = x357 & n995 ;
  assign n4963 = ( n1104 & n4961 ) | ( n1104 & n4962 ) | ( n4961 & n4962 ) ;
  assign n4964 = ( n1119 & n4961 ) | ( n1119 & n4962 ) | ( n4961 & n4962 ) ;
  assign n4965 = ( ~n1126 & n4961 ) | ( ~n1126 & n4962 ) | ( n4961 & n4962 ) ;
  assign n4966 = ( ~n1115 & n4964 ) | ( ~n1115 & n4965 ) | ( n4964 & n4965 ) ;
  assign n4967 = ( ~n975 & n4963 ) | ( ~n975 & n4966 ) | ( n4963 & n4966 ) ;
  assign n4968 = ( n1154 & n4963 ) | ( n1154 & n4966 ) | ( n4963 & n4966 ) ;
  assign n4969 = ( ~x409 & n4967 ) | ( ~x409 & n4968 ) | ( n4967 & n4968 ) ;
  assign n4970 = ( x281 & n4967 ) | ( x281 & n4968 ) | ( n4967 & n4968 ) ;
  assign n4971 = ( n656 & n4969 ) | ( n656 & n4970 ) | ( n4969 & n4970 ) ;
  assign n4972 = n4960 | n4971 ;
  assign n4973 = x228 & n1767 ;
  assign n4974 = x228 & ~n1771 ;
  assign n4975 = ( ~n1751 & n4973 ) | ( ~n1751 & n4974 ) | ( n4973 & n4974 ) ;
  assign n4976 = ( ~n1787 & n4973 ) | ( ~n1787 & n4974 ) | ( n4973 & n4974 ) ;
  assign n4977 = ( n1794 & n4973 ) | ( n1794 & n4974 ) | ( n4973 & n4974 ) ;
  assign n4978 = ( n1783 & n4976 ) | ( n1783 & n4977 ) | ( n4976 & n4977 ) ;
  assign n4979 = ( n1643 & n4975 ) | ( n1643 & n4978 ) | ( n4975 & n4978 ) ;
  assign n4980 = ( ~n1822 & n4975 ) | ( ~n1822 & n4978 ) | ( n4975 & n4978 ) ;
  assign n4981 = ( ~n1324 & n4979 ) | ( ~n1324 & n4980 ) | ( n4979 & n4980 ) ;
  assign n4982 = x100 & ~n1767 ;
  assign n4983 = x100 & n1771 ;
  assign n4984 = ( n1751 & n4982 ) | ( n1751 & n4983 ) | ( n4982 & n4983 ) ;
  assign n4985 = ( n1787 & n4982 ) | ( n1787 & n4983 ) | ( n4982 & n4983 ) ;
  assign n4986 = ( ~n1794 & n4982 ) | ( ~n1794 & n4983 ) | ( n4982 & n4983 ) ;
  assign n4987 = ( ~n1783 & n4985 ) | ( ~n1783 & n4986 ) | ( n4985 & n4986 ) ;
  assign n4988 = ( ~n1643 & n4984 ) | ( ~n1643 & n4987 ) | ( n4984 & n4987 ) ;
  assign n4989 = ( n1822 & n4984 ) | ( n1822 & n4987 ) | ( n4984 & n4987 ) ;
  assign n4990 = ( n1324 & n4988 ) | ( n1324 & n4989 ) | ( n4988 & n4989 ) ;
  assign n4991 = n4981 | n4990 ;
  assign n4992 = x484 & n991 ;
  assign n4993 = x484 & ~n995 ;
  assign n4994 = ( ~n1104 & n4992 ) | ( ~n1104 & n4993 ) | ( n4992 & n4993 ) ;
  assign n4995 = ( ~n1119 & n4992 ) | ( ~n1119 & n4993 ) | ( n4992 & n4993 ) ;
  assign n4996 = ( n1126 & n4992 ) | ( n1126 & n4993 ) | ( n4992 & n4993 ) ;
  assign n4997 = ( n1115 & n4995 ) | ( n1115 & n4996 ) | ( n4995 & n4996 ) ;
  assign n4998 = ( n975 & n4994 ) | ( n975 & n4997 ) | ( n4994 & n4997 ) ;
  assign n4999 = ( ~n1154 & n4994 ) | ( ~n1154 & n4997 ) | ( n4994 & n4997 ) ;
  assign n5000 = ( x409 & n4998 ) | ( x409 & n4999 ) | ( n4998 & n4999 ) ;
  assign n5001 = ( ~x281 & n4998 ) | ( ~x281 & n4999 ) | ( n4998 & n4999 ) ;
  assign n5002 = ( ~n656 & n5000 ) | ( ~n656 & n5001 ) | ( n5000 & n5001 ) ;
  assign n5003 = x356 & ~n991 ;
  assign n5004 = x356 & n995 ;
  assign n5005 = ( n1104 & n5003 ) | ( n1104 & n5004 ) | ( n5003 & n5004 ) ;
  assign n5006 = ( n1119 & n5003 ) | ( n1119 & n5004 ) | ( n5003 & n5004 ) ;
  assign n5007 = ( ~n1126 & n5003 ) | ( ~n1126 & n5004 ) | ( n5003 & n5004 ) ;
  assign n5008 = ( ~n1115 & n5006 ) | ( ~n1115 & n5007 ) | ( n5006 & n5007 ) ;
  assign n5009 = ( ~n975 & n5005 ) | ( ~n975 & n5008 ) | ( n5005 & n5008 ) ;
  assign n5010 = ( n1154 & n5005 ) | ( n1154 & n5008 ) | ( n5005 & n5008 ) ;
  assign n5011 = ( ~x409 & n5009 ) | ( ~x409 & n5010 ) | ( n5009 & n5010 ) ;
  assign n5012 = ( x281 & n5009 ) | ( x281 & n5010 ) | ( n5009 & n5010 ) ;
  assign n5013 = ( n656 & n5011 ) | ( n656 & n5012 ) | ( n5011 & n5012 ) ;
  assign n5014 = n5002 | n5013 ;
  assign n5015 = n4991 & ~n5014 ;
  assign n5016 = ( n4949 & ~n4972 ) | ( n4949 & n5015 ) | ( ~n4972 & n5015 ) ;
  assign n5017 = ~n4930 & n5016 ;
  assign n5018 = ~n4909 & n4928 ;
  assign n5019 = ~n4886 & n5018 ;
  assign n5020 = ~n4949 & n4972 ;
  assign n5021 = ~n4991 & n5014 ;
  assign n5022 = n5020 | n5021 ;
  assign n5023 = n4930 | n5022 ;
  assign n5024 = ~n5019 & n5023 ;
  assign n5025 = x227 & n1767 ;
  assign n5026 = x227 & ~n1771 ;
  assign n5027 = ( ~n1751 & n5025 ) | ( ~n1751 & n5026 ) | ( n5025 & n5026 ) ;
  assign n5028 = ( ~n1787 & n5025 ) | ( ~n1787 & n5026 ) | ( n5025 & n5026 ) ;
  assign n5029 = ( n1794 & n5025 ) | ( n1794 & n5026 ) | ( n5025 & n5026 ) ;
  assign n5030 = ( n1783 & n5028 ) | ( n1783 & n5029 ) | ( n5028 & n5029 ) ;
  assign n5031 = ( n1643 & n5027 ) | ( n1643 & n5030 ) | ( n5027 & n5030 ) ;
  assign n5032 = ( ~n1822 & n5027 ) | ( ~n1822 & n5030 ) | ( n5027 & n5030 ) ;
  assign n5033 = ( ~n1324 & n5031 ) | ( ~n1324 & n5032 ) | ( n5031 & n5032 ) ;
  assign n5034 = x99 & ~n1767 ;
  assign n5035 = x99 & n1771 ;
  assign n5036 = ( n1751 & n5034 ) | ( n1751 & n5035 ) | ( n5034 & n5035 ) ;
  assign n5037 = ( n1787 & n5034 ) | ( n1787 & n5035 ) | ( n5034 & n5035 ) ;
  assign n5038 = ( ~n1794 & n5034 ) | ( ~n1794 & n5035 ) | ( n5034 & n5035 ) ;
  assign n5039 = ( ~n1783 & n5037 ) | ( ~n1783 & n5038 ) | ( n5037 & n5038 ) ;
  assign n5040 = ( ~n1643 & n5036 ) | ( ~n1643 & n5039 ) | ( n5036 & n5039 ) ;
  assign n5041 = ( n1822 & n5036 ) | ( n1822 & n5039 ) | ( n5036 & n5039 ) ;
  assign n5042 = ( n1324 & n5040 ) | ( n1324 & n5041 ) | ( n5040 & n5041 ) ;
  assign n5043 = n5033 | n5042 ;
  assign n5044 = x483 & n991 ;
  assign n5045 = x483 & ~n995 ;
  assign n5046 = ( ~n1104 & n5044 ) | ( ~n1104 & n5045 ) | ( n5044 & n5045 ) ;
  assign n5047 = ( ~n1119 & n5044 ) | ( ~n1119 & n5045 ) | ( n5044 & n5045 ) ;
  assign n5048 = ( n1126 & n5044 ) | ( n1126 & n5045 ) | ( n5044 & n5045 ) ;
  assign n5049 = ( n1115 & n5047 ) | ( n1115 & n5048 ) | ( n5047 & n5048 ) ;
  assign n5050 = ( n975 & n5046 ) | ( n975 & n5049 ) | ( n5046 & n5049 ) ;
  assign n5051 = ( ~n1154 & n5046 ) | ( ~n1154 & n5049 ) | ( n5046 & n5049 ) ;
  assign n5052 = ( x409 & n5050 ) | ( x409 & n5051 ) | ( n5050 & n5051 ) ;
  assign n5053 = ( ~x281 & n5050 ) | ( ~x281 & n5051 ) | ( n5050 & n5051 ) ;
  assign n5054 = ( ~n656 & n5052 ) | ( ~n656 & n5053 ) | ( n5052 & n5053 ) ;
  assign n5055 = x355 & ~n991 ;
  assign n5056 = x355 & n995 ;
  assign n5057 = ( n1104 & n5055 ) | ( n1104 & n5056 ) | ( n5055 & n5056 ) ;
  assign n5058 = ( n1119 & n5055 ) | ( n1119 & n5056 ) | ( n5055 & n5056 ) ;
  assign n5059 = ( ~n1126 & n5055 ) | ( ~n1126 & n5056 ) | ( n5055 & n5056 ) ;
  assign n5060 = ( ~n1115 & n5058 ) | ( ~n1115 & n5059 ) | ( n5058 & n5059 ) ;
  assign n5061 = ( ~n975 & n5057 ) | ( ~n975 & n5060 ) | ( n5057 & n5060 ) ;
  assign n5062 = ( n1154 & n5057 ) | ( n1154 & n5060 ) | ( n5057 & n5060 ) ;
  assign n5063 = ( ~x409 & n5061 ) | ( ~x409 & n5062 ) | ( n5061 & n5062 ) ;
  assign n5064 = ( x281 & n5061 ) | ( x281 & n5062 ) | ( n5061 & n5062 ) ;
  assign n5065 = ( n656 & n5063 ) | ( n656 & n5064 ) | ( n5063 & n5064 ) ;
  assign n5066 = n5054 | n5065 ;
  assign n5067 = x482 & n991 ;
  assign n5068 = x482 & ~n995 ;
  assign n5069 = ( ~n1104 & n5067 ) | ( ~n1104 & n5068 ) | ( n5067 & n5068 ) ;
  assign n5070 = ( ~n1119 & n5067 ) | ( ~n1119 & n5068 ) | ( n5067 & n5068 ) ;
  assign n5071 = ( n1126 & n5067 ) | ( n1126 & n5068 ) | ( n5067 & n5068 ) ;
  assign n5072 = ( n1115 & n5070 ) | ( n1115 & n5071 ) | ( n5070 & n5071 ) ;
  assign n5073 = ( n975 & n5069 ) | ( n975 & n5072 ) | ( n5069 & n5072 ) ;
  assign n5074 = ( ~n1154 & n5069 ) | ( ~n1154 & n5072 ) | ( n5069 & n5072 ) ;
  assign n5075 = ( x409 & n5073 ) | ( x409 & n5074 ) | ( n5073 & n5074 ) ;
  assign n5076 = ( ~x281 & n5073 ) | ( ~x281 & n5074 ) | ( n5073 & n5074 ) ;
  assign n5077 = ( ~n656 & n5075 ) | ( ~n656 & n5076 ) | ( n5075 & n5076 ) ;
  assign n5078 = x354 & ~n991 ;
  assign n5079 = x354 & n995 ;
  assign n5080 = ( n1104 & n5078 ) | ( n1104 & n5079 ) | ( n5078 & n5079 ) ;
  assign n5081 = ( n1119 & n5078 ) | ( n1119 & n5079 ) | ( n5078 & n5079 ) ;
  assign n5082 = ( ~n1126 & n5078 ) | ( ~n1126 & n5079 ) | ( n5078 & n5079 ) ;
  assign n5083 = ( ~n1115 & n5081 ) | ( ~n1115 & n5082 ) | ( n5081 & n5082 ) ;
  assign n5084 = ( ~n975 & n5080 ) | ( ~n975 & n5083 ) | ( n5080 & n5083 ) ;
  assign n5085 = ( n1154 & n5080 ) | ( n1154 & n5083 ) | ( n5080 & n5083 ) ;
  assign n5086 = ( ~x409 & n5084 ) | ( ~x409 & n5085 ) | ( n5084 & n5085 ) ;
  assign n5087 = ( x281 & n5084 ) | ( x281 & n5085 ) | ( n5084 & n5085 ) ;
  assign n5088 = ( n656 & n5086 ) | ( n656 & n5087 ) | ( n5086 & n5087 ) ;
  assign n5089 = n5077 | n5088 ;
  assign n5090 = x226 & n1767 ;
  assign n5091 = x226 & ~n1771 ;
  assign n5092 = ( ~n1751 & n5090 ) | ( ~n1751 & n5091 ) | ( n5090 & n5091 ) ;
  assign n5093 = ( ~n1787 & n5090 ) | ( ~n1787 & n5091 ) | ( n5090 & n5091 ) ;
  assign n5094 = ( n1794 & n5090 ) | ( n1794 & n5091 ) | ( n5090 & n5091 ) ;
  assign n5095 = ( n1783 & n5093 ) | ( n1783 & n5094 ) | ( n5093 & n5094 ) ;
  assign n5096 = ( n1643 & n5092 ) | ( n1643 & n5095 ) | ( n5092 & n5095 ) ;
  assign n5097 = ( ~n1822 & n5092 ) | ( ~n1822 & n5095 ) | ( n5092 & n5095 ) ;
  assign n5098 = ( ~n1324 & n5096 ) | ( ~n1324 & n5097 ) | ( n5096 & n5097 ) ;
  assign n5099 = x98 & ~n1767 ;
  assign n5100 = x98 & n1771 ;
  assign n5101 = ( n1751 & n5099 ) | ( n1751 & n5100 ) | ( n5099 & n5100 ) ;
  assign n5102 = ( n1787 & n5099 ) | ( n1787 & n5100 ) | ( n5099 & n5100 ) ;
  assign n5103 = ( ~n1794 & n5099 ) | ( ~n1794 & n5100 ) | ( n5099 & n5100 ) ;
  assign n5104 = ( ~n1783 & n5102 ) | ( ~n1783 & n5103 ) | ( n5102 & n5103 ) ;
  assign n5105 = ( ~n1643 & n5101 ) | ( ~n1643 & n5104 ) | ( n5101 & n5104 ) ;
  assign n5106 = ( n1822 & n5101 ) | ( n1822 & n5104 ) | ( n5101 & n5104 ) ;
  assign n5107 = ( n1324 & n5105 ) | ( n1324 & n5106 ) | ( n5105 & n5106 ) ;
  assign n5108 = n5098 | n5107 ;
  assign n5109 = n5089 & ~n5108 ;
  assign n5110 = x225 & n1767 ;
  assign n5111 = x225 & ~n1771 ;
  assign n5112 = ( ~n1751 & n5110 ) | ( ~n1751 & n5111 ) | ( n5110 & n5111 ) ;
  assign n5113 = ( ~n1787 & n5110 ) | ( ~n1787 & n5111 ) | ( n5110 & n5111 ) ;
  assign n5114 = ( n1794 & n5110 ) | ( n1794 & n5111 ) | ( n5110 & n5111 ) ;
  assign n5115 = ( n1783 & n5113 ) | ( n1783 & n5114 ) | ( n5113 & n5114 ) ;
  assign n5116 = ( n1643 & n5112 ) | ( n1643 & n5115 ) | ( n5112 & n5115 ) ;
  assign n5117 = ( ~n1822 & n5112 ) | ( ~n1822 & n5115 ) | ( n5112 & n5115 ) ;
  assign n5118 = ( ~n1324 & n5116 ) | ( ~n1324 & n5117 ) | ( n5116 & n5117 ) ;
  assign n5119 = x97 & ~n1767 ;
  assign n5120 = x97 & n1771 ;
  assign n5121 = ( n1751 & n5119 ) | ( n1751 & n5120 ) | ( n5119 & n5120 ) ;
  assign n5122 = ( n1787 & n5119 ) | ( n1787 & n5120 ) | ( n5119 & n5120 ) ;
  assign n5123 = ( ~n1794 & n5119 ) | ( ~n1794 & n5120 ) | ( n5119 & n5120 ) ;
  assign n5124 = ( ~n1783 & n5122 ) | ( ~n1783 & n5123 ) | ( n5122 & n5123 ) ;
  assign n5125 = ( ~n1643 & n5121 ) | ( ~n1643 & n5124 ) | ( n5121 & n5124 ) ;
  assign n5126 = ( n1822 & n5121 ) | ( n1822 & n5124 ) | ( n5121 & n5124 ) ;
  assign n5127 = ( n1324 & n5125 ) | ( n1324 & n5126 ) | ( n5125 & n5126 ) ;
  assign n5128 = n5118 | n5127 ;
  assign n5129 = x481 & n991 ;
  assign n5130 = x481 & ~n995 ;
  assign n5131 = ( ~n1104 & n5129 ) | ( ~n1104 & n5130 ) | ( n5129 & n5130 ) ;
  assign n5132 = ( ~n1119 & n5129 ) | ( ~n1119 & n5130 ) | ( n5129 & n5130 ) ;
  assign n5133 = ( n1126 & n5129 ) | ( n1126 & n5130 ) | ( n5129 & n5130 ) ;
  assign n5134 = ( n1115 & n5132 ) | ( n1115 & n5133 ) | ( n5132 & n5133 ) ;
  assign n5135 = ( n975 & n5131 ) | ( n975 & n5134 ) | ( n5131 & n5134 ) ;
  assign n5136 = ( ~n1154 & n5131 ) | ( ~n1154 & n5134 ) | ( n5131 & n5134 ) ;
  assign n5137 = ( x409 & n5135 ) | ( x409 & n5136 ) | ( n5135 & n5136 ) ;
  assign n5138 = ( ~x281 & n5135 ) | ( ~x281 & n5136 ) | ( n5135 & n5136 ) ;
  assign n5139 = ( ~n656 & n5137 ) | ( ~n656 & n5138 ) | ( n5137 & n5138 ) ;
  assign n5140 = x353 & ~n991 ;
  assign n5141 = x353 & n995 ;
  assign n5142 = ( n1104 & n5140 ) | ( n1104 & n5141 ) | ( n5140 & n5141 ) ;
  assign n5143 = ( n1119 & n5140 ) | ( n1119 & n5141 ) | ( n5140 & n5141 ) ;
  assign n5144 = ( ~n1126 & n5140 ) | ( ~n1126 & n5141 ) | ( n5140 & n5141 ) ;
  assign n5145 = ( ~n1115 & n5143 ) | ( ~n1115 & n5144 ) | ( n5143 & n5144 ) ;
  assign n5146 = ( ~n975 & n5142 ) | ( ~n975 & n5145 ) | ( n5142 & n5145 ) ;
  assign n5147 = ( n1154 & n5142 ) | ( n1154 & n5145 ) | ( n5142 & n5145 ) ;
  assign n5148 = ( ~x409 & n5146 ) | ( ~x409 & n5147 ) | ( n5146 & n5147 ) ;
  assign n5149 = ( x281 & n5146 ) | ( x281 & n5147 ) | ( n5146 & n5147 ) ;
  assign n5150 = ( n656 & n5148 ) | ( n656 & n5149 ) | ( n5148 & n5149 ) ;
  assign n5151 = n5139 | n5150 ;
  assign n5152 = x480 & n991 ;
  assign n5153 = x480 & ~n995 ;
  assign n5154 = ( ~n1104 & n5152 ) | ( ~n1104 & n5153 ) | ( n5152 & n5153 ) ;
  assign n5155 = ( ~n1119 & n5152 ) | ( ~n1119 & n5153 ) | ( n5152 & n5153 ) ;
  assign n5156 = ( n1126 & n5152 ) | ( n1126 & n5153 ) | ( n5152 & n5153 ) ;
  assign n5157 = ( n1115 & n5155 ) | ( n1115 & n5156 ) | ( n5155 & n5156 ) ;
  assign n5158 = ( n975 & n5154 ) | ( n975 & n5157 ) | ( n5154 & n5157 ) ;
  assign n5159 = ( ~n1154 & n5154 ) | ( ~n1154 & n5157 ) | ( n5154 & n5157 ) ;
  assign n5160 = ( x409 & n5158 ) | ( x409 & n5159 ) | ( n5158 & n5159 ) ;
  assign n5161 = ( ~x281 & n5158 ) | ( ~x281 & n5159 ) | ( n5158 & n5159 ) ;
  assign n5162 = ( ~n656 & n5160 ) | ( ~n656 & n5161 ) | ( n5160 & n5161 ) ;
  assign n5163 = x352 & ~n991 ;
  assign n5164 = x352 & n995 ;
  assign n5165 = ( n1104 & n5163 ) | ( n1104 & n5164 ) | ( n5163 & n5164 ) ;
  assign n5166 = ( n1119 & n5163 ) | ( n1119 & n5164 ) | ( n5163 & n5164 ) ;
  assign n5167 = ( ~n1126 & n5163 ) | ( ~n1126 & n5164 ) | ( n5163 & n5164 ) ;
  assign n5168 = ( ~n1115 & n5166 ) | ( ~n1115 & n5167 ) | ( n5166 & n5167 ) ;
  assign n5169 = ( ~n975 & n5165 ) | ( ~n975 & n5168 ) | ( n5165 & n5168 ) ;
  assign n5170 = ( n1154 & n5165 ) | ( n1154 & n5168 ) | ( n5165 & n5168 ) ;
  assign n5171 = ( ~x409 & n5169 ) | ( ~x409 & n5170 ) | ( n5169 & n5170 ) ;
  assign n5172 = ( x281 & n5169 ) | ( x281 & n5170 ) | ( n5169 & n5170 ) ;
  assign n5173 = ( n656 & n5171 ) | ( n656 & n5172 ) | ( n5171 & n5172 ) ;
  assign n5174 = n5162 | n5173 ;
  assign n5175 = x224 & n1767 ;
  assign n5176 = x224 & ~n1771 ;
  assign n5177 = ( ~n1751 & n5175 ) | ( ~n1751 & n5176 ) | ( n5175 & n5176 ) ;
  assign n5178 = ( ~n1787 & n5175 ) | ( ~n1787 & n5176 ) | ( n5175 & n5176 ) ;
  assign n5179 = ( n1794 & n5175 ) | ( n1794 & n5176 ) | ( n5175 & n5176 ) ;
  assign n5180 = ( n1783 & n5178 ) | ( n1783 & n5179 ) | ( n5178 & n5179 ) ;
  assign n5181 = ( n1643 & n5177 ) | ( n1643 & n5180 ) | ( n5177 & n5180 ) ;
  assign n5182 = ( ~n1822 & n5177 ) | ( ~n1822 & n5180 ) | ( n5177 & n5180 ) ;
  assign n5183 = ( ~n1324 & n5181 ) | ( ~n1324 & n5182 ) | ( n5181 & n5182 ) ;
  assign n5184 = x96 & ~n1767 ;
  assign n5185 = x96 & n1771 ;
  assign n5186 = ( n1751 & n5184 ) | ( n1751 & n5185 ) | ( n5184 & n5185 ) ;
  assign n5187 = ( n1787 & n5184 ) | ( n1787 & n5185 ) | ( n5184 & n5185 ) ;
  assign n5188 = ( ~n1794 & n5184 ) | ( ~n1794 & n5185 ) | ( n5184 & n5185 ) ;
  assign n5189 = ( ~n1783 & n5187 ) | ( ~n1783 & n5188 ) | ( n5187 & n5188 ) ;
  assign n5190 = ( ~n1643 & n5186 ) | ( ~n1643 & n5189 ) | ( n5186 & n5189 ) ;
  assign n5191 = ( n1822 & n5186 ) | ( n1822 & n5189 ) | ( n5186 & n5189 ) ;
  assign n5192 = ( n1324 & n5190 ) | ( n1324 & n5191 ) | ( n5190 & n5191 ) ;
  assign n5193 = n5183 | n5192 ;
  assign n5194 = ~n5174 & n5193 ;
  assign n5195 = ( n5128 & ~n5151 ) | ( n5128 & n5194 ) | ( ~n5151 & n5194 ) ;
  assign n5196 = ~n5089 & n5108 ;
  assign n5197 = ~n5109 & n5196 ;
  assign n5198 = ( ~n5109 & n5195 ) | ( ~n5109 & n5197 ) | ( n5195 & n5197 ) ;
  assign n5199 = ( n5043 & ~n5066 ) | ( n5043 & n5198 ) | ( ~n5066 & n5198 ) ;
  assign n5200 = ( n5019 & ~n5024 ) | ( n5019 & n5199 ) | ( ~n5024 & n5199 ) ;
  assign n5201 = n5017 | n5200 ;
  assign n5202 = ~n5128 & n5151 ;
  assign n5203 = n4541 & ~n4564 ;
  assign n5204 = ~n5202 & n5203 ;
  assign n5205 = n4671 & ~n4694 ;
  assign n5206 = ( n4588 & ~n4607 ) | ( n4588 & n4651 ) | ( ~n4607 & n4651 ) ;
  assign n5207 = ( ~n4588 & n4607 ) | ( ~n4588 & n4628 ) | ( n4607 & n4628 ) ;
  assign n5208 = ( n5205 & ~n5206 ) | ( n5205 & n5207 ) | ( ~n5206 & n5207 ) ;
  assign n5209 = ~n4565 & n5208 ;
  assign n5210 = ( ~n5202 & n5204 ) | ( ~n5202 & n5209 ) | ( n5204 & n5209 ) ;
  assign n5211 = ~n5043 & n5066 ;
  assign n5212 = n5109 | n5211 ;
  assign n5213 = n5174 & ~n5193 ;
  assign n5214 = n5212 | n5213 ;
  assign n5215 = n5023 | n5214 ;
  assign n5216 = ( n5023 & ~n5199 ) | ( n5023 & n5215 ) | ( ~n5199 & n5215 ) ;
  assign n5217 = n5017 | n5019 ;
  assign n5218 = n5216 & ~n5217 ;
  assign n5219 = ( n5201 & n5210 ) | ( n5201 & ~n5218 ) | ( n5210 & ~n5218 ) ;
  assign n5220 = ( ~n5201 & n5202 ) | ( ~n5201 & n5218 ) | ( n5202 & n5218 ) ;
  assign n5221 = ( n4885 & ~n5219 ) | ( n4885 & n5220 ) | ( ~n5219 & n5220 ) ;
  assign n5222 = ( n4115 & ~n4159 ) | ( n4115 & n5221 ) | ( ~n4159 & n5221 ) ;
  assign n5223 = n4334 & ~n4517 ;
  assign n5224 = ( n4514 & n4517 ) | ( n4514 & ~n5223 ) | ( n4517 & ~n5223 ) ;
  assign n5225 = n4246 & ~n4698 ;
  assign n5226 = ( n4520 & n4698 ) | ( n4520 & ~n5225 ) | ( n4698 & ~n5225 ) ;
  assign n5227 = n5224 | n5226 ;
  assign n5228 = ( n4884 & n5202 ) | ( n4884 & ~n5210 ) | ( n5202 & ~n5210 ) ;
  assign n5229 = ~n4697 & n4880 ;
  assign n5230 = ( ~n5202 & n5210 ) | ( ~n5202 & n5229 ) | ( n5210 & n5229 ) ;
  assign n5231 = ( n5227 & ~n5228 ) | ( n5227 & n5230 ) | ( ~n5228 & n5230 ) ;
  assign n5232 = n4115 & ~n4159 ;
  assign n5233 = ( ~n4115 & n4159 ) | ( ~n4115 & n5017 ) | ( n4159 & n5017 ) ;
  assign n5234 = ( n5200 & ~n5232 ) | ( n5200 & n5233 ) | ( ~n5232 & n5233 ) ;
  assign n5235 = ( ~n4115 & n4159 ) | ( ~n4115 & n5217 ) | ( n4159 & n5217 ) ;
  assign n5236 = ( n5216 & n5232 ) | ( n5216 & ~n5235 ) | ( n5232 & ~n5235 ) ;
  assign n5237 = ( n5231 & n5234 ) | ( n5231 & ~n5236 ) | ( n5234 & ~n5236 ) ;
  assign n5238 = ~n4485 & n4508 ;
  assign n5239 = x191 & n1767 ;
  assign n5240 = x191 & ~n1771 ;
  assign n5241 = ( ~n1751 & n5239 ) | ( ~n1751 & n5240 ) | ( n5239 & n5240 ) ;
  assign n5242 = ( ~n1787 & n5239 ) | ( ~n1787 & n5240 ) | ( n5239 & n5240 ) ;
  assign n5243 = ( n1794 & n5239 ) | ( n1794 & n5240 ) | ( n5239 & n5240 ) ;
  assign n5244 = ( n1783 & n5242 ) | ( n1783 & n5243 ) | ( n5242 & n5243 ) ;
  assign n5245 = ( n1643 & n5241 ) | ( n1643 & n5244 ) | ( n5241 & n5244 ) ;
  assign n5246 = ( ~n1822 & n5241 ) | ( ~n1822 & n5244 ) | ( n5241 & n5244 ) ;
  assign n5247 = ( ~n1324 & n5245 ) | ( ~n1324 & n5246 ) | ( n5245 & n5246 ) ;
  assign n5248 = x63 & ~n1767 ;
  assign n5249 = x63 & n1771 ;
  assign n5250 = ( n1751 & n5248 ) | ( n1751 & n5249 ) | ( n5248 & n5249 ) ;
  assign n5251 = ( n1787 & n5248 ) | ( n1787 & n5249 ) | ( n5248 & n5249 ) ;
  assign n5252 = ( ~n1794 & n5248 ) | ( ~n1794 & n5249 ) | ( n5248 & n5249 ) ;
  assign n5253 = ( ~n1783 & n5251 ) | ( ~n1783 & n5252 ) | ( n5251 & n5252 ) ;
  assign n5254 = ( ~n1643 & n5250 ) | ( ~n1643 & n5253 ) | ( n5250 & n5253 ) ;
  assign n5255 = ( n1822 & n5250 ) | ( n1822 & n5253 ) | ( n5250 & n5253 ) ;
  assign n5256 = ( n1324 & n5254 ) | ( n1324 & n5255 ) | ( n5254 & n5255 ) ;
  assign n5257 = n5247 | n5256 ;
  assign n5258 = x447 & n991 ;
  assign n5259 = x447 & ~n995 ;
  assign n5260 = ( ~n1104 & n5258 ) | ( ~n1104 & n5259 ) | ( n5258 & n5259 ) ;
  assign n5261 = ( ~n1119 & n5258 ) | ( ~n1119 & n5259 ) | ( n5258 & n5259 ) ;
  assign n5262 = ( n1126 & n5258 ) | ( n1126 & n5259 ) | ( n5258 & n5259 ) ;
  assign n5263 = ( n1115 & n5261 ) | ( n1115 & n5262 ) | ( n5261 & n5262 ) ;
  assign n5264 = ( n975 & n5260 ) | ( n975 & n5263 ) | ( n5260 & n5263 ) ;
  assign n5265 = ( ~n1154 & n5260 ) | ( ~n1154 & n5263 ) | ( n5260 & n5263 ) ;
  assign n5266 = ( x409 & n5264 ) | ( x409 & n5265 ) | ( n5264 & n5265 ) ;
  assign n5267 = ( ~x281 & n5264 ) | ( ~x281 & n5265 ) | ( n5264 & n5265 ) ;
  assign n5268 = ( ~n656 & n5266 ) | ( ~n656 & n5267 ) | ( n5266 & n5267 ) ;
  assign n5269 = x319 & ~n991 ;
  assign n5270 = x319 & n995 ;
  assign n5271 = ( n1104 & n5269 ) | ( n1104 & n5270 ) | ( n5269 & n5270 ) ;
  assign n5272 = ( n1119 & n5269 ) | ( n1119 & n5270 ) | ( n5269 & n5270 ) ;
  assign n5273 = ( ~n1126 & n5269 ) | ( ~n1126 & n5270 ) | ( n5269 & n5270 ) ;
  assign n5274 = ( ~n1115 & n5272 ) | ( ~n1115 & n5273 ) | ( n5272 & n5273 ) ;
  assign n5275 = ( ~n975 & n5271 ) | ( ~n975 & n5274 ) | ( n5271 & n5274 ) ;
  assign n5276 = ( n1154 & n5271 ) | ( n1154 & n5274 ) | ( n5271 & n5274 ) ;
  assign n5277 = ( ~x409 & n5275 ) | ( ~x409 & n5276 ) | ( n5275 & n5276 ) ;
  assign n5278 = ( x281 & n5275 ) | ( x281 & n5276 ) | ( n5275 & n5276 ) ;
  assign n5279 = ( n656 & n5277 ) | ( n656 & n5278 ) | ( n5277 & n5278 ) ;
  assign n5280 = n5268 | n5279 ;
  assign n5281 = ~n5257 & n5280 ;
  assign n5282 = x446 & n991 ;
  assign n5283 = x446 & ~n995 ;
  assign n5284 = ( ~n1104 & n5282 ) | ( ~n1104 & n5283 ) | ( n5282 & n5283 ) ;
  assign n5285 = ( ~n1119 & n5282 ) | ( ~n1119 & n5283 ) | ( n5282 & n5283 ) ;
  assign n5286 = ( n1126 & n5282 ) | ( n1126 & n5283 ) | ( n5282 & n5283 ) ;
  assign n5287 = ( n1115 & n5285 ) | ( n1115 & n5286 ) | ( n5285 & n5286 ) ;
  assign n5288 = ( n975 & n5284 ) | ( n975 & n5287 ) | ( n5284 & n5287 ) ;
  assign n5289 = ( ~n1154 & n5284 ) | ( ~n1154 & n5287 ) | ( n5284 & n5287 ) ;
  assign n5290 = ( x409 & n5288 ) | ( x409 & n5289 ) | ( n5288 & n5289 ) ;
  assign n5291 = ( ~x281 & n5288 ) | ( ~x281 & n5289 ) | ( n5288 & n5289 ) ;
  assign n5292 = ( ~n656 & n5290 ) | ( ~n656 & n5291 ) | ( n5290 & n5291 ) ;
  assign n5293 = x318 & ~n991 ;
  assign n5294 = x318 & n995 ;
  assign n5295 = ( n1104 & n5293 ) | ( n1104 & n5294 ) | ( n5293 & n5294 ) ;
  assign n5296 = ( n1119 & n5293 ) | ( n1119 & n5294 ) | ( n5293 & n5294 ) ;
  assign n5297 = ( ~n1126 & n5293 ) | ( ~n1126 & n5294 ) | ( n5293 & n5294 ) ;
  assign n5298 = ( ~n1115 & n5296 ) | ( ~n1115 & n5297 ) | ( n5296 & n5297 ) ;
  assign n5299 = ( ~n975 & n5295 ) | ( ~n975 & n5298 ) | ( n5295 & n5298 ) ;
  assign n5300 = ( n1154 & n5295 ) | ( n1154 & n5298 ) | ( n5295 & n5298 ) ;
  assign n5301 = ( ~x409 & n5299 ) | ( ~x409 & n5300 ) | ( n5299 & n5300 ) ;
  assign n5302 = ( x281 & n5299 ) | ( x281 & n5300 ) | ( n5299 & n5300 ) ;
  assign n5303 = ( n656 & n5301 ) | ( n656 & n5302 ) | ( n5301 & n5302 ) ;
  assign n5304 = n5292 | n5303 ;
  assign n5305 = x190 & n1767 ;
  assign n5306 = x190 & ~n1771 ;
  assign n5307 = ( ~n1751 & n5305 ) | ( ~n1751 & n5306 ) | ( n5305 & n5306 ) ;
  assign n5308 = ( ~n1787 & n5305 ) | ( ~n1787 & n5306 ) | ( n5305 & n5306 ) ;
  assign n5309 = ( n1794 & n5305 ) | ( n1794 & n5306 ) | ( n5305 & n5306 ) ;
  assign n5310 = ( n1783 & n5308 ) | ( n1783 & n5309 ) | ( n5308 & n5309 ) ;
  assign n5311 = ( n1643 & n5307 ) | ( n1643 & n5310 ) | ( n5307 & n5310 ) ;
  assign n5312 = ( ~n1822 & n5307 ) | ( ~n1822 & n5310 ) | ( n5307 & n5310 ) ;
  assign n5313 = ( ~n1324 & n5311 ) | ( ~n1324 & n5312 ) | ( n5311 & n5312 ) ;
  assign n5314 = x62 & ~n1767 ;
  assign n5315 = x62 & n1771 ;
  assign n5316 = ( n1751 & n5314 ) | ( n1751 & n5315 ) | ( n5314 & n5315 ) ;
  assign n5317 = ( n1787 & n5314 ) | ( n1787 & n5315 ) | ( n5314 & n5315 ) ;
  assign n5318 = ( ~n1794 & n5314 ) | ( ~n1794 & n5315 ) | ( n5314 & n5315 ) ;
  assign n5319 = ( ~n1783 & n5317 ) | ( ~n1783 & n5318 ) | ( n5317 & n5318 ) ;
  assign n5320 = ( ~n1643 & n5316 ) | ( ~n1643 & n5319 ) | ( n5316 & n5319 ) ;
  assign n5321 = ( n1822 & n5316 ) | ( n1822 & n5319 ) | ( n5316 & n5319 ) ;
  assign n5322 = ( n1324 & n5320 ) | ( n1324 & n5321 ) | ( n5320 & n5321 ) ;
  assign n5323 = n5313 | n5322 ;
  assign n5324 = n5304 & ~n5323 ;
  assign n5325 = n5281 | n5324 ;
  assign n5326 = x189 & n1767 ;
  assign n5327 = x189 & ~n1771 ;
  assign n5328 = ( ~n1751 & n5326 ) | ( ~n1751 & n5327 ) | ( n5326 & n5327 ) ;
  assign n5329 = ( ~n1787 & n5326 ) | ( ~n1787 & n5327 ) | ( n5326 & n5327 ) ;
  assign n5330 = ( n1794 & n5326 ) | ( n1794 & n5327 ) | ( n5326 & n5327 ) ;
  assign n5331 = ( n1783 & n5329 ) | ( n1783 & n5330 ) | ( n5329 & n5330 ) ;
  assign n5332 = ( n1643 & n5328 ) | ( n1643 & n5331 ) | ( n5328 & n5331 ) ;
  assign n5333 = ( ~n1822 & n5328 ) | ( ~n1822 & n5331 ) | ( n5328 & n5331 ) ;
  assign n5334 = ( ~n1324 & n5332 ) | ( ~n1324 & n5333 ) | ( n5332 & n5333 ) ;
  assign n5335 = x61 & ~n1767 ;
  assign n5336 = x61 & n1771 ;
  assign n5337 = ( n1751 & n5335 ) | ( n1751 & n5336 ) | ( n5335 & n5336 ) ;
  assign n5338 = ( n1787 & n5335 ) | ( n1787 & n5336 ) | ( n5335 & n5336 ) ;
  assign n5339 = ( ~n1794 & n5335 ) | ( ~n1794 & n5336 ) | ( n5335 & n5336 ) ;
  assign n5340 = ( ~n1783 & n5338 ) | ( ~n1783 & n5339 ) | ( n5338 & n5339 ) ;
  assign n5341 = ( ~n1643 & n5337 ) | ( ~n1643 & n5340 ) | ( n5337 & n5340 ) ;
  assign n5342 = ( n1822 & n5337 ) | ( n1822 & n5340 ) | ( n5337 & n5340 ) ;
  assign n5343 = ( n1324 & n5341 ) | ( n1324 & n5342 ) | ( n5341 & n5342 ) ;
  assign n5344 = n5334 | n5343 ;
  assign n5345 = x445 & n991 ;
  assign n5346 = x445 & ~n995 ;
  assign n5347 = ( ~n1104 & n5345 ) | ( ~n1104 & n5346 ) | ( n5345 & n5346 ) ;
  assign n5348 = ( ~n1119 & n5345 ) | ( ~n1119 & n5346 ) | ( n5345 & n5346 ) ;
  assign n5349 = ( n1126 & n5345 ) | ( n1126 & n5346 ) | ( n5345 & n5346 ) ;
  assign n5350 = ( n1115 & n5348 ) | ( n1115 & n5349 ) | ( n5348 & n5349 ) ;
  assign n5351 = ( n975 & n5347 ) | ( n975 & n5350 ) | ( n5347 & n5350 ) ;
  assign n5352 = ( ~n1154 & n5347 ) | ( ~n1154 & n5350 ) | ( n5347 & n5350 ) ;
  assign n5353 = ( x409 & n5351 ) | ( x409 & n5352 ) | ( n5351 & n5352 ) ;
  assign n5354 = ( ~x281 & n5351 ) | ( ~x281 & n5352 ) | ( n5351 & n5352 ) ;
  assign n5355 = ( ~n656 & n5353 ) | ( ~n656 & n5354 ) | ( n5353 & n5354 ) ;
  assign n5356 = x317 & ~n991 ;
  assign n5357 = x317 & n995 ;
  assign n5358 = ( n1104 & n5356 ) | ( n1104 & n5357 ) | ( n5356 & n5357 ) ;
  assign n5359 = ( n1119 & n5356 ) | ( n1119 & n5357 ) | ( n5356 & n5357 ) ;
  assign n5360 = ( ~n1126 & n5356 ) | ( ~n1126 & n5357 ) | ( n5356 & n5357 ) ;
  assign n5361 = ( ~n1115 & n5359 ) | ( ~n1115 & n5360 ) | ( n5359 & n5360 ) ;
  assign n5362 = ( ~n975 & n5358 ) | ( ~n975 & n5361 ) | ( n5358 & n5361 ) ;
  assign n5363 = ( n1154 & n5358 ) | ( n1154 & n5361 ) | ( n5358 & n5361 ) ;
  assign n5364 = ( ~x409 & n5362 ) | ( ~x409 & n5363 ) | ( n5362 & n5363 ) ;
  assign n5365 = ( x281 & n5362 ) | ( x281 & n5363 ) | ( n5362 & n5363 ) ;
  assign n5366 = ( n656 & n5364 ) | ( n656 & n5365 ) | ( n5364 & n5365 ) ;
  assign n5367 = n5355 | n5366 ;
  assign n5368 = ~n5344 & n5367 ;
  assign n5369 = x188 & n1767 ;
  assign n5370 = x188 & ~n1771 ;
  assign n5371 = ( ~n1751 & n5369 ) | ( ~n1751 & n5370 ) | ( n5369 & n5370 ) ;
  assign n5372 = ( ~n1787 & n5369 ) | ( ~n1787 & n5370 ) | ( n5369 & n5370 ) ;
  assign n5373 = ( n1794 & n5369 ) | ( n1794 & n5370 ) | ( n5369 & n5370 ) ;
  assign n5374 = ( n1783 & n5372 ) | ( n1783 & n5373 ) | ( n5372 & n5373 ) ;
  assign n5375 = ( n1643 & n5371 ) | ( n1643 & n5374 ) | ( n5371 & n5374 ) ;
  assign n5376 = ( ~n1822 & n5371 ) | ( ~n1822 & n5374 ) | ( n5371 & n5374 ) ;
  assign n5377 = ( ~n1324 & n5375 ) | ( ~n1324 & n5376 ) | ( n5375 & n5376 ) ;
  assign n5378 = x60 & ~n1767 ;
  assign n5379 = x60 & n1771 ;
  assign n5380 = ( n1751 & n5378 ) | ( n1751 & n5379 ) | ( n5378 & n5379 ) ;
  assign n5381 = ( n1787 & n5378 ) | ( n1787 & n5379 ) | ( n5378 & n5379 ) ;
  assign n5382 = ( ~n1794 & n5378 ) | ( ~n1794 & n5379 ) | ( n5378 & n5379 ) ;
  assign n5383 = ( ~n1783 & n5381 ) | ( ~n1783 & n5382 ) | ( n5381 & n5382 ) ;
  assign n5384 = ( ~n1643 & n5380 ) | ( ~n1643 & n5383 ) | ( n5380 & n5383 ) ;
  assign n5385 = ( n1822 & n5380 ) | ( n1822 & n5383 ) | ( n5380 & n5383 ) ;
  assign n5386 = ( n1324 & n5384 ) | ( n1324 & n5385 ) | ( n5384 & n5385 ) ;
  assign n5387 = n5377 | n5386 ;
  assign n5388 = x444 & n991 ;
  assign n5389 = x444 & ~n995 ;
  assign n5390 = ( ~n1104 & n5388 ) | ( ~n1104 & n5389 ) | ( n5388 & n5389 ) ;
  assign n5391 = ( ~n1119 & n5388 ) | ( ~n1119 & n5389 ) | ( n5388 & n5389 ) ;
  assign n5392 = ( n1126 & n5388 ) | ( n1126 & n5389 ) | ( n5388 & n5389 ) ;
  assign n5393 = ( n1115 & n5391 ) | ( n1115 & n5392 ) | ( n5391 & n5392 ) ;
  assign n5394 = ( n975 & n5390 ) | ( n975 & n5393 ) | ( n5390 & n5393 ) ;
  assign n5395 = ( ~n1154 & n5390 ) | ( ~n1154 & n5393 ) | ( n5390 & n5393 ) ;
  assign n5396 = ( x409 & n5394 ) | ( x409 & n5395 ) | ( n5394 & n5395 ) ;
  assign n5397 = ( ~x281 & n5394 ) | ( ~x281 & n5395 ) | ( n5394 & n5395 ) ;
  assign n5398 = ( ~n656 & n5396 ) | ( ~n656 & n5397 ) | ( n5396 & n5397 ) ;
  assign n5399 = x316 & ~n991 ;
  assign n5400 = x316 & n995 ;
  assign n5401 = ( n1104 & n5399 ) | ( n1104 & n5400 ) | ( n5399 & n5400 ) ;
  assign n5402 = ( n1119 & n5399 ) | ( n1119 & n5400 ) | ( n5399 & n5400 ) ;
  assign n5403 = ( ~n1126 & n5399 ) | ( ~n1126 & n5400 ) | ( n5399 & n5400 ) ;
  assign n5404 = ( ~n1115 & n5402 ) | ( ~n1115 & n5403 ) | ( n5402 & n5403 ) ;
  assign n5405 = ( ~n975 & n5401 ) | ( ~n975 & n5404 ) | ( n5401 & n5404 ) ;
  assign n5406 = ( n1154 & n5401 ) | ( n1154 & n5404 ) | ( n5401 & n5404 ) ;
  assign n5407 = ( ~x409 & n5405 ) | ( ~x409 & n5406 ) | ( n5405 & n5406 ) ;
  assign n5408 = ( x281 & n5405 ) | ( x281 & n5406 ) | ( n5405 & n5406 ) ;
  assign n5409 = ( n656 & n5407 ) | ( n656 & n5408 ) | ( n5407 & n5408 ) ;
  assign n5410 = n5398 | n5409 ;
  assign n5411 = ~n5387 & n5410 ;
  assign n5412 = n5368 | n5411 ;
  assign n5413 = n5325 | n5412 ;
  assign n5414 = x187 & n1767 ;
  assign n5415 = x187 & ~n1771 ;
  assign n5416 = ( ~n1751 & n5414 ) | ( ~n1751 & n5415 ) | ( n5414 & n5415 ) ;
  assign n5417 = ( ~n1787 & n5414 ) | ( ~n1787 & n5415 ) | ( n5414 & n5415 ) ;
  assign n5418 = ( n1794 & n5414 ) | ( n1794 & n5415 ) | ( n5414 & n5415 ) ;
  assign n5419 = ( n1783 & n5417 ) | ( n1783 & n5418 ) | ( n5417 & n5418 ) ;
  assign n5420 = ( n1643 & n5416 ) | ( n1643 & n5419 ) | ( n5416 & n5419 ) ;
  assign n5421 = ( ~n1822 & n5416 ) | ( ~n1822 & n5419 ) | ( n5416 & n5419 ) ;
  assign n5422 = ( ~n1324 & n5420 ) | ( ~n1324 & n5421 ) | ( n5420 & n5421 ) ;
  assign n5423 = x59 & ~n1767 ;
  assign n5424 = x59 & n1771 ;
  assign n5425 = ( n1751 & n5423 ) | ( n1751 & n5424 ) | ( n5423 & n5424 ) ;
  assign n5426 = ( n1787 & n5423 ) | ( n1787 & n5424 ) | ( n5423 & n5424 ) ;
  assign n5427 = ( ~n1794 & n5423 ) | ( ~n1794 & n5424 ) | ( n5423 & n5424 ) ;
  assign n5428 = ( ~n1783 & n5426 ) | ( ~n1783 & n5427 ) | ( n5426 & n5427 ) ;
  assign n5429 = ( ~n1643 & n5425 ) | ( ~n1643 & n5428 ) | ( n5425 & n5428 ) ;
  assign n5430 = ( n1822 & n5425 ) | ( n1822 & n5428 ) | ( n5425 & n5428 ) ;
  assign n5431 = ( n1324 & n5429 ) | ( n1324 & n5430 ) | ( n5429 & n5430 ) ;
  assign n5432 = n5422 | n5431 ;
  assign n5433 = x443 & n991 ;
  assign n5434 = x443 & ~n995 ;
  assign n5435 = ( ~n1104 & n5433 ) | ( ~n1104 & n5434 ) | ( n5433 & n5434 ) ;
  assign n5436 = ( ~n1119 & n5433 ) | ( ~n1119 & n5434 ) | ( n5433 & n5434 ) ;
  assign n5437 = ( n1126 & n5433 ) | ( n1126 & n5434 ) | ( n5433 & n5434 ) ;
  assign n5438 = ( n1115 & n5436 ) | ( n1115 & n5437 ) | ( n5436 & n5437 ) ;
  assign n5439 = ( n975 & n5435 ) | ( n975 & n5438 ) | ( n5435 & n5438 ) ;
  assign n5440 = ( ~n1154 & n5435 ) | ( ~n1154 & n5438 ) | ( n5435 & n5438 ) ;
  assign n5441 = ( x409 & n5439 ) | ( x409 & n5440 ) | ( n5439 & n5440 ) ;
  assign n5442 = ( ~x281 & n5439 ) | ( ~x281 & n5440 ) | ( n5439 & n5440 ) ;
  assign n5443 = ( ~n656 & n5441 ) | ( ~n656 & n5442 ) | ( n5441 & n5442 ) ;
  assign n5444 = x315 & ~n991 ;
  assign n5445 = x315 & n995 ;
  assign n5446 = ( n1104 & n5444 ) | ( n1104 & n5445 ) | ( n5444 & n5445 ) ;
  assign n5447 = ( n1119 & n5444 ) | ( n1119 & n5445 ) | ( n5444 & n5445 ) ;
  assign n5448 = ( ~n1126 & n5444 ) | ( ~n1126 & n5445 ) | ( n5444 & n5445 ) ;
  assign n5449 = ( ~n1115 & n5447 ) | ( ~n1115 & n5448 ) | ( n5447 & n5448 ) ;
  assign n5450 = ( ~n975 & n5446 ) | ( ~n975 & n5449 ) | ( n5446 & n5449 ) ;
  assign n5451 = ( n1154 & n5446 ) | ( n1154 & n5449 ) | ( n5446 & n5449 ) ;
  assign n5452 = ( ~x409 & n5450 ) | ( ~x409 & n5451 ) | ( n5450 & n5451 ) ;
  assign n5453 = ( x281 & n5450 ) | ( x281 & n5451 ) | ( n5450 & n5451 ) ;
  assign n5454 = ( n656 & n5452 ) | ( n656 & n5453 ) | ( n5452 & n5453 ) ;
  assign n5455 = n5443 | n5454 ;
  assign n5456 = ~n5432 & n5455 ;
  assign n5457 = x186 & n1767 ;
  assign n5458 = x186 & ~n1771 ;
  assign n5459 = ( ~n1751 & n5457 ) | ( ~n1751 & n5458 ) | ( n5457 & n5458 ) ;
  assign n5460 = ( ~n1787 & n5457 ) | ( ~n1787 & n5458 ) | ( n5457 & n5458 ) ;
  assign n5461 = ( n1794 & n5457 ) | ( n1794 & n5458 ) | ( n5457 & n5458 ) ;
  assign n5462 = ( n1783 & n5460 ) | ( n1783 & n5461 ) | ( n5460 & n5461 ) ;
  assign n5463 = ( n1643 & n5459 ) | ( n1643 & n5462 ) | ( n5459 & n5462 ) ;
  assign n5464 = ( ~n1822 & n5459 ) | ( ~n1822 & n5462 ) | ( n5459 & n5462 ) ;
  assign n5465 = ( ~n1324 & n5463 ) | ( ~n1324 & n5464 ) | ( n5463 & n5464 ) ;
  assign n5466 = x58 & ~n1767 ;
  assign n5467 = x58 & n1771 ;
  assign n5468 = ( n1751 & n5466 ) | ( n1751 & n5467 ) | ( n5466 & n5467 ) ;
  assign n5469 = ( n1787 & n5466 ) | ( n1787 & n5467 ) | ( n5466 & n5467 ) ;
  assign n5470 = ( ~n1794 & n5466 ) | ( ~n1794 & n5467 ) | ( n5466 & n5467 ) ;
  assign n5471 = ( ~n1783 & n5469 ) | ( ~n1783 & n5470 ) | ( n5469 & n5470 ) ;
  assign n5472 = ( ~n1643 & n5468 ) | ( ~n1643 & n5471 ) | ( n5468 & n5471 ) ;
  assign n5473 = ( n1822 & n5468 ) | ( n1822 & n5471 ) | ( n5468 & n5471 ) ;
  assign n5474 = ( n1324 & n5472 ) | ( n1324 & n5473 ) | ( n5472 & n5473 ) ;
  assign n5475 = n5465 | n5474 ;
  assign n5476 = x442 & n991 ;
  assign n5477 = x442 & ~n995 ;
  assign n5478 = ( ~n1104 & n5476 ) | ( ~n1104 & n5477 ) | ( n5476 & n5477 ) ;
  assign n5479 = ( ~n1119 & n5476 ) | ( ~n1119 & n5477 ) | ( n5476 & n5477 ) ;
  assign n5480 = ( n1126 & n5476 ) | ( n1126 & n5477 ) | ( n5476 & n5477 ) ;
  assign n5481 = ( n1115 & n5479 ) | ( n1115 & n5480 ) | ( n5479 & n5480 ) ;
  assign n5482 = ( n975 & n5478 ) | ( n975 & n5481 ) | ( n5478 & n5481 ) ;
  assign n5483 = ( ~n1154 & n5478 ) | ( ~n1154 & n5481 ) | ( n5478 & n5481 ) ;
  assign n5484 = ( x409 & n5482 ) | ( x409 & n5483 ) | ( n5482 & n5483 ) ;
  assign n5485 = ( ~x281 & n5482 ) | ( ~x281 & n5483 ) | ( n5482 & n5483 ) ;
  assign n5486 = ( ~n656 & n5484 ) | ( ~n656 & n5485 ) | ( n5484 & n5485 ) ;
  assign n5487 = x314 & ~n991 ;
  assign n5488 = x314 & n995 ;
  assign n5489 = ( n1104 & n5487 ) | ( n1104 & n5488 ) | ( n5487 & n5488 ) ;
  assign n5490 = ( n1119 & n5487 ) | ( n1119 & n5488 ) | ( n5487 & n5488 ) ;
  assign n5491 = ( ~n1126 & n5487 ) | ( ~n1126 & n5488 ) | ( n5487 & n5488 ) ;
  assign n5492 = ( ~n1115 & n5490 ) | ( ~n1115 & n5491 ) | ( n5490 & n5491 ) ;
  assign n5493 = ( ~n975 & n5489 ) | ( ~n975 & n5492 ) | ( n5489 & n5492 ) ;
  assign n5494 = ( n1154 & n5489 ) | ( n1154 & n5492 ) | ( n5489 & n5492 ) ;
  assign n5495 = ( ~x409 & n5493 ) | ( ~x409 & n5494 ) | ( n5493 & n5494 ) ;
  assign n5496 = ( x281 & n5493 ) | ( x281 & n5494 ) | ( n5493 & n5494 ) ;
  assign n5497 = ( n656 & n5495 ) | ( n656 & n5496 ) | ( n5495 & n5496 ) ;
  assign n5498 = n5486 | n5497 ;
  assign n5499 = ~n5475 & n5498 ;
  assign n5500 = n5456 | n5499 ;
  assign n5501 = x185 & n1767 ;
  assign n5502 = x185 & ~n1771 ;
  assign n5503 = ( ~n1751 & n5501 ) | ( ~n1751 & n5502 ) | ( n5501 & n5502 ) ;
  assign n5504 = ( ~n1787 & n5501 ) | ( ~n1787 & n5502 ) | ( n5501 & n5502 ) ;
  assign n5505 = ( n1794 & n5501 ) | ( n1794 & n5502 ) | ( n5501 & n5502 ) ;
  assign n5506 = ( n1783 & n5504 ) | ( n1783 & n5505 ) | ( n5504 & n5505 ) ;
  assign n5507 = ( n1643 & n5503 ) | ( n1643 & n5506 ) | ( n5503 & n5506 ) ;
  assign n5508 = ( ~n1822 & n5503 ) | ( ~n1822 & n5506 ) | ( n5503 & n5506 ) ;
  assign n5509 = ( ~n1324 & n5507 ) | ( ~n1324 & n5508 ) | ( n5507 & n5508 ) ;
  assign n5510 = x57 & ~n1767 ;
  assign n5511 = x57 & n1771 ;
  assign n5512 = ( n1751 & n5510 ) | ( n1751 & n5511 ) | ( n5510 & n5511 ) ;
  assign n5513 = ( n1787 & n5510 ) | ( n1787 & n5511 ) | ( n5510 & n5511 ) ;
  assign n5514 = ( ~n1794 & n5510 ) | ( ~n1794 & n5511 ) | ( n5510 & n5511 ) ;
  assign n5515 = ( ~n1783 & n5513 ) | ( ~n1783 & n5514 ) | ( n5513 & n5514 ) ;
  assign n5516 = ( ~n1643 & n5512 ) | ( ~n1643 & n5515 ) | ( n5512 & n5515 ) ;
  assign n5517 = ( n1822 & n5512 ) | ( n1822 & n5515 ) | ( n5512 & n5515 ) ;
  assign n5518 = ( n1324 & n5516 ) | ( n1324 & n5517 ) | ( n5516 & n5517 ) ;
  assign n5519 = n5509 | n5518 ;
  assign n5520 = x441 & n991 ;
  assign n5521 = x441 & ~n995 ;
  assign n5522 = ( ~n1104 & n5520 ) | ( ~n1104 & n5521 ) | ( n5520 & n5521 ) ;
  assign n5523 = ( ~n1119 & n5520 ) | ( ~n1119 & n5521 ) | ( n5520 & n5521 ) ;
  assign n5524 = ( n1126 & n5520 ) | ( n1126 & n5521 ) | ( n5520 & n5521 ) ;
  assign n5525 = ( n1115 & n5523 ) | ( n1115 & n5524 ) | ( n5523 & n5524 ) ;
  assign n5526 = ( n975 & n5522 ) | ( n975 & n5525 ) | ( n5522 & n5525 ) ;
  assign n5527 = ( ~n1154 & n5522 ) | ( ~n1154 & n5525 ) | ( n5522 & n5525 ) ;
  assign n5528 = ( x409 & n5526 ) | ( x409 & n5527 ) | ( n5526 & n5527 ) ;
  assign n5529 = ( ~x281 & n5526 ) | ( ~x281 & n5527 ) | ( n5526 & n5527 ) ;
  assign n5530 = ( ~n656 & n5528 ) | ( ~n656 & n5529 ) | ( n5528 & n5529 ) ;
  assign n5531 = x313 & ~n991 ;
  assign n5532 = x313 & n995 ;
  assign n5533 = ( n1104 & n5531 ) | ( n1104 & n5532 ) | ( n5531 & n5532 ) ;
  assign n5534 = ( n1119 & n5531 ) | ( n1119 & n5532 ) | ( n5531 & n5532 ) ;
  assign n5535 = ( ~n1126 & n5531 ) | ( ~n1126 & n5532 ) | ( n5531 & n5532 ) ;
  assign n5536 = ( ~n1115 & n5534 ) | ( ~n1115 & n5535 ) | ( n5534 & n5535 ) ;
  assign n5537 = ( ~n975 & n5533 ) | ( ~n975 & n5536 ) | ( n5533 & n5536 ) ;
  assign n5538 = ( n1154 & n5533 ) | ( n1154 & n5536 ) | ( n5533 & n5536 ) ;
  assign n5539 = ( ~x409 & n5537 ) | ( ~x409 & n5538 ) | ( n5537 & n5538 ) ;
  assign n5540 = ( x281 & n5537 ) | ( x281 & n5538 ) | ( n5537 & n5538 ) ;
  assign n5541 = ( n656 & n5539 ) | ( n656 & n5540 ) | ( n5539 & n5540 ) ;
  assign n5542 = n5530 | n5541 ;
  assign n5543 = ~n5519 & n5542 ;
  assign n5544 = x184 & n1767 ;
  assign n5545 = x184 & ~n1771 ;
  assign n5546 = ( ~n1751 & n5544 ) | ( ~n1751 & n5545 ) | ( n5544 & n5545 ) ;
  assign n5547 = ( ~n1787 & n5544 ) | ( ~n1787 & n5545 ) | ( n5544 & n5545 ) ;
  assign n5548 = ( n1794 & n5544 ) | ( n1794 & n5545 ) | ( n5544 & n5545 ) ;
  assign n5549 = ( n1783 & n5547 ) | ( n1783 & n5548 ) | ( n5547 & n5548 ) ;
  assign n5550 = ( n1643 & n5546 ) | ( n1643 & n5549 ) | ( n5546 & n5549 ) ;
  assign n5551 = ( ~n1822 & n5546 ) | ( ~n1822 & n5549 ) | ( n5546 & n5549 ) ;
  assign n5552 = ( ~n1324 & n5550 ) | ( ~n1324 & n5551 ) | ( n5550 & n5551 ) ;
  assign n5553 = x56 & ~n1767 ;
  assign n5554 = x56 & n1771 ;
  assign n5555 = ( n1751 & n5553 ) | ( n1751 & n5554 ) | ( n5553 & n5554 ) ;
  assign n5556 = ( n1787 & n5553 ) | ( n1787 & n5554 ) | ( n5553 & n5554 ) ;
  assign n5557 = ( ~n1794 & n5553 ) | ( ~n1794 & n5554 ) | ( n5553 & n5554 ) ;
  assign n5558 = ( ~n1783 & n5556 ) | ( ~n1783 & n5557 ) | ( n5556 & n5557 ) ;
  assign n5559 = ( ~n1643 & n5555 ) | ( ~n1643 & n5558 ) | ( n5555 & n5558 ) ;
  assign n5560 = ( n1822 & n5555 ) | ( n1822 & n5558 ) | ( n5555 & n5558 ) ;
  assign n5561 = ( n1324 & n5559 ) | ( n1324 & n5560 ) | ( n5559 & n5560 ) ;
  assign n5562 = n5552 | n5561 ;
  assign n5563 = x440 & n991 ;
  assign n5564 = x440 & ~n995 ;
  assign n5565 = ( ~n1104 & n5563 ) | ( ~n1104 & n5564 ) | ( n5563 & n5564 ) ;
  assign n5566 = ( ~n1119 & n5563 ) | ( ~n1119 & n5564 ) | ( n5563 & n5564 ) ;
  assign n5567 = ( n1126 & n5563 ) | ( n1126 & n5564 ) | ( n5563 & n5564 ) ;
  assign n5568 = ( n1115 & n5566 ) | ( n1115 & n5567 ) | ( n5566 & n5567 ) ;
  assign n5569 = ( n975 & n5565 ) | ( n975 & n5568 ) | ( n5565 & n5568 ) ;
  assign n5570 = ( ~n1154 & n5565 ) | ( ~n1154 & n5568 ) | ( n5565 & n5568 ) ;
  assign n5571 = ( x409 & n5569 ) | ( x409 & n5570 ) | ( n5569 & n5570 ) ;
  assign n5572 = ( ~x281 & n5569 ) | ( ~x281 & n5570 ) | ( n5569 & n5570 ) ;
  assign n5573 = ( ~n656 & n5571 ) | ( ~n656 & n5572 ) | ( n5571 & n5572 ) ;
  assign n5574 = x312 & ~n991 ;
  assign n5575 = x312 & n995 ;
  assign n5576 = ( n1104 & n5574 ) | ( n1104 & n5575 ) | ( n5574 & n5575 ) ;
  assign n5577 = ( n1119 & n5574 ) | ( n1119 & n5575 ) | ( n5574 & n5575 ) ;
  assign n5578 = ( ~n1126 & n5574 ) | ( ~n1126 & n5575 ) | ( n5574 & n5575 ) ;
  assign n5579 = ( ~n1115 & n5577 ) | ( ~n1115 & n5578 ) | ( n5577 & n5578 ) ;
  assign n5580 = ( ~n975 & n5576 ) | ( ~n975 & n5579 ) | ( n5576 & n5579 ) ;
  assign n5581 = ( n1154 & n5576 ) | ( n1154 & n5579 ) | ( n5576 & n5579 ) ;
  assign n5582 = ( ~x409 & n5580 ) | ( ~x409 & n5581 ) | ( n5580 & n5581 ) ;
  assign n5583 = ( x281 & n5580 ) | ( x281 & n5581 ) | ( n5580 & n5581 ) ;
  assign n5584 = ( n656 & n5582 ) | ( n656 & n5583 ) | ( n5582 & n5583 ) ;
  assign n5585 = n5573 | n5584 ;
  assign n5586 = ~n5562 & n5585 ;
  assign n5587 = n5543 | n5586 ;
  assign n5588 = n5500 | n5587 ;
  assign n5589 = n5413 | n5588 ;
  assign n5590 = n5387 & ~n5410 ;
  assign n5591 = ( n5344 & ~n5367 ) | ( n5344 & n5590 ) | ( ~n5367 & n5590 ) ;
  assign n5592 = ~n5325 & n5591 ;
  assign n5593 = ~n5304 & n5323 ;
  assign n5594 = ~n5281 & n5593 ;
  assign n5595 = n5592 | n5594 ;
  assign n5596 = n5589 & ~n5595 ;
  assign n5597 = n5257 & ~n5280 ;
  assign n5598 = n5562 & ~n5585 ;
  assign n5599 = ( n5519 & ~n5542 ) | ( n5519 & n5598 ) | ( ~n5542 & n5598 ) ;
  assign n5600 = n5475 & ~n5498 ;
  assign n5601 = ~n5499 & n5600 ;
  assign n5602 = ( ~n5499 & n5599 ) | ( ~n5499 & n5601 ) | ( n5599 & n5601 ) ;
  assign n5603 = ( n5432 & ~n5455 ) | ( n5432 & n5602 ) | ( ~n5455 & n5602 ) ;
  assign n5604 = n5413 & ~n5597 ;
  assign n5605 = ( n5597 & n5603 ) | ( n5597 & ~n5604 ) | ( n5603 & ~n5604 ) ;
  assign n5606 = n5596 & ~n5605 ;
  assign n5607 = x199 & n1767 ;
  assign n5608 = x199 & ~n1771 ;
  assign n5609 = ( ~n1751 & n5607 ) | ( ~n1751 & n5608 ) | ( n5607 & n5608 ) ;
  assign n5610 = ( ~n1787 & n5607 ) | ( ~n1787 & n5608 ) | ( n5607 & n5608 ) ;
  assign n5611 = ( n1794 & n5607 ) | ( n1794 & n5608 ) | ( n5607 & n5608 ) ;
  assign n5612 = ( n1783 & n5610 ) | ( n1783 & n5611 ) | ( n5610 & n5611 ) ;
  assign n5613 = ( n1643 & n5609 ) | ( n1643 & n5612 ) | ( n5609 & n5612 ) ;
  assign n5614 = ( ~n1822 & n5609 ) | ( ~n1822 & n5612 ) | ( n5609 & n5612 ) ;
  assign n5615 = ( ~n1324 & n5613 ) | ( ~n1324 & n5614 ) | ( n5613 & n5614 ) ;
  assign n5616 = x71 & ~n1767 ;
  assign n5617 = x71 & n1771 ;
  assign n5618 = ( n1751 & n5616 ) | ( n1751 & n5617 ) | ( n5616 & n5617 ) ;
  assign n5619 = ( n1787 & n5616 ) | ( n1787 & n5617 ) | ( n5616 & n5617 ) ;
  assign n5620 = ( ~n1794 & n5616 ) | ( ~n1794 & n5617 ) | ( n5616 & n5617 ) ;
  assign n5621 = ( ~n1783 & n5619 ) | ( ~n1783 & n5620 ) | ( n5619 & n5620 ) ;
  assign n5622 = ( ~n1643 & n5618 ) | ( ~n1643 & n5621 ) | ( n5618 & n5621 ) ;
  assign n5623 = ( n1822 & n5618 ) | ( n1822 & n5621 ) | ( n5618 & n5621 ) ;
  assign n5624 = ( n1324 & n5622 ) | ( n1324 & n5623 ) | ( n5622 & n5623 ) ;
  assign n5625 = n5615 | n5624 ;
  assign n5626 = x455 & n991 ;
  assign n5627 = x455 & ~n995 ;
  assign n5628 = ( ~n1104 & n5626 ) | ( ~n1104 & n5627 ) | ( n5626 & n5627 ) ;
  assign n5629 = ( ~n1119 & n5626 ) | ( ~n1119 & n5627 ) | ( n5626 & n5627 ) ;
  assign n5630 = ( n1126 & n5626 ) | ( n1126 & n5627 ) | ( n5626 & n5627 ) ;
  assign n5631 = ( n1115 & n5629 ) | ( n1115 & n5630 ) | ( n5629 & n5630 ) ;
  assign n5632 = ( n975 & n5628 ) | ( n975 & n5631 ) | ( n5628 & n5631 ) ;
  assign n5633 = ( ~n1154 & n5628 ) | ( ~n1154 & n5631 ) | ( n5628 & n5631 ) ;
  assign n5634 = ( x409 & n5632 ) | ( x409 & n5633 ) | ( n5632 & n5633 ) ;
  assign n5635 = ( ~x281 & n5632 ) | ( ~x281 & n5633 ) | ( n5632 & n5633 ) ;
  assign n5636 = ( ~n656 & n5634 ) | ( ~n656 & n5635 ) | ( n5634 & n5635 ) ;
  assign n5637 = x327 & ~n991 ;
  assign n5638 = x327 & n995 ;
  assign n5639 = ( n1104 & n5637 ) | ( n1104 & n5638 ) | ( n5637 & n5638 ) ;
  assign n5640 = ( n1119 & n5637 ) | ( n1119 & n5638 ) | ( n5637 & n5638 ) ;
  assign n5641 = ( ~n1126 & n5637 ) | ( ~n1126 & n5638 ) | ( n5637 & n5638 ) ;
  assign n5642 = ( ~n1115 & n5640 ) | ( ~n1115 & n5641 ) | ( n5640 & n5641 ) ;
  assign n5643 = ( ~n975 & n5639 ) | ( ~n975 & n5642 ) | ( n5639 & n5642 ) ;
  assign n5644 = ( n1154 & n5639 ) | ( n1154 & n5642 ) | ( n5639 & n5642 ) ;
  assign n5645 = ( ~x409 & n5643 ) | ( ~x409 & n5644 ) | ( n5643 & n5644 ) ;
  assign n5646 = ( x281 & n5643 ) | ( x281 & n5644 ) | ( n5643 & n5644 ) ;
  assign n5647 = ( n656 & n5645 ) | ( n656 & n5646 ) | ( n5645 & n5646 ) ;
  assign n5648 = n5636 | n5647 ;
  assign n5649 = ~n5625 & n5648 ;
  assign n5650 = x454 & n991 ;
  assign n5651 = x454 & ~n995 ;
  assign n5652 = ( ~n1104 & n5650 ) | ( ~n1104 & n5651 ) | ( n5650 & n5651 ) ;
  assign n5653 = ( ~n1119 & n5650 ) | ( ~n1119 & n5651 ) | ( n5650 & n5651 ) ;
  assign n5654 = ( n1126 & n5650 ) | ( n1126 & n5651 ) | ( n5650 & n5651 ) ;
  assign n5655 = ( n1115 & n5653 ) | ( n1115 & n5654 ) | ( n5653 & n5654 ) ;
  assign n5656 = ( n975 & n5652 ) | ( n975 & n5655 ) | ( n5652 & n5655 ) ;
  assign n5657 = ( ~n1154 & n5652 ) | ( ~n1154 & n5655 ) | ( n5652 & n5655 ) ;
  assign n5658 = ( x409 & n5656 ) | ( x409 & n5657 ) | ( n5656 & n5657 ) ;
  assign n5659 = ( ~x281 & n5656 ) | ( ~x281 & n5657 ) | ( n5656 & n5657 ) ;
  assign n5660 = ( ~n656 & n5658 ) | ( ~n656 & n5659 ) | ( n5658 & n5659 ) ;
  assign n5661 = x326 & ~n991 ;
  assign n5662 = x326 & n995 ;
  assign n5663 = ( n1104 & n5661 ) | ( n1104 & n5662 ) | ( n5661 & n5662 ) ;
  assign n5664 = ( n1119 & n5661 ) | ( n1119 & n5662 ) | ( n5661 & n5662 ) ;
  assign n5665 = ( ~n1126 & n5661 ) | ( ~n1126 & n5662 ) | ( n5661 & n5662 ) ;
  assign n5666 = ( ~n1115 & n5664 ) | ( ~n1115 & n5665 ) | ( n5664 & n5665 ) ;
  assign n5667 = ( ~n975 & n5663 ) | ( ~n975 & n5666 ) | ( n5663 & n5666 ) ;
  assign n5668 = ( n1154 & n5663 ) | ( n1154 & n5666 ) | ( n5663 & n5666 ) ;
  assign n5669 = ( ~x409 & n5667 ) | ( ~x409 & n5668 ) | ( n5667 & n5668 ) ;
  assign n5670 = ( x281 & n5667 ) | ( x281 & n5668 ) | ( n5667 & n5668 ) ;
  assign n5671 = ( n656 & n5669 ) | ( n656 & n5670 ) | ( n5669 & n5670 ) ;
  assign n5672 = n5660 | n5671 ;
  assign n5673 = x198 & n1767 ;
  assign n5674 = x198 & ~n1771 ;
  assign n5675 = ( ~n1751 & n5673 ) | ( ~n1751 & n5674 ) | ( n5673 & n5674 ) ;
  assign n5676 = ( ~n1787 & n5673 ) | ( ~n1787 & n5674 ) | ( n5673 & n5674 ) ;
  assign n5677 = ( n1794 & n5673 ) | ( n1794 & n5674 ) | ( n5673 & n5674 ) ;
  assign n5678 = ( n1783 & n5676 ) | ( n1783 & n5677 ) | ( n5676 & n5677 ) ;
  assign n5679 = ( n1643 & n5675 ) | ( n1643 & n5678 ) | ( n5675 & n5678 ) ;
  assign n5680 = ( ~n1822 & n5675 ) | ( ~n1822 & n5678 ) | ( n5675 & n5678 ) ;
  assign n5681 = ( ~n1324 & n5679 ) | ( ~n1324 & n5680 ) | ( n5679 & n5680 ) ;
  assign n5682 = x70 & ~n1767 ;
  assign n5683 = x70 & n1771 ;
  assign n5684 = ( n1751 & n5682 ) | ( n1751 & n5683 ) | ( n5682 & n5683 ) ;
  assign n5685 = ( n1787 & n5682 ) | ( n1787 & n5683 ) | ( n5682 & n5683 ) ;
  assign n5686 = ( ~n1794 & n5682 ) | ( ~n1794 & n5683 ) | ( n5682 & n5683 ) ;
  assign n5687 = ( ~n1783 & n5685 ) | ( ~n1783 & n5686 ) | ( n5685 & n5686 ) ;
  assign n5688 = ( ~n1643 & n5684 ) | ( ~n1643 & n5687 ) | ( n5684 & n5687 ) ;
  assign n5689 = ( n1822 & n5684 ) | ( n1822 & n5687 ) | ( n5684 & n5687 ) ;
  assign n5690 = ( n1324 & n5688 ) | ( n1324 & n5689 ) | ( n5688 & n5689 ) ;
  assign n5691 = n5681 | n5690 ;
  assign n5692 = ~n5672 & n5691 ;
  assign n5693 = ~n5649 & n5692 ;
  assign n5694 = n5672 & ~n5691 ;
  assign n5695 = n5649 | n5694 ;
  assign n5696 = x197 & n1767 ;
  assign n5697 = x197 & ~n1771 ;
  assign n5698 = ( ~n1751 & n5696 ) | ( ~n1751 & n5697 ) | ( n5696 & n5697 ) ;
  assign n5699 = ( ~n1787 & n5696 ) | ( ~n1787 & n5697 ) | ( n5696 & n5697 ) ;
  assign n5700 = ( n1794 & n5696 ) | ( n1794 & n5697 ) | ( n5696 & n5697 ) ;
  assign n5701 = ( n1783 & n5699 ) | ( n1783 & n5700 ) | ( n5699 & n5700 ) ;
  assign n5702 = ( n1643 & n5698 ) | ( n1643 & n5701 ) | ( n5698 & n5701 ) ;
  assign n5703 = ( ~n1822 & n5698 ) | ( ~n1822 & n5701 ) | ( n5698 & n5701 ) ;
  assign n5704 = ( ~n1324 & n5702 ) | ( ~n1324 & n5703 ) | ( n5702 & n5703 ) ;
  assign n5705 = x69 & ~n1767 ;
  assign n5706 = x69 & n1771 ;
  assign n5707 = ( n1751 & n5705 ) | ( n1751 & n5706 ) | ( n5705 & n5706 ) ;
  assign n5708 = ( n1787 & n5705 ) | ( n1787 & n5706 ) | ( n5705 & n5706 ) ;
  assign n5709 = ( ~n1794 & n5705 ) | ( ~n1794 & n5706 ) | ( n5705 & n5706 ) ;
  assign n5710 = ( ~n1783 & n5708 ) | ( ~n1783 & n5709 ) | ( n5708 & n5709 ) ;
  assign n5711 = ( ~n1643 & n5707 ) | ( ~n1643 & n5710 ) | ( n5707 & n5710 ) ;
  assign n5712 = ( n1822 & n5707 ) | ( n1822 & n5710 ) | ( n5707 & n5710 ) ;
  assign n5713 = ( n1324 & n5711 ) | ( n1324 & n5712 ) | ( n5711 & n5712 ) ;
  assign n5714 = n5704 | n5713 ;
  assign n5715 = x453 & n991 ;
  assign n5716 = x453 & ~n995 ;
  assign n5717 = ( ~n1104 & n5715 ) | ( ~n1104 & n5716 ) | ( n5715 & n5716 ) ;
  assign n5718 = ( ~n1119 & n5715 ) | ( ~n1119 & n5716 ) | ( n5715 & n5716 ) ;
  assign n5719 = ( n1126 & n5715 ) | ( n1126 & n5716 ) | ( n5715 & n5716 ) ;
  assign n5720 = ( n1115 & n5718 ) | ( n1115 & n5719 ) | ( n5718 & n5719 ) ;
  assign n5721 = ( n975 & n5717 ) | ( n975 & n5720 ) | ( n5717 & n5720 ) ;
  assign n5722 = ( ~n1154 & n5717 ) | ( ~n1154 & n5720 ) | ( n5717 & n5720 ) ;
  assign n5723 = ( x409 & n5721 ) | ( x409 & n5722 ) | ( n5721 & n5722 ) ;
  assign n5724 = ( ~x281 & n5721 ) | ( ~x281 & n5722 ) | ( n5721 & n5722 ) ;
  assign n5725 = ( ~n656 & n5723 ) | ( ~n656 & n5724 ) | ( n5723 & n5724 ) ;
  assign n5726 = x325 & ~n991 ;
  assign n5727 = x325 & n995 ;
  assign n5728 = ( n1104 & n5726 ) | ( n1104 & n5727 ) | ( n5726 & n5727 ) ;
  assign n5729 = ( n1119 & n5726 ) | ( n1119 & n5727 ) | ( n5726 & n5727 ) ;
  assign n5730 = ( ~n1126 & n5726 ) | ( ~n1126 & n5727 ) | ( n5726 & n5727 ) ;
  assign n5731 = ( ~n1115 & n5729 ) | ( ~n1115 & n5730 ) | ( n5729 & n5730 ) ;
  assign n5732 = ( ~n975 & n5728 ) | ( ~n975 & n5731 ) | ( n5728 & n5731 ) ;
  assign n5733 = ( n1154 & n5728 ) | ( n1154 & n5731 ) | ( n5728 & n5731 ) ;
  assign n5734 = ( ~x409 & n5732 ) | ( ~x409 & n5733 ) | ( n5732 & n5733 ) ;
  assign n5735 = ( x281 & n5732 ) | ( x281 & n5733 ) | ( n5732 & n5733 ) ;
  assign n5736 = ( n656 & n5734 ) | ( n656 & n5735 ) | ( n5734 & n5735 ) ;
  assign n5737 = n5725 | n5736 ;
  assign n5738 = ~n5714 & n5737 ;
  assign n5739 = x196 & n1767 ;
  assign n5740 = x196 & ~n1771 ;
  assign n5741 = ( ~n1751 & n5739 ) | ( ~n1751 & n5740 ) | ( n5739 & n5740 ) ;
  assign n5742 = ( ~n1787 & n5739 ) | ( ~n1787 & n5740 ) | ( n5739 & n5740 ) ;
  assign n5743 = ( n1794 & n5739 ) | ( n1794 & n5740 ) | ( n5739 & n5740 ) ;
  assign n5744 = ( n1783 & n5742 ) | ( n1783 & n5743 ) | ( n5742 & n5743 ) ;
  assign n5745 = ( n1643 & n5741 ) | ( n1643 & n5744 ) | ( n5741 & n5744 ) ;
  assign n5746 = ( ~n1822 & n5741 ) | ( ~n1822 & n5744 ) | ( n5741 & n5744 ) ;
  assign n5747 = ( ~n1324 & n5745 ) | ( ~n1324 & n5746 ) | ( n5745 & n5746 ) ;
  assign n5748 = x68 & ~n1767 ;
  assign n5749 = x68 & n1771 ;
  assign n5750 = ( n1751 & n5748 ) | ( n1751 & n5749 ) | ( n5748 & n5749 ) ;
  assign n5751 = ( n1787 & n5748 ) | ( n1787 & n5749 ) | ( n5748 & n5749 ) ;
  assign n5752 = ( ~n1794 & n5748 ) | ( ~n1794 & n5749 ) | ( n5748 & n5749 ) ;
  assign n5753 = ( ~n1783 & n5751 ) | ( ~n1783 & n5752 ) | ( n5751 & n5752 ) ;
  assign n5754 = ( ~n1643 & n5750 ) | ( ~n1643 & n5753 ) | ( n5750 & n5753 ) ;
  assign n5755 = ( n1822 & n5750 ) | ( n1822 & n5753 ) | ( n5750 & n5753 ) ;
  assign n5756 = ( n1324 & n5754 ) | ( n1324 & n5755 ) | ( n5754 & n5755 ) ;
  assign n5757 = n5747 | n5756 ;
  assign n5758 = x452 & n991 ;
  assign n5759 = x452 & ~n995 ;
  assign n5760 = ( ~n1104 & n5758 ) | ( ~n1104 & n5759 ) | ( n5758 & n5759 ) ;
  assign n5761 = ( ~n1119 & n5758 ) | ( ~n1119 & n5759 ) | ( n5758 & n5759 ) ;
  assign n5762 = ( n1126 & n5758 ) | ( n1126 & n5759 ) | ( n5758 & n5759 ) ;
  assign n5763 = ( n1115 & n5761 ) | ( n1115 & n5762 ) | ( n5761 & n5762 ) ;
  assign n5764 = ( n975 & n5760 ) | ( n975 & n5763 ) | ( n5760 & n5763 ) ;
  assign n5765 = ( ~n1154 & n5760 ) | ( ~n1154 & n5763 ) | ( n5760 & n5763 ) ;
  assign n5766 = ( x409 & n5764 ) | ( x409 & n5765 ) | ( n5764 & n5765 ) ;
  assign n5767 = ( ~x281 & n5764 ) | ( ~x281 & n5765 ) | ( n5764 & n5765 ) ;
  assign n5768 = ( ~n656 & n5766 ) | ( ~n656 & n5767 ) | ( n5766 & n5767 ) ;
  assign n5769 = x324 & ~n991 ;
  assign n5770 = x324 & n995 ;
  assign n5771 = ( n1104 & n5769 ) | ( n1104 & n5770 ) | ( n5769 & n5770 ) ;
  assign n5772 = ( n1119 & n5769 ) | ( n1119 & n5770 ) | ( n5769 & n5770 ) ;
  assign n5773 = ( ~n1126 & n5769 ) | ( ~n1126 & n5770 ) | ( n5769 & n5770 ) ;
  assign n5774 = ( ~n1115 & n5772 ) | ( ~n1115 & n5773 ) | ( n5772 & n5773 ) ;
  assign n5775 = ( ~n975 & n5771 ) | ( ~n975 & n5774 ) | ( n5771 & n5774 ) ;
  assign n5776 = ( n1154 & n5771 ) | ( n1154 & n5774 ) | ( n5771 & n5774 ) ;
  assign n5777 = ( ~x409 & n5775 ) | ( ~x409 & n5776 ) | ( n5775 & n5776 ) ;
  assign n5778 = ( x281 & n5775 ) | ( x281 & n5776 ) | ( n5775 & n5776 ) ;
  assign n5779 = ( n656 & n5777 ) | ( n656 & n5778 ) | ( n5777 & n5778 ) ;
  assign n5780 = n5768 | n5779 ;
  assign n5781 = ~n5757 & n5780 ;
  assign n5782 = n5738 | n5781 ;
  assign n5783 = n5695 | n5782 ;
  assign n5784 = x195 & n1767 ;
  assign n5785 = x195 & ~n1771 ;
  assign n5786 = ( ~n1751 & n5784 ) | ( ~n1751 & n5785 ) | ( n5784 & n5785 ) ;
  assign n5787 = ( ~n1787 & n5784 ) | ( ~n1787 & n5785 ) | ( n5784 & n5785 ) ;
  assign n5788 = ( n1794 & n5784 ) | ( n1794 & n5785 ) | ( n5784 & n5785 ) ;
  assign n5789 = ( n1783 & n5787 ) | ( n1783 & n5788 ) | ( n5787 & n5788 ) ;
  assign n5790 = ( n1643 & n5786 ) | ( n1643 & n5789 ) | ( n5786 & n5789 ) ;
  assign n5791 = ( ~n1822 & n5786 ) | ( ~n1822 & n5789 ) | ( n5786 & n5789 ) ;
  assign n5792 = ( ~n1324 & n5790 ) | ( ~n1324 & n5791 ) | ( n5790 & n5791 ) ;
  assign n5793 = x67 & ~n1767 ;
  assign n5794 = x67 & n1771 ;
  assign n5795 = ( n1751 & n5793 ) | ( n1751 & n5794 ) | ( n5793 & n5794 ) ;
  assign n5796 = ( n1787 & n5793 ) | ( n1787 & n5794 ) | ( n5793 & n5794 ) ;
  assign n5797 = ( ~n1794 & n5793 ) | ( ~n1794 & n5794 ) | ( n5793 & n5794 ) ;
  assign n5798 = ( ~n1783 & n5796 ) | ( ~n1783 & n5797 ) | ( n5796 & n5797 ) ;
  assign n5799 = ( ~n1643 & n5795 ) | ( ~n1643 & n5798 ) | ( n5795 & n5798 ) ;
  assign n5800 = ( n1822 & n5795 ) | ( n1822 & n5798 ) | ( n5795 & n5798 ) ;
  assign n5801 = ( n1324 & n5799 ) | ( n1324 & n5800 ) | ( n5799 & n5800 ) ;
  assign n5802 = n5792 | n5801 ;
  assign n5803 = x451 & n991 ;
  assign n5804 = x451 & ~n995 ;
  assign n5805 = ( ~n1104 & n5803 ) | ( ~n1104 & n5804 ) | ( n5803 & n5804 ) ;
  assign n5806 = ( ~n1119 & n5803 ) | ( ~n1119 & n5804 ) | ( n5803 & n5804 ) ;
  assign n5807 = ( n1126 & n5803 ) | ( n1126 & n5804 ) | ( n5803 & n5804 ) ;
  assign n5808 = ( n1115 & n5806 ) | ( n1115 & n5807 ) | ( n5806 & n5807 ) ;
  assign n5809 = ( n975 & n5805 ) | ( n975 & n5808 ) | ( n5805 & n5808 ) ;
  assign n5810 = ( ~n1154 & n5805 ) | ( ~n1154 & n5808 ) | ( n5805 & n5808 ) ;
  assign n5811 = ( x409 & n5809 ) | ( x409 & n5810 ) | ( n5809 & n5810 ) ;
  assign n5812 = ( ~x281 & n5809 ) | ( ~x281 & n5810 ) | ( n5809 & n5810 ) ;
  assign n5813 = ( ~n656 & n5811 ) | ( ~n656 & n5812 ) | ( n5811 & n5812 ) ;
  assign n5814 = x323 & ~n991 ;
  assign n5815 = x323 & n995 ;
  assign n5816 = ( n1104 & n5814 ) | ( n1104 & n5815 ) | ( n5814 & n5815 ) ;
  assign n5817 = ( n1119 & n5814 ) | ( n1119 & n5815 ) | ( n5814 & n5815 ) ;
  assign n5818 = ( ~n1126 & n5814 ) | ( ~n1126 & n5815 ) | ( n5814 & n5815 ) ;
  assign n5819 = ( ~n1115 & n5817 ) | ( ~n1115 & n5818 ) | ( n5817 & n5818 ) ;
  assign n5820 = ( ~n975 & n5816 ) | ( ~n975 & n5819 ) | ( n5816 & n5819 ) ;
  assign n5821 = ( n1154 & n5816 ) | ( n1154 & n5819 ) | ( n5816 & n5819 ) ;
  assign n5822 = ( ~x409 & n5820 ) | ( ~x409 & n5821 ) | ( n5820 & n5821 ) ;
  assign n5823 = ( x281 & n5820 ) | ( x281 & n5821 ) | ( n5820 & n5821 ) ;
  assign n5824 = ( n656 & n5822 ) | ( n656 & n5823 ) | ( n5822 & n5823 ) ;
  assign n5825 = n5813 | n5824 ;
  assign n5826 = ~n5802 & n5825 ;
  assign n5827 = x450 & n991 ;
  assign n5828 = x450 & ~n995 ;
  assign n5829 = ( ~n1104 & n5827 ) | ( ~n1104 & n5828 ) | ( n5827 & n5828 ) ;
  assign n5830 = ( ~n1119 & n5827 ) | ( ~n1119 & n5828 ) | ( n5827 & n5828 ) ;
  assign n5831 = ( n1126 & n5827 ) | ( n1126 & n5828 ) | ( n5827 & n5828 ) ;
  assign n5832 = ( n1115 & n5830 ) | ( n1115 & n5831 ) | ( n5830 & n5831 ) ;
  assign n5833 = ( n975 & n5829 ) | ( n975 & n5832 ) | ( n5829 & n5832 ) ;
  assign n5834 = ( ~n1154 & n5829 ) | ( ~n1154 & n5832 ) | ( n5829 & n5832 ) ;
  assign n5835 = ( x409 & n5833 ) | ( x409 & n5834 ) | ( n5833 & n5834 ) ;
  assign n5836 = ( ~x281 & n5833 ) | ( ~x281 & n5834 ) | ( n5833 & n5834 ) ;
  assign n5837 = ( ~n656 & n5835 ) | ( ~n656 & n5836 ) | ( n5835 & n5836 ) ;
  assign n5838 = x322 & ~n991 ;
  assign n5839 = x322 & n995 ;
  assign n5840 = ( n1104 & n5838 ) | ( n1104 & n5839 ) | ( n5838 & n5839 ) ;
  assign n5841 = ( n1119 & n5838 ) | ( n1119 & n5839 ) | ( n5838 & n5839 ) ;
  assign n5842 = ( ~n1126 & n5838 ) | ( ~n1126 & n5839 ) | ( n5838 & n5839 ) ;
  assign n5843 = ( ~n1115 & n5841 ) | ( ~n1115 & n5842 ) | ( n5841 & n5842 ) ;
  assign n5844 = ( ~n975 & n5840 ) | ( ~n975 & n5843 ) | ( n5840 & n5843 ) ;
  assign n5845 = ( n1154 & n5840 ) | ( n1154 & n5843 ) | ( n5840 & n5843 ) ;
  assign n5846 = ( ~x409 & n5844 ) | ( ~x409 & n5845 ) | ( n5844 & n5845 ) ;
  assign n5847 = ( x281 & n5844 ) | ( x281 & n5845 ) | ( n5844 & n5845 ) ;
  assign n5848 = ( n656 & n5846 ) | ( n656 & n5847 ) | ( n5846 & n5847 ) ;
  assign n5849 = n5837 | n5848 ;
  assign n5850 = x194 & n1767 ;
  assign n5851 = x194 & ~n1771 ;
  assign n5852 = ( ~n1751 & n5850 ) | ( ~n1751 & n5851 ) | ( n5850 & n5851 ) ;
  assign n5853 = ( ~n1787 & n5850 ) | ( ~n1787 & n5851 ) | ( n5850 & n5851 ) ;
  assign n5854 = ( n1794 & n5850 ) | ( n1794 & n5851 ) | ( n5850 & n5851 ) ;
  assign n5855 = ( n1783 & n5853 ) | ( n1783 & n5854 ) | ( n5853 & n5854 ) ;
  assign n5856 = ( n1643 & n5852 ) | ( n1643 & n5855 ) | ( n5852 & n5855 ) ;
  assign n5857 = ( ~n1822 & n5852 ) | ( ~n1822 & n5855 ) | ( n5852 & n5855 ) ;
  assign n5858 = ( ~n1324 & n5856 ) | ( ~n1324 & n5857 ) | ( n5856 & n5857 ) ;
  assign n5859 = x66 & ~n1767 ;
  assign n5860 = x66 & n1771 ;
  assign n5861 = ( n1751 & n5859 ) | ( n1751 & n5860 ) | ( n5859 & n5860 ) ;
  assign n5862 = ( n1787 & n5859 ) | ( n1787 & n5860 ) | ( n5859 & n5860 ) ;
  assign n5863 = ( ~n1794 & n5859 ) | ( ~n1794 & n5860 ) | ( n5859 & n5860 ) ;
  assign n5864 = ( ~n1783 & n5862 ) | ( ~n1783 & n5863 ) | ( n5862 & n5863 ) ;
  assign n5865 = ( ~n1643 & n5861 ) | ( ~n1643 & n5864 ) | ( n5861 & n5864 ) ;
  assign n5866 = ( n1822 & n5861 ) | ( n1822 & n5864 ) | ( n5861 & n5864 ) ;
  assign n5867 = ( n1324 & n5865 ) | ( n1324 & n5866 ) | ( n5865 & n5866 ) ;
  assign n5868 = n5858 | n5867 ;
  assign n5869 = n5849 & ~n5868 ;
  assign n5870 = n5826 | n5869 ;
  assign n5871 = x193 & n1767 ;
  assign n5872 = x193 & ~n1771 ;
  assign n5873 = ( ~n1751 & n5871 ) | ( ~n1751 & n5872 ) | ( n5871 & n5872 ) ;
  assign n5874 = ( ~n1787 & n5871 ) | ( ~n1787 & n5872 ) | ( n5871 & n5872 ) ;
  assign n5875 = ( n1794 & n5871 ) | ( n1794 & n5872 ) | ( n5871 & n5872 ) ;
  assign n5876 = ( n1783 & n5874 ) | ( n1783 & n5875 ) | ( n5874 & n5875 ) ;
  assign n5877 = ( n1643 & n5873 ) | ( n1643 & n5876 ) | ( n5873 & n5876 ) ;
  assign n5878 = ( ~n1822 & n5873 ) | ( ~n1822 & n5876 ) | ( n5873 & n5876 ) ;
  assign n5879 = ( ~n1324 & n5877 ) | ( ~n1324 & n5878 ) | ( n5877 & n5878 ) ;
  assign n5880 = x65 & ~n1767 ;
  assign n5881 = x65 & n1771 ;
  assign n5882 = ( n1751 & n5880 ) | ( n1751 & n5881 ) | ( n5880 & n5881 ) ;
  assign n5883 = ( n1787 & n5880 ) | ( n1787 & n5881 ) | ( n5880 & n5881 ) ;
  assign n5884 = ( ~n1794 & n5880 ) | ( ~n1794 & n5881 ) | ( n5880 & n5881 ) ;
  assign n5885 = ( ~n1783 & n5883 ) | ( ~n1783 & n5884 ) | ( n5883 & n5884 ) ;
  assign n5886 = ( ~n1643 & n5882 ) | ( ~n1643 & n5885 ) | ( n5882 & n5885 ) ;
  assign n5887 = ( n1822 & n5882 ) | ( n1822 & n5885 ) | ( n5882 & n5885 ) ;
  assign n5888 = ( n1324 & n5886 ) | ( n1324 & n5887 ) | ( n5886 & n5887 ) ;
  assign n5889 = n5879 | n5888 ;
  assign n5890 = x449 & n991 ;
  assign n5891 = x449 & ~n995 ;
  assign n5892 = ( ~n1104 & n5890 ) | ( ~n1104 & n5891 ) | ( n5890 & n5891 ) ;
  assign n5893 = ( ~n1119 & n5890 ) | ( ~n1119 & n5891 ) | ( n5890 & n5891 ) ;
  assign n5894 = ( n1126 & n5890 ) | ( n1126 & n5891 ) | ( n5890 & n5891 ) ;
  assign n5895 = ( n1115 & n5893 ) | ( n1115 & n5894 ) | ( n5893 & n5894 ) ;
  assign n5896 = ( n975 & n5892 ) | ( n975 & n5895 ) | ( n5892 & n5895 ) ;
  assign n5897 = ( ~n1154 & n5892 ) | ( ~n1154 & n5895 ) | ( n5892 & n5895 ) ;
  assign n5898 = ( x409 & n5896 ) | ( x409 & n5897 ) | ( n5896 & n5897 ) ;
  assign n5899 = ( ~x281 & n5896 ) | ( ~x281 & n5897 ) | ( n5896 & n5897 ) ;
  assign n5900 = ( ~n656 & n5898 ) | ( ~n656 & n5899 ) | ( n5898 & n5899 ) ;
  assign n5901 = x321 & ~n991 ;
  assign n5902 = x321 & n995 ;
  assign n5903 = ( n1104 & n5901 ) | ( n1104 & n5902 ) | ( n5901 & n5902 ) ;
  assign n5904 = ( n1119 & n5901 ) | ( n1119 & n5902 ) | ( n5901 & n5902 ) ;
  assign n5905 = ( ~n1126 & n5901 ) | ( ~n1126 & n5902 ) | ( n5901 & n5902 ) ;
  assign n5906 = ( ~n1115 & n5904 ) | ( ~n1115 & n5905 ) | ( n5904 & n5905 ) ;
  assign n5907 = ( ~n975 & n5903 ) | ( ~n975 & n5906 ) | ( n5903 & n5906 ) ;
  assign n5908 = ( n1154 & n5903 ) | ( n1154 & n5906 ) | ( n5903 & n5906 ) ;
  assign n5909 = ( ~x409 & n5907 ) | ( ~x409 & n5908 ) | ( n5907 & n5908 ) ;
  assign n5910 = ( x281 & n5907 ) | ( x281 & n5908 ) | ( n5907 & n5908 ) ;
  assign n5911 = ( n656 & n5909 ) | ( n656 & n5910 ) | ( n5909 & n5910 ) ;
  assign n5912 = n5900 | n5911 ;
  assign n5913 = ~n5889 & n5912 ;
  assign n5914 = x448 & n991 ;
  assign n5915 = x448 & ~n995 ;
  assign n5916 = ( ~n1104 & n5914 ) | ( ~n1104 & n5915 ) | ( n5914 & n5915 ) ;
  assign n5917 = ( ~n1119 & n5914 ) | ( ~n1119 & n5915 ) | ( n5914 & n5915 ) ;
  assign n5918 = ( n1126 & n5914 ) | ( n1126 & n5915 ) | ( n5914 & n5915 ) ;
  assign n5919 = ( n1115 & n5917 ) | ( n1115 & n5918 ) | ( n5917 & n5918 ) ;
  assign n5920 = ( n975 & n5916 ) | ( n975 & n5919 ) | ( n5916 & n5919 ) ;
  assign n5921 = ( ~n1154 & n5916 ) | ( ~n1154 & n5919 ) | ( n5916 & n5919 ) ;
  assign n5922 = ( x409 & n5920 ) | ( x409 & n5921 ) | ( n5920 & n5921 ) ;
  assign n5923 = ( ~x281 & n5920 ) | ( ~x281 & n5921 ) | ( n5920 & n5921 ) ;
  assign n5924 = ( ~n656 & n5922 ) | ( ~n656 & n5923 ) | ( n5922 & n5923 ) ;
  assign n5925 = x320 & ~n991 ;
  assign n5926 = x320 & n995 ;
  assign n5927 = ( n1104 & n5925 ) | ( n1104 & n5926 ) | ( n5925 & n5926 ) ;
  assign n5928 = ( n1119 & n5925 ) | ( n1119 & n5926 ) | ( n5925 & n5926 ) ;
  assign n5929 = ( ~n1126 & n5925 ) | ( ~n1126 & n5926 ) | ( n5925 & n5926 ) ;
  assign n5930 = ( ~n1115 & n5928 ) | ( ~n1115 & n5929 ) | ( n5928 & n5929 ) ;
  assign n5931 = ( ~n975 & n5927 ) | ( ~n975 & n5930 ) | ( n5927 & n5930 ) ;
  assign n5932 = ( n1154 & n5927 ) | ( n1154 & n5930 ) | ( n5927 & n5930 ) ;
  assign n5933 = ( ~x409 & n5931 ) | ( ~x409 & n5932 ) | ( n5931 & n5932 ) ;
  assign n5934 = ( x281 & n5931 ) | ( x281 & n5932 ) | ( n5931 & n5932 ) ;
  assign n5935 = ( n656 & n5933 ) | ( n656 & n5934 ) | ( n5933 & n5934 ) ;
  assign n5936 = n5924 | n5935 ;
  assign n5937 = x192 & n1767 ;
  assign n5938 = x192 & ~n1771 ;
  assign n5939 = ( ~n1751 & n5937 ) | ( ~n1751 & n5938 ) | ( n5937 & n5938 ) ;
  assign n5940 = ( ~n1787 & n5937 ) | ( ~n1787 & n5938 ) | ( n5937 & n5938 ) ;
  assign n5941 = ( n1794 & n5937 ) | ( n1794 & n5938 ) | ( n5937 & n5938 ) ;
  assign n5942 = ( n1783 & n5940 ) | ( n1783 & n5941 ) | ( n5940 & n5941 ) ;
  assign n5943 = ( n1643 & n5939 ) | ( n1643 & n5942 ) | ( n5939 & n5942 ) ;
  assign n5944 = ( ~n1822 & n5939 ) | ( ~n1822 & n5942 ) | ( n5939 & n5942 ) ;
  assign n5945 = ( ~n1324 & n5943 ) | ( ~n1324 & n5944 ) | ( n5943 & n5944 ) ;
  assign n5946 = x64 & ~n1767 ;
  assign n5947 = x64 & n1771 ;
  assign n5948 = ( n1751 & n5946 ) | ( n1751 & n5947 ) | ( n5946 & n5947 ) ;
  assign n5949 = ( n1787 & n5946 ) | ( n1787 & n5947 ) | ( n5946 & n5947 ) ;
  assign n5950 = ( ~n1794 & n5946 ) | ( ~n1794 & n5947 ) | ( n5946 & n5947 ) ;
  assign n5951 = ( ~n1783 & n5949 ) | ( ~n1783 & n5950 ) | ( n5949 & n5950 ) ;
  assign n5952 = ( ~n1643 & n5948 ) | ( ~n1643 & n5951 ) | ( n5948 & n5951 ) ;
  assign n5953 = ( n1822 & n5948 ) | ( n1822 & n5951 ) | ( n5948 & n5951 ) ;
  assign n5954 = ( n1324 & n5952 ) | ( n1324 & n5953 ) | ( n5952 & n5953 ) ;
  assign n5955 = n5945 | n5954 ;
  assign n5956 = n5936 & ~n5955 ;
  assign n5957 = n5913 | n5956 ;
  assign n5958 = n5870 | n5957 ;
  assign n5959 = n5783 | n5958 ;
  assign n5960 = ~n5936 & n5955 ;
  assign n5961 = ( n5889 & ~n5912 ) | ( n5889 & n5960 ) | ( ~n5912 & n5960 ) ;
  assign n5962 = ~n5849 & n5868 ;
  assign n5963 = ~n5869 & n5962 ;
  assign n5964 = ( ~n5869 & n5961 ) | ( ~n5869 & n5963 ) | ( n5961 & n5963 ) ;
  assign n5965 = ( n5802 & ~n5825 ) | ( n5802 & n5964 ) | ( ~n5825 & n5964 ) ;
  assign n5966 = ( n5783 & n5959 ) | ( n5783 & ~n5965 ) | ( n5959 & ~n5965 ) ;
  assign n5967 = ~n5693 & n5966 ;
  assign n5968 = x207 & n1767 ;
  assign n5969 = x207 & ~n1771 ;
  assign n5970 = ( ~n1751 & n5968 ) | ( ~n1751 & n5969 ) | ( n5968 & n5969 ) ;
  assign n5971 = ( ~n1787 & n5968 ) | ( ~n1787 & n5969 ) | ( n5968 & n5969 ) ;
  assign n5972 = ( n1794 & n5968 ) | ( n1794 & n5969 ) | ( n5968 & n5969 ) ;
  assign n5973 = ( n1783 & n5971 ) | ( n1783 & n5972 ) | ( n5971 & n5972 ) ;
  assign n5974 = ( n1643 & n5970 ) | ( n1643 & n5973 ) | ( n5970 & n5973 ) ;
  assign n5975 = ( ~n1822 & n5970 ) | ( ~n1822 & n5973 ) | ( n5970 & n5973 ) ;
  assign n5976 = ( ~n1324 & n5974 ) | ( ~n1324 & n5975 ) | ( n5974 & n5975 ) ;
  assign n5977 = x79 & ~n1767 ;
  assign n5978 = x79 & n1771 ;
  assign n5979 = ( n1751 & n5977 ) | ( n1751 & n5978 ) | ( n5977 & n5978 ) ;
  assign n5980 = ( n1787 & n5977 ) | ( n1787 & n5978 ) | ( n5977 & n5978 ) ;
  assign n5981 = ( ~n1794 & n5977 ) | ( ~n1794 & n5978 ) | ( n5977 & n5978 ) ;
  assign n5982 = ( ~n1783 & n5980 ) | ( ~n1783 & n5981 ) | ( n5980 & n5981 ) ;
  assign n5983 = ( ~n1643 & n5979 ) | ( ~n1643 & n5982 ) | ( n5979 & n5982 ) ;
  assign n5984 = ( n1822 & n5979 ) | ( n1822 & n5982 ) | ( n5979 & n5982 ) ;
  assign n5985 = ( n1324 & n5983 ) | ( n1324 & n5984 ) | ( n5983 & n5984 ) ;
  assign n5986 = n5976 | n5985 ;
  assign n5987 = x463 & n991 ;
  assign n5988 = x463 & ~n995 ;
  assign n5989 = ( ~n1104 & n5987 ) | ( ~n1104 & n5988 ) | ( n5987 & n5988 ) ;
  assign n5990 = ( ~n1119 & n5987 ) | ( ~n1119 & n5988 ) | ( n5987 & n5988 ) ;
  assign n5991 = ( n1126 & n5987 ) | ( n1126 & n5988 ) | ( n5987 & n5988 ) ;
  assign n5992 = ( n1115 & n5990 ) | ( n1115 & n5991 ) | ( n5990 & n5991 ) ;
  assign n5993 = ( n975 & n5989 ) | ( n975 & n5992 ) | ( n5989 & n5992 ) ;
  assign n5994 = ( ~n1154 & n5989 ) | ( ~n1154 & n5992 ) | ( n5989 & n5992 ) ;
  assign n5995 = ( x409 & n5993 ) | ( x409 & n5994 ) | ( n5993 & n5994 ) ;
  assign n5996 = ( ~x281 & n5993 ) | ( ~x281 & n5994 ) | ( n5993 & n5994 ) ;
  assign n5997 = ( ~n656 & n5995 ) | ( ~n656 & n5996 ) | ( n5995 & n5996 ) ;
  assign n5998 = x335 & ~n991 ;
  assign n5999 = x335 & n995 ;
  assign n6000 = ( n1104 & n5998 ) | ( n1104 & n5999 ) | ( n5998 & n5999 ) ;
  assign n6001 = ( n1119 & n5998 ) | ( n1119 & n5999 ) | ( n5998 & n5999 ) ;
  assign n6002 = ( ~n1126 & n5998 ) | ( ~n1126 & n5999 ) | ( n5998 & n5999 ) ;
  assign n6003 = ( ~n1115 & n6001 ) | ( ~n1115 & n6002 ) | ( n6001 & n6002 ) ;
  assign n6004 = ( ~n975 & n6000 ) | ( ~n975 & n6003 ) | ( n6000 & n6003 ) ;
  assign n6005 = ( n1154 & n6000 ) | ( n1154 & n6003 ) | ( n6000 & n6003 ) ;
  assign n6006 = ( ~x409 & n6004 ) | ( ~x409 & n6005 ) | ( n6004 & n6005 ) ;
  assign n6007 = ( x281 & n6004 ) | ( x281 & n6005 ) | ( n6004 & n6005 ) ;
  assign n6008 = ( n656 & n6006 ) | ( n656 & n6007 ) | ( n6006 & n6007 ) ;
  assign n6009 = n5997 | n6008 ;
  assign n6010 = ~n5986 & n6009 ;
  assign n6011 = x462 & n991 ;
  assign n6012 = x462 & ~n995 ;
  assign n6013 = ( ~n1104 & n6011 ) | ( ~n1104 & n6012 ) | ( n6011 & n6012 ) ;
  assign n6014 = ( ~n1119 & n6011 ) | ( ~n1119 & n6012 ) | ( n6011 & n6012 ) ;
  assign n6015 = ( n1126 & n6011 ) | ( n1126 & n6012 ) | ( n6011 & n6012 ) ;
  assign n6016 = ( n1115 & n6014 ) | ( n1115 & n6015 ) | ( n6014 & n6015 ) ;
  assign n6017 = ( n975 & n6013 ) | ( n975 & n6016 ) | ( n6013 & n6016 ) ;
  assign n6018 = ( ~n1154 & n6013 ) | ( ~n1154 & n6016 ) | ( n6013 & n6016 ) ;
  assign n6019 = ( x409 & n6017 ) | ( x409 & n6018 ) | ( n6017 & n6018 ) ;
  assign n6020 = ( ~x281 & n6017 ) | ( ~x281 & n6018 ) | ( n6017 & n6018 ) ;
  assign n6021 = ( ~n656 & n6019 ) | ( ~n656 & n6020 ) | ( n6019 & n6020 ) ;
  assign n6022 = x334 & ~n991 ;
  assign n6023 = x334 & n995 ;
  assign n6024 = ( n1104 & n6022 ) | ( n1104 & n6023 ) | ( n6022 & n6023 ) ;
  assign n6025 = ( n1119 & n6022 ) | ( n1119 & n6023 ) | ( n6022 & n6023 ) ;
  assign n6026 = ( ~n1126 & n6022 ) | ( ~n1126 & n6023 ) | ( n6022 & n6023 ) ;
  assign n6027 = ( ~n1115 & n6025 ) | ( ~n1115 & n6026 ) | ( n6025 & n6026 ) ;
  assign n6028 = ( ~n975 & n6024 ) | ( ~n975 & n6027 ) | ( n6024 & n6027 ) ;
  assign n6029 = ( n1154 & n6024 ) | ( n1154 & n6027 ) | ( n6024 & n6027 ) ;
  assign n6030 = ( ~x409 & n6028 ) | ( ~x409 & n6029 ) | ( n6028 & n6029 ) ;
  assign n6031 = ( x281 & n6028 ) | ( x281 & n6029 ) | ( n6028 & n6029 ) ;
  assign n6032 = ( n656 & n6030 ) | ( n656 & n6031 ) | ( n6030 & n6031 ) ;
  assign n6033 = n6021 | n6032 ;
  assign n6034 = x206 & n1767 ;
  assign n6035 = x206 & ~n1771 ;
  assign n6036 = ( ~n1751 & n6034 ) | ( ~n1751 & n6035 ) | ( n6034 & n6035 ) ;
  assign n6037 = ( ~n1787 & n6034 ) | ( ~n1787 & n6035 ) | ( n6034 & n6035 ) ;
  assign n6038 = ( n1794 & n6034 ) | ( n1794 & n6035 ) | ( n6034 & n6035 ) ;
  assign n6039 = ( n1783 & n6037 ) | ( n1783 & n6038 ) | ( n6037 & n6038 ) ;
  assign n6040 = ( n1643 & n6036 ) | ( n1643 & n6039 ) | ( n6036 & n6039 ) ;
  assign n6041 = ( ~n1822 & n6036 ) | ( ~n1822 & n6039 ) | ( n6036 & n6039 ) ;
  assign n6042 = ( ~n1324 & n6040 ) | ( ~n1324 & n6041 ) | ( n6040 & n6041 ) ;
  assign n6043 = x78 & ~n1767 ;
  assign n6044 = x78 & n1771 ;
  assign n6045 = ( n1751 & n6043 ) | ( n1751 & n6044 ) | ( n6043 & n6044 ) ;
  assign n6046 = ( n1787 & n6043 ) | ( n1787 & n6044 ) | ( n6043 & n6044 ) ;
  assign n6047 = ( ~n1794 & n6043 ) | ( ~n1794 & n6044 ) | ( n6043 & n6044 ) ;
  assign n6048 = ( ~n1783 & n6046 ) | ( ~n1783 & n6047 ) | ( n6046 & n6047 ) ;
  assign n6049 = ( ~n1643 & n6045 ) | ( ~n1643 & n6048 ) | ( n6045 & n6048 ) ;
  assign n6050 = ( n1822 & n6045 ) | ( n1822 & n6048 ) | ( n6045 & n6048 ) ;
  assign n6051 = ( n1324 & n6049 ) | ( n1324 & n6050 ) | ( n6049 & n6050 ) ;
  assign n6052 = n6042 | n6051 ;
  assign n6053 = n6033 & ~n6052 ;
  assign n6054 = n6010 | n6053 ;
  assign n6055 = x205 & n1767 ;
  assign n6056 = x205 & ~n1771 ;
  assign n6057 = ( ~n1751 & n6055 ) | ( ~n1751 & n6056 ) | ( n6055 & n6056 ) ;
  assign n6058 = ( ~n1787 & n6055 ) | ( ~n1787 & n6056 ) | ( n6055 & n6056 ) ;
  assign n6059 = ( n1794 & n6055 ) | ( n1794 & n6056 ) | ( n6055 & n6056 ) ;
  assign n6060 = ( n1783 & n6058 ) | ( n1783 & n6059 ) | ( n6058 & n6059 ) ;
  assign n6061 = ( n1643 & n6057 ) | ( n1643 & n6060 ) | ( n6057 & n6060 ) ;
  assign n6062 = ( ~n1822 & n6057 ) | ( ~n1822 & n6060 ) | ( n6057 & n6060 ) ;
  assign n6063 = ( ~n1324 & n6061 ) | ( ~n1324 & n6062 ) | ( n6061 & n6062 ) ;
  assign n6064 = x77 & ~n1767 ;
  assign n6065 = x77 & n1771 ;
  assign n6066 = ( n1751 & n6064 ) | ( n1751 & n6065 ) | ( n6064 & n6065 ) ;
  assign n6067 = ( n1787 & n6064 ) | ( n1787 & n6065 ) | ( n6064 & n6065 ) ;
  assign n6068 = ( ~n1794 & n6064 ) | ( ~n1794 & n6065 ) | ( n6064 & n6065 ) ;
  assign n6069 = ( ~n1783 & n6067 ) | ( ~n1783 & n6068 ) | ( n6067 & n6068 ) ;
  assign n6070 = ( ~n1643 & n6066 ) | ( ~n1643 & n6069 ) | ( n6066 & n6069 ) ;
  assign n6071 = ( n1822 & n6066 ) | ( n1822 & n6069 ) | ( n6066 & n6069 ) ;
  assign n6072 = ( n1324 & n6070 ) | ( n1324 & n6071 ) | ( n6070 & n6071 ) ;
  assign n6073 = n6063 | n6072 ;
  assign n6074 = x461 & n991 ;
  assign n6075 = x461 & ~n995 ;
  assign n6076 = ( ~n1104 & n6074 ) | ( ~n1104 & n6075 ) | ( n6074 & n6075 ) ;
  assign n6077 = ( ~n1119 & n6074 ) | ( ~n1119 & n6075 ) | ( n6074 & n6075 ) ;
  assign n6078 = ( n1126 & n6074 ) | ( n1126 & n6075 ) | ( n6074 & n6075 ) ;
  assign n6079 = ( n1115 & n6077 ) | ( n1115 & n6078 ) | ( n6077 & n6078 ) ;
  assign n6080 = ( n975 & n6076 ) | ( n975 & n6079 ) | ( n6076 & n6079 ) ;
  assign n6081 = ( ~n1154 & n6076 ) | ( ~n1154 & n6079 ) | ( n6076 & n6079 ) ;
  assign n6082 = ( x409 & n6080 ) | ( x409 & n6081 ) | ( n6080 & n6081 ) ;
  assign n6083 = ( ~x281 & n6080 ) | ( ~x281 & n6081 ) | ( n6080 & n6081 ) ;
  assign n6084 = ( ~n656 & n6082 ) | ( ~n656 & n6083 ) | ( n6082 & n6083 ) ;
  assign n6085 = x333 & ~n991 ;
  assign n6086 = x333 & n995 ;
  assign n6087 = ( n1104 & n6085 ) | ( n1104 & n6086 ) | ( n6085 & n6086 ) ;
  assign n6088 = ( n1119 & n6085 ) | ( n1119 & n6086 ) | ( n6085 & n6086 ) ;
  assign n6089 = ( ~n1126 & n6085 ) | ( ~n1126 & n6086 ) | ( n6085 & n6086 ) ;
  assign n6090 = ( ~n1115 & n6088 ) | ( ~n1115 & n6089 ) | ( n6088 & n6089 ) ;
  assign n6091 = ( ~n975 & n6087 ) | ( ~n975 & n6090 ) | ( n6087 & n6090 ) ;
  assign n6092 = ( n1154 & n6087 ) | ( n1154 & n6090 ) | ( n6087 & n6090 ) ;
  assign n6093 = ( ~x409 & n6091 ) | ( ~x409 & n6092 ) | ( n6091 & n6092 ) ;
  assign n6094 = ( x281 & n6091 ) | ( x281 & n6092 ) | ( n6091 & n6092 ) ;
  assign n6095 = ( n656 & n6093 ) | ( n656 & n6094 ) | ( n6093 & n6094 ) ;
  assign n6096 = n6084 | n6095 ;
  assign n6097 = ~n6073 & n6096 ;
  assign n6098 = x204 & n1767 ;
  assign n6099 = x204 & ~n1771 ;
  assign n6100 = ( ~n1751 & n6098 ) | ( ~n1751 & n6099 ) | ( n6098 & n6099 ) ;
  assign n6101 = ( ~n1787 & n6098 ) | ( ~n1787 & n6099 ) | ( n6098 & n6099 ) ;
  assign n6102 = ( n1794 & n6098 ) | ( n1794 & n6099 ) | ( n6098 & n6099 ) ;
  assign n6103 = ( n1783 & n6101 ) | ( n1783 & n6102 ) | ( n6101 & n6102 ) ;
  assign n6104 = ( n1643 & n6100 ) | ( n1643 & n6103 ) | ( n6100 & n6103 ) ;
  assign n6105 = ( ~n1822 & n6100 ) | ( ~n1822 & n6103 ) | ( n6100 & n6103 ) ;
  assign n6106 = ( ~n1324 & n6104 ) | ( ~n1324 & n6105 ) | ( n6104 & n6105 ) ;
  assign n6107 = x76 & ~n1767 ;
  assign n6108 = x76 & n1771 ;
  assign n6109 = ( n1751 & n6107 ) | ( n1751 & n6108 ) | ( n6107 & n6108 ) ;
  assign n6110 = ( n1787 & n6107 ) | ( n1787 & n6108 ) | ( n6107 & n6108 ) ;
  assign n6111 = ( ~n1794 & n6107 ) | ( ~n1794 & n6108 ) | ( n6107 & n6108 ) ;
  assign n6112 = ( ~n1783 & n6110 ) | ( ~n1783 & n6111 ) | ( n6110 & n6111 ) ;
  assign n6113 = ( ~n1643 & n6109 ) | ( ~n1643 & n6112 ) | ( n6109 & n6112 ) ;
  assign n6114 = ( n1822 & n6109 ) | ( n1822 & n6112 ) | ( n6109 & n6112 ) ;
  assign n6115 = ( n1324 & n6113 ) | ( n1324 & n6114 ) | ( n6113 & n6114 ) ;
  assign n6116 = n6106 | n6115 ;
  assign n6117 = x460 & n991 ;
  assign n6118 = x460 & ~n995 ;
  assign n6119 = ( ~n1104 & n6117 ) | ( ~n1104 & n6118 ) | ( n6117 & n6118 ) ;
  assign n6120 = ( ~n1119 & n6117 ) | ( ~n1119 & n6118 ) | ( n6117 & n6118 ) ;
  assign n6121 = ( n1126 & n6117 ) | ( n1126 & n6118 ) | ( n6117 & n6118 ) ;
  assign n6122 = ( n1115 & n6120 ) | ( n1115 & n6121 ) | ( n6120 & n6121 ) ;
  assign n6123 = ( n975 & n6119 ) | ( n975 & n6122 ) | ( n6119 & n6122 ) ;
  assign n6124 = ( ~n1154 & n6119 ) | ( ~n1154 & n6122 ) | ( n6119 & n6122 ) ;
  assign n6125 = ( x409 & n6123 ) | ( x409 & n6124 ) | ( n6123 & n6124 ) ;
  assign n6126 = ( ~x281 & n6123 ) | ( ~x281 & n6124 ) | ( n6123 & n6124 ) ;
  assign n6127 = ( ~n656 & n6125 ) | ( ~n656 & n6126 ) | ( n6125 & n6126 ) ;
  assign n6128 = x332 & ~n991 ;
  assign n6129 = x332 & n995 ;
  assign n6130 = ( n1104 & n6128 ) | ( n1104 & n6129 ) | ( n6128 & n6129 ) ;
  assign n6131 = ( n1119 & n6128 ) | ( n1119 & n6129 ) | ( n6128 & n6129 ) ;
  assign n6132 = ( ~n1126 & n6128 ) | ( ~n1126 & n6129 ) | ( n6128 & n6129 ) ;
  assign n6133 = ( ~n1115 & n6131 ) | ( ~n1115 & n6132 ) | ( n6131 & n6132 ) ;
  assign n6134 = ( ~n975 & n6130 ) | ( ~n975 & n6133 ) | ( n6130 & n6133 ) ;
  assign n6135 = ( n1154 & n6130 ) | ( n1154 & n6133 ) | ( n6130 & n6133 ) ;
  assign n6136 = ( ~x409 & n6134 ) | ( ~x409 & n6135 ) | ( n6134 & n6135 ) ;
  assign n6137 = ( x281 & n6134 ) | ( x281 & n6135 ) | ( n6134 & n6135 ) ;
  assign n6138 = ( n656 & n6136 ) | ( n656 & n6137 ) | ( n6136 & n6137 ) ;
  assign n6139 = n6127 | n6138 ;
  assign n6140 = ~n6116 & n6139 ;
  assign n6141 = n6097 | n6140 ;
  assign n6142 = n6054 | n6141 ;
  assign n6143 = x203 & n1767 ;
  assign n6144 = x203 & ~n1771 ;
  assign n6145 = ( ~n1751 & n6143 ) | ( ~n1751 & n6144 ) | ( n6143 & n6144 ) ;
  assign n6146 = ( ~n1787 & n6143 ) | ( ~n1787 & n6144 ) | ( n6143 & n6144 ) ;
  assign n6147 = ( n1794 & n6143 ) | ( n1794 & n6144 ) | ( n6143 & n6144 ) ;
  assign n6148 = ( n1783 & n6146 ) | ( n1783 & n6147 ) | ( n6146 & n6147 ) ;
  assign n6149 = ( n1643 & n6145 ) | ( n1643 & n6148 ) | ( n6145 & n6148 ) ;
  assign n6150 = ( ~n1822 & n6145 ) | ( ~n1822 & n6148 ) | ( n6145 & n6148 ) ;
  assign n6151 = ( ~n1324 & n6149 ) | ( ~n1324 & n6150 ) | ( n6149 & n6150 ) ;
  assign n6152 = x75 & ~n1767 ;
  assign n6153 = x75 & n1771 ;
  assign n6154 = ( n1751 & n6152 ) | ( n1751 & n6153 ) | ( n6152 & n6153 ) ;
  assign n6155 = ( n1787 & n6152 ) | ( n1787 & n6153 ) | ( n6152 & n6153 ) ;
  assign n6156 = ( ~n1794 & n6152 ) | ( ~n1794 & n6153 ) | ( n6152 & n6153 ) ;
  assign n6157 = ( ~n1783 & n6155 ) | ( ~n1783 & n6156 ) | ( n6155 & n6156 ) ;
  assign n6158 = ( ~n1643 & n6154 ) | ( ~n1643 & n6157 ) | ( n6154 & n6157 ) ;
  assign n6159 = ( n1822 & n6154 ) | ( n1822 & n6157 ) | ( n6154 & n6157 ) ;
  assign n6160 = ( n1324 & n6158 ) | ( n1324 & n6159 ) | ( n6158 & n6159 ) ;
  assign n6161 = n6151 | n6160 ;
  assign n6162 = x459 & n991 ;
  assign n6163 = x459 & ~n995 ;
  assign n6164 = ( ~n1104 & n6162 ) | ( ~n1104 & n6163 ) | ( n6162 & n6163 ) ;
  assign n6165 = ( ~n1119 & n6162 ) | ( ~n1119 & n6163 ) | ( n6162 & n6163 ) ;
  assign n6166 = ( n1126 & n6162 ) | ( n1126 & n6163 ) | ( n6162 & n6163 ) ;
  assign n6167 = ( n1115 & n6165 ) | ( n1115 & n6166 ) | ( n6165 & n6166 ) ;
  assign n6168 = ( n975 & n6164 ) | ( n975 & n6167 ) | ( n6164 & n6167 ) ;
  assign n6169 = ( ~n1154 & n6164 ) | ( ~n1154 & n6167 ) | ( n6164 & n6167 ) ;
  assign n6170 = ( x409 & n6168 ) | ( x409 & n6169 ) | ( n6168 & n6169 ) ;
  assign n6171 = ( ~x281 & n6168 ) | ( ~x281 & n6169 ) | ( n6168 & n6169 ) ;
  assign n6172 = ( ~n656 & n6170 ) | ( ~n656 & n6171 ) | ( n6170 & n6171 ) ;
  assign n6173 = x331 & ~n991 ;
  assign n6174 = x331 & n995 ;
  assign n6175 = ( n1104 & n6173 ) | ( n1104 & n6174 ) | ( n6173 & n6174 ) ;
  assign n6176 = ( n1119 & n6173 ) | ( n1119 & n6174 ) | ( n6173 & n6174 ) ;
  assign n6177 = ( ~n1126 & n6173 ) | ( ~n1126 & n6174 ) | ( n6173 & n6174 ) ;
  assign n6178 = ( ~n1115 & n6176 ) | ( ~n1115 & n6177 ) | ( n6176 & n6177 ) ;
  assign n6179 = ( ~n975 & n6175 ) | ( ~n975 & n6178 ) | ( n6175 & n6178 ) ;
  assign n6180 = ( n1154 & n6175 ) | ( n1154 & n6178 ) | ( n6175 & n6178 ) ;
  assign n6181 = ( ~x409 & n6179 ) | ( ~x409 & n6180 ) | ( n6179 & n6180 ) ;
  assign n6182 = ( x281 & n6179 ) | ( x281 & n6180 ) | ( n6179 & n6180 ) ;
  assign n6183 = ( n656 & n6181 ) | ( n656 & n6182 ) | ( n6181 & n6182 ) ;
  assign n6184 = n6172 | n6183 ;
  assign n6185 = ~n6161 & n6184 ;
  assign n6186 = x458 & n991 ;
  assign n6187 = x458 & ~n995 ;
  assign n6188 = ( ~n1104 & n6186 ) | ( ~n1104 & n6187 ) | ( n6186 & n6187 ) ;
  assign n6189 = ( ~n1119 & n6186 ) | ( ~n1119 & n6187 ) | ( n6186 & n6187 ) ;
  assign n6190 = ( n1126 & n6186 ) | ( n1126 & n6187 ) | ( n6186 & n6187 ) ;
  assign n6191 = ( n1115 & n6189 ) | ( n1115 & n6190 ) | ( n6189 & n6190 ) ;
  assign n6192 = ( n975 & n6188 ) | ( n975 & n6191 ) | ( n6188 & n6191 ) ;
  assign n6193 = ( ~n1154 & n6188 ) | ( ~n1154 & n6191 ) | ( n6188 & n6191 ) ;
  assign n6194 = ( x409 & n6192 ) | ( x409 & n6193 ) | ( n6192 & n6193 ) ;
  assign n6195 = ( ~x281 & n6192 ) | ( ~x281 & n6193 ) | ( n6192 & n6193 ) ;
  assign n6196 = ( ~n656 & n6194 ) | ( ~n656 & n6195 ) | ( n6194 & n6195 ) ;
  assign n6197 = x330 & ~n991 ;
  assign n6198 = x330 & n995 ;
  assign n6199 = ( n1104 & n6197 ) | ( n1104 & n6198 ) | ( n6197 & n6198 ) ;
  assign n6200 = ( n1119 & n6197 ) | ( n1119 & n6198 ) | ( n6197 & n6198 ) ;
  assign n6201 = ( ~n1126 & n6197 ) | ( ~n1126 & n6198 ) | ( n6197 & n6198 ) ;
  assign n6202 = ( ~n1115 & n6200 ) | ( ~n1115 & n6201 ) | ( n6200 & n6201 ) ;
  assign n6203 = ( ~n975 & n6199 ) | ( ~n975 & n6202 ) | ( n6199 & n6202 ) ;
  assign n6204 = ( n1154 & n6199 ) | ( n1154 & n6202 ) | ( n6199 & n6202 ) ;
  assign n6205 = ( ~x409 & n6203 ) | ( ~x409 & n6204 ) | ( n6203 & n6204 ) ;
  assign n6206 = ( x281 & n6203 ) | ( x281 & n6204 ) | ( n6203 & n6204 ) ;
  assign n6207 = ( n656 & n6205 ) | ( n656 & n6206 ) | ( n6205 & n6206 ) ;
  assign n6208 = n6196 | n6207 ;
  assign n6209 = x202 & n1767 ;
  assign n6210 = x202 & ~n1771 ;
  assign n6211 = ( ~n1751 & n6209 ) | ( ~n1751 & n6210 ) | ( n6209 & n6210 ) ;
  assign n6212 = ( ~n1787 & n6209 ) | ( ~n1787 & n6210 ) | ( n6209 & n6210 ) ;
  assign n6213 = ( n1794 & n6209 ) | ( n1794 & n6210 ) | ( n6209 & n6210 ) ;
  assign n6214 = ( n1783 & n6212 ) | ( n1783 & n6213 ) | ( n6212 & n6213 ) ;
  assign n6215 = ( n1643 & n6211 ) | ( n1643 & n6214 ) | ( n6211 & n6214 ) ;
  assign n6216 = ( ~n1822 & n6211 ) | ( ~n1822 & n6214 ) | ( n6211 & n6214 ) ;
  assign n6217 = ( ~n1324 & n6215 ) | ( ~n1324 & n6216 ) | ( n6215 & n6216 ) ;
  assign n6218 = x74 & ~n1767 ;
  assign n6219 = x74 & n1771 ;
  assign n6220 = ( n1751 & n6218 ) | ( n1751 & n6219 ) | ( n6218 & n6219 ) ;
  assign n6221 = ( n1787 & n6218 ) | ( n1787 & n6219 ) | ( n6218 & n6219 ) ;
  assign n6222 = ( ~n1794 & n6218 ) | ( ~n1794 & n6219 ) | ( n6218 & n6219 ) ;
  assign n6223 = ( ~n1783 & n6221 ) | ( ~n1783 & n6222 ) | ( n6221 & n6222 ) ;
  assign n6224 = ( ~n1643 & n6220 ) | ( ~n1643 & n6223 ) | ( n6220 & n6223 ) ;
  assign n6225 = ( n1822 & n6220 ) | ( n1822 & n6223 ) | ( n6220 & n6223 ) ;
  assign n6226 = ( n1324 & n6224 ) | ( n1324 & n6225 ) | ( n6224 & n6225 ) ;
  assign n6227 = n6217 | n6226 ;
  assign n6228 = n6208 & ~n6227 ;
  assign n6229 = n6185 | n6228 ;
  assign n6230 = x201 & n1767 ;
  assign n6231 = x201 & ~n1771 ;
  assign n6232 = ( ~n1751 & n6230 ) | ( ~n1751 & n6231 ) | ( n6230 & n6231 ) ;
  assign n6233 = ( ~n1787 & n6230 ) | ( ~n1787 & n6231 ) | ( n6230 & n6231 ) ;
  assign n6234 = ( n1794 & n6230 ) | ( n1794 & n6231 ) | ( n6230 & n6231 ) ;
  assign n6235 = ( n1783 & n6233 ) | ( n1783 & n6234 ) | ( n6233 & n6234 ) ;
  assign n6236 = ( n1643 & n6232 ) | ( n1643 & n6235 ) | ( n6232 & n6235 ) ;
  assign n6237 = ( ~n1822 & n6232 ) | ( ~n1822 & n6235 ) | ( n6232 & n6235 ) ;
  assign n6238 = ( ~n1324 & n6236 ) | ( ~n1324 & n6237 ) | ( n6236 & n6237 ) ;
  assign n6239 = x73 & ~n1767 ;
  assign n6240 = x73 & n1771 ;
  assign n6241 = ( n1751 & n6239 ) | ( n1751 & n6240 ) | ( n6239 & n6240 ) ;
  assign n6242 = ( n1787 & n6239 ) | ( n1787 & n6240 ) | ( n6239 & n6240 ) ;
  assign n6243 = ( ~n1794 & n6239 ) | ( ~n1794 & n6240 ) | ( n6239 & n6240 ) ;
  assign n6244 = ( ~n1783 & n6242 ) | ( ~n1783 & n6243 ) | ( n6242 & n6243 ) ;
  assign n6245 = ( ~n1643 & n6241 ) | ( ~n1643 & n6244 ) | ( n6241 & n6244 ) ;
  assign n6246 = ( n1822 & n6241 ) | ( n1822 & n6244 ) | ( n6241 & n6244 ) ;
  assign n6247 = ( n1324 & n6245 ) | ( n1324 & n6246 ) | ( n6245 & n6246 ) ;
  assign n6248 = n6238 | n6247 ;
  assign n6249 = x457 & n991 ;
  assign n6250 = x457 & ~n995 ;
  assign n6251 = ( ~n1104 & n6249 ) | ( ~n1104 & n6250 ) | ( n6249 & n6250 ) ;
  assign n6252 = ( ~n1119 & n6249 ) | ( ~n1119 & n6250 ) | ( n6249 & n6250 ) ;
  assign n6253 = ( n1126 & n6249 ) | ( n1126 & n6250 ) | ( n6249 & n6250 ) ;
  assign n6254 = ( n1115 & n6252 ) | ( n1115 & n6253 ) | ( n6252 & n6253 ) ;
  assign n6255 = ( n975 & n6251 ) | ( n975 & n6254 ) | ( n6251 & n6254 ) ;
  assign n6256 = ( ~n1154 & n6251 ) | ( ~n1154 & n6254 ) | ( n6251 & n6254 ) ;
  assign n6257 = ( x409 & n6255 ) | ( x409 & n6256 ) | ( n6255 & n6256 ) ;
  assign n6258 = ( ~x281 & n6255 ) | ( ~x281 & n6256 ) | ( n6255 & n6256 ) ;
  assign n6259 = ( ~n656 & n6257 ) | ( ~n656 & n6258 ) | ( n6257 & n6258 ) ;
  assign n6260 = x329 & ~n991 ;
  assign n6261 = x329 & n995 ;
  assign n6262 = ( n1104 & n6260 ) | ( n1104 & n6261 ) | ( n6260 & n6261 ) ;
  assign n6263 = ( n1119 & n6260 ) | ( n1119 & n6261 ) | ( n6260 & n6261 ) ;
  assign n6264 = ( ~n1126 & n6260 ) | ( ~n1126 & n6261 ) | ( n6260 & n6261 ) ;
  assign n6265 = ( ~n1115 & n6263 ) | ( ~n1115 & n6264 ) | ( n6263 & n6264 ) ;
  assign n6266 = ( ~n975 & n6262 ) | ( ~n975 & n6265 ) | ( n6262 & n6265 ) ;
  assign n6267 = ( n1154 & n6262 ) | ( n1154 & n6265 ) | ( n6262 & n6265 ) ;
  assign n6268 = ( ~x409 & n6266 ) | ( ~x409 & n6267 ) | ( n6266 & n6267 ) ;
  assign n6269 = ( x281 & n6266 ) | ( x281 & n6267 ) | ( n6266 & n6267 ) ;
  assign n6270 = ( n656 & n6268 ) | ( n656 & n6269 ) | ( n6268 & n6269 ) ;
  assign n6271 = n6259 | n6270 ;
  assign n6272 = ~n6248 & n6271 ;
  assign n6273 = x456 & n991 ;
  assign n6274 = x456 & ~n995 ;
  assign n6275 = ( ~n1104 & n6273 ) | ( ~n1104 & n6274 ) | ( n6273 & n6274 ) ;
  assign n6276 = ( ~n1119 & n6273 ) | ( ~n1119 & n6274 ) | ( n6273 & n6274 ) ;
  assign n6277 = ( n1126 & n6273 ) | ( n1126 & n6274 ) | ( n6273 & n6274 ) ;
  assign n6278 = ( n1115 & n6276 ) | ( n1115 & n6277 ) | ( n6276 & n6277 ) ;
  assign n6279 = ( n975 & n6275 ) | ( n975 & n6278 ) | ( n6275 & n6278 ) ;
  assign n6280 = ( ~n1154 & n6275 ) | ( ~n1154 & n6278 ) | ( n6275 & n6278 ) ;
  assign n6281 = ( x409 & n6279 ) | ( x409 & n6280 ) | ( n6279 & n6280 ) ;
  assign n6282 = ( ~x281 & n6279 ) | ( ~x281 & n6280 ) | ( n6279 & n6280 ) ;
  assign n6283 = ( ~n656 & n6281 ) | ( ~n656 & n6282 ) | ( n6281 & n6282 ) ;
  assign n6284 = x328 & ~n991 ;
  assign n6285 = x328 & n995 ;
  assign n6286 = ( n1104 & n6284 ) | ( n1104 & n6285 ) | ( n6284 & n6285 ) ;
  assign n6287 = ( n1119 & n6284 ) | ( n1119 & n6285 ) | ( n6284 & n6285 ) ;
  assign n6288 = ( ~n1126 & n6284 ) | ( ~n1126 & n6285 ) | ( n6284 & n6285 ) ;
  assign n6289 = ( ~n1115 & n6287 ) | ( ~n1115 & n6288 ) | ( n6287 & n6288 ) ;
  assign n6290 = ( ~n975 & n6286 ) | ( ~n975 & n6289 ) | ( n6286 & n6289 ) ;
  assign n6291 = ( n1154 & n6286 ) | ( n1154 & n6289 ) | ( n6286 & n6289 ) ;
  assign n6292 = ( ~x409 & n6290 ) | ( ~x409 & n6291 ) | ( n6290 & n6291 ) ;
  assign n6293 = ( x281 & n6290 ) | ( x281 & n6291 ) | ( n6290 & n6291 ) ;
  assign n6294 = ( n656 & n6292 ) | ( n656 & n6293 ) | ( n6292 & n6293 ) ;
  assign n6295 = n6283 | n6294 ;
  assign n6296 = x200 & n1767 ;
  assign n6297 = x200 & ~n1771 ;
  assign n6298 = ( ~n1751 & n6296 ) | ( ~n1751 & n6297 ) | ( n6296 & n6297 ) ;
  assign n6299 = ( ~n1787 & n6296 ) | ( ~n1787 & n6297 ) | ( n6296 & n6297 ) ;
  assign n6300 = ( n1794 & n6296 ) | ( n1794 & n6297 ) | ( n6296 & n6297 ) ;
  assign n6301 = ( n1783 & n6299 ) | ( n1783 & n6300 ) | ( n6299 & n6300 ) ;
  assign n6302 = ( n1643 & n6298 ) | ( n1643 & n6301 ) | ( n6298 & n6301 ) ;
  assign n6303 = ( ~n1822 & n6298 ) | ( ~n1822 & n6301 ) | ( n6298 & n6301 ) ;
  assign n6304 = ( ~n1324 & n6302 ) | ( ~n1324 & n6303 ) | ( n6302 & n6303 ) ;
  assign n6305 = x72 & ~n1767 ;
  assign n6306 = x72 & n1771 ;
  assign n6307 = ( n1751 & n6305 ) | ( n1751 & n6306 ) | ( n6305 & n6306 ) ;
  assign n6308 = ( n1787 & n6305 ) | ( n1787 & n6306 ) | ( n6305 & n6306 ) ;
  assign n6309 = ( ~n1794 & n6305 ) | ( ~n1794 & n6306 ) | ( n6305 & n6306 ) ;
  assign n6310 = ( ~n1783 & n6308 ) | ( ~n1783 & n6309 ) | ( n6308 & n6309 ) ;
  assign n6311 = ( ~n1643 & n6307 ) | ( ~n1643 & n6310 ) | ( n6307 & n6310 ) ;
  assign n6312 = ( n1822 & n6307 ) | ( n1822 & n6310 ) | ( n6307 & n6310 ) ;
  assign n6313 = ( n1324 & n6311 ) | ( n1324 & n6312 ) | ( n6311 & n6312 ) ;
  assign n6314 = n6304 | n6313 ;
  assign n6315 = n6295 & ~n6314 ;
  assign n6316 = n6272 | n6315 ;
  assign n6317 = n6229 | n6316 ;
  assign n6318 = n5625 & ~n5648 ;
  assign n6319 = n5695 & ~n6318 ;
  assign n6320 = n5757 & ~n5780 ;
  assign n6321 = ( n5714 & ~n5737 ) | ( n5714 & n6320 ) | ( ~n5737 & n6320 ) ;
  assign n6322 = ( n6318 & ~n6319 ) | ( n6318 & n6321 ) | ( ~n6319 & n6321 ) ;
  assign n6323 = ~n6317 & n6322 ;
  assign n6324 = ~n6295 & n6314 ;
  assign n6325 = ( n6248 & ~n6271 ) | ( n6248 & n6324 ) | ( ~n6271 & n6324 ) ;
  assign n6326 = ~n6208 & n6227 ;
  assign n6327 = ~n6228 & n6326 ;
  assign n6328 = ( ~n6228 & n6325 ) | ( ~n6228 & n6327 ) | ( n6325 & n6327 ) ;
  assign n6329 = ( n6161 & ~n6184 ) | ( n6161 & n6328 ) | ( ~n6184 & n6328 ) ;
  assign n6330 = ~n6142 & n6329 ;
  assign n6331 = ( ~n6142 & n6323 ) | ( ~n6142 & n6330 ) | ( n6323 & n6330 ) ;
  assign n6332 = n6142 | n6317 ;
  assign n6333 = ( n6142 & ~n6329 ) | ( n6142 & n6332 ) | ( ~n6329 & n6332 ) ;
  assign n6334 = ( n5967 & ~n6331 ) | ( n5967 & n6333 ) | ( ~n6331 & n6333 ) ;
  assign n6335 = ~n5693 & n5783 ;
  assign n6336 = ( n5693 & n5965 ) | ( n5693 & ~n6335 ) | ( n5965 & ~n6335 ) ;
  assign n6337 = ( n6331 & ~n6333 ) | ( n6331 & n6336 ) | ( ~n6333 & n6336 ) ;
  assign n6338 = ( n5606 & n6334 ) | ( n5606 & ~n6337 ) | ( n6334 & ~n6337 ) ;
  assign n6339 = n6116 & ~n6139 ;
  assign n6340 = ( n6073 & ~n6096 ) | ( n6073 & n6339 ) | ( ~n6096 & n6339 ) ;
  assign n6341 = ~n6054 & n6340 ;
  assign n6342 = n5986 & ~n6009 ;
  assign n6343 = ~n5238 & n6342 ;
  assign n6344 = ~n6033 & n6052 ;
  assign n6345 = ~n6010 & n6344 ;
  assign n6346 = ( ~n5238 & n6343 ) | ( ~n5238 & n6345 ) | ( n6343 & n6345 ) ;
  assign n6347 = n5238 & ~n6343 ;
  assign n6348 = ( n6341 & n6346 ) | ( n6341 & ~n6347 ) | ( n6346 & ~n6347 ) ;
  assign n6349 = ( n5238 & n6338 ) | ( n5238 & ~n6348 ) | ( n6338 & ~n6348 ) ;
  assign n6350 = ~n5413 & n5603 ;
  assign n6351 = n5594 | n5597 ;
  assign n6352 = n5592 | n6351 ;
  assign n6353 = n6350 | n6352 ;
  assign n6354 = ~n5693 & n5695 ;
  assign n6355 = ( n5693 & n6321 ) | ( n5693 & ~n6354 ) | ( n6321 & ~n6354 ) ;
  assign n6356 = ~n6317 & n6318 ;
  assign n6357 = ( ~n6317 & n6355 ) | ( ~n6317 & n6356 ) | ( n6355 & n6356 ) ;
  assign n6358 = ( n5966 & n6317 ) | ( n5966 & ~n6357 ) | ( n6317 & ~n6357 ) ;
  assign n6359 = ~n5783 & n5965 ;
  assign n6360 = ( ~n6317 & n6357 ) | ( ~n6317 & n6359 ) | ( n6357 & n6359 ) ;
  assign n6361 = ( n6353 & ~n6358 ) | ( n6353 & n6360 ) | ( ~n6358 & n6360 ) ;
  assign n6362 = n6142 & ~n6345 ;
  assign n6363 = ( n6329 & n6345 ) | ( n6329 & ~n6362 ) | ( n6345 & ~n6362 ) ;
  assign n6364 = ( ~n5238 & n6341 ) | ( ~n5238 & n6343 ) | ( n6341 & n6343 ) ;
  assign n6365 = ( ~n5238 & n6363 ) | ( ~n5238 & n6364 ) | ( n6363 & n6364 ) ;
  assign n6366 = ( n6347 & n6362 ) | ( n6347 & ~n6364 ) | ( n6362 & ~n6364 ) ;
  assign n6367 = ( n6361 & n6365 ) | ( n6361 & ~n6366 ) | ( n6365 & ~n6366 ) ;
  assign n6368 = x183 & n1767 ;
  assign n6369 = x183 & ~n1771 ;
  assign n6370 = ( ~n1751 & n6368 ) | ( ~n1751 & n6369 ) | ( n6368 & n6369 ) ;
  assign n6371 = ( ~n1787 & n6368 ) | ( ~n1787 & n6369 ) | ( n6368 & n6369 ) ;
  assign n6372 = ( n1794 & n6368 ) | ( n1794 & n6369 ) | ( n6368 & n6369 ) ;
  assign n6373 = ( n1783 & n6371 ) | ( n1783 & n6372 ) | ( n6371 & n6372 ) ;
  assign n6374 = ( n1643 & n6370 ) | ( n1643 & n6373 ) | ( n6370 & n6373 ) ;
  assign n6375 = ( ~n1822 & n6370 ) | ( ~n1822 & n6373 ) | ( n6370 & n6373 ) ;
  assign n6376 = ( ~n1324 & n6374 ) | ( ~n1324 & n6375 ) | ( n6374 & n6375 ) ;
  assign n6377 = x55 & ~n1767 ;
  assign n6378 = x55 & n1771 ;
  assign n6379 = ( n1751 & n6377 ) | ( n1751 & n6378 ) | ( n6377 & n6378 ) ;
  assign n6380 = ( n1787 & n6377 ) | ( n1787 & n6378 ) | ( n6377 & n6378 ) ;
  assign n6381 = ( ~n1794 & n6377 ) | ( ~n1794 & n6378 ) | ( n6377 & n6378 ) ;
  assign n6382 = ( ~n1783 & n6380 ) | ( ~n1783 & n6381 ) | ( n6380 & n6381 ) ;
  assign n6383 = ( ~n1643 & n6379 ) | ( ~n1643 & n6382 ) | ( n6379 & n6382 ) ;
  assign n6384 = ( n1822 & n6379 ) | ( n1822 & n6382 ) | ( n6379 & n6382 ) ;
  assign n6385 = ( n1324 & n6383 ) | ( n1324 & n6384 ) | ( n6383 & n6384 ) ;
  assign n6386 = n6376 | n6385 ;
  assign n6387 = x439 & n991 ;
  assign n6388 = x439 & ~n995 ;
  assign n6389 = ( ~n1104 & n6387 ) | ( ~n1104 & n6388 ) | ( n6387 & n6388 ) ;
  assign n6390 = ( ~n1119 & n6387 ) | ( ~n1119 & n6388 ) | ( n6387 & n6388 ) ;
  assign n6391 = ( n1126 & n6387 ) | ( n1126 & n6388 ) | ( n6387 & n6388 ) ;
  assign n6392 = ( n1115 & n6390 ) | ( n1115 & n6391 ) | ( n6390 & n6391 ) ;
  assign n6393 = ( n975 & n6389 ) | ( n975 & n6392 ) | ( n6389 & n6392 ) ;
  assign n6394 = ( ~n1154 & n6389 ) | ( ~n1154 & n6392 ) | ( n6389 & n6392 ) ;
  assign n6395 = ( x409 & n6393 ) | ( x409 & n6394 ) | ( n6393 & n6394 ) ;
  assign n6396 = ( ~x281 & n6393 ) | ( ~x281 & n6394 ) | ( n6393 & n6394 ) ;
  assign n6397 = ( ~n656 & n6395 ) | ( ~n656 & n6396 ) | ( n6395 & n6396 ) ;
  assign n6398 = x311 & ~n991 ;
  assign n6399 = x311 & n995 ;
  assign n6400 = ( n1104 & n6398 ) | ( n1104 & n6399 ) | ( n6398 & n6399 ) ;
  assign n6401 = ( n1119 & n6398 ) | ( n1119 & n6399 ) | ( n6398 & n6399 ) ;
  assign n6402 = ( ~n1126 & n6398 ) | ( ~n1126 & n6399 ) | ( n6398 & n6399 ) ;
  assign n6403 = ( ~n1115 & n6401 ) | ( ~n1115 & n6402 ) | ( n6401 & n6402 ) ;
  assign n6404 = ( ~n975 & n6400 ) | ( ~n975 & n6403 ) | ( n6400 & n6403 ) ;
  assign n6405 = ( n1154 & n6400 ) | ( n1154 & n6403 ) | ( n6400 & n6403 ) ;
  assign n6406 = ( ~x409 & n6404 ) | ( ~x409 & n6405 ) | ( n6404 & n6405 ) ;
  assign n6407 = ( x281 & n6404 ) | ( x281 & n6405 ) | ( n6404 & n6405 ) ;
  assign n6408 = ( n656 & n6406 ) | ( n656 & n6407 ) | ( n6406 & n6407 ) ;
  assign n6409 = n6397 | n6408 ;
  assign n6410 = ~n6386 & n6409 ;
  assign n6411 = x438 & n991 ;
  assign n6412 = x438 & ~n995 ;
  assign n6413 = ( ~n1104 & n6411 ) | ( ~n1104 & n6412 ) | ( n6411 & n6412 ) ;
  assign n6414 = ( ~n1119 & n6411 ) | ( ~n1119 & n6412 ) | ( n6411 & n6412 ) ;
  assign n6415 = ( n1126 & n6411 ) | ( n1126 & n6412 ) | ( n6411 & n6412 ) ;
  assign n6416 = ( n1115 & n6414 ) | ( n1115 & n6415 ) | ( n6414 & n6415 ) ;
  assign n6417 = ( n975 & n6413 ) | ( n975 & n6416 ) | ( n6413 & n6416 ) ;
  assign n6418 = ( ~n1154 & n6413 ) | ( ~n1154 & n6416 ) | ( n6413 & n6416 ) ;
  assign n6419 = ( x409 & n6417 ) | ( x409 & n6418 ) | ( n6417 & n6418 ) ;
  assign n6420 = ( ~x281 & n6417 ) | ( ~x281 & n6418 ) | ( n6417 & n6418 ) ;
  assign n6421 = ( ~n656 & n6419 ) | ( ~n656 & n6420 ) | ( n6419 & n6420 ) ;
  assign n6422 = x310 & ~n991 ;
  assign n6423 = x310 & n995 ;
  assign n6424 = ( n1104 & n6422 ) | ( n1104 & n6423 ) | ( n6422 & n6423 ) ;
  assign n6425 = ( n1119 & n6422 ) | ( n1119 & n6423 ) | ( n6422 & n6423 ) ;
  assign n6426 = ( ~n1126 & n6422 ) | ( ~n1126 & n6423 ) | ( n6422 & n6423 ) ;
  assign n6427 = ( ~n1115 & n6425 ) | ( ~n1115 & n6426 ) | ( n6425 & n6426 ) ;
  assign n6428 = ( ~n975 & n6424 ) | ( ~n975 & n6427 ) | ( n6424 & n6427 ) ;
  assign n6429 = ( n1154 & n6424 ) | ( n1154 & n6427 ) | ( n6424 & n6427 ) ;
  assign n6430 = ( ~x409 & n6428 ) | ( ~x409 & n6429 ) | ( n6428 & n6429 ) ;
  assign n6431 = ( x281 & n6428 ) | ( x281 & n6429 ) | ( n6428 & n6429 ) ;
  assign n6432 = ( n656 & n6430 ) | ( n656 & n6431 ) | ( n6430 & n6431 ) ;
  assign n6433 = n6421 | n6432 ;
  assign n6434 = x182 & n1767 ;
  assign n6435 = x182 & ~n1771 ;
  assign n6436 = ( ~n1751 & n6434 ) | ( ~n1751 & n6435 ) | ( n6434 & n6435 ) ;
  assign n6437 = ( ~n1787 & n6434 ) | ( ~n1787 & n6435 ) | ( n6434 & n6435 ) ;
  assign n6438 = ( n1794 & n6434 ) | ( n1794 & n6435 ) | ( n6434 & n6435 ) ;
  assign n6439 = ( n1783 & n6437 ) | ( n1783 & n6438 ) | ( n6437 & n6438 ) ;
  assign n6440 = ( n1643 & n6436 ) | ( n1643 & n6439 ) | ( n6436 & n6439 ) ;
  assign n6441 = ( ~n1822 & n6436 ) | ( ~n1822 & n6439 ) | ( n6436 & n6439 ) ;
  assign n6442 = ( ~n1324 & n6440 ) | ( ~n1324 & n6441 ) | ( n6440 & n6441 ) ;
  assign n6443 = x54 & ~n1767 ;
  assign n6444 = x54 & n1771 ;
  assign n6445 = ( n1751 & n6443 ) | ( n1751 & n6444 ) | ( n6443 & n6444 ) ;
  assign n6446 = ( n1787 & n6443 ) | ( n1787 & n6444 ) | ( n6443 & n6444 ) ;
  assign n6447 = ( ~n1794 & n6443 ) | ( ~n1794 & n6444 ) | ( n6443 & n6444 ) ;
  assign n6448 = ( ~n1783 & n6446 ) | ( ~n1783 & n6447 ) | ( n6446 & n6447 ) ;
  assign n6449 = ( ~n1643 & n6445 ) | ( ~n1643 & n6448 ) | ( n6445 & n6448 ) ;
  assign n6450 = ( n1822 & n6445 ) | ( n1822 & n6448 ) | ( n6445 & n6448 ) ;
  assign n6451 = ( n1324 & n6449 ) | ( n1324 & n6450 ) | ( n6449 & n6450 ) ;
  assign n6452 = n6442 | n6451 ;
  assign n6453 = n6433 & ~n6452 ;
  assign n6454 = n6410 | n6453 ;
  assign n6455 = x181 & n1767 ;
  assign n6456 = x181 & ~n1771 ;
  assign n6457 = ( ~n1751 & n6455 ) | ( ~n1751 & n6456 ) | ( n6455 & n6456 ) ;
  assign n6458 = ( ~n1787 & n6455 ) | ( ~n1787 & n6456 ) | ( n6455 & n6456 ) ;
  assign n6459 = ( n1794 & n6455 ) | ( n1794 & n6456 ) | ( n6455 & n6456 ) ;
  assign n6460 = ( n1783 & n6458 ) | ( n1783 & n6459 ) | ( n6458 & n6459 ) ;
  assign n6461 = ( n1643 & n6457 ) | ( n1643 & n6460 ) | ( n6457 & n6460 ) ;
  assign n6462 = ( ~n1822 & n6457 ) | ( ~n1822 & n6460 ) | ( n6457 & n6460 ) ;
  assign n6463 = ( ~n1324 & n6461 ) | ( ~n1324 & n6462 ) | ( n6461 & n6462 ) ;
  assign n6464 = x53 & ~n1767 ;
  assign n6465 = x53 & n1771 ;
  assign n6466 = ( n1751 & n6464 ) | ( n1751 & n6465 ) | ( n6464 & n6465 ) ;
  assign n6467 = ( n1787 & n6464 ) | ( n1787 & n6465 ) | ( n6464 & n6465 ) ;
  assign n6468 = ( ~n1794 & n6464 ) | ( ~n1794 & n6465 ) | ( n6464 & n6465 ) ;
  assign n6469 = ( ~n1783 & n6467 ) | ( ~n1783 & n6468 ) | ( n6467 & n6468 ) ;
  assign n6470 = ( ~n1643 & n6466 ) | ( ~n1643 & n6469 ) | ( n6466 & n6469 ) ;
  assign n6471 = ( n1822 & n6466 ) | ( n1822 & n6469 ) | ( n6466 & n6469 ) ;
  assign n6472 = ( n1324 & n6470 ) | ( n1324 & n6471 ) | ( n6470 & n6471 ) ;
  assign n6473 = n6463 | n6472 ;
  assign n6474 = x437 & n991 ;
  assign n6475 = x437 & ~n995 ;
  assign n6476 = ( ~n1104 & n6474 ) | ( ~n1104 & n6475 ) | ( n6474 & n6475 ) ;
  assign n6477 = ( ~n1119 & n6474 ) | ( ~n1119 & n6475 ) | ( n6474 & n6475 ) ;
  assign n6478 = ( n1126 & n6474 ) | ( n1126 & n6475 ) | ( n6474 & n6475 ) ;
  assign n6479 = ( n1115 & n6477 ) | ( n1115 & n6478 ) | ( n6477 & n6478 ) ;
  assign n6480 = ( n975 & n6476 ) | ( n975 & n6479 ) | ( n6476 & n6479 ) ;
  assign n6481 = ( ~n1154 & n6476 ) | ( ~n1154 & n6479 ) | ( n6476 & n6479 ) ;
  assign n6482 = ( x409 & n6480 ) | ( x409 & n6481 ) | ( n6480 & n6481 ) ;
  assign n6483 = ( ~x281 & n6480 ) | ( ~x281 & n6481 ) | ( n6480 & n6481 ) ;
  assign n6484 = ( ~n656 & n6482 ) | ( ~n656 & n6483 ) | ( n6482 & n6483 ) ;
  assign n6485 = x309 & ~n991 ;
  assign n6486 = x309 & n995 ;
  assign n6487 = ( n1104 & n6485 ) | ( n1104 & n6486 ) | ( n6485 & n6486 ) ;
  assign n6488 = ( n1119 & n6485 ) | ( n1119 & n6486 ) | ( n6485 & n6486 ) ;
  assign n6489 = ( ~n1126 & n6485 ) | ( ~n1126 & n6486 ) | ( n6485 & n6486 ) ;
  assign n6490 = ( ~n1115 & n6488 ) | ( ~n1115 & n6489 ) | ( n6488 & n6489 ) ;
  assign n6491 = ( ~n975 & n6487 ) | ( ~n975 & n6490 ) | ( n6487 & n6490 ) ;
  assign n6492 = ( n1154 & n6487 ) | ( n1154 & n6490 ) | ( n6487 & n6490 ) ;
  assign n6493 = ( ~x409 & n6491 ) | ( ~x409 & n6492 ) | ( n6491 & n6492 ) ;
  assign n6494 = ( x281 & n6491 ) | ( x281 & n6492 ) | ( n6491 & n6492 ) ;
  assign n6495 = ( n656 & n6493 ) | ( n656 & n6494 ) | ( n6493 & n6494 ) ;
  assign n6496 = n6484 | n6495 ;
  assign n6497 = ~n6473 & n6496 ;
  assign n6498 = x436 & n991 ;
  assign n6499 = x436 & ~n995 ;
  assign n6500 = ( ~n1104 & n6498 ) | ( ~n1104 & n6499 ) | ( n6498 & n6499 ) ;
  assign n6501 = ( ~n1119 & n6498 ) | ( ~n1119 & n6499 ) | ( n6498 & n6499 ) ;
  assign n6502 = ( n1126 & n6498 ) | ( n1126 & n6499 ) | ( n6498 & n6499 ) ;
  assign n6503 = ( n1115 & n6501 ) | ( n1115 & n6502 ) | ( n6501 & n6502 ) ;
  assign n6504 = ( n975 & n6500 ) | ( n975 & n6503 ) | ( n6500 & n6503 ) ;
  assign n6505 = ( ~n1154 & n6500 ) | ( ~n1154 & n6503 ) | ( n6500 & n6503 ) ;
  assign n6506 = ( x409 & n6504 ) | ( x409 & n6505 ) | ( n6504 & n6505 ) ;
  assign n6507 = ( ~x281 & n6504 ) | ( ~x281 & n6505 ) | ( n6504 & n6505 ) ;
  assign n6508 = ( ~n656 & n6506 ) | ( ~n656 & n6507 ) | ( n6506 & n6507 ) ;
  assign n6509 = x308 & ~n991 ;
  assign n6510 = x308 & n995 ;
  assign n6511 = ( n1104 & n6509 ) | ( n1104 & n6510 ) | ( n6509 & n6510 ) ;
  assign n6512 = ( n1119 & n6509 ) | ( n1119 & n6510 ) | ( n6509 & n6510 ) ;
  assign n6513 = ( ~n1126 & n6509 ) | ( ~n1126 & n6510 ) | ( n6509 & n6510 ) ;
  assign n6514 = ( ~n1115 & n6512 ) | ( ~n1115 & n6513 ) | ( n6512 & n6513 ) ;
  assign n6515 = ( ~n975 & n6511 ) | ( ~n975 & n6514 ) | ( n6511 & n6514 ) ;
  assign n6516 = ( n1154 & n6511 ) | ( n1154 & n6514 ) | ( n6511 & n6514 ) ;
  assign n6517 = ( ~x409 & n6515 ) | ( ~x409 & n6516 ) | ( n6515 & n6516 ) ;
  assign n6518 = ( x281 & n6515 ) | ( x281 & n6516 ) | ( n6515 & n6516 ) ;
  assign n6519 = ( n656 & n6517 ) | ( n656 & n6518 ) | ( n6517 & n6518 ) ;
  assign n6520 = n6508 | n6519 ;
  assign n6521 = x180 & n1767 ;
  assign n6522 = x180 & ~n1771 ;
  assign n6523 = ( ~n1751 & n6521 ) | ( ~n1751 & n6522 ) | ( n6521 & n6522 ) ;
  assign n6524 = ( ~n1787 & n6521 ) | ( ~n1787 & n6522 ) | ( n6521 & n6522 ) ;
  assign n6525 = ( n1794 & n6521 ) | ( n1794 & n6522 ) | ( n6521 & n6522 ) ;
  assign n6526 = ( n1783 & n6524 ) | ( n1783 & n6525 ) | ( n6524 & n6525 ) ;
  assign n6527 = ( n1643 & n6523 ) | ( n1643 & n6526 ) | ( n6523 & n6526 ) ;
  assign n6528 = ( ~n1822 & n6523 ) | ( ~n1822 & n6526 ) | ( n6523 & n6526 ) ;
  assign n6529 = ( ~n1324 & n6527 ) | ( ~n1324 & n6528 ) | ( n6527 & n6528 ) ;
  assign n6530 = x52 & ~n1767 ;
  assign n6531 = x52 & n1771 ;
  assign n6532 = ( n1751 & n6530 ) | ( n1751 & n6531 ) | ( n6530 & n6531 ) ;
  assign n6533 = ( n1787 & n6530 ) | ( n1787 & n6531 ) | ( n6530 & n6531 ) ;
  assign n6534 = ( ~n1794 & n6530 ) | ( ~n1794 & n6531 ) | ( n6530 & n6531 ) ;
  assign n6535 = ( ~n1783 & n6533 ) | ( ~n1783 & n6534 ) | ( n6533 & n6534 ) ;
  assign n6536 = ( ~n1643 & n6532 ) | ( ~n1643 & n6535 ) | ( n6532 & n6535 ) ;
  assign n6537 = ( n1822 & n6532 ) | ( n1822 & n6535 ) | ( n6532 & n6535 ) ;
  assign n6538 = ( n1324 & n6536 ) | ( n1324 & n6537 ) | ( n6536 & n6537 ) ;
  assign n6539 = n6529 | n6538 ;
  assign n6540 = n6520 & ~n6539 ;
  assign n6541 = n6497 | n6540 ;
  assign n6542 = n6454 | n6541 ;
  assign n6543 = x177 & n1767 ;
  assign n6544 = x177 & ~n1771 ;
  assign n6545 = ( ~n1751 & n6543 ) | ( ~n1751 & n6544 ) | ( n6543 & n6544 ) ;
  assign n6546 = ( ~n1787 & n6543 ) | ( ~n1787 & n6544 ) | ( n6543 & n6544 ) ;
  assign n6547 = ( n1794 & n6543 ) | ( n1794 & n6544 ) | ( n6543 & n6544 ) ;
  assign n6548 = ( n1783 & n6546 ) | ( n1783 & n6547 ) | ( n6546 & n6547 ) ;
  assign n6549 = ( n1643 & n6545 ) | ( n1643 & n6548 ) | ( n6545 & n6548 ) ;
  assign n6550 = ( ~n1822 & n6545 ) | ( ~n1822 & n6548 ) | ( n6545 & n6548 ) ;
  assign n6551 = ( ~n1324 & n6549 ) | ( ~n1324 & n6550 ) | ( n6549 & n6550 ) ;
  assign n6552 = x49 & ~n1767 ;
  assign n6553 = x49 & n1771 ;
  assign n6554 = ( n1751 & n6552 ) | ( n1751 & n6553 ) | ( n6552 & n6553 ) ;
  assign n6555 = ( n1787 & n6552 ) | ( n1787 & n6553 ) | ( n6552 & n6553 ) ;
  assign n6556 = ( ~n1794 & n6552 ) | ( ~n1794 & n6553 ) | ( n6552 & n6553 ) ;
  assign n6557 = ( ~n1783 & n6555 ) | ( ~n1783 & n6556 ) | ( n6555 & n6556 ) ;
  assign n6558 = ( ~n1643 & n6554 ) | ( ~n1643 & n6557 ) | ( n6554 & n6557 ) ;
  assign n6559 = ( n1822 & n6554 ) | ( n1822 & n6557 ) | ( n6554 & n6557 ) ;
  assign n6560 = ( n1324 & n6558 ) | ( n1324 & n6559 ) | ( n6558 & n6559 ) ;
  assign n6561 = n6551 | n6560 ;
  assign n6562 = x433 & n991 ;
  assign n6563 = x433 & ~n995 ;
  assign n6564 = ( ~n1104 & n6562 ) | ( ~n1104 & n6563 ) | ( n6562 & n6563 ) ;
  assign n6565 = ( ~n1119 & n6562 ) | ( ~n1119 & n6563 ) | ( n6562 & n6563 ) ;
  assign n6566 = ( n1126 & n6562 ) | ( n1126 & n6563 ) | ( n6562 & n6563 ) ;
  assign n6567 = ( n1115 & n6565 ) | ( n1115 & n6566 ) | ( n6565 & n6566 ) ;
  assign n6568 = ( n975 & n6564 ) | ( n975 & n6567 ) | ( n6564 & n6567 ) ;
  assign n6569 = ( ~n1154 & n6564 ) | ( ~n1154 & n6567 ) | ( n6564 & n6567 ) ;
  assign n6570 = ( x409 & n6568 ) | ( x409 & n6569 ) | ( n6568 & n6569 ) ;
  assign n6571 = ( ~x281 & n6568 ) | ( ~x281 & n6569 ) | ( n6568 & n6569 ) ;
  assign n6572 = ( ~n656 & n6570 ) | ( ~n656 & n6571 ) | ( n6570 & n6571 ) ;
  assign n6573 = x305 & ~n991 ;
  assign n6574 = x305 & n995 ;
  assign n6575 = ( n1104 & n6573 ) | ( n1104 & n6574 ) | ( n6573 & n6574 ) ;
  assign n6576 = ( n1119 & n6573 ) | ( n1119 & n6574 ) | ( n6573 & n6574 ) ;
  assign n6577 = ( ~n1126 & n6573 ) | ( ~n1126 & n6574 ) | ( n6573 & n6574 ) ;
  assign n6578 = ( ~n1115 & n6576 ) | ( ~n1115 & n6577 ) | ( n6576 & n6577 ) ;
  assign n6579 = ( ~n975 & n6575 ) | ( ~n975 & n6578 ) | ( n6575 & n6578 ) ;
  assign n6580 = ( n1154 & n6575 ) | ( n1154 & n6578 ) | ( n6575 & n6578 ) ;
  assign n6581 = ( ~x409 & n6579 ) | ( ~x409 & n6580 ) | ( n6579 & n6580 ) ;
  assign n6582 = ( x281 & n6579 ) | ( x281 & n6580 ) | ( n6579 & n6580 ) ;
  assign n6583 = ( n656 & n6581 ) | ( n656 & n6582 ) | ( n6581 & n6582 ) ;
  assign n6584 = n6572 | n6583 ;
  assign n6585 = ~n6561 & n6584 ;
  assign n6586 = x179 & n1767 ;
  assign n6587 = x179 & ~n1771 ;
  assign n6588 = ( ~n1751 & n6586 ) | ( ~n1751 & n6587 ) | ( n6586 & n6587 ) ;
  assign n6589 = ( ~n1787 & n6586 ) | ( ~n1787 & n6587 ) | ( n6586 & n6587 ) ;
  assign n6590 = ( n1794 & n6586 ) | ( n1794 & n6587 ) | ( n6586 & n6587 ) ;
  assign n6591 = ( n1783 & n6589 ) | ( n1783 & n6590 ) | ( n6589 & n6590 ) ;
  assign n6592 = ( n1643 & n6588 ) | ( n1643 & n6591 ) | ( n6588 & n6591 ) ;
  assign n6593 = ( ~n1822 & n6588 ) | ( ~n1822 & n6591 ) | ( n6588 & n6591 ) ;
  assign n6594 = ( ~n1324 & n6592 ) | ( ~n1324 & n6593 ) | ( n6592 & n6593 ) ;
  assign n6595 = x51 & ~n1767 ;
  assign n6596 = x51 & n1771 ;
  assign n6597 = ( n1751 & n6595 ) | ( n1751 & n6596 ) | ( n6595 & n6596 ) ;
  assign n6598 = ( n1787 & n6595 ) | ( n1787 & n6596 ) | ( n6595 & n6596 ) ;
  assign n6599 = ( ~n1794 & n6595 ) | ( ~n1794 & n6596 ) | ( n6595 & n6596 ) ;
  assign n6600 = ( ~n1783 & n6598 ) | ( ~n1783 & n6599 ) | ( n6598 & n6599 ) ;
  assign n6601 = ( ~n1643 & n6597 ) | ( ~n1643 & n6600 ) | ( n6597 & n6600 ) ;
  assign n6602 = ( n1822 & n6597 ) | ( n1822 & n6600 ) | ( n6597 & n6600 ) ;
  assign n6603 = ( n1324 & n6601 ) | ( n1324 & n6602 ) | ( n6601 & n6602 ) ;
  assign n6604 = n6594 | n6603 ;
  assign n6605 = x435 & n991 ;
  assign n6606 = x435 & ~n995 ;
  assign n6607 = ( ~n1104 & n6605 ) | ( ~n1104 & n6606 ) | ( n6605 & n6606 ) ;
  assign n6608 = ( ~n1119 & n6605 ) | ( ~n1119 & n6606 ) | ( n6605 & n6606 ) ;
  assign n6609 = ( n1126 & n6605 ) | ( n1126 & n6606 ) | ( n6605 & n6606 ) ;
  assign n6610 = ( n1115 & n6608 ) | ( n1115 & n6609 ) | ( n6608 & n6609 ) ;
  assign n6611 = ( n975 & n6607 ) | ( n975 & n6610 ) | ( n6607 & n6610 ) ;
  assign n6612 = ( ~n1154 & n6607 ) | ( ~n1154 & n6610 ) | ( n6607 & n6610 ) ;
  assign n6613 = ( x409 & n6611 ) | ( x409 & n6612 ) | ( n6611 & n6612 ) ;
  assign n6614 = ( ~x281 & n6611 ) | ( ~x281 & n6612 ) | ( n6611 & n6612 ) ;
  assign n6615 = ( ~n656 & n6613 ) | ( ~n656 & n6614 ) | ( n6613 & n6614 ) ;
  assign n6616 = x307 & ~n991 ;
  assign n6617 = x307 & n995 ;
  assign n6618 = ( n1104 & n6616 ) | ( n1104 & n6617 ) | ( n6616 & n6617 ) ;
  assign n6619 = ( n1119 & n6616 ) | ( n1119 & n6617 ) | ( n6616 & n6617 ) ;
  assign n6620 = ( ~n1126 & n6616 ) | ( ~n1126 & n6617 ) | ( n6616 & n6617 ) ;
  assign n6621 = ( ~n1115 & n6619 ) | ( ~n1115 & n6620 ) | ( n6619 & n6620 ) ;
  assign n6622 = ( ~n975 & n6618 ) | ( ~n975 & n6621 ) | ( n6618 & n6621 ) ;
  assign n6623 = ( n1154 & n6618 ) | ( n1154 & n6621 ) | ( n6618 & n6621 ) ;
  assign n6624 = ( ~x409 & n6622 ) | ( ~x409 & n6623 ) | ( n6622 & n6623 ) ;
  assign n6625 = ( x281 & n6622 ) | ( x281 & n6623 ) | ( n6622 & n6623 ) ;
  assign n6626 = ( n656 & n6624 ) | ( n656 & n6625 ) | ( n6624 & n6625 ) ;
  assign n6627 = n6615 | n6626 ;
  assign n6628 = ~n6604 & n6627 ;
  assign n6629 = x434 & n991 ;
  assign n6630 = x434 & ~n995 ;
  assign n6631 = ( ~n1104 & n6629 ) | ( ~n1104 & n6630 ) | ( n6629 & n6630 ) ;
  assign n6632 = ( ~n1119 & n6629 ) | ( ~n1119 & n6630 ) | ( n6629 & n6630 ) ;
  assign n6633 = ( n1126 & n6629 ) | ( n1126 & n6630 ) | ( n6629 & n6630 ) ;
  assign n6634 = ( n1115 & n6632 ) | ( n1115 & n6633 ) | ( n6632 & n6633 ) ;
  assign n6635 = ( n975 & n6631 ) | ( n975 & n6634 ) | ( n6631 & n6634 ) ;
  assign n6636 = ( ~n1154 & n6631 ) | ( ~n1154 & n6634 ) | ( n6631 & n6634 ) ;
  assign n6637 = ( x409 & n6635 ) | ( x409 & n6636 ) | ( n6635 & n6636 ) ;
  assign n6638 = ( ~x281 & n6635 ) | ( ~x281 & n6636 ) | ( n6635 & n6636 ) ;
  assign n6639 = ( ~n656 & n6637 ) | ( ~n656 & n6638 ) | ( n6637 & n6638 ) ;
  assign n6640 = x306 & ~n991 ;
  assign n6641 = x306 & n995 ;
  assign n6642 = ( n1104 & n6640 ) | ( n1104 & n6641 ) | ( n6640 & n6641 ) ;
  assign n6643 = ( n1119 & n6640 ) | ( n1119 & n6641 ) | ( n6640 & n6641 ) ;
  assign n6644 = ( ~n1126 & n6640 ) | ( ~n1126 & n6641 ) | ( n6640 & n6641 ) ;
  assign n6645 = ( ~n1115 & n6643 ) | ( ~n1115 & n6644 ) | ( n6643 & n6644 ) ;
  assign n6646 = ( ~n975 & n6642 ) | ( ~n975 & n6645 ) | ( n6642 & n6645 ) ;
  assign n6647 = ( n1154 & n6642 ) | ( n1154 & n6645 ) | ( n6642 & n6645 ) ;
  assign n6648 = ( ~x409 & n6646 ) | ( ~x409 & n6647 ) | ( n6646 & n6647 ) ;
  assign n6649 = ( x281 & n6646 ) | ( x281 & n6647 ) | ( n6646 & n6647 ) ;
  assign n6650 = ( n656 & n6648 ) | ( n656 & n6649 ) | ( n6648 & n6649 ) ;
  assign n6651 = n6639 | n6650 ;
  assign n6652 = x178 & n1767 ;
  assign n6653 = x178 & ~n1771 ;
  assign n6654 = ( ~n1751 & n6652 ) | ( ~n1751 & n6653 ) | ( n6652 & n6653 ) ;
  assign n6655 = ( ~n1787 & n6652 ) | ( ~n1787 & n6653 ) | ( n6652 & n6653 ) ;
  assign n6656 = ( n1794 & n6652 ) | ( n1794 & n6653 ) | ( n6652 & n6653 ) ;
  assign n6657 = ( n1783 & n6655 ) | ( n1783 & n6656 ) | ( n6655 & n6656 ) ;
  assign n6658 = ( n1643 & n6654 ) | ( n1643 & n6657 ) | ( n6654 & n6657 ) ;
  assign n6659 = ( ~n1822 & n6654 ) | ( ~n1822 & n6657 ) | ( n6654 & n6657 ) ;
  assign n6660 = ( ~n1324 & n6658 ) | ( ~n1324 & n6659 ) | ( n6658 & n6659 ) ;
  assign n6661 = x50 & ~n1767 ;
  assign n6662 = x50 & n1771 ;
  assign n6663 = ( n1751 & n6661 ) | ( n1751 & n6662 ) | ( n6661 & n6662 ) ;
  assign n6664 = ( n1787 & n6661 ) | ( n1787 & n6662 ) | ( n6661 & n6662 ) ;
  assign n6665 = ( ~n1794 & n6661 ) | ( ~n1794 & n6662 ) | ( n6661 & n6662 ) ;
  assign n6666 = ( ~n1783 & n6664 ) | ( ~n1783 & n6665 ) | ( n6664 & n6665 ) ;
  assign n6667 = ( ~n1643 & n6663 ) | ( ~n1643 & n6666 ) | ( n6663 & n6666 ) ;
  assign n6668 = ( n1822 & n6663 ) | ( n1822 & n6666 ) | ( n6663 & n6666 ) ;
  assign n6669 = ( n1324 & n6667 ) | ( n1324 & n6668 ) | ( n6667 & n6668 ) ;
  assign n6670 = n6660 | n6669 ;
  assign n6671 = n6651 & ~n6670 ;
  assign n6672 = n6628 | n6671 ;
  assign n6673 = n6585 | n6672 ;
  assign n6674 = ~n6651 & n6670 ;
  assign n6675 = ~n6628 & n6674 ;
  assign n6676 = x432 & n991 ;
  assign n6677 = x432 & ~n995 ;
  assign n6678 = ( ~n1104 & n6676 ) | ( ~n1104 & n6677 ) | ( n6676 & n6677 ) ;
  assign n6679 = ( ~n1119 & n6676 ) | ( ~n1119 & n6677 ) | ( n6676 & n6677 ) ;
  assign n6680 = ( n1126 & n6676 ) | ( n1126 & n6677 ) | ( n6676 & n6677 ) ;
  assign n6681 = ( n1115 & n6679 ) | ( n1115 & n6680 ) | ( n6679 & n6680 ) ;
  assign n6682 = ( n975 & n6678 ) | ( n975 & n6681 ) | ( n6678 & n6681 ) ;
  assign n6683 = ( ~n1154 & n6678 ) | ( ~n1154 & n6681 ) | ( n6678 & n6681 ) ;
  assign n6684 = ( x409 & n6682 ) | ( x409 & n6683 ) | ( n6682 & n6683 ) ;
  assign n6685 = ( ~x281 & n6682 ) | ( ~x281 & n6683 ) | ( n6682 & n6683 ) ;
  assign n6686 = ( ~n656 & n6684 ) | ( ~n656 & n6685 ) | ( n6684 & n6685 ) ;
  assign n6687 = x304 & ~n991 ;
  assign n6688 = x304 & n995 ;
  assign n6689 = ( n1104 & n6687 ) | ( n1104 & n6688 ) | ( n6687 & n6688 ) ;
  assign n6690 = ( n1119 & n6687 ) | ( n1119 & n6688 ) | ( n6687 & n6688 ) ;
  assign n6691 = ( ~n1126 & n6687 ) | ( ~n1126 & n6688 ) | ( n6687 & n6688 ) ;
  assign n6692 = ( ~n1115 & n6690 ) | ( ~n1115 & n6691 ) | ( n6690 & n6691 ) ;
  assign n6693 = ( ~n975 & n6689 ) | ( ~n975 & n6692 ) | ( n6689 & n6692 ) ;
  assign n6694 = ( n1154 & n6689 ) | ( n1154 & n6692 ) | ( n6689 & n6692 ) ;
  assign n6695 = ( ~x409 & n6693 ) | ( ~x409 & n6694 ) | ( n6693 & n6694 ) ;
  assign n6696 = ( x281 & n6693 ) | ( x281 & n6694 ) | ( n6693 & n6694 ) ;
  assign n6697 = ( n656 & n6695 ) | ( n656 & n6696 ) | ( n6695 & n6696 ) ;
  assign n6698 = n6686 | n6697 ;
  assign n6699 = x176 & n1767 ;
  assign n6700 = x176 & ~n1771 ;
  assign n6701 = ( ~n1751 & n6699 ) | ( ~n1751 & n6700 ) | ( n6699 & n6700 ) ;
  assign n6702 = ( ~n1787 & n6699 ) | ( ~n1787 & n6700 ) | ( n6699 & n6700 ) ;
  assign n6703 = ( n1794 & n6699 ) | ( n1794 & n6700 ) | ( n6699 & n6700 ) ;
  assign n6704 = ( n1783 & n6702 ) | ( n1783 & n6703 ) | ( n6702 & n6703 ) ;
  assign n6705 = ( n1643 & n6701 ) | ( n1643 & n6704 ) | ( n6701 & n6704 ) ;
  assign n6706 = ( ~n1822 & n6701 ) | ( ~n1822 & n6704 ) | ( n6701 & n6704 ) ;
  assign n6707 = ( ~n1324 & n6705 ) | ( ~n1324 & n6706 ) | ( n6705 & n6706 ) ;
  assign n6708 = x48 & ~n1767 ;
  assign n6709 = x48 & n1771 ;
  assign n6710 = ( n1751 & n6708 ) | ( n1751 & n6709 ) | ( n6708 & n6709 ) ;
  assign n6711 = ( n1787 & n6708 ) | ( n1787 & n6709 ) | ( n6708 & n6709 ) ;
  assign n6712 = ( ~n1794 & n6708 ) | ( ~n1794 & n6709 ) | ( n6708 & n6709 ) ;
  assign n6713 = ( ~n1783 & n6711 ) | ( ~n1783 & n6712 ) | ( n6711 & n6712 ) ;
  assign n6714 = ( ~n1643 & n6710 ) | ( ~n1643 & n6713 ) | ( n6710 & n6713 ) ;
  assign n6715 = ( n1822 & n6710 ) | ( n1822 & n6713 ) | ( n6710 & n6713 ) ;
  assign n6716 = ( n1324 & n6714 ) | ( n1324 & n6715 ) | ( n6714 & n6715 ) ;
  assign n6717 = n6707 | n6716 ;
  assign n6718 = ~n6698 & n6717 ;
  assign n6719 = n6561 & ~n6584 ;
  assign n6720 = n6718 | n6719 ;
  assign n6721 = n6675 | n6720 ;
  assign n6722 = ( ~n6673 & n6675 ) | ( ~n6673 & n6721 ) | ( n6675 & n6721 ) ;
  assign n6723 = n6604 & ~n6627 ;
  assign n6724 = ~n6542 & n6723 ;
  assign n6725 = ( ~n6542 & n6722 ) | ( ~n6542 & n6724 ) | ( n6722 & n6724 ) ;
  assign n6726 = ~n6520 & n6539 ;
  assign n6727 = ( n6473 & ~n6496 ) | ( n6473 & n6726 ) | ( ~n6496 & n6726 ) ;
  assign n6728 = ~n6433 & n6452 ;
  assign n6729 = ~n6453 & n6728 ;
  assign n6730 = ( ~n6453 & n6727 ) | ( ~n6453 & n6729 ) | ( n6727 & n6729 ) ;
  assign n6731 = ( n6386 & ~n6409 ) | ( n6386 & n6730 ) | ( ~n6409 & n6730 ) ;
  assign n6732 = n6725 | n6731 ;
  assign n6733 = n6542 | n6673 ;
  assign n6734 = n6698 & ~n6717 ;
  assign n6735 = n6733 | n6734 ;
  assign n6736 = ~n6732 & n6735 ;
  assign n6737 = x175 & n1767 ;
  assign n6738 = x175 & ~n1771 ;
  assign n6739 = ( ~n1751 & n6737 ) | ( ~n1751 & n6738 ) | ( n6737 & n6738 ) ;
  assign n6740 = ( ~n1787 & n6737 ) | ( ~n1787 & n6738 ) | ( n6737 & n6738 ) ;
  assign n6741 = ( n1794 & n6737 ) | ( n1794 & n6738 ) | ( n6737 & n6738 ) ;
  assign n6742 = ( n1783 & n6740 ) | ( n1783 & n6741 ) | ( n6740 & n6741 ) ;
  assign n6743 = ( n1643 & n6739 ) | ( n1643 & n6742 ) | ( n6739 & n6742 ) ;
  assign n6744 = ( ~n1822 & n6739 ) | ( ~n1822 & n6742 ) | ( n6739 & n6742 ) ;
  assign n6745 = ( ~n1324 & n6743 ) | ( ~n1324 & n6744 ) | ( n6743 & n6744 ) ;
  assign n6746 = x47 & ~n1767 ;
  assign n6747 = x47 & n1771 ;
  assign n6748 = ( n1751 & n6746 ) | ( n1751 & n6747 ) | ( n6746 & n6747 ) ;
  assign n6749 = ( n1787 & n6746 ) | ( n1787 & n6747 ) | ( n6746 & n6747 ) ;
  assign n6750 = ( ~n1794 & n6746 ) | ( ~n1794 & n6747 ) | ( n6746 & n6747 ) ;
  assign n6751 = ( ~n1783 & n6749 ) | ( ~n1783 & n6750 ) | ( n6749 & n6750 ) ;
  assign n6752 = ( ~n1643 & n6748 ) | ( ~n1643 & n6751 ) | ( n6748 & n6751 ) ;
  assign n6753 = ( n1822 & n6748 ) | ( n1822 & n6751 ) | ( n6748 & n6751 ) ;
  assign n6754 = ( n1324 & n6752 ) | ( n1324 & n6753 ) | ( n6752 & n6753 ) ;
  assign n6755 = n6745 | n6754 ;
  assign n6756 = x431 & n991 ;
  assign n6757 = x431 & ~n995 ;
  assign n6758 = ( ~n1104 & n6756 ) | ( ~n1104 & n6757 ) | ( n6756 & n6757 ) ;
  assign n6759 = ( ~n1119 & n6756 ) | ( ~n1119 & n6757 ) | ( n6756 & n6757 ) ;
  assign n6760 = ( n1126 & n6756 ) | ( n1126 & n6757 ) | ( n6756 & n6757 ) ;
  assign n6761 = ( n1115 & n6759 ) | ( n1115 & n6760 ) | ( n6759 & n6760 ) ;
  assign n6762 = ( n975 & n6758 ) | ( n975 & n6761 ) | ( n6758 & n6761 ) ;
  assign n6763 = ( ~n1154 & n6758 ) | ( ~n1154 & n6761 ) | ( n6758 & n6761 ) ;
  assign n6764 = ( x409 & n6762 ) | ( x409 & n6763 ) | ( n6762 & n6763 ) ;
  assign n6765 = ( ~x281 & n6762 ) | ( ~x281 & n6763 ) | ( n6762 & n6763 ) ;
  assign n6766 = ( ~n656 & n6764 ) | ( ~n656 & n6765 ) | ( n6764 & n6765 ) ;
  assign n6767 = x303 & ~n991 ;
  assign n6768 = x303 & n995 ;
  assign n6769 = ( n1104 & n6767 ) | ( n1104 & n6768 ) | ( n6767 & n6768 ) ;
  assign n6770 = ( n1119 & n6767 ) | ( n1119 & n6768 ) | ( n6767 & n6768 ) ;
  assign n6771 = ( ~n1126 & n6767 ) | ( ~n1126 & n6768 ) | ( n6767 & n6768 ) ;
  assign n6772 = ( ~n1115 & n6770 ) | ( ~n1115 & n6771 ) | ( n6770 & n6771 ) ;
  assign n6773 = ( ~n975 & n6769 ) | ( ~n975 & n6772 ) | ( n6769 & n6772 ) ;
  assign n6774 = ( n1154 & n6769 ) | ( n1154 & n6772 ) | ( n6769 & n6772 ) ;
  assign n6775 = ( ~x409 & n6773 ) | ( ~x409 & n6774 ) | ( n6773 & n6774 ) ;
  assign n6776 = ( x281 & n6773 ) | ( x281 & n6774 ) | ( n6773 & n6774 ) ;
  assign n6777 = ( n656 & n6775 ) | ( n656 & n6776 ) | ( n6775 & n6776 ) ;
  assign n6778 = n6766 | n6777 ;
  assign n6779 = ~n6755 & n6778 ;
  assign n6780 = x430 & n991 ;
  assign n6781 = x430 & ~n995 ;
  assign n6782 = ( ~n1104 & n6780 ) | ( ~n1104 & n6781 ) | ( n6780 & n6781 ) ;
  assign n6783 = ( ~n1119 & n6780 ) | ( ~n1119 & n6781 ) | ( n6780 & n6781 ) ;
  assign n6784 = ( n1126 & n6780 ) | ( n1126 & n6781 ) | ( n6780 & n6781 ) ;
  assign n6785 = ( n1115 & n6783 ) | ( n1115 & n6784 ) | ( n6783 & n6784 ) ;
  assign n6786 = ( n975 & n6782 ) | ( n975 & n6785 ) | ( n6782 & n6785 ) ;
  assign n6787 = ( ~n1154 & n6782 ) | ( ~n1154 & n6785 ) | ( n6782 & n6785 ) ;
  assign n6788 = ( x409 & n6786 ) | ( x409 & n6787 ) | ( n6786 & n6787 ) ;
  assign n6789 = ( ~x281 & n6786 ) | ( ~x281 & n6787 ) | ( n6786 & n6787 ) ;
  assign n6790 = ( ~n656 & n6788 ) | ( ~n656 & n6789 ) | ( n6788 & n6789 ) ;
  assign n6791 = x302 & ~n991 ;
  assign n6792 = x302 & n995 ;
  assign n6793 = ( n1104 & n6791 ) | ( n1104 & n6792 ) | ( n6791 & n6792 ) ;
  assign n6794 = ( n1119 & n6791 ) | ( n1119 & n6792 ) | ( n6791 & n6792 ) ;
  assign n6795 = ( ~n1126 & n6791 ) | ( ~n1126 & n6792 ) | ( n6791 & n6792 ) ;
  assign n6796 = ( ~n1115 & n6794 ) | ( ~n1115 & n6795 ) | ( n6794 & n6795 ) ;
  assign n6797 = ( ~n975 & n6793 ) | ( ~n975 & n6796 ) | ( n6793 & n6796 ) ;
  assign n6798 = ( n1154 & n6793 ) | ( n1154 & n6796 ) | ( n6793 & n6796 ) ;
  assign n6799 = ( ~x409 & n6797 ) | ( ~x409 & n6798 ) | ( n6797 & n6798 ) ;
  assign n6800 = ( x281 & n6797 ) | ( x281 & n6798 ) | ( n6797 & n6798 ) ;
  assign n6801 = ( n656 & n6799 ) | ( n656 & n6800 ) | ( n6799 & n6800 ) ;
  assign n6802 = n6790 | n6801 ;
  assign n6803 = x174 & n1767 ;
  assign n6804 = x174 & ~n1771 ;
  assign n6805 = ( ~n1751 & n6803 ) | ( ~n1751 & n6804 ) | ( n6803 & n6804 ) ;
  assign n6806 = ( ~n1787 & n6803 ) | ( ~n1787 & n6804 ) | ( n6803 & n6804 ) ;
  assign n6807 = ( n1794 & n6803 ) | ( n1794 & n6804 ) | ( n6803 & n6804 ) ;
  assign n6808 = ( n1783 & n6806 ) | ( n1783 & n6807 ) | ( n6806 & n6807 ) ;
  assign n6809 = ( n1643 & n6805 ) | ( n1643 & n6808 ) | ( n6805 & n6808 ) ;
  assign n6810 = ( ~n1822 & n6805 ) | ( ~n1822 & n6808 ) | ( n6805 & n6808 ) ;
  assign n6811 = ( ~n1324 & n6809 ) | ( ~n1324 & n6810 ) | ( n6809 & n6810 ) ;
  assign n6812 = x46 & ~n1767 ;
  assign n6813 = x46 & n1771 ;
  assign n6814 = ( n1751 & n6812 ) | ( n1751 & n6813 ) | ( n6812 & n6813 ) ;
  assign n6815 = ( n1787 & n6812 ) | ( n1787 & n6813 ) | ( n6812 & n6813 ) ;
  assign n6816 = ( ~n1794 & n6812 ) | ( ~n1794 & n6813 ) | ( n6812 & n6813 ) ;
  assign n6817 = ( ~n1783 & n6815 ) | ( ~n1783 & n6816 ) | ( n6815 & n6816 ) ;
  assign n6818 = ( ~n1643 & n6814 ) | ( ~n1643 & n6817 ) | ( n6814 & n6817 ) ;
  assign n6819 = ( n1822 & n6814 ) | ( n1822 & n6817 ) | ( n6814 & n6817 ) ;
  assign n6820 = ( n1324 & n6818 ) | ( n1324 & n6819 ) | ( n6818 & n6819 ) ;
  assign n6821 = n6811 | n6820 ;
  assign n6822 = n6802 & ~n6821 ;
  assign n6823 = n6779 | n6822 ;
  assign n6824 = x172 & n1767 ;
  assign n6825 = x172 & ~n1771 ;
  assign n6826 = ( ~n1751 & n6824 ) | ( ~n1751 & n6825 ) | ( n6824 & n6825 ) ;
  assign n6827 = ( ~n1787 & n6824 ) | ( ~n1787 & n6825 ) | ( n6824 & n6825 ) ;
  assign n6828 = ( n1794 & n6824 ) | ( n1794 & n6825 ) | ( n6824 & n6825 ) ;
  assign n6829 = ( n1783 & n6827 ) | ( n1783 & n6828 ) | ( n6827 & n6828 ) ;
  assign n6830 = ( n1643 & n6826 ) | ( n1643 & n6829 ) | ( n6826 & n6829 ) ;
  assign n6831 = ( ~n1822 & n6826 ) | ( ~n1822 & n6829 ) | ( n6826 & n6829 ) ;
  assign n6832 = ( ~n1324 & n6830 ) | ( ~n1324 & n6831 ) | ( n6830 & n6831 ) ;
  assign n6833 = x44 & ~n1767 ;
  assign n6834 = x44 & n1771 ;
  assign n6835 = ( n1751 & n6833 ) | ( n1751 & n6834 ) | ( n6833 & n6834 ) ;
  assign n6836 = ( n1787 & n6833 ) | ( n1787 & n6834 ) | ( n6833 & n6834 ) ;
  assign n6837 = ( ~n1794 & n6833 ) | ( ~n1794 & n6834 ) | ( n6833 & n6834 ) ;
  assign n6838 = ( ~n1783 & n6836 ) | ( ~n1783 & n6837 ) | ( n6836 & n6837 ) ;
  assign n6839 = ( ~n1643 & n6835 ) | ( ~n1643 & n6838 ) | ( n6835 & n6838 ) ;
  assign n6840 = ( n1822 & n6835 ) | ( n1822 & n6838 ) | ( n6835 & n6838 ) ;
  assign n6841 = ( n1324 & n6839 ) | ( n1324 & n6840 ) | ( n6839 & n6840 ) ;
  assign n6842 = n6832 | n6841 ;
  assign n6843 = x428 & n991 ;
  assign n6844 = x428 & ~n995 ;
  assign n6845 = ( ~n1104 & n6843 ) | ( ~n1104 & n6844 ) | ( n6843 & n6844 ) ;
  assign n6846 = ( ~n1119 & n6843 ) | ( ~n1119 & n6844 ) | ( n6843 & n6844 ) ;
  assign n6847 = ( n1126 & n6843 ) | ( n1126 & n6844 ) | ( n6843 & n6844 ) ;
  assign n6848 = ( n1115 & n6846 ) | ( n1115 & n6847 ) | ( n6846 & n6847 ) ;
  assign n6849 = ( n975 & n6845 ) | ( n975 & n6848 ) | ( n6845 & n6848 ) ;
  assign n6850 = ( ~n1154 & n6845 ) | ( ~n1154 & n6848 ) | ( n6845 & n6848 ) ;
  assign n6851 = ( x409 & n6849 ) | ( x409 & n6850 ) | ( n6849 & n6850 ) ;
  assign n6852 = ( ~x281 & n6849 ) | ( ~x281 & n6850 ) | ( n6849 & n6850 ) ;
  assign n6853 = ( ~n656 & n6851 ) | ( ~n656 & n6852 ) | ( n6851 & n6852 ) ;
  assign n6854 = x300 & ~n991 ;
  assign n6855 = x300 & n995 ;
  assign n6856 = ( n1104 & n6854 ) | ( n1104 & n6855 ) | ( n6854 & n6855 ) ;
  assign n6857 = ( n1119 & n6854 ) | ( n1119 & n6855 ) | ( n6854 & n6855 ) ;
  assign n6858 = ( ~n1126 & n6854 ) | ( ~n1126 & n6855 ) | ( n6854 & n6855 ) ;
  assign n6859 = ( ~n1115 & n6857 ) | ( ~n1115 & n6858 ) | ( n6857 & n6858 ) ;
  assign n6860 = ( ~n975 & n6856 ) | ( ~n975 & n6859 ) | ( n6856 & n6859 ) ;
  assign n6861 = ( n1154 & n6856 ) | ( n1154 & n6859 ) | ( n6856 & n6859 ) ;
  assign n6862 = ( ~x409 & n6860 ) | ( ~x409 & n6861 ) | ( n6860 & n6861 ) ;
  assign n6863 = ( x281 & n6860 ) | ( x281 & n6861 ) | ( n6860 & n6861 ) ;
  assign n6864 = ( n656 & n6862 ) | ( n656 & n6863 ) | ( n6862 & n6863 ) ;
  assign n6865 = n6853 | n6864 ;
  assign n6866 = ~n6842 & n6865 ;
  assign n6867 = x173 & n1767 ;
  assign n6868 = x173 & ~n1771 ;
  assign n6869 = ( ~n1751 & n6867 ) | ( ~n1751 & n6868 ) | ( n6867 & n6868 ) ;
  assign n6870 = ( ~n1787 & n6867 ) | ( ~n1787 & n6868 ) | ( n6867 & n6868 ) ;
  assign n6871 = ( n1794 & n6867 ) | ( n1794 & n6868 ) | ( n6867 & n6868 ) ;
  assign n6872 = ( n1783 & n6870 ) | ( n1783 & n6871 ) | ( n6870 & n6871 ) ;
  assign n6873 = ( n1643 & n6869 ) | ( n1643 & n6872 ) | ( n6869 & n6872 ) ;
  assign n6874 = ( ~n1822 & n6869 ) | ( ~n1822 & n6872 ) | ( n6869 & n6872 ) ;
  assign n6875 = ( ~n1324 & n6873 ) | ( ~n1324 & n6874 ) | ( n6873 & n6874 ) ;
  assign n6876 = x45 & ~n1767 ;
  assign n6877 = x45 & n1771 ;
  assign n6878 = ( n1751 & n6876 ) | ( n1751 & n6877 ) | ( n6876 & n6877 ) ;
  assign n6879 = ( n1787 & n6876 ) | ( n1787 & n6877 ) | ( n6876 & n6877 ) ;
  assign n6880 = ( ~n1794 & n6876 ) | ( ~n1794 & n6877 ) | ( n6876 & n6877 ) ;
  assign n6881 = ( ~n1783 & n6879 ) | ( ~n1783 & n6880 ) | ( n6879 & n6880 ) ;
  assign n6882 = ( ~n1643 & n6878 ) | ( ~n1643 & n6881 ) | ( n6878 & n6881 ) ;
  assign n6883 = ( n1822 & n6878 ) | ( n1822 & n6881 ) | ( n6878 & n6881 ) ;
  assign n6884 = ( n1324 & n6882 ) | ( n1324 & n6883 ) | ( n6882 & n6883 ) ;
  assign n6885 = n6875 | n6884 ;
  assign n6886 = x429 & n991 ;
  assign n6887 = x429 & ~n995 ;
  assign n6888 = ( ~n1104 & n6886 ) | ( ~n1104 & n6887 ) | ( n6886 & n6887 ) ;
  assign n6889 = ( ~n1119 & n6886 ) | ( ~n1119 & n6887 ) | ( n6886 & n6887 ) ;
  assign n6890 = ( n1126 & n6886 ) | ( n1126 & n6887 ) | ( n6886 & n6887 ) ;
  assign n6891 = ( n1115 & n6889 ) | ( n1115 & n6890 ) | ( n6889 & n6890 ) ;
  assign n6892 = ( n975 & n6888 ) | ( n975 & n6891 ) | ( n6888 & n6891 ) ;
  assign n6893 = ( ~n1154 & n6888 ) | ( ~n1154 & n6891 ) | ( n6888 & n6891 ) ;
  assign n6894 = ( x409 & n6892 ) | ( x409 & n6893 ) | ( n6892 & n6893 ) ;
  assign n6895 = ( ~x281 & n6892 ) | ( ~x281 & n6893 ) | ( n6892 & n6893 ) ;
  assign n6896 = ( ~n656 & n6894 ) | ( ~n656 & n6895 ) | ( n6894 & n6895 ) ;
  assign n6897 = x301 & ~n991 ;
  assign n6898 = x301 & n995 ;
  assign n6899 = ( n1104 & n6897 ) | ( n1104 & n6898 ) | ( n6897 & n6898 ) ;
  assign n6900 = ( n1119 & n6897 ) | ( n1119 & n6898 ) | ( n6897 & n6898 ) ;
  assign n6901 = ( ~n1126 & n6897 ) | ( ~n1126 & n6898 ) | ( n6897 & n6898 ) ;
  assign n6902 = ( ~n1115 & n6900 ) | ( ~n1115 & n6901 ) | ( n6900 & n6901 ) ;
  assign n6903 = ( ~n975 & n6899 ) | ( ~n975 & n6902 ) | ( n6899 & n6902 ) ;
  assign n6904 = ( n1154 & n6899 ) | ( n1154 & n6902 ) | ( n6899 & n6902 ) ;
  assign n6905 = ( ~x409 & n6903 ) | ( ~x409 & n6904 ) | ( n6903 & n6904 ) ;
  assign n6906 = ( x281 & n6903 ) | ( x281 & n6904 ) | ( n6903 & n6904 ) ;
  assign n6907 = ( n656 & n6905 ) | ( n656 & n6906 ) | ( n6905 & n6906 ) ;
  assign n6908 = n6896 | n6907 ;
  assign n6909 = ~n6885 & n6908 ;
  assign n6910 = n6866 | n6909 ;
  assign n6911 = n6823 | n6910 ;
  assign n6912 = x170 & n1767 ;
  assign n6913 = x170 & ~n1771 ;
  assign n6914 = ( ~n1751 & n6912 ) | ( ~n1751 & n6913 ) | ( n6912 & n6913 ) ;
  assign n6915 = ( ~n1787 & n6912 ) | ( ~n1787 & n6913 ) | ( n6912 & n6913 ) ;
  assign n6916 = ( n1794 & n6912 ) | ( n1794 & n6913 ) | ( n6912 & n6913 ) ;
  assign n6917 = ( n1783 & n6915 ) | ( n1783 & n6916 ) | ( n6915 & n6916 ) ;
  assign n6918 = ( n1643 & n6914 ) | ( n1643 & n6917 ) | ( n6914 & n6917 ) ;
  assign n6919 = ( ~n1822 & n6914 ) | ( ~n1822 & n6917 ) | ( n6914 & n6917 ) ;
  assign n6920 = ( ~n1324 & n6918 ) | ( ~n1324 & n6919 ) | ( n6918 & n6919 ) ;
  assign n6921 = x42 & ~n1767 ;
  assign n6922 = x42 & n1771 ;
  assign n6923 = ( n1751 & n6921 ) | ( n1751 & n6922 ) | ( n6921 & n6922 ) ;
  assign n6924 = ( n1787 & n6921 ) | ( n1787 & n6922 ) | ( n6921 & n6922 ) ;
  assign n6925 = ( ~n1794 & n6921 ) | ( ~n1794 & n6922 ) | ( n6921 & n6922 ) ;
  assign n6926 = ( ~n1783 & n6924 ) | ( ~n1783 & n6925 ) | ( n6924 & n6925 ) ;
  assign n6927 = ( ~n1643 & n6923 ) | ( ~n1643 & n6926 ) | ( n6923 & n6926 ) ;
  assign n6928 = ( n1822 & n6923 ) | ( n1822 & n6926 ) | ( n6923 & n6926 ) ;
  assign n6929 = ( n1324 & n6927 ) | ( n1324 & n6928 ) | ( n6927 & n6928 ) ;
  assign n6930 = n6920 | n6929 ;
  assign n6931 = x426 & n991 ;
  assign n6932 = x426 & ~n995 ;
  assign n6933 = ( ~n1104 & n6931 ) | ( ~n1104 & n6932 ) | ( n6931 & n6932 ) ;
  assign n6934 = ( ~n1119 & n6931 ) | ( ~n1119 & n6932 ) | ( n6931 & n6932 ) ;
  assign n6935 = ( n1126 & n6931 ) | ( n1126 & n6932 ) | ( n6931 & n6932 ) ;
  assign n6936 = ( n1115 & n6934 ) | ( n1115 & n6935 ) | ( n6934 & n6935 ) ;
  assign n6937 = ( n975 & n6933 ) | ( n975 & n6936 ) | ( n6933 & n6936 ) ;
  assign n6938 = ( ~n1154 & n6933 ) | ( ~n1154 & n6936 ) | ( n6933 & n6936 ) ;
  assign n6939 = ( x409 & n6937 ) | ( x409 & n6938 ) | ( n6937 & n6938 ) ;
  assign n6940 = ( ~x281 & n6937 ) | ( ~x281 & n6938 ) | ( n6937 & n6938 ) ;
  assign n6941 = ( ~n656 & n6939 ) | ( ~n656 & n6940 ) | ( n6939 & n6940 ) ;
  assign n6942 = x298 & ~n991 ;
  assign n6943 = x298 & n995 ;
  assign n6944 = ( n1104 & n6942 ) | ( n1104 & n6943 ) | ( n6942 & n6943 ) ;
  assign n6945 = ( n1119 & n6942 ) | ( n1119 & n6943 ) | ( n6942 & n6943 ) ;
  assign n6946 = ( ~n1126 & n6942 ) | ( ~n1126 & n6943 ) | ( n6942 & n6943 ) ;
  assign n6947 = ( ~n1115 & n6945 ) | ( ~n1115 & n6946 ) | ( n6945 & n6946 ) ;
  assign n6948 = ( ~n975 & n6944 ) | ( ~n975 & n6947 ) | ( n6944 & n6947 ) ;
  assign n6949 = ( n1154 & n6944 ) | ( n1154 & n6947 ) | ( n6944 & n6947 ) ;
  assign n6950 = ( ~x409 & n6948 ) | ( ~x409 & n6949 ) | ( n6948 & n6949 ) ;
  assign n6951 = ( x281 & n6948 ) | ( x281 & n6949 ) | ( n6948 & n6949 ) ;
  assign n6952 = ( n656 & n6950 ) | ( n656 & n6951 ) | ( n6950 & n6951 ) ;
  assign n6953 = n6941 | n6952 ;
  assign n6954 = ~n6930 & n6953 ;
  assign n6955 = x171 & n1767 ;
  assign n6956 = x171 & ~n1771 ;
  assign n6957 = ( ~n1751 & n6955 ) | ( ~n1751 & n6956 ) | ( n6955 & n6956 ) ;
  assign n6958 = ( ~n1787 & n6955 ) | ( ~n1787 & n6956 ) | ( n6955 & n6956 ) ;
  assign n6959 = ( n1794 & n6955 ) | ( n1794 & n6956 ) | ( n6955 & n6956 ) ;
  assign n6960 = ( n1783 & n6958 ) | ( n1783 & n6959 ) | ( n6958 & n6959 ) ;
  assign n6961 = ( n1643 & n6957 ) | ( n1643 & n6960 ) | ( n6957 & n6960 ) ;
  assign n6962 = ( ~n1822 & n6957 ) | ( ~n1822 & n6960 ) | ( n6957 & n6960 ) ;
  assign n6963 = ( ~n1324 & n6961 ) | ( ~n1324 & n6962 ) | ( n6961 & n6962 ) ;
  assign n6964 = x43 & ~n1767 ;
  assign n6965 = x43 & n1771 ;
  assign n6966 = ( n1751 & n6964 ) | ( n1751 & n6965 ) | ( n6964 & n6965 ) ;
  assign n6967 = ( n1787 & n6964 ) | ( n1787 & n6965 ) | ( n6964 & n6965 ) ;
  assign n6968 = ( ~n1794 & n6964 ) | ( ~n1794 & n6965 ) | ( n6964 & n6965 ) ;
  assign n6969 = ( ~n1783 & n6967 ) | ( ~n1783 & n6968 ) | ( n6967 & n6968 ) ;
  assign n6970 = ( ~n1643 & n6966 ) | ( ~n1643 & n6969 ) | ( n6966 & n6969 ) ;
  assign n6971 = ( n1822 & n6966 ) | ( n1822 & n6969 ) | ( n6966 & n6969 ) ;
  assign n6972 = ( n1324 & n6970 ) | ( n1324 & n6971 ) | ( n6970 & n6971 ) ;
  assign n6973 = n6963 | n6972 ;
  assign n6974 = x427 & n991 ;
  assign n6975 = x427 & ~n995 ;
  assign n6976 = ( ~n1104 & n6974 ) | ( ~n1104 & n6975 ) | ( n6974 & n6975 ) ;
  assign n6977 = ( ~n1119 & n6974 ) | ( ~n1119 & n6975 ) | ( n6974 & n6975 ) ;
  assign n6978 = ( n1126 & n6974 ) | ( n1126 & n6975 ) | ( n6974 & n6975 ) ;
  assign n6979 = ( n1115 & n6977 ) | ( n1115 & n6978 ) | ( n6977 & n6978 ) ;
  assign n6980 = ( n975 & n6976 ) | ( n975 & n6979 ) | ( n6976 & n6979 ) ;
  assign n6981 = ( ~n1154 & n6976 ) | ( ~n1154 & n6979 ) | ( n6976 & n6979 ) ;
  assign n6982 = ( x409 & n6980 ) | ( x409 & n6981 ) | ( n6980 & n6981 ) ;
  assign n6983 = ( ~x281 & n6980 ) | ( ~x281 & n6981 ) | ( n6980 & n6981 ) ;
  assign n6984 = ( ~n656 & n6982 ) | ( ~n656 & n6983 ) | ( n6982 & n6983 ) ;
  assign n6985 = x299 & ~n991 ;
  assign n6986 = x299 & n995 ;
  assign n6987 = ( n1104 & n6985 ) | ( n1104 & n6986 ) | ( n6985 & n6986 ) ;
  assign n6988 = ( n1119 & n6985 ) | ( n1119 & n6986 ) | ( n6985 & n6986 ) ;
  assign n6989 = ( ~n1126 & n6985 ) | ( ~n1126 & n6986 ) | ( n6985 & n6986 ) ;
  assign n6990 = ( ~n1115 & n6988 ) | ( ~n1115 & n6989 ) | ( n6988 & n6989 ) ;
  assign n6991 = ( ~n975 & n6987 ) | ( ~n975 & n6990 ) | ( n6987 & n6990 ) ;
  assign n6992 = ( n1154 & n6987 ) | ( n1154 & n6990 ) | ( n6987 & n6990 ) ;
  assign n6993 = ( ~x409 & n6991 ) | ( ~x409 & n6992 ) | ( n6991 & n6992 ) ;
  assign n6994 = ( x281 & n6991 ) | ( x281 & n6992 ) | ( n6991 & n6992 ) ;
  assign n6995 = ( n656 & n6993 ) | ( n656 & n6994 ) | ( n6993 & n6994 ) ;
  assign n6996 = n6984 | n6995 ;
  assign n6997 = ~n6973 & n6996 ;
  assign n6998 = n6954 | n6997 ;
  assign n6999 = x169 & n1767 ;
  assign n7000 = x169 & ~n1771 ;
  assign n7001 = ( ~n1751 & n6999 ) | ( ~n1751 & n7000 ) | ( n6999 & n7000 ) ;
  assign n7002 = ( ~n1787 & n6999 ) | ( ~n1787 & n7000 ) | ( n6999 & n7000 ) ;
  assign n7003 = ( n1794 & n6999 ) | ( n1794 & n7000 ) | ( n6999 & n7000 ) ;
  assign n7004 = ( n1783 & n7002 ) | ( n1783 & n7003 ) | ( n7002 & n7003 ) ;
  assign n7005 = ( n1643 & n7001 ) | ( n1643 & n7004 ) | ( n7001 & n7004 ) ;
  assign n7006 = ( ~n1822 & n7001 ) | ( ~n1822 & n7004 ) | ( n7001 & n7004 ) ;
  assign n7007 = ( ~n1324 & n7005 ) | ( ~n1324 & n7006 ) | ( n7005 & n7006 ) ;
  assign n7008 = x41 & ~n1767 ;
  assign n7009 = x41 & n1771 ;
  assign n7010 = ( n1751 & n7008 ) | ( n1751 & n7009 ) | ( n7008 & n7009 ) ;
  assign n7011 = ( n1787 & n7008 ) | ( n1787 & n7009 ) | ( n7008 & n7009 ) ;
  assign n7012 = ( ~n1794 & n7008 ) | ( ~n1794 & n7009 ) | ( n7008 & n7009 ) ;
  assign n7013 = ( ~n1783 & n7011 ) | ( ~n1783 & n7012 ) | ( n7011 & n7012 ) ;
  assign n7014 = ( ~n1643 & n7010 ) | ( ~n1643 & n7013 ) | ( n7010 & n7013 ) ;
  assign n7015 = ( n1822 & n7010 ) | ( n1822 & n7013 ) | ( n7010 & n7013 ) ;
  assign n7016 = ( n1324 & n7014 ) | ( n1324 & n7015 ) | ( n7014 & n7015 ) ;
  assign n7017 = n7007 | n7016 ;
  assign n7018 = x425 & n991 ;
  assign n7019 = x425 & ~n995 ;
  assign n7020 = ( ~n1104 & n7018 ) | ( ~n1104 & n7019 ) | ( n7018 & n7019 ) ;
  assign n7021 = ( ~n1119 & n7018 ) | ( ~n1119 & n7019 ) | ( n7018 & n7019 ) ;
  assign n7022 = ( n1126 & n7018 ) | ( n1126 & n7019 ) | ( n7018 & n7019 ) ;
  assign n7023 = ( n1115 & n7021 ) | ( n1115 & n7022 ) | ( n7021 & n7022 ) ;
  assign n7024 = ( n975 & n7020 ) | ( n975 & n7023 ) | ( n7020 & n7023 ) ;
  assign n7025 = ( ~n1154 & n7020 ) | ( ~n1154 & n7023 ) | ( n7020 & n7023 ) ;
  assign n7026 = ( x409 & n7024 ) | ( x409 & n7025 ) | ( n7024 & n7025 ) ;
  assign n7027 = ( ~x281 & n7024 ) | ( ~x281 & n7025 ) | ( n7024 & n7025 ) ;
  assign n7028 = ( ~n656 & n7026 ) | ( ~n656 & n7027 ) | ( n7026 & n7027 ) ;
  assign n7029 = x297 & ~n991 ;
  assign n7030 = x297 & n995 ;
  assign n7031 = ( n1104 & n7029 ) | ( n1104 & n7030 ) | ( n7029 & n7030 ) ;
  assign n7032 = ( n1119 & n7029 ) | ( n1119 & n7030 ) | ( n7029 & n7030 ) ;
  assign n7033 = ( ~n1126 & n7029 ) | ( ~n1126 & n7030 ) | ( n7029 & n7030 ) ;
  assign n7034 = ( ~n1115 & n7032 ) | ( ~n1115 & n7033 ) | ( n7032 & n7033 ) ;
  assign n7035 = ( ~n975 & n7031 ) | ( ~n975 & n7034 ) | ( n7031 & n7034 ) ;
  assign n7036 = ( n1154 & n7031 ) | ( n1154 & n7034 ) | ( n7031 & n7034 ) ;
  assign n7037 = ( ~x409 & n7035 ) | ( ~x409 & n7036 ) | ( n7035 & n7036 ) ;
  assign n7038 = ( x281 & n7035 ) | ( x281 & n7036 ) | ( n7035 & n7036 ) ;
  assign n7039 = ( n656 & n7037 ) | ( n656 & n7038 ) | ( n7037 & n7038 ) ;
  assign n7040 = n7028 | n7039 ;
  assign n7041 = ~n7017 & n7040 ;
  assign n7042 = x168 & n1767 ;
  assign n7043 = x168 & ~n1771 ;
  assign n7044 = ( ~n1751 & n7042 ) | ( ~n1751 & n7043 ) | ( n7042 & n7043 ) ;
  assign n7045 = ( ~n1787 & n7042 ) | ( ~n1787 & n7043 ) | ( n7042 & n7043 ) ;
  assign n7046 = ( n1794 & n7042 ) | ( n1794 & n7043 ) | ( n7042 & n7043 ) ;
  assign n7047 = ( n1783 & n7045 ) | ( n1783 & n7046 ) | ( n7045 & n7046 ) ;
  assign n7048 = ( n1643 & n7044 ) | ( n1643 & n7047 ) | ( n7044 & n7047 ) ;
  assign n7049 = ( ~n1822 & n7044 ) | ( ~n1822 & n7047 ) | ( n7044 & n7047 ) ;
  assign n7050 = ( ~n1324 & n7048 ) | ( ~n1324 & n7049 ) | ( n7048 & n7049 ) ;
  assign n7051 = x40 & ~n1767 ;
  assign n7052 = x40 & n1771 ;
  assign n7053 = ( n1751 & n7051 ) | ( n1751 & n7052 ) | ( n7051 & n7052 ) ;
  assign n7054 = ( n1787 & n7051 ) | ( n1787 & n7052 ) | ( n7051 & n7052 ) ;
  assign n7055 = ( ~n1794 & n7051 ) | ( ~n1794 & n7052 ) | ( n7051 & n7052 ) ;
  assign n7056 = ( ~n1783 & n7054 ) | ( ~n1783 & n7055 ) | ( n7054 & n7055 ) ;
  assign n7057 = ( ~n1643 & n7053 ) | ( ~n1643 & n7056 ) | ( n7053 & n7056 ) ;
  assign n7058 = ( n1822 & n7053 ) | ( n1822 & n7056 ) | ( n7053 & n7056 ) ;
  assign n7059 = ( n1324 & n7057 ) | ( n1324 & n7058 ) | ( n7057 & n7058 ) ;
  assign n7060 = n7050 | n7059 ;
  assign n7061 = x424 & n991 ;
  assign n7062 = x424 & ~n995 ;
  assign n7063 = ( ~n1104 & n7061 ) | ( ~n1104 & n7062 ) | ( n7061 & n7062 ) ;
  assign n7064 = ( ~n1119 & n7061 ) | ( ~n1119 & n7062 ) | ( n7061 & n7062 ) ;
  assign n7065 = ( n1126 & n7061 ) | ( n1126 & n7062 ) | ( n7061 & n7062 ) ;
  assign n7066 = ( n1115 & n7064 ) | ( n1115 & n7065 ) | ( n7064 & n7065 ) ;
  assign n7067 = ( n975 & n7063 ) | ( n975 & n7066 ) | ( n7063 & n7066 ) ;
  assign n7068 = ( ~n1154 & n7063 ) | ( ~n1154 & n7066 ) | ( n7063 & n7066 ) ;
  assign n7069 = ( x409 & n7067 ) | ( x409 & n7068 ) | ( n7067 & n7068 ) ;
  assign n7070 = ( ~x281 & n7067 ) | ( ~x281 & n7068 ) | ( n7067 & n7068 ) ;
  assign n7071 = ( ~n656 & n7069 ) | ( ~n656 & n7070 ) | ( n7069 & n7070 ) ;
  assign n7072 = x296 & ~n991 ;
  assign n7073 = x296 & n995 ;
  assign n7074 = ( n1104 & n7072 ) | ( n1104 & n7073 ) | ( n7072 & n7073 ) ;
  assign n7075 = ( n1119 & n7072 ) | ( n1119 & n7073 ) | ( n7072 & n7073 ) ;
  assign n7076 = ( ~n1126 & n7072 ) | ( ~n1126 & n7073 ) | ( n7072 & n7073 ) ;
  assign n7077 = ( ~n1115 & n7075 ) | ( ~n1115 & n7076 ) | ( n7075 & n7076 ) ;
  assign n7078 = ( ~n975 & n7074 ) | ( ~n975 & n7077 ) | ( n7074 & n7077 ) ;
  assign n7079 = ( n1154 & n7074 ) | ( n1154 & n7077 ) | ( n7074 & n7077 ) ;
  assign n7080 = ( ~x409 & n7078 ) | ( ~x409 & n7079 ) | ( n7078 & n7079 ) ;
  assign n7081 = ( x281 & n7078 ) | ( x281 & n7079 ) | ( n7078 & n7079 ) ;
  assign n7082 = ( n656 & n7080 ) | ( n656 & n7081 ) | ( n7080 & n7081 ) ;
  assign n7083 = n7071 | n7082 ;
  assign n7084 = ~n7060 & n7083 ;
  assign n7085 = n7041 | n7084 ;
  assign n7086 = n6998 | n7085 ;
  assign n7087 = n6911 | n7086 ;
  assign n7088 = x416 & n991 ;
  assign n7089 = x416 & ~n995 ;
  assign n7090 = ( ~n1104 & n7088 ) | ( ~n1104 & n7089 ) | ( n7088 & n7089 ) ;
  assign n7091 = ( ~n1119 & n7088 ) | ( ~n1119 & n7089 ) | ( n7088 & n7089 ) ;
  assign n7092 = ( n1126 & n7088 ) | ( n1126 & n7089 ) | ( n7088 & n7089 ) ;
  assign n7093 = ( n1115 & n7091 ) | ( n1115 & n7092 ) | ( n7091 & n7092 ) ;
  assign n7094 = ( n975 & n7090 ) | ( n975 & n7093 ) | ( n7090 & n7093 ) ;
  assign n7095 = ( ~n1154 & n7090 ) | ( ~n1154 & n7093 ) | ( n7090 & n7093 ) ;
  assign n7096 = ( x409 & n7094 ) | ( x409 & n7095 ) | ( n7094 & n7095 ) ;
  assign n7097 = ( ~x281 & n7094 ) | ( ~x281 & n7095 ) | ( n7094 & n7095 ) ;
  assign n7098 = ( ~n656 & n7096 ) | ( ~n656 & n7097 ) | ( n7096 & n7097 ) ;
  assign n7099 = x288 & ~n991 ;
  assign n7100 = x288 & n995 ;
  assign n7101 = ( n1104 & n7099 ) | ( n1104 & n7100 ) | ( n7099 & n7100 ) ;
  assign n7102 = ( n1119 & n7099 ) | ( n1119 & n7100 ) | ( n7099 & n7100 ) ;
  assign n7103 = ( ~n1126 & n7099 ) | ( ~n1126 & n7100 ) | ( n7099 & n7100 ) ;
  assign n7104 = ( ~n1115 & n7102 ) | ( ~n1115 & n7103 ) | ( n7102 & n7103 ) ;
  assign n7105 = ( ~n975 & n7101 ) | ( ~n975 & n7104 ) | ( n7101 & n7104 ) ;
  assign n7106 = ( n1154 & n7101 ) | ( n1154 & n7104 ) | ( n7101 & n7104 ) ;
  assign n7107 = ( ~x409 & n7105 ) | ( ~x409 & n7106 ) | ( n7105 & n7106 ) ;
  assign n7108 = ( x281 & n7105 ) | ( x281 & n7106 ) | ( n7105 & n7106 ) ;
  assign n7109 = ( n656 & n7107 ) | ( n656 & n7108 ) | ( n7107 & n7108 ) ;
  assign n7110 = n7098 | n7109 ;
  assign n7111 = x160 & n1767 ;
  assign n7112 = x160 & ~n1771 ;
  assign n7113 = ( ~n1751 & n7111 ) | ( ~n1751 & n7112 ) | ( n7111 & n7112 ) ;
  assign n7114 = ( ~n1787 & n7111 ) | ( ~n1787 & n7112 ) | ( n7111 & n7112 ) ;
  assign n7115 = ( n1794 & n7111 ) | ( n1794 & n7112 ) | ( n7111 & n7112 ) ;
  assign n7116 = ( n1783 & n7114 ) | ( n1783 & n7115 ) | ( n7114 & n7115 ) ;
  assign n7117 = ( n1643 & n7113 ) | ( n1643 & n7116 ) | ( n7113 & n7116 ) ;
  assign n7118 = ( ~n1822 & n7113 ) | ( ~n1822 & n7116 ) | ( n7113 & n7116 ) ;
  assign n7119 = ( ~n1324 & n7117 ) | ( ~n1324 & n7118 ) | ( n7117 & n7118 ) ;
  assign n7120 = x32 & ~n1767 ;
  assign n7121 = x32 & n1771 ;
  assign n7122 = ( n1751 & n7120 ) | ( n1751 & n7121 ) | ( n7120 & n7121 ) ;
  assign n7123 = ( n1787 & n7120 ) | ( n1787 & n7121 ) | ( n7120 & n7121 ) ;
  assign n7124 = ( ~n1794 & n7120 ) | ( ~n1794 & n7121 ) | ( n7120 & n7121 ) ;
  assign n7125 = ( ~n1783 & n7123 ) | ( ~n1783 & n7124 ) | ( n7123 & n7124 ) ;
  assign n7126 = ( ~n1643 & n7122 ) | ( ~n1643 & n7125 ) | ( n7122 & n7125 ) ;
  assign n7127 = ( n1822 & n7122 ) | ( n1822 & n7125 ) | ( n7122 & n7125 ) ;
  assign n7128 = ( n1324 & n7126 ) | ( n1324 & n7127 ) | ( n7126 & n7127 ) ;
  assign n7129 = n7119 | n7128 ;
  assign n7130 = n7110 & ~n7129 ;
  assign n7131 = x167 & n1767 ;
  assign n7132 = x167 & ~n1771 ;
  assign n7133 = ( ~n1751 & n7131 ) | ( ~n1751 & n7132 ) | ( n7131 & n7132 ) ;
  assign n7134 = ( ~n1787 & n7131 ) | ( ~n1787 & n7132 ) | ( n7131 & n7132 ) ;
  assign n7135 = ( n1794 & n7131 ) | ( n1794 & n7132 ) | ( n7131 & n7132 ) ;
  assign n7136 = ( n1783 & n7134 ) | ( n1783 & n7135 ) | ( n7134 & n7135 ) ;
  assign n7137 = ( n1643 & n7133 ) | ( n1643 & n7136 ) | ( n7133 & n7136 ) ;
  assign n7138 = ( ~n1822 & n7133 ) | ( ~n1822 & n7136 ) | ( n7133 & n7136 ) ;
  assign n7139 = ( ~n1324 & n7137 ) | ( ~n1324 & n7138 ) | ( n7137 & n7138 ) ;
  assign n7140 = x39 & ~n1767 ;
  assign n7141 = x39 & n1771 ;
  assign n7142 = ( n1751 & n7140 ) | ( n1751 & n7141 ) | ( n7140 & n7141 ) ;
  assign n7143 = ( n1787 & n7140 ) | ( n1787 & n7141 ) | ( n7140 & n7141 ) ;
  assign n7144 = ( ~n1794 & n7140 ) | ( ~n1794 & n7141 ) | ( n7140 & n7141 ) ;
  assign n7145 = ( ~n1783 & n7143 ) | ( ~n1783 & n7144 ) | ( n7143 & n7144 ) ;
  assign n7146 = ( ~n1643 & n7142 ) | ( ~n1643 & n7145 ) | ( n7142 & n7145 ) ;
  assign n7147 = ( n1822 & n7142 ) | ( n1822 & n7145 ) | ( n7142 & n7145 ) ;
  assign n7148 = ( n1324 & n7146 ) | ( n1324 & n7147 ) | ( n7146 & n7147 ) ;
  assign n7149 = n7139 | n7148 ;
  assign n7150 = x423 & n991 ;
  assign n7151 = x423 & ~n995 ;
  assign n7152 = ( ~n1104 & n7150 ) | ( ~n1104 & n7151 ) | ( n7150 & n7151 ) ;
  assign n7153 = ( ~n1119 & n7150 ) | ( ~n1119 & n7151 ) | ( n7150 & n7151 ) ;
  assign n7154 = ( n1126 & n7150 ) | ( n1126 & n7151 ) | ( n7150 & n7151 ) ;
  assign n7155 = ( n1115 & n7153 ) | ( n1115 & n7154 ) | ( n7153 & n7154 ) ;
  assign n7156 = ( n975 & n7152 ) | ( n975 & n7155 ) | ( n7152 & n7155 ) ;
  assign n7157 = ( ~n1154 & n7152 ) | ( ~n1154 & n7155 ) | ( n7152 & n7155 ) ;
  assign n7158 = ( x409 & n7156 ) | ( x409 & n7157 ) | ( n7156 & n7157 ) ;
  assign n7159 = ( ~x281 & n7156 ) | ( ~x281 & n7157 ) | ( n7156 & n7157 ) ;
  assign n7160 = ( ~n656 & n7158 ) | ( ~n656 & n7159 ) | ( n7158 & n7159 ) ;
  assign n7161 = x295 & ~n991 ;
  assign n7162 = x295 & n995 ;
  assign n7163 = ( n1104 & n7161 ) | ( n1104 & n7162 ) | ( n7161 & n7162 ) ;
  assign n7164 = ( n1119 & n7161 ) | ( n1119 & n7162 ) | ( n7161 & n7162 ) ;
  assign n7165 = ( ~n1126 & n7161 ) | ( ~n1126 & n7162 ) | ( n7161 & n7162 ) ;
  assign n7166 = ( ~n1115 & n7164 ) | ( ~n1115 & n7165 ) | ( n7164 & n7165 ) ;
  assign n7167 = ( ~n975 & n7163 ) | ( ~n975 & n7166 ) | ( n7163 & n7166 ) ;
  assign n7168 = ( n1154 & n7163 ) | ( n1154 & n7166 ) | ( n7163 & n7166 ) ;
  assign n7169 = ( ~x409 & n7167 ) | ( ~x409 & n7168 ) | ( n7167 & n7168 ) ;
  assign n7170 = ( x281 & n7167 ) | ( x281 & n7168 ) | ( n7167 & n7168 ) ;
  assign n7171 = ( n656 & n7169 ) | ( n656 & n7170 ) | ( n7169 & n7170 ) ;
  assign n7172 = n7160 | n7171 ;
  assign n7173 = ~n7149 & n7172 ;
  assign n7174 = x422 & n991 ;
  assign n7175 = x422 & ~n995 ;
  assign n7176 = ( ~n1104 & n7174 ) | ( ~n1104 & n7175 ) | ( n7174 & n7175 ) ;
  assign n7177 = ( ~n1119 & n7174 ) | ( ~n1119 & n7175 ) | ( n7174 & n7175 ) ;
  assign n7178 = ( n1126 & n7174 ) | ( n1126 & n7175 ) | ( n7174 & n7175 ) ;
  assign n7179 = ( n1115 & n7177 ) | ( n1115 & n7178 ) | ( n7177 & n7178 ) ;
  assign n7180 = ( n975 & n7176 ) | ( n975 & n7179 ) | ( n7176 & n7179 ) ;
  assign n7181 = ( ~n1154 & n7176 ) | ( ~n1154 & n7179 ) | ( n7176 & n7179 ) ;
  assign n7182 = ( x409 & n7180 ) | ( x409 & n7181 ) | ( n7180 & n7181 ) ;
  assign n7183 = ( ~x281 & n7180 ) | ( ~x281 & n7181 ) | ( n7180 & n7181 ) ;
  assign n7184 = ( ~n656 & n7182 ) | ( ~n656 & n7183 ) | ( n7182 & n7183 ) ;
  assign n7185 = x294 & ~n991 ;
  assign n7186 = x294 & n995 ;
  assign n7187 = ( n1104 & n7185 ) | ( n1104 & n7186 ) | ( n7185 & n7186 ) ;
  assign n7188 = ( n1119 & n7185 ) | ( n1119 & n7186 ) | ( n7185 & n7186 ) ;
  assign n7189 = ( ~n1126 & n7185 ) | ( ~n1126 & n7186 ) | ( n7185 & n7186 ) ;
  assign n7190 = ( ~n1115 & n7188 ) | ( ~n1115 & n7189 ) | ( n7188 & n7189 ) ;
  assign n7191 = ( ~n975 & n7187 ) | ( ~n975 & n7190 ) | ( n7187 & n7190 ) ;
  assign n7192 = ( n1154 & n7187 ) | ( n1154 & n7190 ) | ( n7187 & n7190 ) ;
  assign n7193 = ( ~x409 & n7191 ) | ( ~x409 & n7192 ) | ( n7191 & n7192 ) ;
  assign n7194 = ( x281 & n7191 ) | ( x281 & n7192 ) | ( n7191 & n7192 ) ;
  assign n7195 = ( n656 & n7193 ) | ( n656 & n7194 ) | ( n7193 & n7194 ) ;
  assign n7196 = n7184 | n7195 ;
  assign n7197 = x166 & n1767 ;
  assign n7198 = x166 & ~n1771 ;
  assign n7199 = ( ~n1751 & n7197 ) | ( ~n1751 & n7198 ) | ( n7197 & n7198 ) ;
  assign n7200 = ( ~n1787 & n7197 ) | ( ~n1787 & n7198 ) | ( n7197 & n7198 ) ;
  assign n7201 = ( n1794 & n7197 ) | ( n1794 & n7198 ) | ( n7197 & n7198 ) ;
  assign n7202 = ( n1783 & n7200 ) | ( n1783 & n7201 ) | ( n7200 & n7201 ) ;
  assign n7203 = ( n1643 & n7199 ) | ( n1643 & n7202 ) | ( n7199 & n7202 ) ;
  assign n7204 = ( ~n1822 & n7199 ) | ( ~n1822 & n7202 ) | ( n7199 & n7202 ) ;
  assign n7205 = ( ~n1324 & n7203 ) | ( ~n1324 & n7204 ) | ( n7203 & n7204 ) ;
  assign n7206 = x38 & ~n1767 ;
  assign n7207 = x38 & n1771 ;
  assign n7208 = ( n1751 & n7206 ) | ( n1751 & n7207 ) | ( n7206 & n7207 ) ;
  assign n7209 = ( n1787 & n7206 ) | ( n1787 & n7207 ) | ( n7206 & n7207 ) ;
  assign n7210 = ( ~n1794 & n7206 ) | ( ~n1794 & n7207 ) | ( n7206 & n7207 ) ;
  assign n7211 = ( ~n1783 & n7209 ) | ( ~n1783 & n7210 ) | ( n7209 & n7210 ) ;
  assign n7212 = ( ~n1643 & n7208 ) | ( ~n1643 & n7211 ) | ( n7208 & n7211 ) ;
  assign n7213 = ( n1822 & n7208 ) | ( n1822 & n7211 ) | ( n7208 & n7211 ) ;
  assign n7214 = ( n1324 & n7212 ) | ( n1324 & n7213 ) | ( n7212 & n7213 ) ;
  assign n7215 = n7205 | n7214 ;
  assign n7216 = n7196 & ~n7215 ;
  assign n7217 = n7173 | n7216 ;
  assign n7218 = x164 & n1767 ;
  assign n7219 = x164 & ~n1771 ;
  assign n7220 = ( ~n1751 & n7218 ) | ( ~n1751 & n7219 ) | ( n7218 & n7219 ) ;
  assign n7221 = ( ~n1787 & n7218 ) | ( ~n1787 & n7219 ) | ( n7218 & n7219 ) ;
  assign n7222 = ( n1794 & n7218 ) | ( n1794 & n7219 ) | ( n7218 & n7219 ) ;
  assign n7223 = ( n1783 & n7221 ) | ( n1783 & n7222 ) | ( n7221 & n7222 ) ;
  assign n7224 = ( n1643 & n7220 ) | ( n1643 & n7223 ) | ( n7220 & n7223 ) ;
  assign n7225 = ( ~n1822 & n7220 ) | ( ~n1822 & n7223 ) | ( n7220 & n7223 ) ;
  assign n7226 = ( ~n1324 & n7224 ) | ( ~n1324 & n7225 ) | ( n7224 & n7225 ) ;
  assign n7227 = x36 & ~n1767 ;
  assign n7228 = x36 & n1771 ;
  assign n7229 = ( n1751 & n7227 ) | ( n1751 & n7228 ) | ( n7227 & n7228 ) ;
  assign n7230 = ( n1787 & n7227 ) | ( n1787 & n7228 ) | ( n7227 & n7228 ) ;
  assign n7231 = ( ~n1794 & n7227 ) | ( ~n1794 & n7228 ) | ( n7227 & n7228 ) ;
  assign n7232 = ( ~n1783 & n7230 ) | ( ~n1783 & n7231 ) | ( n7230 & n7231 ) ;
  assign n7233 = ( ~n1643 & n7229 ) | ( ~n1643 & n7232 ) | ( n7229 & n7232 ) ;
  assign n7234 = ( n1822 & n7229 ) | ( n1822 & n7232 ) | ( n7229 & n7232 ) ;
  assign n7235 = ( n1324 & n7233 ) | ( n1324 & n7234 ) | ( n7233 & n7234 ) ;
  assign n7236 = n7226 | n7235 ;
  assign n7237 = x420 & n991 ;
  assign n7238 = x420 & ~n995 ;
  assign n7239 = ( ~n1104 & n7237 ) | ( ~n1104 & n7238 ) | ( n7237 & n7238 ) ;
  assign n7240 = ( ~n1119 & n7237 ) | ( ~n1119 & n7238 ) | ( n7237 & n7238 ) ;
  assign n7241 = ( n1126 & n7237 ) | ( n1126 & n7238 ) | ( n7237 & n7238 ) ;
  assign n7242 = ( n1115 & n7240 ) | ( n1115 & n7241 ) | ( n7240 & n7241 ) ;
  assign n7243 = ( n975 & n7239 ) | ( n975 & n7242 ) | ( n7239 & n7242 ) ;
  assign n7244 = ( ~n1154 & n7239 ) | ( ~n1154 & n7242 ) | ( n7239 & n7242 ) ;
  assign n7245 = ( x409 & n7243 ) | ( x409 & n7244 ) | ( n7243 & n7244 ) ;
  assign n7246 = ( ~x281 & n7243 ) | ( ~x281 & n7244 ) | ( n7243 & n7244 ) ;
  assign n7247 = ( ~n656 & n7245 ) | ( ~n656 & n7246 ) | ( n7245 & n7246 ) ;
  assign n7248 = x292 & ~n991 ;
  assign n7249 = x292 & n995 ;
  assign n7250 = ( n1104 & n7248 ) | ( n1104 & n7249 ) | ( n7248 & n7249 ) ;
  assign n7251 = ( n1119 & n7248 ) | ( n1119 & n7249 ) | ( n7248 & n7249 ) ;
  assign n7252 = ( ~n1126 & n7248 ) | ( ~n1126 & n7249 ) | ( n7248 & n7249 ) ;
  assign n7253 = ( ~n1115 & n7251 ) | ( ~n1115 & n7252 ) | ( n7251 & n7252 ) ;
  assign n7254 = ( ~n975 & n7250 ) | ( ~n975 & n7253 ) | ( n7250 & n7253 ) ;
  assign n7255 = ( n1154 & n7250 ) | ( n1154 & n7253 ) | ( n7250 & n7253 ) ;
  assign n7256 = ( ~x409 & n7254 ) | ( ~x409 & n7255 ) | ( n7254 & n7255 ) ;
  assign n7257 = ( x281 & n7254 ) | ( x281 & n7255 ) | ( n7254 & n7255 ) ;
  assign n7258 = ( n656 & n7256 ) | ( n656 & n7257 ) | ( n7256 & n7257 ) ;
  assign n7259 = n7247 | n7258 ;
  assign n7260 = ~n7236 & n7259 ;
  assign n7261 = x165 & n1767 ;
  assign n7262 = x165 & ~n1771 ;
  assign n7263 = ( ~n1751 & n7261 ) | ( ~n1751 & n7262 ) | ( n7261 & n7262 ) ;
  assign n7264 = ( ~n1787 & n7261 ) | ( ~n1787 & n7262 ) | ( n7261 & n7262 ) ;
  assign n7265 = ( n1794 & n7261 ) | ( n1794 & n7262 ) | ( n7261 & n7262 ) ;
  assign n7266 = ( n1783 & n7264 ) | ( n1783 & n7265 ) | ( n7264 & n7265 ) ;
  assign n7267 = ( n1643 & n7263 ) | ( n1643 & n7266 ) | ( n7263 & n7266 ) ;
  assign n7268 = ( ~n1822 & n7263 ) | ( ~n1822 & n7266 ) | ( n7263 & n7266 ) ;
  assign n7269 = ( ~n1324 & n7267 ) | ( ~n1324 & n7268 ) | ( n7267 & n7268 ) ;
  assign n7270 = x37 & ~n1767 ;
  assign n7271 = x37 & n1771 ;
  assign n7272 = ( n1751 & n7270 ) | ( n1751 & n7271 ) | ( n7270 & n7271 ) ;
  assign n7273 = ( n1787 & n7270 ) | ( n1787 & n7271 ) | ( n7270 & n7271 ) ;
  assign n7274 = ( ~n1794 & n7270 ) | ( ~n1794 & n7271 ) | ( n7270 & n7271 ) ;
  assign n7275 = ( ~n1783 & n7273 ) | ( ~n1783 & n7274 ) | ( n7273 & n7274 ) ;
  assign n7276 = ( ~n1643 & n7272 ) | ( ~n1643 & n7275 ) | ( n7272 & n7275 ) ;
  assign n7277 = ( n1822 & n7272 ) | ( n1822 & n7275 ) | ( n7272 & n7275 ) ;
  assign n7278 = ( n1324 & n7276 ) | ( n1324 & n7277 ) | ( n7276 & n7277 ) ;
  assign n7279 = n7269 | n7278 ;
  assign n7280 = x421 & n991 ;
  assign n7281 = x421 & ~n995 ;
  assign n7282 = ( ~n1104 & n7280 ) | ( ~n1104 & n7281 ) | ( n7280 & n7281 ) ;
  assign n7283 = ( ~n1119 & n7280 ) | ( ~n1119 & n7281 ) | ( n7280 & n7281 ) ;
  assign n7284 = ( n1126 & n7280 ) | ( n1126 & n7281 ) | ( n7280 & n7281 ) ;
  assign n7285 = ( n1115 & n7283 ) | ( n1115 & n7284 ) | ( n7283 & n7284 ) ;
  assign n7286 = ( n975 & n7282 ) | ( n975 & n7285 ) | ( n7282 & n7285 ) ;
  assign n7287 = ( ~n1154 & n7282 ) | ( ~n1154 & n7285 ) | ( n7282 & n7285 ) ;
  assign n7288 = ( x409 & n7286 ) | ( x409 & n7287 ) | ( n7286 & n7287 ) ;
  assign n7289 = ( ~x281 & n7286 ) | ( ~x281 & n7287 ) | ( n7286 & n7287 ) ;
  assign n7290 = ( ~n656 & n7288 ) | ( ~n656 & n7289 ) | ( n7288 & n7289 ) ;
  assign n7291 = x293 & ~n991 ;
  assign n7292 = x293 & n995 ;
  assign n7293 = ( n1104 & n7291 ) | ( n1104 & n7292 ) | ( n7291 & n7292 ) ;
  assign n7294 = ( n1119 & n7291 ) | ( n1119 & n7292 ) | ( n7291 & n7292 ) ;
  assign n7295 = ( ~n1126 & n7291 ) | ( ~n1126 & n7292 ) | ( n7291 & n7292 ) ;
  assign n7296 = ( ~n1115 & n7294 ) | ( ~n1115 & n7295 ) | ( n7294 & n7295 ) ;
  assign n7297 = ( ~n975 & n7293 ) | ( ~n975 & n7296 ) | ( n7293 & n7296 ) ;
  assign n7298 = ( n1154 & n7293 ) | ( n1154 & n7296 ) | ( n7293 & n7296 ) ;
  assign n7299 = ( ~x409 & n7297 ) | ( ~x409 & n7298 ) | ( n7297 & n7298 ) ;
  assign n7300 = ( x281 & n7297 ) | ( x281 & n7298 ) | ( n7297 & n7298 ) ;
  assign n7301 = ( n656 & n7299 ) | ( n656 & n7300 ) | ( n7299 & n7300 ) ;
  assign n7302 = n7290 | n7301 ;
  assign n7303 = ~n7279 & n7302 ;
  assign n7304 = n7260 | n7303 ;
  assign n7305 = n7217 | n7304 ;
  assign n7306 = x161 & n1767 ;
  assign n7307 = x161 & ~n1771 ;
  assign n7308 = ( ~n1751 & n7306 ) | ( ~n1751 & n7307 ) | ( n7306 & n7307 ) ;
  assign n7309 = ( ~n1787 & n7306 ) | ( ~n1787 & n7307 ) | ( n7306 & n7307 ) ;
  assign n7310 = ( n1794 & n7306 ) | ( n1794 & n7307 ) | ( n7306 & n7307 ) ;
  assign n7311 = ( n1783 & n7309 ) | ( n1783 & n7310 ) | ( n7309 & n7310 ) ;
  assign n7312 = ( n1643 & n7308 ) | ( n1643 & n7311 ) | ( n7308 & n7311 ) ;
  assign n7313 = ( ~n1822 & n7308 ) | ( ~n1822 & n7311 ) | ( n7308 & n7311 ) ;
  assign n7314 = ( ~n1324 & n7312 ) | ( ~n1324 & n7313 ) | ( n7312 & n7313 ) ;
  assign n7315 = x33 & ~n1767 ;
  assign n7316 = x33 & n1771 ;
  assign n7317 = ( n1751 & n7315 ) | ( n1751 & n7316 ) | ( n7315 & n7316 ) ;
  assign n7318 = ( n1787 & n7315 ) | ( n1787 & n7316 ) | ( n7315 & n7316 ) ;
  assign n7319 = ( ~n1794 & n7315 ) | ( ~n1794 & n7316 ) | ( n7315 & n7316 ) ;
  assign n7320 = ( ~n1783 & n7318 ) | ( ~n1783 & n7319 ) | ( n7318 & n7319 ) ;
  assign n7321 = ( ~n1643 & n7317 ) | ( ~n1643 & n7320 ) | ( n7317 & n7320 ) ;
  assign n7322 = ( n1822 & n7317 ) | ( n1822 & n7320 ) | ( n7317 & n7320 ) ;
  assign n7323 = ( n1324 & n7321 ) | ( n1324 & n7322 ) | ( n7321 & n7322 ) ;
  assign n7324 = n7314 | n7323 ;
  assign n7325 = x417 & n991 ;
  assign n7326 = x417 & ~n995 ;
  assign n7327 = ( ~n1104 & n7325 ) | ( ~n1104 & n7326 ) | ( n7325 & n7326 ) ;
  assign n7328 = ( ~n1119 & n7325 ) | ( ~n1119 & n7326 ) | ( n7325 & n7326 ) ;
  assign n7329 = ( n1126 & n7325 ) | ( n1126 & n7326 ) | ( n7325 & n7326 ) ;
  assign n7330 = ( n1115 & n7328 ) | ( n1115 & n7329 ) | ( n7328 & n7329 ) ;
  assign n7331 = ( n975 & n7327 ) | ( n975 & n7330 ) | ( n7327 & n7330 ) ;
  assign n7332 = ( ~n1154 & n7327 ) | ( ~n1154 & n7330 ) | ( n7327 & n7330 ) ;
  assign n7333 = ( x409 & n7331 ) | ( x409 & n7332 ) | ( n7331 & n7332 ) ;
  assign n7334 = ( ~x281 & n7331 ) | ( ~x281 & n7332 ) | ( n7331 & n7332 ) ;
  assign n7335 = ( ~n656 & n7333 ) | ( ~n656 & n7334 ) | ( n7333 & n7334 ) ;
  assign n7336 = x289 & ~n991 ;
  assign n7337 = x289 & n995 ;
  assign n7338 = ( n1104 & n7336 ) | ( n1104 & n7337 ) | ( n7336 & n7337 ) ;
  assign n7339 = ( n1119 & n7336 ) | ( n1119 & n7337 ) | ( n7336 & n7337 ) ;
  assign n7340 = ( ~n1126 & n7336 ) | ( ~n1126 & n7337 ) | ( n7336 & n7337 ) ;
  assign n7341 = ( ~n1115 & n7339 ) | ( ~n1115 & n7340 ) | ( n7339 & n7340 ) ;
  assign n7342 = ( ~n975 & n7338 ) | ( ~n975 & n7341 ) | ( n7338 & n7341 ) ;
  assign n7343 = ( n1154 & n7338 ) | ( n1154 & n7341 ) | ( n7338 & n7341 ) ;
  assign n7344 = ( ~x409 & n7342 ) | ( ~x409 & n7343 ) | ( n7342 & n7343 ) ;
  assign n7345 = ( x281 & n7342 ) | ( x281 & n7343 ) | ( n7342 & n7343 ) ;
  assign n7346 = ( n656 & n7344 ) | ( n656 & n7345 ) | ( n7344 & n7345 ) ;
  assign n7347 = n7335 | n7346 ;
  assign n7348 = ~n7324 & n7347 ;
  assign n7349 = x163 & n1767 ;
  assign n7350 = x163 & ~n1771 ;
  assign n7351 = ( ~n1751 & n7349 ) | ( ~n1751 & n7350 ) | ( n7349 & n7350 ) ;
  assign n7352 = ( ~n1787 & n7349 ) | ( ~n1787 & n7350 ) | ( n7349 & n7350 ) ;
  assign n7353 = ( n1794 & n7349 ) | ( n1794 & n7350 ) | ( n7349 & n7350 ) ;
  assign n7354 = ( n1783 & n7352 ) | ( n1783 & n7353 ) | ( n7352 & n7353 ) ;
  assign n7355 = ( n1643 & n7351 ) | ( n1643 & n7354 ) | ( n7351 & n7354 ) ;
  assign n7356 = ( ~n1822 & n7351 ) | ( ~n1822 & n7354 ) | ( n7351 & n7354 ) ;
  assign n7357 = ( ~n1324 & n7355 ) | ( ~n1324 & n7356 ) | ( n7355 & n7356 ) ;
  assign n7358 = x35 & ~n1767 ;
  assign n7359 = x35 & n1771 ;
  assign n7360 = ( n1751 & n7358 ) | ( n1751 & n7359 ) | ( n7358 & n7359 ) ;
  assign n7361 = ( n1787 & n7358 ) | ( n1787 & n7359 ) | ( n7358 & n7359 ) ;
  assign n7362 = ( ~n1794 & n7358 ) | ( ~n1794 & n7359 ) | ( n7358 & n7359 ) ;
  assign n7363 = ( ~n1783 & n7361 ) | ( ~n1783 & n7362 ) | ( n7361 & n7362 ) ;
  assign n7364 = ( ~n1643 & n7360 ) | ( ~n1643 & n7363 ) | ( n7360 & n7363 ) ;
  assign n7365 = ( n1822 & n7360 ) | ( n1822 & n7363 ) | ( n7360 & n7363 ) ;
  assign n7366 = ( n1324 & n7364 ) | ( n1324 & n7365 ) | ( n7364 & n7365 ) ;
  assign n7367 = n7357 | n7366 ;
  assign n7368 = x419 & n991 ;
  assign n7369 = x419 & ~n995 ;
  assign n7370 = ( ~n1104 & n7368 ) | ( ~n1104 & n7369 ) | ( n7368 & n7369 ) ;
  assign n7371 = ( ~n1119 & n7368 ) | ( ~n1119 & n7369 ) | ( n7368 & n7369 ) ;
  assign n7372 = ( n1126 & n7368 ) | ( n1126 & n7369 ) | ( n7368 & n7369 ) ;
  assign n7373 = ( n1115 & n7371 ) | ( n1115 & n7372 ) | ( n7371 & n7372 ) ;
  assign n7374 = ( n975 & n7370 ) | ( n975 & n7373 ) | ( n7370 & n7373 ) ;
  assign n7375 = ( ~n1154 & n7370 ) | ( ~n1154 & n7373 ) | ( n7370 & n7373 ) ;
  assign n7376 = ( x409 & n7374 ) | ( x409 & n7375 ) | ( n7374 & n7375 ) ;
  assign n7377 = ( ~x281 & n7374 ) | ( ~x281 & n7375 ) | ( n7374 & n7375 ) ;
  assign n7378 = ( ~n656 & n7376 ) | ( ~n656 & n7377 ) | ( n7376 & n7377 ) ;
  assign n7379 = x291 & ~n991 ;
  assign n7380 = x291 & n995 ;
  assign n7381 = ( n1104 & n7379 ) | ( n1104 & n7380 ) | ( n7379 & n7380 ) ;
  assign n7382 = ( n1119 & n7379 ) | ( n1119 & n7380 ) | ( n7379 & n7380 ) ;
  assign n7383 = ( ~n1126 & n7379 ) | ( ~n1126 & n7380 ) | ( n7379 & n7380 ) ;
  assign n7384 = ( ~n1115 & n7382 ) | ( ~n1115 & n7383 ) | ( n7382 & n7383 ) ;
  assign n7385 = ( ~n975 & n7381 ) | ( ~n975 & n7384 ) | ( n7381 & n7384 ) ;
  assign n7386 = ( n1154 & n7381 ) | ( n1154 & n7384 ) | ( n7381 & n7384 ) ;
  assign n7387 = ( ~x409 & n7385 ) | ( ~x409 & n7386 ) | ( n7385 & n7386 ) ;
  assign n7388 = ( x281 & n7385 ) | ( x281 & n7386 ) | ( n7385 & n7386 ) ;
  assign n7389 = ( n656 & n7387 ) | ( n656 & n7388 ) | ( n7387 & n7388 ) ;
  assign n7390 = n7378 | n7389 ;
  assign n7391 = ~n7367 & n7390 ;
  assign n7392 = x418 & n991 ;
  assign n7393 = x418 & ~n995 ;
  assign n7394 = ( ~n1104 & n7392 ) | ( ~n1104 & n7393 ) | ( n7392 & n7393 ) ;
  assign n7395 = ( ~n1119 & n7392 ) | ( ~n1119 & n7393 ) | ( n7392 & n7393 ) ;
  assign n7396 = ( n1126 & n7392 ) | ( n1126 & n7393 ) | ( n7392 & n7393 ) ;
  assign n7397 = ( n1115 & n7395 ) | ( n1115 & n7396 ) | ( n7395 & n7396 ) ;
  assign n7398 = ( n975 & n7394 ) | ( n975 & n7397 ) | ( n7394 & n7397 ) ;
  assign n7399 = ( ~n1154 & n7394 ) | ( ~n1154 & n7397 ) | ( n7394 & n7397 ) ;
  assign n7400 = ( x409 & n7398 ) | ( x409 & n7399 ) | ( n7398 & n7399 ) ;
  assign n7401 = ( ~x281 & n7398 ) | ( ~x281 & n7399 ) | ( n7398 & n7399 ) ;
  assign n7402 = ( ~n656 & n7400 ) | ( ~n656 & n7401 ) | ( n7400 & n7401 ) ;
  assign n7403 = x290 & ~n991 ;
  assign n7404 = x290 & n995 ;
  assign n7405 = ( n1104 & n7403 ) | ( n1104 & n7404 ) | ( n7403 & n7404 ) ;
  assign n7406 = ( n1119 & n7403 ) | ( n1119 & n7404 ) | ( n7403 & n7404 ) ;
  assign n7407 = ( ~n1126 & n7403 ) | ( ~n1126 & n7404 ) | ( n7403 & n7404 ) ;
  assign n7408 = ( ~n1115 & n7406 ) | ( ~n1115 & n7407 ) | ( n7406 & n7407 ) ;
  assign n7409 = ( ~n975 & n7405 ) | ( ~n975 & n7408 ) | ( n7405 & n7408 ) ;
  assign n7410 = ( n1154 & n7405 ) | ( n1154 & n7408 ) | ( n7405 & n7408 ) ;
  assign n7411 = ( ~x409 & n7409 ) | ( ~x409 & n7410 ) | ( n7409 & n7410 ) ;
  assign n7412 = ( x281 & n7409 ) | ( x281 & n7410 ) | ( n7409 & n7410 ) ;
  assign n7413 = ( n656 & n7411 ) | ( n656 & n7412 ) | ( n7411 & n7412 ) ;
  assign n7414 = n7402 | n7413 ;
  assign n7415 = x162 & n1767 ;
  assign n7416 = x162 & ~n1771 ;
  assign n7417 = ( ~n1751 & n7415 ) | ( ~n1751 & n7416 ) | ( n7415 & n7416 ) ;
  assign n7418 = ( ~n1787 & n7415 ) | ( ~n1787 & n7416 ) | ( n7415 & n7416 ) ;
  assign n7419 = ( n1794 & n7415 ) | ( n1794 & n7416 ) | ( n7415 & n7416 ) ;
  assign n7420 = ( n1783 & n7418 ) | ( n1783 & n7419 ) | ( n7418 & n7419 ) ;
  assign n7421 = ( n1643 & n7417 ) | ( n1643 & n7420 ) | ( n7417 & n7420 ) ;
  assign n7422 = ( ~n1822 & n7417 ) | ( ~n1822 & n7420 ) | ( n7417 & n7420 ) ;
  assign n7423 = ( ~n1324 & n7421 ) | ( ~n1324 & n7422 ) | ( n7421 & n7422 ) ;
  assign n7424 = x34 & ~n1767 ;
  assign n7425 = x34 & n1771 ;
  assign n7426 = ( n1751 & n7424 ) | ( n1751 & n7425 ) | ( n7424 & n7425 ) ;
  assign n7427 = ( n1787 & n7424 ) | ( n1787 & n7425 ) | ( n7424 & n7425 ) ;
  assign n7428 = ( ~n1794 & n7424 ) | ( ~n1794 & n7425 ) | ( n7424 & n7425 ) ;
  assign n7429 = ( ~n1783 & n7427 ) | ( ~n1783 & n7428 ) | ( n7427 & n7428 ) ;
  assign n7430 = ( ~n1643 & n7426 ) | ( ~n1643 & n7429 ) | ( n7426 & n7429 ) ;
  assign n7431 = ( n1822 & n7426 ) | ( n1822 & n7429 ) | ( n7426 & n7429 ) ;
  assign n7432 = ( n1324 & n7430 ) | ( n1324 & n7431 ) | ( n7430 & n7431 ) ;
  assign n7433 = n7423 | n7432 ;
  assign n7434 = n7414 & ~n7433 ;
  assign n7435 = n7391 | n7434 ;
  assign n7436 = n7348 | n7435 ;
  assign n7437 = n7305 | n7436 ;
  assign n7438 = n7130 | n7437 ;
  assign n7439 = x159 & n1767 ;
  assign n7440 = x159 & ~n1771 ;
  assign n7441 = ( ~n1751 & n7439 ) | ( ~n1751 & n7440 ) | ( n7439 & n7440 ) ;
  assign n7442 = ( ~n1787 & n7439 ) | ( ~n1787 & n7440 ) | ( n7439 & n7440 ) ;
  assign n7443 = ( n1794 & n7439 ) | ( n1794 & n7440 ) | ( n7439 & n7440 ) ;
  assign n7444 = ( n1783 & n7442 ) | ( n1783 & n7443 ) | ( n7442 & n7443 ) ;
  assign n7445 = ( n1643 & n7441 ) | ( n1643 & n7444 ) | ( n7441 & n7444 ) ;
  assign n7446 = ( ~n1822 & n7441 ) | ( ~n1822 & n7444 ) | ( n7441 & n7444 ) ;
  assign n7447 = ( ~n1324 & n7445 ) | ( ~n1324 & n7446 ) | ( n7445 & n7446 ) ;
  assign n7448 = x31 & ~n1767 ;
  assign n7449 = x31 & n1771 ;
  assign n7450 = ( n1751 & n7448 ) | ( n1751 & n7449 ) | ( n7448 & n7449 ) ;
  assign n7451 = ( n1787 & n7448 ) | ( n1787 & n7449 ) | ( n7448 & n7449 ) ;
  assign n7452 = ( ~n1794 & n7448 ) | ( ~n1794 & n7449 ) | ( n7448 & n7449 ) ;
  assign n7453 = ( ~n1783 & n7451 ) | ( ~n1783 & n7452 ) | ( n7451 & n7452 ) ;
  assign n7454 = ( ~n1643 & n7450 ) | ( ~n1643 & n7453 ) | ( n7450 & n7453 ) ;
  assign n7455 = ( n1822 & n7450 ) | ( n1822 & n7453 ) | ( n7450 & n7453 ) ;
  assign n7456 = ( n1324 & n7454 ) | ( n1324 & n7455 ) | ( n7454 & n7455 ) ;
  assign n7457 = n7447 | n7456 ;
  assign n7458 = x415 & n991 ;
  assign n7459 = x415 & ~n995 ;
  assign n7460 = ( ~n1104 & n7458 ) | ( ~n1104 & n7459 ) | ( n7458 & n7459 ) ;
  assign n7461 = ( ~n1119 & n7458 ) | ( ~n1119 & n7459 ) | ( n7458 & n7459 ) ;
  assign n7462 = ( n1126 & n7458 ) | ( n1126 & n7459 ) | ( n7458 & n7459 ) ;
  assign n7463 = ( n1115 & n7461 ) | ( n1115 & n7462 ) | ( n7461 & n7462 ) ;
  assign n7464 = ( n975 & n7460 ) | ( n975 & n7463 ) | ( n7460 & n7463 ) ;
  assign n7465 = ( ~n1154 & n7460 ) | ( ~n1154 & n7463 ) | ( n7460 & n7463 ) ;
  assign n7466 = ( x409 & n7464 ) | ( x409 & n7465 ) | ( n7464 & n7465 ) ;
  assign n7467 = ( ~x281 & n7464 ) | ( ~x281 & n7465 ) | ( n7464 & n7465 ) ;
  assign n7468 = ( ~n656 & n7466 ) | ( ~n656 & n7467 ) | ( n7466 & n7467 ) ;
  assign n7469 = x287 & ~n991 ;
  assign n7470 = x287 & n995 ;
  assign n7471 = ( n1104 & n7469 ) | ( n1104 & n7470 ) | ( n7469 & n7470 ) ;
  assign n7472 = ( n1119 & n7469 ) | ( n1119 & n7470 ) | ( n7469 & n7470 ) ;
  assign n7473 = ( ~n1126 & n7469 ) | ( ~n1126 & n7470 ) | ( n7469 & n7470 ) ;
  assign n7474 = ( ~n1115 & n7472 ) | ( ~n1115 & n7473 ) | ( n7472 & n7473 ) ;
  assign n7475 = ( ~n975 & n7471 ) | ( ~n975 & n7474 ) | ( n7471 & n7474 ) ;
  assign n7476 = ( n1154 & n7471 ) | ( n1154 & n7474 ) | ( n7471 & n7474 ) ;
  assign n7477 = ( ~x409 & n7475 ) | ( ~x409 & n7476 ) | ( n7475 & n7476 ) ;
  assign n7478 = ( x281 & n7475 ) | ( x281 & n7476 ) | ( n7475 & n7476 ) ;
  assign n7479 = ( n656 & n7477 ) | ( n656 & n7478 ) | ( n7477 & n7478 ) ;
  assign n7480 = n7468 | n7479 ;
  assign n7481 = n7457 & ~n7480 ;
  assign n7482 = ~n7457 & n7480 ;
  assign n7483 = x158 & n1767 ;
  assign n7484 = x158 & ~n1771 ;
  assign n7485 = ( ~n1751 & n7483 ) | ( ~n1751 & n7484 ) | ( n7483 & n7484 ) ;
  assign n7486 = ( ~n1787 & n7483 ) | ( ~n1787 & n7484 ) | ( n7483 & n7484 ) ;
  assign n7487 = ( n1794 & n7483 ) | ( n1794 & n7484 ) | ( n7483 & n7484 ) ;
  assign n7488 = ( n1783 & n7486 ) | ( n1783 & n7487 ) | ( n7486 & n7487 ) ;
  assign n7489 = ( n1643 & n7485 ) | ( n1643 & n7488 ) | ( n7485 & n7488 ) ;
  assign n7490 = ( ~n1822 & n7485 ) | ( ~n1822 & n7488 ) | ( n7485 & n7488 ) ;
  assign n7491 = ( ~n1324 & n7489 ) | ( ~n1324 & n7490 ) | ( n7489 & n7490 ) ;
  assign n7492 = x30 & ~n1767 ;
  assign n7493 = x30 & n1771 ;
  assign n7494 = ( n1751 & n7492 ) | ( n1751 & n7493 ) | ( n7492 & n7493 ) ;
  assign n7495 = ( n1787 & n7492 ) | ( n1787 & n7493 ) | ( n7492 & n7493 ) ;
  assign n7496 = ( ~n1794 & n7492 ) | ( ~n1794 & n7493 ) | ( n7492 & n7493 ) ;
  assign n7497 = ( ~n1783 & n7495 ) | ( ~n1783 & n7496 ) | ( n7495 & n7496 ) ;
  assign n7498 = ( ~n1643 & n7494 ) | ( ~n1643 & n7497 ) | ( n7494 & n7497 ) ;
  assign n7499 = ( n1822 & n7494 ) | ( n1822 & n7497 ) | ( n7494 & n7497 ) ;
  assign n7500 = ( n1324 & n7498 ) | ( n1324 & n7499 ) | ( n7498 & n7499 ) ;
  assign n7501 = n7491 | n7500 ;
  assign n7502 = x414 & n991 ;
  assign n7503 = x414 & ~n995 ;
  assign n7504 = ( ~n1104 & n7502 ) | ( ~n1104 & n7503 ) | ( n7502 & n7503 ) ;
  assign n7505 = ( ~n1119 & n7502 ) | ( ~n1119 & n7503 ) | ( n7502 & n7503 ) ;
  assign n7506 = ( n1126 & n7502 ) | ( n1126 & n7503 ) | ( n7502 & n7503 ) ;
  assign n7507 = ( n1115 & n7505 ) | ( n1115 & n7506 ) | ( n7505 & n7506 ) ;
  assign n7508 = ( n975 & n7504 ) | ( n975 & n7507 ) | ( n7504 & n7507 ) ;
  assign n7509 = ( ~n1154 & n7504 ) | ( ~n1154 & n7507 ) | ( n7504 & n7507 ) ;
  assign n7510 = ( x409 & n7508 ) | ( x409 & n7509 ) | ( n7508 & n7509 ) ;
  assign n7511 = ( ~x281 & n7508 ) | ( ~x281 & n7509 ) | ( n7508 & n7509 ) ;
  assign n7512 = ( ~n656 & n7510 ) | ( ~n656 & n7511 ) | ( n7510 & n7511 ) ;
  assign n7513 = x286 & ~n991 ;
  assign n7514 = x286 & n995 ;
  assign n7515 = ( n1104 & n7513 ) | ( n1104 & n7514 ) | ( n7513 & n7514 ) ;
  assign n7516 = ( n1119 & n7513 ) | ( n1119 & n7514 ) | ( n7513 & n7514 ) ;
  assign n7517 = ( ~n1126 & n7513 ) | ( ~n1126 & n7514 ) | ( n7513 & n7514 ) ;
  assign n7518 = ( ~n1115 & n7516 ) | ( ~n1115 & n7517 ) | ( n7516 & n7517 ) ;
  assign n7519 = ( ~n975 & n7515 ) | ( ~n975 & n7518 ) | ( n7515 & n7518 ) ;
  assign n7520 = ( n1154 & n7515 ) | ( n1154 & n7518 ) | ( n7515 & n7518 ) ;
  assign n7521 = ( ~x409 & n7519 ) | ( ~x409 & n7520 ) | ( n7519 & n7520 ) ;
  assign n7522 = ( x281 & n7519 ) | ( x281 & n7520 ) | ( n7519 & n7520 ) ;
  assign n7523 = ( n656 & n7521 ) | ( n656 & n7522 ) | ( n7521 & n7522 ) ;
  assign n7524 = n7512 | n7523 ;
  assign n7525 = n7501 & ~n7524 ;
  assign n7526 = ~n7501 & n7524 ;
  assign n7527 = ~n7525 & n7526 ;
  assign n7528 = n7482 | n7527 ;
  assign n7529 = x157 & n1767 ;
  assign n7530 = x157 & ~n1771 ;
  assign n7531 = ( ~n1751 & n7529 ) | ( ~n1751 & n7530 ) | ( n7529 & n7530 ) ;
  assign n7532 = ( ~n1787 & n7529 ) | ( ~n1787 & n7530 ) | ( n7529 & n7530 ) ;
  assign n7533 = ( n1794 & n7529 ) | ( n1794 & n7530 ) | ( n7529 & n7530 ) ;
  assign n7534 = ( n1783 & n7532 ) | ( n1783 & n7533 ) | ( n7532 & n7533 ) ;
  assign n7535 = ( n1643 & n7531 ) | ( n1643 & n7534 ) | ( n7531 & n7534 ) ;
  assign n7536 = ( ~n1822 & n7531 ) | ( ~n1822 & n7534 ) | ( n7531 & n7534 ) ;
  assign n7537 = ( ~n1324 & n7535 ) | ( ~n1324 & n7536 ) | ( n7535 & n7536 ) ;
  assign n7538 = x29 & ~n1767 ;
  assign n7539 = x29 & n1771 ;
  assign n7540 = ( n1751 & n7538 ) | ( n1751 & n7539 ) | ( n7538 & n7539 ) ;
  assign n7541 = ( n1787 & n7538 ) | ( n1787 & n7539 ) | ( n7538 & n7539 ) ;
  assign n7542 = ( ~n1794 & n7538 ) | ( ~n1794 & n7539 ) | ( n7538 & n7539 ) ;
  assign n7543 = ( ~n1783 & n7541 ) | ( ~n1783 & n7542 ) | ( n7541 & n7542 ) ;
  assign n7544 = ( ~n1643 & n7540 ) | ( ~n1643 & n7543 ) | ( n7540 & n7543 ) ;
  assign n7545 = ( n1822 & n7540 ) | ( n1822 & n7543 ) | ( n7540 & n7543 ) ;
  assign n7546 = ( n1324 & n7544 ) | ( n1324 & n7545 ) | ( n7544 & n7545 ) ;
  assign n7547 = n7537 | n7546 ;
  assign n7548 = x413 & n991 ;
  assign n7549 = x413 & ~n995 ;
  assign n7550 = ( ~n1104 & n7548 ) | ( ~n1104 & n7549 ) | ( n7548 & n7549 ) ;
  assign n7551 = ( ~n1119 & n7548 ) | ( ~n1119 & n7549 ) | ( n7548 & n7549 ) ;
  assign n7552 = ( n1126 & n7548 ) | ( n1126 & n7549 ) | ( n7548 & n7549 ) ;
  assign n7553 = ( n1115 & n7551 ) | ( n1115 & n7552 ) | ( n7551 & n7552 ) ;
  assign n7554 = ( n975 & n7550 ) | ( n975 & n7553 ) | ( n7550 & n7553 ) ;
  assign n7555 = ( ~n1154 & n7550 ) | ( ~n1154 & n7553 ) | ( n7550 & n7553 ) ;
  assign n7556 = ( x409 & n7554 ) | ( x409 & n7555 ) | ( n7554 & n7555 ) ;
  assign n7557 = ( ~x281 & n7554 ) | ( ~x281 & n7555 ) | ( n7554 & n7555 ) ;
  assign n7558 = ( ~n656 & n7556 ) | ( ~n656 & n7557 ) | ( n7556 & n7557 ) ;
  assign n7559 = x285 & ~n991 ;
  assign n7560 = x285 & n995 ;
  assign n7561 = ( n1104 & n7559 ) | ( n1104 & n7560 ) | ( n7559 & n7560 ) ;
  assign n7562 = ( n1119 & n7559 ) | ( n1119 & n7560 ) | ( n7559 & n7560 ) ;
  assign n7563 = ( ~n1126 & n7559 ) | ( ~n1126 & n7560 ) | ( n7559 & n7560 ) ;
  assign n7564 = ( ~n1115 & n7562 ) | ( ~n1115 & n7563 ) | ( n7562 & n7563 ) ;
  assign n7565 = ( ~n975 & n7561 ) | ( ~n975 & n7564 ) | ( n7561 & n7564 ) ;
  assign n7566 = ( n1154 & n7561 ) | ( n1154 & n7564 ) | ( n7561 & n7564 ) ;
  assign n7567 = ( ~x409 & n7565 ) | ( ~x409 & n7566 ) | ( n7565 & n7566 ) ;
  assign n7568 = ( x281 & n7565 ) | ( x281 & n7566 ) | ( n7565 & n7566 ) ;
  assign n7569 = ( n656 & n7567 ) | ( n656 & n7568 ) | ( n7567 & n7568 ) ;
  assign n7570 = n7558 | n7569 ;
  assign n7571 = ~n7547 & n7570 ;
  assign n7572 = x156 & n1767 ;
  assign n7573 = x156 & ~n1771 ;
  assign n7574 = ( ~n1751 & n7572 ) | ( ~n1751 & n7573 ) | ( n7572 & n7573 ) ;
  assign n7575 = ( ~n1787 & n7572 ) | ( ~n1787 & n7573 ) | ( n7572 & n7573 ) ;
  assign n7576 = ( n1794 & n7572 ) | ( n1794 & n7573 ) | ( n7572 & n7573 ) ;
  assign n7577 = ( n1783 & n7575 ) | ( n1783 & n7576 ) | ( n7575 & n7576 ) ;
  assign n7578 = ( n1643 & n7574 ) | ( n1643 & n7577 ) | ( n7574 & n7577 ) ;
  assign n7579 = ( ~n1822 & n7574 ) | ( ~n1822 & n7577 ) | ( n7574 & n7577 ) ;
  assign n7580 = ( ~n1324 & n7578 ) | ( ~n1324 & n7579 ) | ( n7578 & n7579 ) ;
  assign n7581 = x28 & ~n1767 ;
  assign n7582 = x28 & n1771 ;
  assign n7583 = ( n1751 & n7581 ) | ( n1751 & n7582 ) | ( n7581 & n7582 ) ;
  assign n7584 = ( n1787 & n7581 ) | ( n1787 & n7582 ) | ( n7581 & n7582 ) ;
  assign n7585 = ( ~n1794 & n7581 ) | ( ~n1794 & n7582 ) | ( n7581 & n7582 ) ;
  assign n7586 = ( ~n1783 & n7584 ) | ( ~n1783 & n7585 ) | ( n7584 & n7585 ) ;
  assign n7587 = ( ~n1643 & n7583 ) | ( ~n1643 & n7586 ) | ( n7583 & n7586 ) ;
  assign n7588 = ( n1822 & n7583 ) | ( n1822 & n7586 ) | ( n7583 & n7586 ) ;
  assign n7589 = ( n1324 & n7587 ) | ( n1324 & n7588 ) | ( n7587 & n7588 ) ;
  assign n7590 = n7580 | n7589 ;
  assign n7591 = x412 & n991 ;
  assign n7592 = x412 & ~n995 ;
  assign n7593 = ( ~n1104 & n7591 ) | ( ~n1104 & n7592 ) | ( n7591 & n7592 ) ;
  assign n7594 = ( ~n1119 & n7591 ) | ( ~n1119 & n7592 ) | ( n7591 & n7592 ) ;
  assign n7595 = ( n1126 & n7591 ) | ( n1126 & n7592 ) | ( n7591 & n7592 ) ;
  assign n7596 = ( n1115 & n7594 ) | ( n1115 & n7595 ) | ( n7594 & n7595 ) ;
  assign n7597 = ( n975 & n7593 ) | ( n975 & n7596 ) | ( n7593 & n7596 ) ;
  assign n7598 = ( ~n1154 & n7593 ) | ( ~n1154 & n7596 ) | ( n7593 & n7596 ) ;
  assign n7599 = ( x409 & n7597 ) | ( x409 & n7598 ) | ( n7597 & n7598 ) ;
  assign n7600 = ( ~x281 & n7597 ) | ( ~x281 & n7598 ) | ( n7597 & n7598 ) ;
  assign n7601 = ( ~n656 & n7599 ) | ( ~n656 & n7600 ) | ( n7599 & n7600 ) ;
  assign n7602 = x284 & ~n991 ;
  assign n7603 = x284 & n995 ;
  assign n7604 = ( n1104 & n7602 ) | ( n1104 & n7603 ) | ( n7602 & n7603 ) ;
  assign n7605 = ( n1119 & n7602 ) | ( n1119 & n7603 ) | ( n7602 & n7603 ) ;
  assign n7606 = ( ~n1126 & n7602 ) | ( ~n1126 & n7603 ) | ( n7602 & n7603 ) ;
  assign n7607 = ( ~n1115 & n7605 ) | ( ~n1115 & n7606 ) | ( n7605 & n7606 ) ;
  assign n7608 = ( ~n975 & n7604 ) | ( ~n975 & n7607 ) | ( n7604 & n7607 ) ;
  assign n7609 = ( n1154 & n7604 ) | ( n1154 & n7607 ) | ( n7604 & n7607 ) ;
  assign n7610 = ( ~x409 & n7608 ) | ( ~x409 & n7609 ) | ( n7608 & n7609 ) ;
  assign n7611 = ( x281 & n7608 ) | ( x281 & n7609 ) | ( n7608 & n7609 ) ;
  assign n7612 = ( n656 & n7610 ) | ( n656 & n7611 ) | ( n7610 & n7611 ) ;
  assign n7613 = n7601 | n7612 ;
  assign n7614 = n7590 & ~n7613 ;
  assign n7615 = ~n7571 & n7614 ;
  assign n7616 = x155 & n1767 ;
  assign n7617 = x155 & ~n1771 ;
  assign n7618 = ( ~n1751 & n7616 ) | ( ~n1751 & n7617 ) | ( n7616 & n7617 ) ;
  assign n7619 = ( ~n1787 & n7616 ) | ( ~n1787 & n7617 ) | ( n7616 & n7617 ) ;
  assign n7620 = ( n1794 & n7616 ) | ( n1794 & n7617 ) | ( n7616 & n7617 ) ;
  assign n7621 = ( n1783 & n7619 ) | ( n1783 & n7620 ) | ( n7619 & n7620 ) ;
  assign n7622 = ( n1643 & n7618 ) | ( n1643 & n7621 ) | ( n7618 & n7621 ) ;
  assign n7623 = ( ~n1822 & n7618 ) | ( ~n1822 & n7621 ) | ( n7618 & n7621 ) ;
  assign n7624 = ( ~n1324 & n7622 ) | ( ~n1324 & n7623 ) | ( n7622 & n7623 ) ;
  assign n7625 = x27 & ~n1767 ;
  assign n7626 = x27 & n1771 ;
  assign n7627 = ( n1751 & n7625 ) | ( n1751 & n7626 ) | ( n7625 & n7626 ) ;
  assign n7628 = ( n1787 & n7625 ) | ( n1787 & n7626 ) | ( n7625 & n7626 ) ;
  assign n7629 = ( ~n1794 & n7625 ) | ( ~n1794 & n7626 ) | ( n7625 & n7626 ) ;
  assign n7630 = ( ~n1783 & n7628 ) | ( ~n1783 & n7629 ) | ( n7628 & n7629 ) ;
  assign n7631 = ( ~n1643 & n7627 ) | ( ~n1643 & n7630 ) | ( n7627 & n7630 ) ;
  assign n7632 = ( n1822 & n7627 ) | ( n1822 & n7630 ) | ( n7627 & n7630 ) ;
  assign n7633 = ( n1324 & n7631 ) | ( n1324 & n7632 ) | ( n7631 & n7632 ) ;
  assign n7634 = n7624 | n7633 ;
  assign n7635 = x411 & n991 ;
  assign n7636 = x411 & ~n995 ;
  assign n7637 = ( ~n1104 & n7635 ) | ( ~n1104 & n7636 ) | ( n7635 & n7636 ) ;
  assign n7638 = ( ~n1119 & n7635 ) | ( ~n1119 & n7636 ) | ( n7635 & n7636 ) ;
  assign n7639 = ( n1126 & n7635 ) | ( n1126 & n7636 ) | ( n7635 & n7636 ) ;
  assign n7640 = ( n1115 & n7638 ) | ( n1115 & n7639 ) | ( n7638 & n7639 ) ;
  assign n7641 = ( n975 & n7637 ) | ( n975 & n7640 ) | ( n7637 & n7640 ) ;
  assign n7642 = ( ~n1154 & n7637 ) | ( ~n1154 & n7640 ) | ( n7637 & n7640 ) ;
  assign n7643 = ( x409 & n7641 ) | ( x409 & n7642 ) | ( n7641 & n7642 ) ;
  assign n7644 = ( ~x281 & n7641 ) | ( ~x281 & n7642 ) | ( n7641 & n7642 ) ;
  assign n7645 = ( ~n656 & n7643 ) | ( ~n656 & n7644 ) | ( n7643 & n7644 ) ;
  assign n7646 = x283 & ~n991 ;
  assign n7647 = x283 & n995 ;
  assign n7648 = ( n1104 & n7646 ) | ( n1104 & n7647 ) | ( n7646 & n7647 ) ;
  assign n7649 = ( n1119 & n7646 ) | ( n1119 & n7647 ) | ( n7646 & n7647 ) ;
  assign n7650 = ( ~n1126 & n7646 ) | ( ~n1126 & n7647 ) | ( n7646 & n7647 ) ;
  assign n7651 = ( ~n1115 & n7649 ) | ( ~n1115 & n7650 ) | ( n7649 & n7650 ) ;
  assign n7652 = ( ~n975 & n7648 ) | ( ~n975 & n7651 ) | ( n7648 & n7651 ) ;
  assign n7653 = ( n1154 & n7648 ) | ( n1154 & n7651 ) | ( n7648 & n7651 ) ;
  assign n7654 = ( ~x409 & n7652 ) | ( ~x409 & n7653 ) | ( n7652 & n7653 ) ;
  assign n7655 = ( x281 & n7652 ) | ( x281 & n7653 ) | ( n7652 & n7653 ) ;
  assign n7656 = ( n656 & n7654 ) | ( n656 & n7655 ) | ( n7654 & n7655 ) ;
  assign n7657 = n7645 | n7656 ;
  assign n7658 = x154 & n1767 ;
  assign n7659 = x154 & ~n1771 ;
  assign n7660 = ( ~n1751 & n7658 ) | ( ~n1751 & n7659 ) | ( n7658 & n7659 ) ;
  assign n7661 = ( ~n1787 & n7658 ) | ( ~n1787 & n7659 ) | ( n7658 & n7659 ) ;
  assign n7662 = ( n1794 & n7658 ) | ( n1794 & n7659 ) | ( n7658 & n7659 ) ;
  assign n7663 = ( n1783 & n7661 ) | ( n1783 & n7662 ) | ( n7661 & n7662 ) ;
  assign n7664 = ( n1643 & n7660 ) | ( n1643 & n7663 ) | ( n7660 & n7663 ) ;
  assign n7665 = ( ~n1822 & n7660 ) | ( ~n1822 & n7663 ) | ( n7660 & n7663 ) ;
  assign n7666 = ( ~n1324 & n7664 ) | ( ~n1324 & n7665 ) | ( n7664 & n7665 ) ;
  assign n7667 = x26 & ~n1767 ;
  assign n7668 = x26 & n1771 ;
  assign n7669 = ( n1751 & n7667 ) | ( n1751 & n7668 ) | ( n7667 & n7668 ) ;
  assign n7670 = ( n1787 & n7667 ) | ( n1787 & n7668 ) | ( n7667 & n7668 ) ;
  assign n7671 = ( ~n1794 & n7667 ) | ( ~n1794 & n7668 ) | ( n7667 & n7668 ) ;
  assign n7672 = ( ~n1783 & n7670 ) | ( ~n1783 & n7671 ) | ( n7670 & n7671 ) ;
  assign n7673 = ( ~n1643 & n7669 ) | ( ~n1643 & n7672 ) | ( n7669 & n7672 ) ;
  assign n7674 = ( n1822 & n7669 ) | ( n1822 & n7672 ) | ( n7669 & n7672 ) ;
  assign n7675 = ( n1324 & n7673 ) | ( n1324 & n7674 ) | ( n7673 & n7674 ) ;
  assign n7676 = n7666 | n7675 ;
  assign n7677 = x410 & n991 ;
  assign n7678 = x410 & ~n995 ;
  assign n7679 = ( ~n1104 & n7677 ) | ( ~n1104 & n7678 ) | ( n7677 & n7678 ) ;
  assign n7680 = ( ~n1119 & n7677 ) | ( ~n1119 & n7678 ) | ( n7677 & n7678 ) ;
  assign n7681 = ( n1126 & n7677 ) | ( n1126 & n7678 ) | ( n7677 & n7678 ) ;
  assign n7682 = ( n1115 & n7680 ) | ( n1115 & n7681 ) | ( n7680 & n7681 ) ;
  assign n7683 = ( n975 & n7679 ) | ( n975 & n7682 ) | ( n7679 & n7682 ) ;
  assign n7684 = ( ~n1154 & n7679 ) | ( ~n1154 & n7682 ) | ( n7679 & n7682 ) ;
  assign n7685 = ( x409 & n7683 ) | ( x409 & n7684 ) | ( n7683 & n7684 ) ;
  assign n7686 = ( ~x281 & n7683 ) | ( ~x281 & n7684 ) | ( n7683 & n7684 ) ;
  assign n7687 = ( ~n656 & n7685 ) | ( ~n656 & n7686 ) | ( n7685 & n7686 ) ;
  assign n7688 = x282 & ~n991 ;
  assign n7689 = x282 & n995 ;
  assign n7690 = ( n1104 & n7688 ) | ( n1104 & n7689 ) | ( n7688 & n7689 ) ;
  assign n7691 = ( n1119 & n7688 ) | ( n1119 & n7689 ) | ( n7688 & n7689 ) ;
  assign n7692 = ( ~n1126 & n7688 ) | ( ~n1126 & n7689 ) | ( n7688 & n7689 ) ;
  assign n7693 = ( ~n1115 & n7691 ) | ( ~n1115 & n7692 ) | ( n7691 & n7692 ) ;
  assign n7694 = ( ~n975 & n7690 ) | ( ~n975 & n7693 ) | ( n7690 & n7693 ) ;
  assign n7695 = ( n1154 & n7690 ) | ( n1154 & n7693 ) | ( n7690 & n7693 ) ;
  assign n7696 = ( ~x409 & n7694 ) | ( ~x409 & n7695 ) | ( n7694 & n7695 ) ;
  assign n7697 = ( x281 & n7694 ) | ( x281 & n7695 ) | ( n7694 & n7695 ) ;
  assign n7698 = ( n656 & n7696 ) | ( n656 & n7697 ) | ( n7696 & n7697 ) ;
  assign n7699 = n7687 | n7698 ;
  assign n7700 = ~n7676 & n7699 ;
  assign n7701 = ( ~n7634 & n7657 ) | ( ~n7634 & n7700 ) | ( n7657 & n7700 ) ;
  assign n7702 = ~n7590 & n7613 ;
  assign n7703 = n7571 | n7702 ;
  assign n7704 = ( ~n7615 & n7701 ) | ( ~n7615 & n7703 ) | ( n7701 & n7703 ) ;
  assign n7705 = ~n7482 & n7525 ;
  assign n7706 = n7547 & ~n7570 ;
  assign n7707 = ~n7526 & n7706 ;
  assign n7708 = ( ~n7482 & n7705 ) | ( ~n7482 & n7707 ) | ( n7705 & n7707 ) ;
  assign n7709 = ( n7528 & n7704 ) | ( n7528 & ~n7708 ) | ( n7704 & ~n7708 ) ;
  assign n7710 = ( n7438 & ~n7481 ) | ( n7438 & n7709 ) | ( ~n7481 & n7709 ) ;
  assign n7711 = n7438 | n7710 ;
  assign n7712 = ~n7414 & n7433 ;
  assign n7713 = ~n7391 & n7712 ;
  assign n7714 = ~n7110 & n7129 ;
  assign n7715 = n7324 & ~n7347 ;
  assign n7716 = n7714 | n7715 ;
  assign n7717 = n7713 | n7716 ;
  assign n7718 = ( ~n7436 & n7713 ) | ( ~n7436 & n7717 ) | ( n7713 & n7717 ) ;
  assign n7719 = n7367 & ~n7390 ;
  assign n7720 = ~n7305 & n7719 ;
  assign n7721 = ( ~n7305 & n7718 ) | ( ~n7305 & n7720 ) | ( n7718 & n7720 ) ;
  assign n7722 = n7149 & ~n7172 ;
  assign n7723 = n7236 & ~n7259 ;
  assign n7724 = ( n7196 & ~n7215 ) | ( n7196 & n7302 ) | ( ~n7215 & n7302 ) ;
  assign n7725 = ( ~n7196 & n7215 ) | ( ~n7196 & n7279 ) | ( n7215 & n7279 ) ;
  assign n7726 = ( n7723 & ~n7724 ) | ( n7723 & n7725 ) | ( ~n7724 & n7725 ) ;
  assign n7727 = n7173 & ~n7722 ;
  assign n7728 = ( n7722 & n7726 ) | ( n7722 & ~n7727 ) | ( n7726 & ~n7727 ) ;
  assign n7729 = ~n7087 & n7728 ;
  assign n7730 = ( ~n7087 & n7721 ) | ( ~n7087 & n7729 ) | ( n7721 & n7729 ) ;
  assign n7731 = ( n7087 & n7711 ) | ( n7087 & ~n7730 ) | ( n7711 & ~n7730 ) ;
  assign n7732 = n6755 & ~n6778 ;
  assign n7733 = ~n6734 & n7732 ;
  assign n7734 = ~n6733 & n7733 ;
  assign n7735 = n7060 & ~n7083 ;
  assign n7736 = ( n7017 & ~n7040 ) | ( n7017 & n7735 ) | ( ~n7040 & n7735 ) ;
  assign n7737 = n6930 & ~n6953 ;
  assign n7738 = ~n6954 & n7737 ;
  assign n7739 = ( ~n6954 & n7736 ) | ( ~n6954 & n7738 ) | ( n7736 & n7738 ) ;
  assign n7740 = ( n6973 & ~n6996 ) | ( n6973 & n7739 ) | ( ~n6996 & n7739 ) ;
  assign n7741 = ~n6911 & n7740 ;
  assign n7742 = n6842 & ~n6865 ;
  assign n7743 = ( n6885 & ~n6908 ) | ( n6885 & n7742 ) | ( ~n6908 & n7742 ) ;
  assign n7744 = ~n6823 & n7743 ;
  assign n7745 = ~n6802 & n6821 ;
  assign n7746 = ~n6779 & n7745 ;
  assign n7747 = n7744 | n7746 ;
  assign n7748 = n7741 | n7747 ;
  assign n7749 = ( ~n6735 & n7734 ) | ( ~n6735 & n7748 ) | ( n7734 & n7748 ) ;
  assign n7750 = n6732 | n7749 ;
  assign n7751 = ( n6736 & n7731 ) | ( n6736 & ~n7750 ) | ( n7731 & ~n7750 ) ;
  assign n7752 = ( n6349 & ~n6367 ) | ( n6349 & n7751 ) | ( ~n6367 & n7751 ) ;
  assign n7753 = ( n5222 & ~n5237 ) | ( n5222 & n7752 ) | ( ~n5237 & n7752 ) ;
  assign n7754 = ( ~n4094 & n4109 ) | ( ~n4094 & n7753 ) | ( n4109 & n7753 ) ;
  assign n7755 = n6732 | n7734 ;
  assign n7756 = n7721 | n7728 ;
  assign n7757 = n7481 | n7705 ;
  assign n7758 = ~n7634 & n7657 ;
  assign n7759 = n7676 & ~n7699 ;
  assign n7760 = ~n7758 & n7759 ;
  assign n7761 = n7634 & ~n7657 ;
  assign n7762 = ~n7702 & n7761 ;
  assign n7763 = ( ~n7702 & n7760 ) | ( ~n7702 & n7762 ) | ( n7760 & n7762 ) ;
  assign n7764 = n7615 | n7706 ;
  assign n7765 = ( ~n7571 & n7763 ) | ( ~n7571 & n7764 ) | ( n7763 & n7764 ) ;
  assign n7766 = ~n7481 & n7482 ;
  assign n7767 = ( ~n7481 & n7527 ) | ( ~n7481 & n7766 ) | ( n7527 & n7766 ) ;
  assign n7768 = ( n7757 & n7765 ) | ( n7757 & ~n7767 ) | ( n7765 & ~n7767 ) ;
  assign n7769 = ~n7438 & n7768 ;
  assign n7770 = n7756 | n7769 ;
  assign n7771 = n7087 & ~n7747 ;
  assign n7772 = ~n7741 & n7771 ;
  assign n7773 = ( n7748 & n7770 ) | ( n7748 & ~n7772 ) | ( n7770 & ~n7772 ) ;
  assign n7774 = ( ~n6736 & n7755 ) | ( ~n6736 & n7773 ) | ( n7755 & n7773 ) ;
  assign n7775 = ( ~n6349 & n6367 ) | ( ~n6349 & n7774 ) | ( n6367 & n7774 ) ;
  assign n7776 = ( ~n5222 & n5237 ) | ( ~n5222 & n7775 ) | ( n5237 & n7775 ) ;
  assign n7777 = ( n4094 & ~n4109 ) | ( n4094 & n7776 ) | ( ~n4109 & n7776 ) ;
  assign n7778 = ( n3007 & ~n7754 ) | ( n3007 & n7777 ) | ( ~n7754 & n7777 ) ;
  assign n7779 = n1170 & ~n7778 ;
  assign n7780 = n1834 & n7778 ;
  assign n7781 = n7779 | n7780 ;
  assign n7782 = ( ~n4094 & n4109 ) | ( ~n4094 & n5222 ) | ( n4109 & n5222 ) ;
  assign n7783 = ( n4094 & ~n4109 ) | ( n4094 & n5237 ) | ( ~n4109 & n5237 ) ;
  assign n7784 = ( n7752 & n7782 ) | ( n7752 & ~n7783 ) | ( n7782 & ~n7783 ) ;
  assign n7785 = n1193 & n7784 ;
  assign n7786 = ( n7775 & ~n7782 ) | ( n7775 & n7783 ) | ( ~n7782 & n7783 ) ;
  assign n7787 = n1193 & ~n7786 ;
  assign n7788 = ( ~n3007 & n7785 ) | ( ~n3007 & n7787 ) | ( n7785 & n7787 ) ;
  assign n7789 = n1855 & ~n7784 ;
  assign n7790 = n1855 & n7786 ;
  assign n7791 = ( n3007 & n7789 ) | ( n3007 & n7790 ) | ( n7789 & n7790 ) ;
  assign n7792 = n7788 | n7791 ;
  assign n7793 = n1970 & n7784 ;
  assign n7794 = n1970 & ~n7786 ;
  assign n7795 = ( ~n3007 & n7793 ) | ( ~n3007 & n7794 ) | ( n7793 & n7794 ) ;
  assign n7796 = n1990 & ~n7784 ;
  assign n7797 = n1990 & n7786 ;
  assign n7798 = ( n3007 & n7796 ) | ( n3007 & n7797 ) | ( n7796 & n7797 ) ;
  assign n7799 = n7795 | n7798 ;
  assign n7800 = n1923 & n7784 ;
  assign n7801 = n1923 & ~n7786 ;
  assign n7802 = ( ~n3007 & n7800 ) | ( ~n3007 & n7801 ) | ( n7800 & n7801 ) ;
  assign n7803 = n1900 & ~n7784 ;
  assign n7804 = n1900 & n7786 ;
  assign n7805 = ( n3007 & n7803 ) | ( n3007 & n7804 ) | ( n7803 & n7804 ) ;
  assign n7806 = n7802 | n7805 ;
  assign n7807 = n1881 & n7784 ;
  assign n7808 = n1881 & ~n7786 ;
  assign n7809 = ( ~n3007 & n7807 ) | ( ~n3007 & n7808 ) | ( n7807 & n7808 ) ;
  assign n7810 = n1943 & ~n7784 ;
  assign n7811 = n1943 & n7786 ;
  assign n7812 = ( n3007 & n7810 ) | ( n3007 & n7811 ) | ( n7810 & n7811 ) ;
  assign n7813 = n7809 | n7812 ;
  assign n7814 = n2173 & n7784 ;
  assign n7815 = n2173 & ~n7786 ;
  assign n7816 = ( ~n3007 & n7814 ) | ( ~n3007 & n7815 ) | ( n7814 & n7815 ) ;
  assign n7817 = n2148 & ~n7784 ;
  assign n7818 = n2148 & n7786 ;
  assign n7819 = ( n3007 & n7817 ) | ( n3007 & n7818 ) | ( n7817 & n7818 ) ;
  assign n7820 = n7816 | n7819 ;
  assign n7821 = n2129 & n7784 ;
  assign n7822 = n2129 & ~n7786 ;
  assign n7823 = ( ~n3007 & n7821 ) | ( ~n3007 & n7822 ) | ( n7821 & n7822 ) ;
  assign n7824 = n2106 & ~n7784 ;
  assign n7825 = n2106 & n7786 ;
  assign n7826 = ( n3007 & n7824 ) | ( n3007 & n7825 ) | ( n7824 & n7825 ) ;
  assign n7827 = n7823 | n7826 ;
  assign n7828 = n2063 & n7784 ;
  assign n7829 = n2063 & ~n7786 ;
  assign n7830 = ( ~n3007 & n7828 ) | ( ~n3007 & n7829 ) | ( n7828 & n7829 ) ;
  assign n7831 = n2040 & ~n7784 ;
  assign n7832 = n2040 & n7786 ;
  assign n7833 = ( n3007 & n7831 ) | ( n3007 & n7832 ) | ( n7831 & n7832 ) ;
  assign n7834 = n7830 | n7833 ;
  assign n7835 = n2021 & n7784 ;
  assign n7836 = n2021 & ~n7786 ;
  assign n7837 = ( ~n3007 & n7835 ) | ( ~n3007 & n7836 ) | ( n7835 & n7836 ) ;
  assign n7838 = n2083 & ~n7784 ;
  assign n7839 = n2083 & n7786 ;
  assign n7840 = ( n3007 & n7838 ) | ( n3007 & n7839 ) | ( n7838 & n7839 ) ;
  assign n7841 = n7837 | n7840 ;
  assign n7842 = n2537 & n7784 ;
  assign n7843 = n2537 & ~n7786 ;
  assign n7844 = ( ~n3007 & n7842 ) | ( ~n3007 & n7843 ) | ( n7842 & n7843 ) ;
  assign n7845 = n2557 & ~n7784 ;
  assign n7846 = n2557 & n7786 ;
  assign n7847 = ( n3007 & n7845 ) | ( n3007 & n7846 ) | ( n7845 & n7846 ) ;
  assign n7848 = n7844 | n7847 ;
  assign n7849 = n2353 & n7784 ;
  assign n7850 = n2353 & ~n7786 ;
  assign n7851 = ( ~n3007 & n7849 ) | ( ~n3007 & n7850 ) | ( n7849 & n7850 ) ;
  assign n7852 = n2330 & ~n7784 ;
  assign n7853 = n2330 & n7786 ;
  assign n7854 = ( n3007 & n7852 ) | ( n3007 & n7853 ) | ( n7852 & n7853 ) ;
  assign n7855 = n7851 | n7854 ;
  assign n7856 = n2311 & n7784 ;
  assign n7857 = n2311 & ~n7786 ;
  assign n7858 = ( ~n3007 & n7856 ) | ( ~n3007 & n7857 ) | ( n7856 & n7857 ) ;
  assign n7859 = n2288 & ~n7784 ;
  assign n7860 = n2288 & n7786 ;
  assign n7861 = ( n3007 & n7859 ) | ( n3007 & n7860 ) | ( n7859 & n7860 ) ;
  assign n7862 = n7858 | n7861 ;
  assign n7863 = n2267 & n7784 ;
  assign n7864 = n2267 & ~n7786 ;
  assign n7865 = ( ~n3007 & n7863 ) | ( ~n3007 & n7864 ) | ( n7863 & n7864 ) ;
  assign n7866 = n2244 & ~n7784 ;
  assign n7867 = n2244 & n7786 ;
  assign n7868 = ( n3007 & n7866 ) | ( n3007 & n7867 ) | ( n7866 & n7867 ) ;
  assign n7869 = n7865 | n7868 ;
  assign n7870 = n2224 & n7784 ;
  assign n7871 = n2224 & ~n7786 ;
  assign n7872 = ( ~n3007 & n7870 ) | ( ~n3007 & n7871 ) | ( n7870 & n7871 ) ;
  assign n7873 = n2201 & ~n7784 ;
  assign n7874 = n2201 & n7786 ;
  assign n7875 = ( n3007 & n7873 ) | ( n3007 & n7874 ) | ( n7873 & n7874 ) ;
  assign n7876 = n7872 | n7875 ;
  assign n7877 = n2466 & n7784 ;
  assign n7878 = n2466 & ~n7786 ;
  assign n7879 = ( ~n3007 & n7877 ) | ( ~n3007 & n7878 ) | ( n7877 & n7878 ) ;
  assign n7880 = n2443 & ~n7784 ;
  assign n7881 = n2443 & n7786 ;
  assign n7882 = ( n3007 & n7880 ) | ( n3007 & n7881 ) | ( n7880 & n7881 ) ;
  assign n7883 = n7879 | n7882 ;
  assign n7884 = n2423 & n7784 ;
  assign n7885 = n2423 & ~n7786 ;
  assign n7886 = ( ~n3007 & n7884 ) | ( ~n3007 & n7885 ) | ( n7884 & n7885 ) ;
  assign n7887 = n2400 & ~n7784 ;
  assign n7888 = n2400 & n7786 ;
  assign n7889 = ( n3007 & n7887 ) | ( n3007 & n7888 ) | ( n7887 & n7888 ) ;
  assign n7890 = n7886 | n7889 ;
  assign n7891 = n2381 & n7784 ;
  assign n7892 = n2381 & ~n7786 ;
  assign n7893 = ( ~n3007 & n7891 ) | ( ~n3007 & n7892 ) | ( n7891 & n7892 ) ;
  assign n7894 = n2492 & ~n7784 ;
  assign n7895 = n2492 & n7786 ;
  assign n7896 = ( n3007 & n7894 ) | ( n3007 & n7895 ) | ( n7894 & n7895 ) ;
  assign n7897 = n7893 | n7896 ;
  assign n7898 = n2928 & n7784 ;
  assign n7899 = n2928 & ~n7786 ;
  assign n7900 = ( ~n3007 & n7898 ) | ( ~n3007 & n7899 ) | ( n7898 & n7899 ) ;
  assign n7901 = n2948 & ~n7784 ;
  assign n7902 = n2948 & n7786 ;
  assign n7903 = ( n3007 & n7901 ) | ( n3007 & n7902 ) | ( n7901 & n7902 ) ;
  assign n7904 = n7900 | n7903 ;
  assign n7905 = n2744 & n7784 ;
  assign n7906 = n2744 & ~n7786 ;
  assign n7907 = ( ~n3007 & n7905 ) | ( ~n3007 & n7906 ) | ( n7905 & n7906 ) ;
  assign n7908 = n2721 & ~n7784 ;
  assign n7909 = n2721 & n7786 ;
  assign n7910 = ( n3007 & n7908 ) | ( n3007 & n7909 ) | ( n7908 & n7909 ) ;
  assign n7911 = n7907 | n7910 ;
  assign n7912 = n2702 & n7784 ;
  assign n7913 = n2702 & ~n7786 ;
  assign n7914 = ( ~n3007 & n7912 ) | ( ~n3007 & n7913 ) | ( n7912 & n7913 ) ;
  assign n7915 = n2679 & ~n7784 ;
  assign n7916 = n2679 & n7786 ;
  assign n7917 = ( n3007 & n7915 ) | ( n3007 & n7916 ) | ( n7915 & n7916 ) ;
  assign n7918 = n7914 | n7917 ;
  assign n7919 = n2658 & n7784 ;
  assign n7920 = n2658 & ~n7786 ;
  assign n7921 = ( ~n3007 & n7919 ) | ( ~n3007 & n7920 ) | ( n7919 & n7920 ) ;
  assign n7922 = n2635 & ~n7784 ;
  assign n7923 = n2635 & n7786 ;
  assign n7924 = ( n3007 & n7922 ) | ( n3007 & n7923 ) | ( n7922 & n7923 ) ;
  assign n7925 = n7921 | n7924 ;
  assign n7926 = n2615 & n7784 ;
  assign n7927 = n2615 & ~n7786 ;
  assign n7928 = ( ~n3007 & n7926 ) | ( ~n3007 & n7927 ) | ( n7926 & n7927 ) ;
  assign n7929 = n2592 & ~n7784 ;
  assign n7930 = n2592 & n7786 ;
  assign n7931 = ( n3007 & n7929 ) | ( n3007 & n7930 ) | ( n7929 & n7930 ) ;
  assign n7932 = n7928 | n7931 ;
  assign n7933 = n2857 & n7784 ;
  assign n7934 = n2857 & ~n7786 ;
  assign n7935 = ( ~n3007 & n7933 ) | ( ~n3007 & n7934 ) | ( n7933 & n7934 ) ;
  assign n7936 = n2834 & ~n7784 ;
  assign n7937 = n2834 & n7786 ;
  assign n7938 = ( n3007 & n7936 ) | ( n3007 & n7937 ) | ( n7936 & n7937 ) ;
  assign n7939 = n7935 | n7938 ;
  assign n7940 = n2814 & n7784 ;
  assign n7941 = n2814 & ~n7786 ;
  assign n7942 = ( ~n3007 & n7940 ) | ( ~n3007 & n7941 ) | ( n7940 & n7941 ) ;
  assign n7943 = n2791 & ~n7784 ;
  assign n7944 = n2791 & n7786 ;
  assign n7945 = ( n3007 & n7943 ) | ( n3007 & n7944 ) | ( n7943 & n7944 ) ;
  assign n7946 = n7942 | n7945 ;
  assign n7947 = n2772 & n7784 ;
  assign n7948 = n2772 & ~n7786 ;
  assign n7949 = ( ~n3007 & n7947 ) | ( ~n3007 & n7948 ) | ( n7947 & n7948 ) ;
  assign n7950 = n2883 & ~n7784 ;
  assign n7951 = n2883 & n7786 ;
  assign n7952 = ( n3007 & n7950 ) | ( n3007 & n7951 ) | ( n7950 & n7951 ) ;
  assign n7953 = n7949 | n7952 ;
  assign n7954 = n3006 & n7784 ;
  assign n7955 = n3006 & ~n7786 ;
  assign n7956 = ( ~n3007 & n7954 ) | ( ~n3007 & n7955 ) | ( n7954 & n7955 ) ;
  assign n7957 = n2983 & ~n7784 ;
  assign n7958 = n2983 & n7786 ;
  assign n7959 = ( n3007 & n7957 ) | ( n3007 & n7958 ) | ( n7957 & n7958 ) ;
  assign n7960 = n7956 | n7959 ;
  assign n7961 = n7699 & n7784 ;
  assign n7962 = n7699 & ~n7786 ;
  assign n7963 = ( ~n3007 & n7961 ) | ( ~n3007 & n7962 ) | ( n7961 & n7962 ) ;
  assign n7964 = n7676 & ~n7784 ;
  assign n7965 = n7676 & n7786 ;
  assign n7966 = ( n3007 & n7964 ) | ( n3007 & n7965 ) | ( n7964 & n7965 ) ;
  assign n7967 = n7963 | n7966 ;
  assign n7968 = n7657 & n7784 ;
  assign n7969 = n7657 & ~n7786 ;
  assign n7970 = ( ~n3007 & n7968 ) | ( ~n3007 & n7969 ) | ( n7968 & n7969 ) ;
  assign n7971 = n7634 & ~n7784 ;
  assign n7972 = n7634 & n7786 ;
  assign n7973 = ( n3007 & n7971 ) | ( n3007 & n7972 ) | ( n7971 & n7972 ) ;
  assign n7974 = n7970 | n7973 ;
  assign n7975 = n7613 & n7784 ;
  assign n7976 = n7613 & ~n7786 ;
  assign n7977 = ( ~n3007 & n7975 ) | ( ~n3007 & n7976 ) | ( n7975 & n7976 ) ;
  assign n7978 = n7590 & ~n7784 ;
  assign n7979 = n7590 & n7786 ;
  assign n7980 = ( n3007 & n7978 ) | ( n3007 & n7979 ) | ( n7978 & n7979 ) ;
  assign n7981 = n7977 | n7980 ;
  assign n7982 = n7570 & n7784 ;
  assign n7983 = n7570 & ~n7786 ;
  assign n7984 = ( ~n3007 & n7982 ) | ( ~n3007 & n7983 ) | ( n7982 & n7983 ) ;
  assign n7985 = n7547 & ~n7784 ;
  assign n7986 = n7547 & n7786 ;
  assign n7987 = ( n3007 & n7985 ) | ( n3007 & n7986 ) | ( n7985 & n7986 ) ;
  assign n7988 = n7984 | n7987 ;
  assign n7989 = n7524 & n7784 ;
  assign n7990 = n7524 & ~n7786 ;
  assign n7991 = ( ~n3007 & n7989 ) | ( ~n3007 & n7990 ) | ( n7989 & n7990 ) ;
  assign n7992 = n7501 & ~n7784 ;
  assign n7993 = n7501 & n7786 ;
  assign n7994 = ( n3007 & n7992 ) | ( n3007 & n7993 ) | ( n7992 & n7993 ) ;
  assign n7995 = n7991 | n7994 ;
  assign n7996 = n7480 & n7784 ;
  assign n7997 = n7480 & ~n7786 ;
  assign n7998 = ( ~n3007 & n7996 ) | ( ~n3007 & n7997 ) | ( n7996 & n7997 ) ;
  assign n7999 = n7457 & ~n7784 ;
  assign n8000 = n7457 & n7786 ;
  assign n8001 = ( n3007 & n7999 ) | ( n3007 & n8000 ) | ( n7999 & n8000 ) ;
  assign n8002 = n7998 | n8001 ;
  assign n8003 = n7110 & n7784 ;
  assign n8004 = n7110 & ~n7786 ;
  assign n8005 = ( ~n3007 & n8003 ) | ( ~n3007 & n8004 ) | ( n8003 & n8004 ) ;
  assign n8006 = n7129 & ~n7784 ;
  assign n8007 = n7129 & n7786 ;
  assign n8008 = ( n3007 & n8006 ) | ( n3007 & n8007 ) | ( n8006 & n8007 ) ;
  assign n8009 = n8005 | n8008 ;
  assign n8010 = n7347 & n7784 ;
  assign n8011 = n7347 & ~n7786 ;
  assign n8012 = ( ~n3007 & n8010 ) | ( ~n3007 & n8011 ) | ( n8010 & n8011 ) ;
  assign n8013 = n7324 & ~n7784 ;
  assign n8014 = n7324 & n7786 ;
  assign n8015 = ( n3007 & n8013 ) | ( n3007 & n8014 ) | ( n8013 & n8014 ) ;
  assign n8016 = n8012 | n8015 ;
  assign n8017 = n7414 & n7784 ;
  assign n8018 = n7414 & ~n7786 ;
  assign n8019 = ( ~n3007 & n8017 ) | ( ~n3007 & n8018 ) | ( n8017 & n8018 ) ;
  assign n8020 = n7433 & ~n7784 ;
  assign n8021 = n7433 & n7786 ;
  assign n8022 = ( n3007 & n8020 ) | ( n3007 & n8021 ) | ( n8020 & n8021 ) ;
  assign n8023 = n8019 | n8022 ;
  assign n8024 = n7390 & n7784 ;
  assign n8025 = n7390 & ~n7786 ;
  assign n8026 = ( ~n3007 & n8024 ) | ( ~n3007 & n8025 ) | ( n8024 & n8025 ) ;
  assign n8027 = n7367 & ~n7784 ;
  assign n8028 = n7367 & n7786 ;
  assign n8029 = ( n3007 & n8027 ) | ( n3007 & n8028 ) | ( n8027 & n8028 ) ;
  assign n8030 = n8026 | n8029 ;
  assign n8031 = n7259 & n7784 ;
  assign n8032 = n7259 & ~n7786 ;
  assign n8033 = ( ~n3007 & n8031 ) | ( ~n3007 & n8032 ) | ( n8031 & n8032 ) ;
  assign n8034 = n7236 & ~n7784 ;
  assign n8035 = n7236 & n7786 ;
  assign n8036 = ( n3007 & n8034 ) | ( n3007 & n8035 ) | ( n8034 & n8035 ) ;
  assign n8037 = n8033 | n8036 ;
  assign n8038 = n7302 & n7784 ;
  assign n8039 = n7302 & ~n7786 ;
  assign n8040 = ( ~n3007 & n8038 ) | ( ~n3007 & n8039 ) | ( n8038 & n8039 ) ;
  assign n8041 = n7279 & ~n7784 ;
  assign n8042 = n7279 & n7786 ;
  assign n8043 = ( n3007 & n8041 ) | ( n3007 & n8042 ) | ( n8041 & n8042 ) ;
  assign n8044 = n8040 | n8043 ;
  assign n8045 = n7196 & n7784 ;
  assign n8046 = n7196 & ~n7786 ;
  assign n8047 = ( ~n3007 & n8045 ) | ( ~n3007 & n8046 ) | ( n8045 & n8046 ) ;
  assign n8048 = n7215 & ~n7784 ;
  assign n8049 = n7215 & n7786 ;
  assign n8050 = ( n3007 & n8048 ) | ( n3007 & n8049 ) | ( n8048 & n8049 ) ;
  assign n8051 = n8047 | n8050 ;
  assign n8052 = n7172 & n7784 ;
  assign n8053 = n7172 & ~n7786 ;
  assign n8054 = ( ~n3007 & n8052 ) | ( ~n3007 & n8053 ) | ( n8052 & n8053 ) ;
  assign n8055 = n7149 & ~n7784 ;
  assign n8056 = n7149 & n7786 ;
  assign n8057 = ( n3007 & n8055 ) | ( n3007 & n8056 ) | ( n8055 & n8056 ) ;
  assign n8058 = n8054 | n8057 ;
  assign n8059 = n7083 & n7784 ;
  assign n8060 = n7083 & ~n7786 ;
  assign n8061 = ( ~n3007 & n8059 ) | ( ~n3007 & n8060 ) | ( n8059 & n8060 ) ;
  assign n8062 = n7060 & ~n7784 ;
  assign n8063 = n7060 & n7786 ;
  assign n8064 = ( n3007 & n8062 ) | ( n3007 & n8063 ) | ( n8062 & n8063 ) ;
  assign n8065 = n8061 | n8064 ;
  assign n8066 = n7040 & n7784 ;
  assign n8067 = n7040 & ~n7786 ;
  assign n8068 = ( ~n3007 & n8066 ) | ( ~n3007 & n8067 ) | ( n8066 & n8067 ) ;
  assign n8069 = n7017 & ~n7784 ;
  assign n8070 = n7017 & n7786 ;
  assign n8071 = ( n3007 & n8069 ) | ( n3007 & n8070 ) | ( n8069 & n8070 ) ;
  assign n8072 = n8068 | n8071 ;
  assign n8073 = n6953 & n7784 ;
  assign n8074 = n6953 & ~n7786 ;
  assign n8075 = ( ~n3007 & n8073 ) | ( ~n3007 & n8074 ) | ( n8073 & n8074 ) ;
  assign n8076 = n6930 & ~n7784 ;
  assign n8077 = n6930 & n7786 ;
  assign n8078 = ( n3007 & n8076 ) | ( n3007 & n8077 ) | ( n8076 & n8077 ) ;
  assign n8079 = n8075 | n8078 ;
  assign n8080 = n6996 & n7784 ;
  assign n8081 = n6996 & ~n7786 ;
  assign n8082 = ( ~n3007 & n8080 ) | ( ~n3007 & n8081 ) | ( n8080 & n8081 ) ;
  assign n8083 = n6973 & ~n7784 ;
  assign n8084 = n6973 & n7786 ;
  assign n8085 = ( n3007 & n8083 ) | ( n3007 & n8084 ) | ( n8083 & n8084 ) ;
  assign n8086 = n8082 | n8085 ;
  assign n8087 = n6865 & n7784 ;
  assign n8088 = n6865 & ~n7786 ;
  assign n8089 = ( ~n3007 & n8087 ) | ( ~n3007 & n8088 ) | ( n8087 & n8088 ) ;
  assign n8090 = n6842 & ~n7784 ;
  assign n8091 = n6842 & n7786 ;
  assign n8092 = ( n3007 & n8090 ) | ( n3007 & n8091 ) | ( n8090 & n8091 ) ;
  assign n8093 = n8089 | n8092 ;
  assign n8094 = n6908 & n7784 ;
  assign n8095 = n6908 & ~n7786 ;
  assign n8096 = ( ~n3007 & n8094 ) | ( ~n3007 & n8095 ) | ( n8094 & n8095 ) ;
  assign n8097 = n6885 & ~n7784 ;
  assign n8098 = n6885 & n7786 ;
  assign n8099 = ( n3007 & n8097 ) | ( n3007 & n8098 ) | ( n8097 & n8098 ) ;
  assign n8100 = n8096 | n8099 ;
  assign n8101 = n6802 & n7784 ;
  assign n8102 = n6802 & ~n7786 ;
  assign n8103 = ( ~n3007 & n8101 ) | ( ~n3007 & n8102 ) | ( n8101 & n8102 ) ;
  assign n8104 = n6821 & ~n7784 ;
  assign n8105 = n6821 & n7786 ;
  assign n8106 = ( n3007 & n8104 ) | ( n3007 & n8105 ) | ( n8104 & n8105 ) ;
  assign n8107 = n8103 | n8106 ;
  assign n8108 = n6778 & n7784 ;
  assign n8109 = n6778 & ~n7786 ;
  assign n8110 = ( ~n3007 & n8108 ) | ( ~n3007 & n8109 ) | ( n8108 & n8109 ) ;
  assign n8111 = n6755 & ~n7784 ;
  assign n8112 = n6755 & n7786 ;
  assign n8113 = ( n3007 & n8111 ) | ( n3007 & n8112 ) | ( n8111 & n8112 ) ;
  assign n8114 = n8110 | n8113 ;
  assign n8115 = n6698 & n7784 ;
  assign n8116 = n6698 & ~n7786 ;
  assign n8117 = ( ~n3007 & n8115 ) | ( ~n3007 & n8116 ) | ( n8115 & n8116 ) ;
  assign n8118 = n6717 & ~n7784 ;
  assign n8119 = n6717 & n7786 ;
  assign n8120 = ( n3007 & n8118 ) | ( n3007 & n8119 ) | ( n8118 & n8119 ) ;
  assign n8121 = n8117 | n8120 ;
  assign n8122 = n6584 & n7784 ;
  assign n8123 = n6584 & ~n7786 ;
  assign n8124 = ( ~n3007 & n8122 ) | ( ~n3007 & n8123 ) | ( n8122 & n8123 ) ;
  assign n8125 = n6561 & ~n7784 ;
  assign n8126 = n6561 & n7786 ;
  assign n8127 = ( n3007 & n8125 ) | ( n3007 & n8126 ) | ( n8125 & n8126 ) ;
  assign n8128 = n8124 | n8127 ;
  assign n8129 = n6651 & n7784 ;
  assign n8130 = n6651 & ~n7786 ;
  assign n8131 = ( ~n3007 & n8129 ) | ( ~n3007 & n8130 ) | ( n8129 & n8130 ) ;
  assign n8132 = n6670 & ~n7784 ;
  assign n8133 = n6670 & n7786 ;
  assign n8134 = ( n3007 & n8132 ) | ( n3007 & n8133 ) | ( n8132 & n8133 ) ;
  assign n8135 = n8131 | n8134 ;
  assign n8136 = n6627 & n7784 ;
  assign n8137 = n6627 & ~n7786 ;
  assign n8138 = ( ~n3007 & n8136 ) | ( ~n3007 & n8137 ) | ( n8136 & n8137 ) ;
  assign n8139 = n6604 & ~n7784 ;
  assign n8140 = n6604 & n7786 ;
  assign n8141 = ( n3007 & n8139 ) | ( n3007 & n8140 ) | ( n8139 & n8140 ) ;
  assign n8142 = n8138 | n8141 ;
  assign n8143 = n6520 & n7784 ;
  assign n8144 = n6520 & ~n7786 ;
  assign n8145 = ( ~n3007 & n8143 ) | ( ~n3007 & n8144 ) | ( n8143 & n8144 ) ;
  assign n8146 = n6539 & ~n7784 ;
  assign n8147 = n6539 & n7786 ;
  assign n8148 = ( n3007 & n8146 ) | ( n3007 & n8147 ) | ( n8146 & n8147 ) ;
  assign n8149 = n8145 | n8148 ;
  assign n8150 = n6496 & n7784 ;
  assign n8151 = n6496 & ~n7786 ;
  assign n8152 = ( ~n3007 & n8150 ) | ( ~n3007 & n8151 ) | ( n8150 & n8151 ) ;
  assign n8153 = n6473 & ~n7784 ;
  assign n8154 = n6473 & n7786 ;
  assign n8155 = ( n3007 & n8153 ) | ( n3007 & n8154 ) | ( n8153 & n8154 ) ;
  assign n8156 = n8152 | n8155 ;
  assign n8157 = n6433 & n7784 ;
  assign n8158 = n6433 & ~n7786 ;
  assign n8159 = ( ~n3007 & n8157 ) | ( ~n3007 & n8158 ) | ( n8157 & n8158 ) ;
  assign n8160 = n6452 & ~n7784 ;
  assign n8161 = n6452 & n7786 ;
  assign n8162 = ( n3007 & n8160 ) | ( n3007 & n8161 ) | ( n8160 & n8161 ) ;
  assign n8163 = n8159 | n8162 ;
  assign n8164 = n6409 & n7784 ;
  assign n8165 = n6409 & ~n7786 ;
  assign n8166 = ( ~n3007 & n8164 ) | ( ~n3007 & n8165 ) | ( n8164 & n8165 ) ;
  assign n8167 = n6386 & ~n7784 ;
  assign n8168 = n6386 & n7786 ;
  assign n8169 = ( n3007 & n8167 ) | ( n3007 & n8168 ) | ( n8167 & n8168 ) ;
  assign n8170 = n8166 | n8169 ;
  assign n8171 = n5585 & n7784 ;
  assign n8172 = n5585 & ~n7786 ;
  assign n8173 = ( ~n3007 & n8171 ) | ( ~n3007 & n8172 ) | ( n8171 & n8172 ) ;
  assign n8174 = n5562 & ~n7784 ;
  assign n8175 = n5562 & n7786 ;
  assign n8176 = ( n3007 & n8174 ) | ( n3007 & n8175 ) | ( n8174 & n8175 ) ;
  assign n8177 = n8173 | n8176 ;
  assign n8178 = n5542 & n7784 ;
  assign n8179 = n5542 & ~n7786 ;
  assign n8180 = ( ~n3007 & n8178 ) | ( ~n3007 & n8179 ) | ( n8178 & n8179 ) ;
  assign n8181 = n5519 & ~n7784 ;
  assign n8182 = n5519 & n7786 ;
  assign n8183 = ( n3007 & n8181 ) | ( n3007 & n8182 ) | ( n8181 & n8182 ) ;
  assign n8184 = n8180 | n8183 ;
  assign n8185 = n5498 & n7784 ;
  assign n8186 = n5498 & ~n7786 ;
  assign n8187 = ( ~n3007 & n8185 ) | ( ~n3007 & n8186 ) | ( n8185 & n8186 ) ;
  assign n8188 = n5475 & ~n7784 ;
  assign n8189 = n5475 & n7786 ;
  assign n8190 = ( n3007 & n8188 ) | ( n3007 & n8189 ) | ( n8188 & n8189 ) ;
  assign n8191 = n8187 | n8190 ;
  assign n8192 = n5455 & n7784 ;
  assign n8193 = n5455 & ~n7786 ;
  assign n8194 = ( ~n3007 & n8192 ) | ( ~n3007 & n8193 ) | ( n8192 & n8193 ) ;
  assign n8195 = n5432 & ~n7784 ;
  assign n8196 = n5432 & n7786 ;
  assign n8197 = ( n3007 & n8195 ) | ( n3007 & n8196 ) | ( n8195 & n8196 ) ;
  assign n8198 = n8194 | n8197 ;
  assign n8199 = n5410 & n7784 ;
  assign n8200 = n5410 & ~n7786 ;
  assign n8201 = ( ~n3007 & n8199 ) | ( ~n3007 & n8200 ) | ( n8199 & n8200 ) ;
  assign n8202 = n5387 & ~n7784 ;
  assign n8203 = n5387 & n7786 ;
  assign n8204 = ( n3007 & n8202 ) | ( n3007 & n8203 ) | ( n8202 & n8203 ) ;
  assign n8205 = n8201 | n8204 ;
  assign n8206 = n5367 & n7784 ;
  assign n8207 = n5367 & ~n7786 ;
  assign n8208 = ( ~n3007 & n8206 ) | ( ~n3007 & n8207 ) | ( n8206 & n8207 ) ;
  assign n8209 = n5344 & ~n7784 ;
  assign n8210 = n5344 & n7786 ;
  assign n8211 = ( n3007 & n8209 ) | ( n3007 & n8210 ) | ( n8209 & n8210 ) ;
  assign n8212 = n8208 | n8211 ;
  assign n8213 = n5304 & n7784 ;
  assign n8214 = n5304 & ~n7786 ;
  assign n8215 = ( ~n3007 & n8213 ) | ( ~n3007 & n8214 ) | ( n8213 & n8214 ) ;
  assign n8216 = n5323 & ~n7784 ;
  assign n8217 = n5323 & n7786 ;
  assign n8218 = ( n3007 & n8216 ) | ( n3007 & n8217 ) | ( n8216 & n8217 ) ;
  assign n8219 = n8215 | n8218 ;
  assign n8220 = n5280 & n7784 ;
  assign n8221 = n5280 & ~n7786 ;
  assign n8222 = ( ~n3007 & n8220 ) | ( ~n3007 & n8221 ) | ( n8220 & n8221 ) ;
  assign n8223 = n5257 & ~n7784 ;
  assign n8224 = n5257 & n7786 ;
  assign n8225 = ( n3007 & n8223 ) | ( n3007 & n8224 ) | ( n8223 & n8224 ) ;
  assign n8226 = n8222 | n8225 ;
  assign n8227 = n5936 & n7784 ;
  assign n8228 = n5936 & ~n7786 ;
  assign n8229 = ( ~n3007 & n8227 ) | ( ~n3007 & n8228 ) | ( n8227 & n8228 ) ;
  assign n8230 = n5955 & ~n7784 ;
  assign n8231 = n5955 & n7786 ;
  assign n8232 = ( n3007 & n8230 ) | ( n3007 & n8231 ) | ( n8230 & n8231 ) ;
  assign n8233 = n8229 | n8232 ;
  assign n8234 = n5912 & n7784 ;
  assign n8235 = n5912 & ~n7786 ;
  assign n8236 = ( ~n3007 & n8234 ) | ( ~n3007 & n8235 ) | ( n8234 & n8235 ) ;
  assign n8237 = n5889 & ~n7784 ;
  assign n8238 = n5889 & n7786 ;
  assign n8239 = ( n3007 & n8237 ) | ( n3007 & n8238 ) | ( n8237 & n8238 ) ;
  assign n8240 = n8236 | n8239 ;
  assign n8241 = n5849 & n7784 ;
  assign n8242 = n5849 & ~n7786 ;
  assign n8243 = ( ~n3007 & n8241 ) | ( ~n3007 & n8242 ) | ( n8241 & n8242 ) ;
  assign n8244 = n5868 & ~n7784 ;
  assign n8245 = n5868 & n7786 ;
  assign n8246 = ( n3007 & n8244 ) | ( n3007 & n8245 ) | ( n8244 & n8245 ) ;
  assign n8247 = n8243 | n8246 ;
  assign n8248 = n5825 & n7784 ;
  assign n8249 = n5825 & ~n7786 ;
  assign n8250 = ( ~n3007 & n8248 ) | ( ~n3007 & n8249 ) | ( n8248 & n8249 ) ;
  assign n8251 = n5802 & ~n7784 ;
  assign n8252 = n5802 & n7786 ;
  assign n8253 = ( n3007 & n8251 ) | ( n3007 & n8252 ) | ( n8251 & n8252 ) ;
  assign n8254 = n8250 | n8253 ;
  assign n8255 = n5780 & n7784 ;
  assign n8256 = n5780 & ~n7786 ;
  assign n8257 = ( ~n3007 & n8255 ) | ( ~n3007 & n8256 ) | ( n8255 & n8256 ) ;
  assign n8258 = n5757 & ~n7784 ;
  assign n8259 = n5757 & n7786 ;
  assign n8260 = ( n3007 & n8258 ) | ( n3007 & n8259 ) | ( n8258 & n8259 ) ;
  assign n8261 = n8257 | n8260 ;
  assign n8262 = n5737 & n7784 ;
  assign n8263 = n5737 & ~n7786 ;
  assign n8264 = ( ~n3007 & n8262 ) | ( ~n3007 & n8263 ) | ( n8262 & n8263 ) ;
  assign n8265 = n5714 & ~n7784 ;
  assign n8266 = n5714 & n7786 ;
  assign n8267 = ( n3007 & n8265 ) | ( n3007 & n8266 ) | ( n8265 & n8266 ) ;
  assign n8268 = n8264 | n8267 ;
  assign n8269 = n5672 & n7784 ;
  assign n8270 = n5672 & ~n7786 ;
  assign n8271 = ( ~n3007 & n8269 ) | ( ~n3007 & n8270 ) | ( n8269 & n8270 ) ;
  assign n8272 = n5691 & ~n7784 ;
  assign n8273 = n5691 & n7786 ;
  assign n8274 = ( n3007 & n8272 ) | ( n3007 & n8273 ) | ( n8272 & n8273 ) ;
  assign n8275 = n8271 | n8274 ;
  assign n8276 = n5648 & n7784 ;
  assign n8277 = n5648 & ~n7786 ;
  assign n8278 = ( ~n3007 & n8276 ) | ( ~n3007 & n8277 ) | ( n8276 & n8277 ) ;
  assign n8279 = n5625 & ~n7784 ;
  assign n8280 = n5625 & n7786 ;
  assign n8281 = ( n3007 & n8279 ) | ( n3007 & n8280 ) | ( n8279 & n8280 ) ;
  assign n8282 = n8278 | n8281 ;
  assign n8283 = n6295 & n7784 ;
  assign n8284 = n6295 & ~n7786 ;
  assign n8285 = ( ~n3007 & n8283 ) | ( ~n3007 & n8284 ) | ( n8283 & n8284 ) ;
  assign n8286 = n6314 & ~n7784 ;
  assign n8287 = n6314 & n7786 ;
  assign n8288 = ( n3007 & n8286 ) | ( n3007 & n8287 ) | ( n8286 & n8287 ) ;
  assign n8289 = n8285 | n8288 ;
  assign n8290 = n6271 & n7784 ;
  assign n8291 = n6271 & ~n7786 ;
  assign n8292 = ( ~n3007 & n8290 ) | ( ~n3007 & n8291 ) | ( n8290 & n8291 ) ;
  assign n8293 = n6248 & ~n7784 ;
  assign n8294 = n6248 & n7786 ;
  assign n8295 = ( n3007 & n8293 ) | ( n3007 & n8294 ) | ( n8293 & n8294 ) ;
  assign n8296 = n8292 | n8295 ;
  assign n8297 = n6208 & n7784 ;
  assign n8298 = n6208 & ~n7786 ;
  assign n8299 = ( ~n3007 & n8297 ) | ( ~n3007 & n8298 ) | ( n8297 & n8298 ) ;
  assign n8300 = n6227 & ~n7784 ;
  assign n8301 = n6227 & n7786 ;
  assign n8302 = ( n3007 & n8300 ) | ( n3007 & n8301 ) | ( n8300 & n8301 ) ;
  assign n8303 = n8299 | n8302 ;
  assign n8304 = n6184 & n7784 ;
  assign n8305 = n6184 & ~n7786 ;
  assign n8306 = ( ~n3007 & n8304 ) | ( ~n3007 & n8305 ) | ( n8304 & n8305 ) ;
  assign n8307 = n6161 & ~n7784 ;
  assign n8308 = n6161 & n7786 ;
  assign n8309 = ( n3007 & n8307 ) | ( n3007 & n8308 ) | ( n8307 & n8308 ) ;
  assign n8310 = n8306 | n8309 ;
  assign n8311 = n6139 & n7784 ;
  assign n8312 = n6139 & ~n7786 ;
  assign n8313 = ( ~n3007 & n8311 ) | ( ~n3007 & n8312 ) | ( n8311 & n8312 ) ;
  assign n8314 = n6116 & ~n7784 ;
  assign n8315 = n6116 & n7786 ;
  assign n8316 = ( n3007 & n8314 ) | ( n3007 & n8315 ) | ( n8314 & n8315 ) ;
  assign n8317 = n8313 | n8316 ;
  assign n8318 = n6096 & n7784 ;
  assign n8319 = n6096 & ~n7786 ;
  assign n8320 = ( ~n3007 & n8318 ) | ( ~n3007 & n8319 ) | ( n8318 & n8319 ) ;
  assign n8321 = n6073 & ~n7784 ;
  assign n8322 = n6073 & n7786 ;
  assign n8323 = ( n3007 & n8321 ) | ( n3007 & n8322 ) | ( n8321 & n8322 ) ;
  assign n8324 = n8320 | n8323 ;
  assign n8325 = n6033 & n7784 ;
  assign n8326 = n6033 & ~n7786 ;
  assign n8327 = ( ~n3007 & n8325 ) | ( ~n3007 & n8326 ) | ( n8325 & n8326 ) ;
  assign n8328 = n6052 & ~n7784 ;
  assign n8329 = n6052 & n7786 ;
  assign n8330 = ( n3007 & n8328 ) | ( n3007 & n8329 ) | ( n8328 & n8329 ) ;
  assign n8331 = n8327 | n8330 ;
  assign n8332 = n6009 & n7784 ;
  assign n8333 = n6009 & ~n7786 ;
  assign n8334 = ( ~n3007 & n8332 ) | ( ~n3007 & n8333 ) | ( n8332 & n8333 ) ;
  assign n8335 = n5986 & ~n7784 ;
  assign n8336 = n5986 & n7786 ;
  assign n8337 = ( n3007 & n8335 ) | ( n3007 & n8336 ) | ( n8335 & n8336 ) ;
  assign n8338 = n8334 | n8337 ;
  assign n8339 = n4444 & n7784 ;
  assign n8340 = n4444 & ~n7786 ;
  assign n8341 = ( ~n3007 & n8339 ) | ( ~n3007 & n8340 ) | ( n8339 & n8340 ) ;
  assign n8342 = n4463 & ~n7784 ;
  assign n8343 = n4463 & n7786 ;
  assign n8344 = ( n3007 & n8342 ) | ( n3007 & n8343 ) | ( n8342 & n8343 ) ;
  assign n8345 = n8341 | n8344 ;
  assign n8346 = n4508 & n7784 ;
  assign n8347 = n4508 & ~n7786 ;
  assign n8348 = ( ~n3007 & n8346 ) | ( ~n3007 & n8347 ) | ( n8346 & n8347 ) ;
  assign n8349 = n4485 & ~n7784 ;
  assign n8350 = n4485 & n7786 ;
  assign n8351 = ( n3007 & n8349 ) | ( n3007 & n8350 ) | ( n8349 & n8350 ) ;
  assign n8352 = n8348 | n8351 ;
  assign n8353 = n4400 & n7784 ;
  assign n8354 = n4400 & ~n7786 ;
  assign n8355 = ( ~n3007 & n8353 ) | ( ~n3007 & n8354 ) | ( n8353 & n8354 ) ;
  assign n8356 = n4419 & ~n7784 ;
  assign n8357 = n4419 & n7786 ;
  assign n8358 = ( n3007 & n8356 ) | ( n3007 & n8357 ) | ( n8356 & n8357 ) ;
  assign n8359 = n8355 | n8358 ;
  assign n8360 = n4376 & n7784 ;
  assign n8361 = n4376 & ~n7786 ;
  assign n8362 = ( ~n3007 & n8360 ) | ( ~n3007 & n8361 ) | ( n8360 & n8361 ) ;
  assign n8363 = n4353 & ~n7784 ;
  assign n8364 = n4353 & n7786 ;
  assign n8365 = ( n3007 & n8363 ) | ( n3007 & n8364 ) | ( n8363 & n8364 ) ;
  assign n8366 = n8362 | n8365 ;
  assign n8367 = n4331 & n7784 ;
  assign n8368 = n4331 & ~n7786 ;
  assign n8369 = ( ~n3007 & n8367 ) | ( ~n3007 & n8368 ) | ( n8367 & n8368 ) ;
  assign n8370 = n4308 & ~n7784 ;
  assign n8371 = n4308 & n7786 ;
  assign n8372 = ( n3007 & n8370 ) | ( n3007 & n8371 ) | ( n8370 & n8371 ) ;
  assign n8373 = n8369 | n8372 ;
  assign n8374 = n4288 & n7784 ;
  assign n8375 = n4288 & ~n7786 ;
  assign n8376 = ( ~n3007 & n8374 ) | ( ~n3007 & n8375 ) | ( n8374 & n8375 ) ;
  assign n8377 = n4265 & ~n7784 ;
  assign n8378 = n4265 & n7786 ;
  assign n8379 = ( n3007 & n8377 ) | ( n3007 & n8378 ) | ( n8377 & n8378 ) ;
  assign n8380 = n8376 | n8379 ;
  assign n8381 = n4225 & n7784 ;
  assign n8382 = n4225 & ~n7786 ;
  assign n8383 = ( ~n3007 & n8381 ) | ( ~n3007 & n8382 ) | ( n8381 & n8382 ) ;
  assign n8384 = n4244 & ~n7784 ;
  assign n8385 = n4244 & n7786 ;
  assign n8386 = ( n3007 & n8384 ) | ( n3007 & n8385 ) | ( n8384 & n8385 ) ;
  assign n8387 = n8383 | n8386 ;
  assign n8388 = n4201 & n7784 ;
  assign n8389 = n4201 & ~n7786 ;
  assign n8390 = ( ~n3007 & n8388 ) | ( ~n3007 & n8389 ) | ( n8388 & n8389 ) ;
  assign n8391 = n4178 & ~n7784 ;
  assign n8392 = n4178 & n7786 ;
  assign n8393 = ( n3007 & n8391 ) | ( n3007 & n8392 ) | ( n8391 & n8392 ) ;
  assign n8394 = n8390 | n8393 ;
  assign n8395 = n4851 & n7784 ;
  assign n8396 = n4851 & ~n7786 ;
  assign n8397 = ( ~n3007 & n8395 ) | ( ~n3007 & n8396 ) | ( n8395 & n8396 ) ;
  assign n8398 = n4870 & ~n7784 ;
  assign n8399 = n4870 & n7786 ;
  assign n8400 = ( n3007 & n8398 ) | ( n3007 & n8399 ) | ( n8398 & n8399 ) ;
  assign n8401 = n8397 | n8400 ;
  assign n8402 = n4827 & n7784 ;
  assign n8403 = n4827 & ~n7786 ;
  assign n8404 = ( ~n3007 & n8402 ) | ( ~n3007 & n8403 ) | ( n8402 & n8403 ) ;
  assign n8405 = n4804 & ~n7784 ;
  assign n8406 = n4804 & n7786 ;
  assign n8407 = ( n3007 & n8405 ) | ( n3007 & n8406 ) | ( n8405 & n8406 ) ;
  assign n8408 = n8404 | n8407 ;
  assign n8409 = n4764 & n7784 ;
  assign n8410 = n4764 & ~n7786 ;
  assign n8411 = ( ~n3007 & n8409 ) | ( ~n3007 & n8410 ) | ( n8409 & n8410 ) ;
  assign n8412 = n4783 & ~n7784 ;
  assign n8413 = n4783 & n7786 ;
  assign n8414 = ( n3007 & n8412 ) | ( n3007 & n8413 ) | ( n8412 & n8413 ) ;
  assign n8415 = n8411 | n8414 ;
  assign n8416 = n4740 & n7784 ;
  assign n8417 = n4740 & ~n7786 ;
  assign n8418 = ( ~n3007 & n8416 ) | ( ~n3007 & n8417 ) | ( n8416 & n8417 ) ;
  assign n8419 = n4717 & ~n7784 ;
  assign n8420 = n4717 & n7786 ;
  assign n8421 = ( n3007 & n8419 ) | ( n3007 & n8420 ) | ( n8419 & n8420 ) ;
  assign n8422 = n8418 | n8421 ;
  assign n8423 = n4694 & n7784 ;
  assign n8424 = n4694 & ~n7786 ;
  assign n8425 = ( ~n3007 & n8423 ) | ( ~n3007 & n8424 ) | ( n8423 & n8424 ) ;
  assign n8426 = n4671 & ~n7784 ;
  assign n8427 = n4671 & n7786 ;
  assign n8428 = ( n3007 & n8426 ) | ( n3007 & n8427 ) | ( n8426 & n8427 ) ;
  assign n8429 = n8425 | n8428 ;
  assign n8430 = n4651 & n7784 ;
  assign n8431 = n4651 & ~n7786 ;
  assign n8432 = ( ~n3007 & n8430 ) | ( ~n3007 & n8431 ) | ( n8430 & n8431 ) ;
  assign n8433 = n4628 & ~n7784 ;
  assign n8434 = n4628 & n7786 ;
  assign n8435 = ( n3007 & n8433 ) | ( n3007 & n8434 ) | ( n8433 & n8434 ) ;
  assign n8436 = n8432 | n8435 ;
  assign n8437 = n4588 & n7784 ;
  assign n8438 = n4588 & ~n7786 ;
  assign n8439 = ( ~n3007 & n8437 ) | ( ~n3007 & n8438 ) | ( n8437 & n8438 ) ;
  assign n8440 = n4607 & ~n7784 ;
  assign n8441 = n4607 & n7786 ;
  assign n8442 = ( n3007 & n8440 ) | ( n3007 & n8441 ) | ( n8440 & n8441 ) ;
  assign n8443 = n8439 | n8442 ;
  assign n8444 = n4564 & n7784 ;
  assign n8445 = n4564 & ~n7786 ;
  assign n8446 = ( ~n3007 & n8444 ) | ( ~n3007 & n8445 ) | ( n8444 & n8445 ) ;
  assign n8447 = n4541 & ~n7784 ;
  assign n8448 = n4541 & n7786 ;
  assign n8449 = ( n3007 & n8447 ) | ( n3007 & n8448 ) | ( n8447 & n8448 ) ;
  assign n8450 = n8446 | n8449 ;
  assign n8451 = n5174 & n7784 ;
  assign n8452 = n5174 & ~n7786 ;
  assign n8453 = ( ~n3007 & n8451 ) | ( ~n3007 & n8452 ) | ( n8451 & n8452 ) ;
  assign n8454 = n5193 & ~n7784 ;
  assign n8455 = n5193 & n7786 ;
  assign n8456 = ( n3007 & n8454 ) | ( n3007 & n8455 ) | ( n8454 & n8455 ) ;
  assign n8457 = n8453 | n8456 ;
  assign n8458 = n5151 & n7784 ;
  assign n8459 = n5151 & ~n7786 ;
  assign n8460 = ( ~n3007 & n8458 ) | ( ~n3007 & n8459 ) | ( n8458 & n8459 ) ;
  assign n8461 = n5128 & ~n7784 ;
  assign n8462 = n5128 & n7786 ;
  assign n8463 = ( n3007 & n8461 ) | ( n3007 & n8462 ) | ( n8461 & n8462 ) ;
  assign n8464 = n8460 | n8463 ;
  assign n8465 = n5089 & n7784 ;
  assign n8466 = n5089 & ~n7786 ;
  assign n8467 = ( ~n3007 & n8465 ) | ( ~n3007 & n8466 ) | ( n8465 & n8466 ) ;
  assign n8468 = n5108 & ~n7784 ;
  assign n8469 = n5108 & n7786 ;
  assign n8470 = ( n3007 & n8468 ) | ( n3007 & n8469 ) | ( n8468 & n8469 ) ;
  assign n8471 = n8467 | n8470 ;
  assign n8472 = n5066 & n7784 ;
  assign n8473 = n5066 & ~n7786 ;
  assign n8474 = ( ~n3007 & n8472 ) | ( ~n3007 & n8473 ) | ( n8472 & n8473 ) ;
  assign n8475 = n5043 & ~n7784 ;
  assign n8476 = n5043 & n7786 ;
  assign n8477 = ( n3007 & n8475 ) | ( n3007 & n8476 ) | ( n8475 & n8476 ) ;
  assign n8478 = n8474 | n8477 ;
  assign n8479 = n5014 & n7784 ;
  assign n8480 = n5014 & ~n7786 ;
  assign n8481 = ( ~n3007 & n8479 ) | ( ~n3007 & n8480 ) | ( n8479 & n8480 ) ;
  assign n8482 = n4991 & ~n7784 ;
  assign n8483 = n4991 & n7786 ;
  assign n8484 = ( n3007 & n8482 ) | ( n3007 & n8483 ) | ( n8482 & n8483 ) ;
  assign n8485 = n8481 | n8484 ;
  assign n8486 = n4972 & n7784 ;
  assign n8487 = n4972 & ~n7786 ;
  assign n8488 = ( ~n3007 & n8486 ) | ( ~n3007 & n8487 ) | ( n8486 & n8487 ) ;
  assign n8489 = n4949 & ~n7784 ;
  assign n8490 = n4949 & n7786 ;
  assign n8491 = ( n3007 & n8489 ) | ( n3007 & n8490 ) | ( n8489 & n8490 ) ;
  assign n8492 = n8488 | n8491 ;
  assign n8493 = n4909 & n7784 ;
  assign n8494 = n4909 & ~n7786 ;
  assign n8495 = ( ~n3007 & n8493 ) | ( ~n3007 & n8494 ) | ( n8493 & n8494 ) ;
  assign n8496 = n4928 & ~n7784 ;
  assign n8497 = n4928 & n7786 ;
  assign n8498 = ( n3007 & n8496 ) | ( n3007 & n8497 ) | ( n8496 & n8497 ) ;
  assign n8499 = n8495 | n8498 ;
  assign n8500 = n4157 & n7784 ;
  assign n8501 = n4157 & ~n7786 ;
  assign n8502 = ( ~n3007 & n8500 ) | ( ~n3007 & n8501 ) | ( n8500 & n8501 ) ;
  assign n8503 = n4134 & ~n7784 ;
  assign n8504 = n4134 & n7786 ;
  assign n8505 = ( n3007 & n8503 ) | ( n3007 & n8504 ) | ( n8503 & n8504 ) ;
  assign n8506 = n8502 | n8505 ;
  assign n8507 = n3335 & n7784 ;
  assign n8508 = n3335 & ~n7786 ;
  assign n8509 = ( ~n3007 & n8507 ) | ( ~n3007 & n8508 ) | ( n8507 & n8508 ) ;
  assign n8510 = n3354 & ~n7784 ;
  assign n8511 = n3354 & n7786 ;
  assign n8512 = ( n3007 & n8510 ) | ( n3007 & n8511 ) | ( n8510 & n8511 ) ;
  assign n8513 = n8509 | n8512 ;
  assign n8514 = n3312 & n7784 ;
  assign n8515 = n3312 & ~n7786 ;
  assign n8516 = ( ~n3007 & n8514 ) | ( ~n3007 & n8515 ) | ( n8514 & n8515 ) ;
  assign n8517 = n3289 & ~n7784 ;
  assign n8518 = n3289 & n7786 ;
  assign n8519 = ( n3007 & n8517 ) | ( n3007 & n8518 ) | ( n8517 & n8518 ) ;
  assign n8520 = n8516 | n8519 ;
  assign n8521 = n3250 & n7784 ;
  assign n8522 = n3250 & ~n7786 ;
  assign n8523 = ( ~n3007 & n8521 ) | ( ~n3007 & n8522 ) | ( n8521 & n8522 ) ;
  assign n8524 = n3269 & ~n7784 ;
  assign n8525 = n3269 & n7786 ;
  assign n8526 = ( n3007 & n8524 ) | ( n3007 & n8525 ) | ( n8524 & n8525 ) ;
  assign n8527 = n8523 | n8526 ;
  assign n8528 = n3227 & n7784 ;
  assign n8529 = n3227 & ~n7786 ;
  assign n8530 = ( ~n3007 & n8528 ) | ( ~n3007 & n8529 ) | ( n8528 & n8529 ) ;
  assign n8531 = n3204 & ~n7784 ;
  assign n8532 = n3204 & n7786 ;
  assign n8533 = ( n3007 & n8531 ) | ( n3007 & n8532 ) | ( n8531 & n8532 ) ;
  assign n8534 = n8530 | n8533 ;
  assign n8535 = n3181 & n7784 ;
  assign n8536 = n3181 & ~n7786 ;
  assign n8537 = ( ~n3007 & n8535 ) | ( ~n3007 & n8536 ) | ( n8535 & n8536 ) ;
  assign n8538 = n3158 & ~n7784 ;
  assign n8539 = n3158 & n7786 ;
  assign n8540 = ( n3007 & n8538 ) | ( n3007 & n8539 ) | ( n8538 & n8539 ) ;
  assign n8541 = n8537 | n8540 ;
  assign n8542 = n3138 & n7784 ;
  assign n8543 = n3138 & ~n7786 ;
  assign n8544 = ( ~n3007 & n8542 ) | ( ~n3007 & n8543 ) | ( n8542 & n8543 ) ;
  assign n8545 = n3115 & ~n7784 ;
  assign n8546 = n3115 & n7786 ;
  assign n8547 = ( n3007 & n8545 ) | ( n3007 & n8546 ) | ( n8545 & n8546 ) ;
  assign n8548 = n8544 | n8547 ;
  assign n8549 = n3073 & n7784 ;
  assign n8550 = n3073 & ~n7786 ;
  assign n8551 = ( ~n3007 & n8549 ) | ( ~n3007 & n8550 ) | ( n8549 & n8550 ) ;
  assign n8552 = n3092 & ~n7784 ;
  assign n8553 = n3092 & n7786 ;
  assign n8554 = ( n3007 & n8552 ) | ( n3007 & n8553 ) | ( n8552 & n8553 ) ;
  assign n8555 = n8551 | n8554 ;
  assign n8556 = n3049 & n7784 ;
  assign n8557 = n3049 & ~n7786 ;
  assign n8558 = ( ~n3007 & n8556 ) | ( ~n3007 & n8557 ) | ( n8556 & n8557 ) ;
  assign n8559 = n3026 & ~n7784 ;
  assign n8560 = n3026 & n7786 ;
  assign n8561 = ( n3007 & n8559 ) | ( n3007 & n8560 ) | ( n8559 & n8560 ) ;
  assign n8562 = n8558 | n8561 ;
  assign n8563 = n3876 & n7784 ;
  assign n8564 = n3876 & ~n7786 ;
  assign n8565 = ( ~n3007 & n8563 ) | ( ~n3007 & n8564 ) | ( n8563 & n8564 ) ;
  assign n8566 = n3895 & ~n7784 ;
  assign n8567 = n3895 & n7786 ;
  assign n8568 = ( n3007 & n8566 ) | ( n3007 & n8567 ) | ( n8566 & n8567 ) ;
  assign n8569 = n8565 | n8568 ;
  assign n8570 = n3853 & n7784 ;
  assign n8571 = n3853 & ~n7786 ;
  assign n8572 = ( ~n3007 & n8570 ) | ( ~n3007 & n8571 ) | ( n8570 & n8571 ) ;
  assign n8573 = n3830 & ~n7784 ;
  assign n8574 = n3830 & n7786 ;
  assign n8575 = ( n3007 & n8573 ) | ( n3007 & n8574 ) | ( n8573 & n8574 ) ;
  assign n8576 = n8572 | n8575 ;
  assign n8577 = n3791 & n7784 ;
  assign n8578 = n3791 & ~n7786 ;
  assign n8579 = ( ~n3007 & n8577 ) | ( ~n3007 & n8578 ) | ( n8577 & n8578 ) ;
  assign n8580 = n3810 & ~n7784 ;
  assign n8581 = n3810 & n7786 ;
  assign n8582 = ( n3007 & n8580 ) | ( n3007 & n8581 ) | ( n8580 & n8581 ) ;
  assign n8583 = n8579 | n8582 ;
  assign n8584 = n3768 & n7784 ;
  assign n8585 = n3768 & ~n7786 ;
  assign n8586 = ( ~n3007 & n8584 ) | ( ~n3007 & n8585 ) | ( n8584 & n8585 ) ;
  assign n8587 = n3745 & ~n7784 ;
  assign n8588 = n3745 & n7786 ;
  assign n8589 = ( n3007 & n8587 ) | ( n3007 & n8588 ) | ( n8587 & n8588 ) ;
  assign n8590 = n8586 | n8589 ;
  assign n8591 = n3713 & n7784 ;
  assign n8592 = n3713 & ~n7786 ;
  assign n8593 = ( ~n3007 & n8591 ) | ( ~n3007 & n8592 ) | ( n8591 & n8592 ) ;
  assign n8594 = n3690 & ~n7784 ;
  assign n8595 = n3690 & n7786 ;
  assign n8596 = ( n3007 & n8594 ) | ( n3007 & n8595 ) | ( n8594 & n8595 ) ;
  assign n8597 = n8593 | n8596 ;
  assign n8598 = n3671 & n7784 ;
  assign n8599 = n3671 & ~n7786 ;
  assign n8600 = ( ~n3007 & n8598 ) | ( ~n3007 & n8599 ) | ( n8598 & n8599 ) ;
  assign n8601 = n3648 & ~n7784 ;
  assign n8602 = n3648 & n7786 ;
  assign n8603 = ( n3007 & n8601 ) | ( n3007 & n8602 ) | ( n8601 & n8602 ) ;
  assign n8604 = n8600 | n8603 ;
  assign n8605 = n3608 & n7784 ;
  assign n8606 = n3608 & ~n7786 ;
  assign n8607 = ( ~n3007 & n8605 ) | ( ~n3007 & n8606 ) | ( n8605 & n8606 ) ;
  assign n8608 = n3627 & ~n7784 ;
  assign n8609 = n3627 & n7786 ;
  assign n8610 = ( n3007 & n8608 ) | ( n3007 & n8609 ) | ( n8608 & n8609 ) ;
  assign n8611 = n8607 | n8610 ;
  assign n8612 = n3584 & n7784 ;
  assign n8613 = n3584 & ~n7786 ;
  assign n8614 = ( ~n3007 & n8612 ) | ( ~n3007 & n8613 ) | ( n8612 & n8613 ) ;
  assign n8615 = n3561 & ~n7784 ;
  assign n8616 = n3561 & n7786 ;
  assign n8617 = ( n3007 & n8615 ) | ( n3007 & n8616 ) | ( n8615 & n8616 ) ;
  assign n8618 = n8614 | n8617 ;
  assign n8619 = n3520 & n7784 ;
  assign n8620 = n3520 & ~n7786 ;
  assign n8621 = ( ~n3007 & n8619 ) | ( ~n3007 & n8620 ) | ( n8619 & n8620 ) ;
  assign n8622 = n3539 & ~n7784 ;
  assign n8623 = n3539 & n7786 ;
  assign n8624 = ( n3007 & n8622 ) | ( n3007 & n8623 ) | ( n8622 & n8623 ) ;
  assign n8625 = n8621 | n8624 ;
  assign n8626 = n3496 & n7784 ;
  assign n8627 = n3496 & ~n7786 ;
  assign n8628 = ( ~n3007 & n8626 ) | ( ~n3007 & n8627 ) | ( n8626 & n8627 ) ;
  assign n8629 = n3473 & ~n7784 ;
  assign n8630 = n3473 & n7786 ;
  assign n8631 = ( n3007 & n8629 ) | ( n3007 & n8630 ) | ( n8629 & n8630 ) ;
  assign n8632 = n8628 | n8631 ;
  assign n8633 = n3433 & n7784 ;
  assign n8634 = n3433 & ~n7786 ;
  assign n8635 = ( ~n3007 & n8633 ) | ( ~n3007 & n8634 ) | ( n8633 & n8634 ) ;
  assign n8636 = n3452 & ~n7784 ;
  assign n8637 = n3452 & n7786 ;
  assign n8638 = ( n3007 & n8636 ) | ( n3007 & n8637 ) | ( n8636 & n8637 ) ;
  assign n8639 = n8635 | n8638 ;
  assign n8640 = n3409 & n7784 ;
  assign n8641 = n3409 & ~n7786 ;
  assign n8642 = ( ~n3007 & n8640 ) | ( ~n3007 & n8641 ) | ( n8640 & n8641 ) ;
  assign n8643 = n3386 & ~n7784 ;
  assign n8644 = n3386 & n7786 ;
  assign n8645 = ( n3007 & n8643 ) | ( n3007 & n8644 ) | ( n8643 & n8644 ) ;
  assign n8646 = n8642 | n8645 ;
  assign n8647 = n4042 & n7784 ;
  assign n8648 = n4042 & ~n7786 ;
  assign n8649 = ( ~n3007 & n8647 ) | ( ~n3007 & n8648 ) | ( n8647 & n8648 ) ;
  assign n8650 = n4019 & ~n7784 ;
  assign n8651 = n4019 & n7786 ;
  assign n8652 = ( n3007 & n8650 ) | ( n3007 & n8651 ) | ( n8650 & n8651 ) ;
  assign n8653 = n8649 | n8652 ;
  assign n8654 = n3998 & n7784 ;
  assign n8655 = n3998 & ~n7786 ;
  assign n8656 = ( ~n3007 & n8654 ) | ( ~n3007 & n8655 ) | ( n8654 & n8655 ) ;
  assign n8657 = n3975 & ~n7784 ;
  assign n8658 = n3975 & n7786 ;
  assign n8659 = ( n3007 & n8657 ) | ( n3007 & n8658 ) | ( n8657 & n8658 ) ;
  assign n8660 = n8656 | n8659 ;
  assign n8661 = n3955 & n7784 ;
  assign n8662 = n3955 & ~n7786 ;
  assign n8663 = ( ~n3007 & n8661 ) | ( ~n3007 & n8662 ) | ( n8661 & n8662 ) ;
  assign n8664 = n3932 & ~n7784 ;
  assign n8665 = n3932 & n7786 ;
  assign n8666 = ( n3007 & n8664 ) | ( n3007 & n8665 ) | ( n8664 & n8665 ) ;
  assign n8667 = n8663 | n8666 ;
  assign n8668 = ~n4074 & n4089 ;
  assign n8669 = ( ~n4074 & n4086 ) | ( ~n4074 & n8668 ) | ( n4086 & n8668 ) ;
  assign n8670 = n4083 | n8669 ;
  assign n8671 = n4076 & ~n8669 ;
  assign n8672 = ( n3913 & n8670 ) | ( n3913 & ~n8671 ) | ( n8670 & ~n8671 ) ;
  assign n8673 = n4096 & ~n8669 ;
  assign n8674 = ( n4108 & ~n8670 ) | ( n4108 & n8673 ) | ( ~n8670 & n8673 ) ;
  assign n8675 = ( n5222 & ~n8672 ) | ( n5222 & n8674 ) | ( ~n8672 & n8674 ) ;
  assign n8676 = ( n5237 & n8672 ) | ( n5237 & ~n8674 ) | ( n8672 & ~n8674 ) ;
  assign n8677 = ( n7752 & n8675 ) | ( n7752 & ~n8676 ) | ( n8675 & ~n8676 ) ;
  assign n8678 = ~n4073 & n8677 ;
  assign n8679 = ( n7775 & ~n8675 ) | ( n7775 & n8676 ) | ( ~n8675 & n8676 ) ;
  assign n8680 = n4073 | n8679 ;
  assign n8681 = ( n3007 & ~n8678 ) | ( n3007 & n8680 ) | ( ~n8678 & n8680 ) ;
  assign n8682 = n4057 & n8681 ;
  assign n8683 = ( x281 & ~x409 ) | ( x281 & n656 ) | ( ~x409 & n656 ) ;
  assign n8684 = ( n1115 & ~n1119 ) | ( n1115 & n1126 ) | ( ~n1119 & n1126 ) ;
  assign n8685 = ( n991 & ~n995 ) | ( n991 & n8684 ) | ( ~n995 & n8684 ) ;
  assign n8686 = ( ~n991 & n995 ) | ( ~n991 & n1104 ) | ( n995 & n1104 ) ;
  assign n8687 = ( n975 & n8685 ) | ( n975 & ~n8686 ) | ( n8685 & ~n8686 ) ;
  assign n8688 = ( n1154 & ~n8685 ) | ( n1154 & n8686 ) | ( ~n8685 & n8686 ) ;
  assign n8689 = ( n8683 & ~n8687 ) | ( n8683 & n8688 ) | ( ~n8687 & n8688 ) ;
  assign n8690 = n7784 & ~n8689 ;
  assign n8691 = n7786 | n8689 ;
  assign n8692 = ( n3007 & ~n8690 ) | ( n3007 & n8691 ) | ( ~n8690 & n8691 ) ;
  assign n8693 = ( n1783 & ~n1787 ) | ( n1783 & n1794 ) | ( ~n1787 & n1794 ) ;
  assign n8694 = ( n1767 & ~n1771 ) | ( n1767 & n8693 ) | ( ~n1771 & n8693 ) ;
  assign n8695 = ( n1751 & ~n1767 ) | ( n1751 & n1771 ) | ( ~n1767 & n1771 ) ;
  assign n8696 = ( n1643 & n8694 ) | ( n1643 & ~n8695 ) | ( n8694 & ~n8695 ) ;
  assign n8697 = ( n1822 & ~n8694 ) | ( n1822 & n8695 ) | ( ~n8694 & n8695 ) ;
  assign n8698 = ( n1324 & ~n8696 ) | ( n1324 & n8697 ) | ( ~n8696 & n8697 ) ;
  assign n8699 = n7784 | n8698 ;
  assign n8700 = n7786 & ~n8698 ;
  assign n8701 = ( n3007 & ~n8699 ) | ( n3007 & n8700 ) | ( ~n8699 & n8700 ) ;
  assign n8702 = n8692 & ~n8701 ;
  assign n8703 = ( n3007 & ~n7784 ) | ( n3007 & n7786 ) | ( ~n7784 & n7786 ) ;
  assign y0 = n7781 ;
  assign y1 = n7792 ;
  assign y2 = n7799 ;
  assign y3 = n7806 ;
  assign y4 = n7813 ;
  assign y5 = n7820 ;
  assign y6 = n7827 ;
  assign y7 = n7834 ;
  assign y8 = n7841 ;
  assign y9 = n7848 ;
  assign y10 = n7855 ;
  assign y11 = n7862 ;
  assign y12 = n7869 ;
  assign y13 = n7876 ;
  assign y14 = n7883 ;
  assign y15 = n7890 ;
  assign y16 = n7897 ;
  assign y17 = n7904 ;
  assign y18 = n7911 ;
  assign y19 = n7918 ;
  assign y20 = n7925 ;
  assign y21 = n7932 ;
  assign y22 = n7939 ;
  assign y23 = n7946 ;
  assign y24 = n7953 ;
  assign y25 = n7960 ;
  assign y26 = n7967 ;
  assign y27 = n7974 ;
  assign y28 = n7981 ;
  assign y29 = n7988 ;
  assign y30 = n7995 ;
  assign y31 = n8002 ;
  assign y32 = n8009 ;
  assign y33 = n8016 ;
  assign y34 = n8023 ;
  assign y35 = n8030 ;
  assign y36 = n8037 ;
  assign y37 = n8044 ;
  assign y38 = n8051 ;
  assign y39 = n8058 ;
  assign y40 = n8065 ;
  assign y41 = n8072 ;
  assign y42 = n8079 ;
  assign y43 = n8086 ;
  assign y44 = n8093 ;
  assign y45 = n8100 ;
  assign y46 = n8107 ;
  assign y47 = n8114 ;
  assign y48 = n8121 ;
  assign y49 = n8128 ;
  assign y50 = n8135 ;
  assign y51 = n8142 ;
  assign y52 = n8149 ;
  assign y53 = n8156 ;
  assign y54 = n8163 ;
  assign y55 = n8170 ;
  assign y56 = n8177 ;
  assign y57 = n8184 ;
  assign y58 = n8191 ;
  assign y59 = n8198 ;
  assign y60 = n8205 ;
  assign y61 = n8212 ;
  assign y62 = n8219 ;
  assign y63 = n8226 ;
  assign y64 = n8233 ;
  assign y65 = n8240 ;
  assign y66 = n8247 ;
  assign y67 = n8254 ;
  assign y68 = n8261 ;
  assign y69 = n8268 ;
  assign y70 = n8275 ;
  assign y71 = n8282 ;
  assign y72 = n8289 ;
  assign y73 = n8296 ;
  assign y74 = n8303 ;
  assign y75 = n8310 ;
  assign y76 = n8317 ;
  assign y77 = n8324 ;
  assign y78 = n8331 ;
  assign y79 = n8338 ;
  assign y80 = n8345 ;
  assign y81 = n8352 ;
  assign y82 = n8359 ;
  assign y83 = n8366 ;
  assign y84 = n8373 ;
  assign y85 = n8380 ;
  assign y86 = n8387 ;
  assign y87 = n8394 ;
  assign y88 = n8401 ;
  assign y89 = n8408 ;
  assign y90 = n8415 ;
  assign y91 = n8422 ;
  assign y92 = n8429 ;
  assign y93 = n8436 ;
  assign y94 = n8443 ;
  assign y95 = n8450 ;
  assign y96 = n8457 ;
  assign y97 = n8464 ;
  assign y98 = n8471 ;
  assign y99 = n8478 ;
  assign y100 = n8485 ;
  assign y101 = n8492 ;
  assign y102 = n8499 ;
  assign y103 = n8506 ;
  assign y104 = n8513 ;
  assign y105 = n8520 ;
  assign y106 = n8527 ;
  assign y107 = n8534 ;
  assign y108 = n8541 ;
  assign y109 = n8548 ;
  assign y110 = n8555 ;
  assign y111 = n8562 ;
  assign y112 = n8569 ;
  assign y113 = n8576 ;
  assign y114 = n8583 ;
  assign y115 = n8590 ;
  assign y116 = n8597 ;
  assign y117 = n8604 ;
  assign y118 = n8611 ;
  assign y119 = n8618 ;
  assign y120 = n8625 ;
  assign y121 = n8632 ;
  assign y122 = n8639 ;
  assign y123 = n8646 ;
  assign y124 = n8653 ;
  assign y125 = n8660 ;
  assign y126 = n8667 ;
  assign y127 = n8682 ;
  assign y128 = ~n8702 ;
  assign y129 = ~n8703 ;
endmodule
