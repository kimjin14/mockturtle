module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 ;
  output y0 ;
  wire n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 ;
  assign n1478 = ~x0 & x1 ;
  assign n1479 = x0 & ~x1 ;
  assign n1480 = n1478 | n1479 ;
  assign n1481 = ~x2 & n1480 ;
  assign n1482 = x2 & ~n1478 ;
  assign n1483 = ~n1479 & n1482 ;
  assign n1484 = n1481 | n1483 ;
  assign n1485 = ~x6 & n1484 ;
  assign n1486 = x3 & ~x4 ;
  assign n1487 = ~x3 & x4 ;
  assign n1488 = n1486 | n1487 ;
  assign n1489 = ~x5 & n1488 ;
  assign n1490 = x5 & ~n1488 ;
  assign n1491 = n1489 | n1490 ;
  assign n1492 = x6 & n1479 ;
  assign n1493 = ( x6 & ~n1482 ) | ( x6 & n1492 ) | ( ~n1482 & n1492 ) ;
  assign n1494 = ~n1481 & n1493 ;
  assign n1495 = n1491 & ~n1494 ;
  assign n1496 = ~n1485 & n1495 ;
  assign n1497 = ~n1491 & n1494 ;
  assign n1498 = ( n1485 & ~n1491 ) | ( n1485 & n1497 ) | ( ~n1491 & n1497 ) ;
  assign n1499 = n1496 | n1498 ;
  assign n1500 = ~x997 & x998 ;
  assign n1501 = x997 & ~x998 ;
  assign n1502 = n1500 | n1501 ;
  assign n1503 = ~x999 & n1502 ;
  assign n1504 = x999 & ~n1502 ;
  assign n1505 = n1503 | n1504 ;
  assign n1506 = n1499 | n1505 ;
  assign n1507 = n1499 & ~n1505 ;
  assign n1508 = ( ~n1499 & n1506 ) | ( ~n1499 & n1507 ) | ( n1506 & n1507 ) ;
  assign n1509 = ~x991 & x992 ;
  assign n1510 = x991 & ~x992 ;
  assign n1511 = n1509 | n1510 ;
  assign n1512 = ~x993 & n1511 ;
  assign n1513 = x993 & ~n1511 ;
  assign n1514 = n1512 | n1513 ;
  assign n1515 = ~x994 & x995 ;
  assign n1516 = x994 & ~x995 ;
  assign n1517 = n1515 | n1516 ;
  assign n1518 = ~x996 & n1517 ;
  assign n1519 = x996 & ~n1517 ;
  assign n1520 = n1518 | n1519 ;
  assign n1521 = n1514 & ~n1520 ;
  assign n1522 = ~n1514 & n1520 ;
  assign n1523 = n1521 | n1522 ;
  assign n1524 = ( x994 & x995 ) | ( x994 & x996 ) | ( x995 & x996 ) ;
  assign n1525 = ( x991 & x992 ) | ( x991 & x993 ) | ( x992 & x993 ) ;
  assign n1526 = n1524 & ~n1525 ;
  assign n1527 = ~n1524 & n1525 ;
  assign n1528 = n1526 | n1527 ;
  assign n1529 = n1514 & n1520 ;
  assign n1530 = n1528 & ~n1529 ;
  assign n1531 = ~n1528 & n1529 ;
  assign n1532 = n1530 | n1531 ;
  assign n1533 = ( n1524 & n1525 ) | ( n1524 & n1529 ) | ( n1525 & n1529 ) ;
  assign n1534 = n1523 & ~n1533 ;
  assign n1535 = ( n1523 & ~n1532 ) | ( n1523 & n1534 ) | ( ~n1532 & n1534 ) ;
  assign n1536 = n1508 & n1535 ;
  assign n1537 = n1491 & n1494 ;
  assign n1538 = ( n1485 & n1491 ) | ( n1485 & n1537 ) | ( n1491 & n1537 ) ;
  assign n1539 = ( x0 & x1 ) | ( x0 & x2 ) | ( x1 & x2 ) ;
  assign n1540 = ( x3 & x4 ) | ( x3 & x5 ) | ( x4 & x5 ) ;
  assign n1541 = ~n1539 & n1540 ;
  assign n1542 = n1539 & ~n1540 ;
  assign n1543 = n1541 | n1542 ;
  assign n1544 = x6 | n1543 ;
  assign n1545 = ( n1484 & n1543 ) | ( n1484 & n1544 ) | ( n1543 & n1544 ) ;
  assign n1546 = n1538 | n1545 ;
  assign n1547 = x6 & n1543 ;
  assign n1548 = n1484 & n1547 ;
  assign n1549 = ( n1538 & n1543 ) | ( n1538 & n1548 ) | ( n1543 & n1548 ) ;
  assign n1550 = n1546 & ~n1549 ;
  assign n1551 = n1499 & n1505 ;
  assign n1552 = n1550 & n1551 ;
  assign n1553 = n1550 | n1551 ;
  assign n1554 = ( x997 & x998 ) | ( x997 & x999 ) | ( x998 & x999 ) ;
  assign n1555 = n1553 & ~n1554 ;
  assign n1556 = ~n1552 & n1555 ;
  assign n1557 = ~n1552 & n1553 ;
  assign n1558 = n1554 & ~n1557 ;
  assign n1559 = n1556 | n1558 ;
  assign n1560 = n1536 & n1559 ;
  assign n1561 = n1523 & n1533 ;
  assign n1562 = n1532 & ~n1561 ;
  assign n1563 = n1536 | n1558 ;
  assign n1564 = n1556 & n1562 ;
  assign n1565 = ( n1562 & n1563 ) | ( n1562 & n1564 ) | ( n1563 & n1564 ) ;
  assign n1566 = n1560 | n1565 ;
  assign n1567 = n1553 & n1554 ;
  assign n1568 = n1539 & n1540 ;
  assign n1569 = n1548 | n1568 ;
  assign n1570 = n1543 | n1568 ;
  assign n1571 = ( n1538 & n1569 ) | ( n1538 & n1570 ) | ( n1569 & n1570 ) ;
  assign n1572 = ~n1552 & n1571 ;
  assign n1573 = ~n1567 & n1572 ;
  assign n1574 = n1552 & ~n1571 ;
  assign n1575 = ( n1567 & ~n1571 ) | ( n1567 & n1574 ) | ( ~n1571 & n1574 ) ;
  assign n1576 = n1573 | n1575 ;
  assign n1577 = n1566 & n1576 ;
  assign n1578 = ~n1523 & n1533 ;
  assign n1579 = ( ~n1532 & n1533 ) | ( ~n1532 & n1578 ) | ( n1533 & n1578 ) ;
  assign n1580 = n1576 & n1579 ;
  assign n1581 = ( n1566 & n1579 ) | ( n1566 & n1580 ) | ( n1579 & n1580 ) ;
  assign n1582 = n1577 | n1581 ;
  assign n1583 = n1552 & n1571 ;
  assign n1584 = ( n1567 & n1571 ) | ( n1567 & n1583 ) | ( n1571 & n1583 ) ;
  assign n1585 = n1582 & n1584 ;
  assign n1586 = n1580 | n1584 ;
  assign n1587 = n1579 | n1584 ;
  assign n1588 = ( n1566 & n1586 ) | ( n1566 & n1587 ) | ( n1586 & n1587 ) ;
  assign n1589 = n1577 | n1588 ;
  assign n1590 = ~n1585 & n1589 ;
  assign n1591 = ~x19 & x20 ;
  assign n1592 = x19 & ~x20 ;
  assign n1593 = n1591 | n1592 ;
  assign n1594 = ~x21 & n1593 ;
  assign n1595 = x21 & ~n1593 ;
  assign n1596 = n1594 | n1595 ;
  assign n1597 = ~x22 & x23 ;
  assign n1598 = x22 & ~x23 ;
  assign n1599 = n1597 | n1598 ;
  assign n1600 = ~x24 & n1599 ;
  assign n1601 = x24 & ~n1599 ;
  assign n1602 = n1600 | n1601 ;
  assign n1603 = n1596 & n1602 ;
  assign n1604 = ( x22 & x23 ) | ( x22 & x24 ) | ( x23 & x24 ) ;
  assign n1605 = ( x19 & x20 ) | ( x19 & x21 ) | ( x20 & x21 ) ;
  assign n1606 = ~n1604 & n1605 ;
  assign n1607 = n1604 & ~n1605 ;
  assign n1608 = n1606 | n1607 ;
  assign n1609 = ~n1603 & n1608 ;
  assign n1610 = n1603 & ~n1608 ;
  assign n1611 = n1609 | n1610 ;
  assign n1612 = n1596 & ~n1602 ;
  assign n1613 = ~n1596 & n1602 ;
  assign n1614 = n1612 | n1613 ;
  assign n1615 = ( n1603 & n1604 ) | ( n1603 & n1605 ) | ( n1604 & n1605 ) ;
  assign n1616 = n1614 & n1615 ;
  assign n1617 = n1611 & ~n1616 ;
  assign n1618 = ( x28 & x29 ) | ( x28 & x30 ) | ( x29 & x30 ) ;
  assign n1619 = ( x25 & x26 ) | ( x25 & x27 ) | ( x26 & x27 ) ;
  assign n1620 = n1618 & ~n1619 ;
  assign n1621 = ~n1618 & n1619 ;
  assign n1622 = n1620 | n1621 ;
  assign n1623 = x25 & ~x26 ;
  assign n1624 = ~x25 & x26 ;
  assign n1625 = n1623 | n1624 ;
  assign n1626 = ~x27 & n1625 ;
  assign n1627 = x27 & ~n1625 ;
  assign n1628 = n1626 | n1627 ;
  assign n1629 = x28 & ~x29 ;
  assign n1630 = ~x28 & x29 ;
  assign n1631 = n1629 | n1630 ;
  assign n1632 = ~x30 & n1631 ;
  assign n1633 = x30 & ~n1631 ;
  assign n1634 = n1632 | n1633 ;
  assign n1635 = n1628 & n1634 ;
  assign n1636 = n1622 & ~n1635 ;
  assign n1637 = ~n1622 & n1635 ;
  assign n1638 = n1636 | n1637 ;
  assign n1639 = ( n1618 & n1619 ) | ( n1618 & n1635 ) | ( n1619 & n1635 ) ;
  assign n1640 = n1638 & n1639 ;
  assign n1641 = n1628 & ~n1634 ;
  assign n1642 = ~n1628 & n1634 ;
  assign n1643 = n1641 | n1642 ;
  assign n1644 = n1614 & n1643 ;
  assign n1645 = ~n1640 & n1644 ;
  assign n1646 = n1639 & n1643 ;
  assign n1647 = n1638 & ~n1646 ;
  assign n1648 = n1611 & n1615 ;
  assign n1649 = ~n1647 & n1648 ;
  assign n1650 = ( n1645 & n1647 ) | ( n1645 & ~n1649 ) | ( n1647 & ~n1649 ) ;
  assign n1651 = n1617 & n1650 ;
  assign n1652 = n1646 | n1648 ;
  assign n1653 = n1638 & n1644 ;
  assign n1654 = ~n1640 & n1653 ;
  assign n1655 = ~n1652 & n1654 ;
  assign n1656 = ~n1614 & n1615 ;
  assign n1657 = ( ~n1611 & n1615 ) | ( ~n1611 & n1656 ) | ( n1615 & n1656 ) ;
  assign n1658 = n1639 & ~n1643 ;
  assign n1659 = ( ~n1638 & n1639 ) | ( ~n1638 & n1658 ) | ( n1639 & n1658 ) ;
  assign n1660 = ( n1655 & n1657 ) | ( n1655 & n1659 ) | ( n1657 & n1659 ) ;
  assign n1661 = n1657 | n1659 ;
  assign n1662 = ( n1651 & n1660 ) | ( n1651 & n1661 ) | ( n1660 & n1661 ) ;
  assign n1663 = ~x7 & x8 ;
  assign n1664 = x7 & ~x8 ;
  assign n1665 = n1663 | n1664 ;
  assign n1666 = ~x9 & n1665 ;
  assign n1667 = x9 & ~n1665 ;
  assign n1668 = n1666 | n1667 ;
  assign n1669 = ~x10 & x11 ;
  assign n1670 = x10 & ~x11 ;
  assign n1671 = n1669 | n1670 ;
  assign n1672 = ~x12 & n1671 ;
  assign n1673 = x12 & ~n1671 ;
  assign n1674 = n1672 | n1673 ;
  assign n1675 = n1668 & n1674 ;
  assign n1676 = ( x10 & x11 ) | ( x10 & x12 ) | ( x11 & x12 ) ;
  assign n1677 = ( x7 & x8 ) | ( x7 & x9 ) | ( x8 & x9 ) ;
  assign n1678 = ~n1676 & n1677 ;
  assign n1679 = n1676 & ~n1677 ;
  assign n1680 = n1678 | n1679 ;
  assign n1681 = ~n1675 & n1680 ;
  assign n1682 = n1675 & ~n1680 ;
  assign n1683 = n1681 | n1682 ;
  assign n1684 = n1668 & ~n1674 ;
  assign n1685 = ~n1668 & n1674 ;
  assign n1686 = n1684 | n1685 ;
  assign n1687 = ( n1675 & n1676 ) | ( n1675 & n1677 ) | ( n1676 & n1677 ) ;
  assign n1688 = n1686 & n1687 ;
  assign n1689 = n1683 & ~n1688 ;
  assign n1690 = ( x16 & x17 ) | ( x16 & x18 ) | ( x17 & x18 ) ;
  assign n1691 = ( x13 & x14 ) | ( x13 & x15 ) | ( x14 & x15 ) ;
  assign n1692 = n1690 & ~n1691 ;
  assign n1693 = ~n1690 & n1691 ;
  assign n1694 = n1692 | n1693 ;
  assign n1695 = x13 & ~x14 ;
  assign n1696 = ~x13 & x14 ;
  assign n1697 = n1695 | n1696 ;
  assign n1698 = ~x15 & n1697 ;
  assign n1699 = x15 & ~n1697 ;
  assign n1700 = n1698 | n1699 ;
  assign n1701 = x16 & ~x17 ;
  assign n1702 = ~x16 & x17 ;
  assign n1703 = n1701 | n1702 ;
  assign n1704 = ~x18 & n1703 ;
  assign n1705 = x18 & ~n1703 ;
  assign n1706 = n1704 | n1705 ;
  assign n1707 = n1700 & n1706 ;
  assign n1708 = n1694 & ~n1707 ;
  assign n1709 = ~n1694 & n1707 ;
  assign n1710 = n1708 | n1709 ;
  assign n1711 = ( n1690 & n1691 ) | ( n1690 & n1707 ) | ( n1691 & n1707 ) ;
  assign n1712 = n1710 & n1711 ;
  assign n1713 = n1700 & ~n1706 ;
  assign n1714 = ~n1700 & n1706 ;
  assign n1715 = n1713 | n1714 ;
  assign n1716 = n1686 & n1715 ;
  assign n1717 = ~n1712 & n1716 ;
  assign n1718 = n1711 & n1715 ;
  assign n1719 = n1710 & ~n1718 ;
  assign n1720 = n1683 & n1687 ;
  assign n1721 = ~n1719 & n1720 ;
  assign n1722 = ( n1717 & n1719 ) | ( n1717 & ~n1721 ) | ( n1719 & ~n1721 ) ;
  assign n1723 = n1689 & n1722 ;
  assign n1724 = n1718 | n1720 ;
  assign n1725 = n1710 & n1716 ;
  assign n1726 = ~n1712 & n1725 ;
  assign n1727 = ~n1724 & n1726 ;
  assign n1728 = ~n1686 & n1687 ;
  assign n1729 = ( ~n1683 & n1687 ) | ( ~n1683 & n1728 ) | ( n1687 & n1728 ) ;
  assign n1730 = n1711 & ~n1715 ;
  assign n1731 = ( ~n1710 & n1711 ) | ( ~n1710 & n1730 ) | ( n1711 & n1730 ) ;
  assign n1732 = ( n1727 & n1729 ) | ( n1727 & n1731 ) | ( n1729 & n1731 ) ;
  assign n1733 = n1729 | n1731 ;
  assign n1734 = ( n1723 & n1732 ) | ( n1723 & n1733 ) | ( n1732 & n1733 ) ;
  assign n1735 = n1662 & n1734 ;
  assign n1736 = n1617 & n1655 ;
  assign n1737 = ( n1617 & ~n1650 ) | ( n1617 & n1736 ) | ( ~n1650 & n1736 ) ;
  assign n1738 = ~n1639 & n1643 ;
  assign n1739 = ( ~n1638 & n1643 ) | ( ~n1638 & n1738 ) | ( n1643 & n1738 ) ;
  assign n1740 = n1614 & ~n1615 ;
  assign n1741 = ( ~n1611 & n1614 ) | ( ~n1611 & n1740 ) | ( n1614 & n1740 ) ;
  assign n1742 = ~n1739 & n1741 ;
  assign n1743 = n1739 & ~n1741 ;
  assign n1744 = n1742 | n1743 ;
  assign n1745 = ~n1711 & n1715 ;
  assign n1746 = ( ~n1710 & n1715 ) | ( ~n1710 & n1745 ) | ( n1715 & n1745 ) ;
  assign n1747 = n1686 & ~n1687 ;
  assign n1748 = ( ~n1683 & n1686 ) | ( ~n1683 & n1747 ) | ( n1686 & n1747 ) ;
  assign n1749 = ~n1746 & n1748 ;
  assign n1750 = n1746 & ~n1748 ;
  assign n1751 = n1749 | n1750 ;
  assign n1752 = n1744 & n1751 ;
  assign n1753 = ( n1617 & n1647 ) | ( n1617 & ~n1648 ) | ( n1647 & ~n1648 ) ;
  assign n1754 = n1617 & n1647 ;
  assign n1755 = ( n1645 & n1753 ) | ( n1645 & n1754 ) | ( n1753 & n1754 ) ;
  assign n1756 = n1650 & ~n1755 ;
  assign n1757 = n1752 | n1756 ;
  assign n1758 = n1737 | n1757 ;
  assign n1759 = n1689 & ~n1727 ;
  assign n1760 = ( n1689 & n1719 ) | ( n1689 & n1720 ) | ( n1719 & n1720 ) ;
  assign n1761 = n1689 | n1719 ;
  assign n1762 = ( ~n1717 & n1760 ) | ( ~n1717 & n1761 ) | ( n1760 & n1761 ) ;
  assign n1763 = n1719 | n1720 ;
  assign n1764 = n1717 & ~n1763 ;
  assign n1765 = ( ~n1719 & n1762 ) | ( ~n1719 & n1764 ) | ( n1762 & n1764 ) ;
  assign n1766 = ( ~n1759 & n1762 ) | ( ~n1759 & n1765 ) | ( n1762 & n1765 ) ;
  assign n1767 = n1758 & n1766 ;
  assign n1768 = n1752 & n1756 ;
  assign n1769 = ( n1737 & n1752 ) | ( n1737 & n1768 ) | ( n1752 & n1768 ) ;
  assign n1770 = n1767 | n1769 ;
  assign n1771 = ~n1729 & n1731 ;
  assign n1772 = n1729 & ~n1731 ;
  assign n1773 = n1771 | n1772 ;
  assign n1774 = n1727 | n1773 ;
  assign n1775 = n1723 | n1774 ;
  assign n1776 = n1727 & n1773 ;
  assign n1777 = ( n1723 & n1773 ) | ( n1723 & n1776 ) | ( n1773 & n1776 ) ;
  assign n1778 = n1775 & ~n1777 ;
  assign n1779 = ~n1657 & n1659 ;
  assign n1780 = n1657 & ~n1659 ;
  assign n1781 = n1779 | n1780 ;
  assign n1782 = n1655 | n1781 ;
  assign n1783 = n1651 | n1782 ;
  assign n1784 = n1655 & n1781 ;
  assign n1785 = ( n1651 & n1781 ) | ( n1651 & n1784 ) | ( n1781 & n1784 ) ;
  assign n1786 = n1783 & ~n1785 ;
  assign n1787 = n1778 | n1786 ;
  assign n1788 = n1770 & n1787 ;
  assign n1789 = n1775 & n1783 ;
  assign n1790 = n1777 | n1785 ;
  assign n1791 = n1789 & ~n1790 ;
  assign n1792 = n1662 & ~n1734 ;
  assign n1793 = ~n1662 & n1734 ;
  assign n1794 = n1792 | n1793 ;
  assign n1795 = n1791 | n1794 ;
  assign n1796 = n1788 | n1795 ;
  assign n1797 = n1787 | n1791 ;
  assign n1798 = ( n1770 & n1791 ) | ( n1770 & n1797 ) | ( n1791 & n1797 ) ;
  assign n1799 = ( n1662 & n1734 ) | ( n1662 & n1798 ) | ( n1734 & n1798 ) ;
  assign n1800 = ( n1735 & n1796 ) | ( n1735 & ~n1799 ) | ( n1796 & ~n1799 ) ;
  assign n1801 = n1590 | n1800 ;
  assign n1802 = n1744 & ~n1751 ;
  assign n1803 = ~n1744 & n1751 ;
  assign n1804 = n1802 | n1803 ;
  assign n1805 = ~n1508 & n1535 ;
  assign n1806 = n1508 & ~n1535 ;
  assign n1807 = n1805 | n1806 ;
  assign n1808 = n1804 & n1807 ;
  assign n1809 = n1758 & ~n1769 ;
  assign n1810 = n1766 & ~n1809 ;
  assign n1811 = ~n1752 & n1758 ;
  assign n1812 = n1758 & ~n1766 ;
  assign n1813 = n1737 | n1756 ;
  assign n1814 = n1766 | n1813 ;
  assign n1815 = ( n1811 & n1812 ) | ( n1811 & ~n1814 ) | ( n1812 & ~n1814 ) ;
  assign n1816 = n1810 | n1815 ;
  assign n1817 = n1808 & n1816 ;
  assign n1818 = n1808 | n1815 ;
  assign n1819 = ( n1536 & ~n1559 ) | ( n1536 & n1562 ) | ( ~n1559 & n1562 ) ;
  assign n1820 = ( ~n1536 & n1559 ) | ( ~n1536 & n1819 ) | ( n1559 & n1819 ) ;
  assign n1821 = ( ~n1562 & n1819 ) | ( ~n1562 & n1820 ) | ( n1819 & n1820 ) ;
  assign n1822 = n1810 & n1821 ;
  assign n1823 = ( n1818 & n1821 ) | ( n1818 & n1822 ) | ( n1821 & n1822 ) ;
  assign n1824 = n1817 | n1823 ;
  assign n1825 = ~n1778 & n1786 ;
  assign n1826 = n1778 & ~n1786 ;
  assign n1827 = n1825 | n1826 ;
  assign n1828 = n1770 & n1827 ;
  assign n1829 = n1770 | n1827 ;
  assign n1830 = ~n1828 & n1829 ;
  assign n1831 = ~n1573 & n1579 ;
  assign n1832 = ~n1575 & n1831 ;
  assign n1833 = n1576 & ~n1579 ;
  assign n1834 = n1832 & ~n1833 ;
  assign n1835 = ( n1566 & n1833 ) | ( n1566 & n1834 ) | ( n1833 & n1834 ) ;
  assign n1836 = ( n1566 & n1833 ) | ( n1566 & ~n1834 ) | ( n1833 & ~n1834 ) ;
  assign n1837 = ( n1834 & ~n1835 ) | ( n1834 & n1836 ) | ( ~n1835 & n1836 ) ;
  assign n1838 = ( n1824 & n1830 ) | ( n1824 & n1837 ) | ( n1830 & n1837 ) ;
  assign n1839 = n1801 & n1838 ;
  assign n1840 = n1662 | n1734 ;
  assign n1841 = n1735 | n1840 ;
  assign n1842 = ( n1735 & n1798 ) | ( n1735 & n1841 ) | ( n1798 & n1841 ) ;
  assign n1843 = n1585 & n1842 ;
  assign n1844 = n1798 & n1840 ;
  assign n1845 = n1584 | n1735 ;
  assign n1846 = ( n1582 & n1735 ) | ( n1582 & n1845 ) | ( n1735 & n1845 ) ;
  assign n1847 = n1844 | n1846 ;
  assign n1848 = n1843 | n1847 ;
  assign n1849 = n1590 & n1800 ;
  assign n1850 = ( n1843 & n1848 ) | ( n1843 & n1849 ) | ( n1848 & n1849 ) ;
  assign n1851 = n1843 | n1848 ;
  assign n1852 = ( n1839 & n1850 ) | ( n1839 & n1851 ) | ( n1850 & n1851 ) ;
  assign n1002 = ~x43 & x44 ;
  assign n1003 = x43 & ~x44 ;
  assign n1004 = n1002 | n1003 ;
  assign n1005 = ~x45 & n1004 ;
  assign n1006 = x45 & ~n1004 ;
  assign n1007 = n1005 | n1006 ;
  assign n1008 = ~x46 & x47 ;
  assign n1009 = x46 & ~x47 ;
  assign n1010 = n1008 | n1009 ;
  assign n1011 = ~x48 & n1010 ;
  assign n1012 = x48 & ~n1010 ;
  assign n1013 = n1011 | n1012 ;
  assign n1014 = n1007 & n1013 ;
  assign n1015 = ( x46 & x47 ) | ( x46 & x48 ) | ( x47 & x48 ) ;
  assign n1016 = ( x43 & x44 ) | ( x43 & x45 ) | ( x44 & x45 ) ;
  assign n1017 = ~n1015 & n1016 ;
  assign n1018 = n1015 & ~n1016 ;
  assign n1019 = n1017 | n1018 ;
  assign n1020 = ~n1014 & n1019 ;
  assign n1021 = n1014 & ~n1019 ;
  assign n1022 = n1020 | n1021 ;
  assign n1023 = n1007 & ~n1013 ;
  assign n1024 = ~n1007 & n1013 ;
  assign n1025 = n1023 | n1024 ;
  assign n1026 = ( n1014 & n1015 ) | ( n1014 & n1016 ) | ( n1015 & n1016 ) ;
  assign n1027 = n1025 & n1026 ;
  assign n1028 = n1022 & ~n1027 ;
  assign n1029 = ( x52 & x53 ) | ( x52 & x54 ) | ( x53 & x54 ) ;
  assign n1030 = ( x49 & x50 ) | ( x49 & x51 ) | ( x50 & x51 ) ;
  assign n1031 = n1029 & ~n1030 ;
  assign n1032 = ~n1029 & n1030 ;
  assign n1033 = n1031 | n1032 ;
  assign n1034 = x49 & ~x50 ;
  assign n1035 = ~x49 & x50 ;
  assign n1036 = n1034 | n1035 ;
  assign n1037 = ~x51 & n1036 ;
  assign n1038 = x51 & ~n1036 ;
  assign n1039 = n1037 | n1038 ;
  assign n1040 = x52 & ~x53 ;
  assign n1041 = ~x52 & x53 ;
  assign n1042 = n1040 | n1041 ;
  assign n1043 = ~x54 & n1042 ;
  assign n1044 = x54 & ~n1042 ;
  assign n1045 = n1043 | n1044 ;
  assign n1046 = n1039 & n1045 ;
  assign n1047 = n1033 & ~n1046 ;
  assign n1048 = ~n1033 & n1046 ;
  assign n1049 = n1047 | n1048 ;
  assign n1050 = ( n1029 & n1030 ) | ( n1029 & n1046 ) | ( n1030 & n1046 ) ;
  assign n1051 = n1049 & n1050 ;
  assign n1052 = n1039 & ~n1045 ;
  assign n1053 = ~n1039 & n1045 ;
  assign n1054 = n1052 | n1053 ;
  assign n1055 = n1025 & n1054 ;
  assign n1056 = ~n1051 & n1055 ;
  assign n1057 = n1050 & n1054 ;
  assign n1058 = n1049 & ~n1057 ;
  assign n1059 = n1022 & n1026 ;
  assign n1060 = ~n1058 & n1059 ;
  assign n1061 = ( n1056 & n1058 ) | ( n1056 & ~n1060 ) | ( n1058 & ~n1060 ) ;
  assign n1062 = n1028 & n1061 ;
  assign n1063 = n1057 | n1059 ;
  assign n1064 = n1049 & n1055 ;
  assign n1065 = ~n1051 & n1064 ;
  assign n1066 = ~n1063 & n1065 ;
  assign n1067 = ~n1025 & n1026 ;
  assign n1068 = ( ~n1022 & n1026 ) | ( ~n1022 & n1067 ) | ( n1026 & n1067 ) ;
  assign n1069 = n1050 & ~n1054 ;
  assign n1070 = ( ~n1049 & n1050 ) | ( ~n1049 & n1069 ) | ( n1050 & n1069 ) ;
  assign n1071 = ( n1066 & n1068 ) | ( n1066 & n1070 ) | ( n1068 & n1070 ) ;
  assign n1072 = n1068 | n1070 ;
  assign n1073 = ( n1062 & n1071 ) | ( n1062 & n1072 ) | ( n1071 & n1072 ) ;
  assign n1074 = ( x34 & x35 ) | ( x34 & x36 ) | ( x35 & x36 ) ;
  assign n1075 = ( x31 & x32 ) | ( x31 & x33 ) | ( x32 & x33 ) ;
  assign n1076 = n1074 & ~n1075 ;
  assign n1077 = ~n1074 & n1075 ;
  assign n1078 = n1076 | n1077 ;
  assign n1079 = ~x31 & x32 ;
  assign n1080 = x31 & ~x32 ;
  assign n1081 = n1079 | n1080 ;
  assign n1082 = ~x33 & n1081 ;
  assign n1083 = x33 & ~n1081 ;
  assign n1084 = n1082 | n1083 ;
  assign n1085 = ~x34 & x35 ;
  assign n1086 = x34 & ~x35 ;
  assign n1087 = n1085 | n1086 ;
  assign n1088 = ~x36 & n1087 ;
  assign n1089 = x36 & ~n1087 ;
  assign n1090 = n1088 | n1089 ;
  assign n1091 = n1084 & n1090 ;
  assign n1092 = n1078 & ~n1091 ;
  assign n1093 = ~n1078 & n1091 ;
  assign n1094 = n1092 | n1093 ;
  assign n1095 = n1084 & ~n1090 ;
  assign n1096 = ~n1084 & n1090 ;
  assign n1097 = n1095 | n1096 ;
  assign n1098 = ( n1074 & n1075 ) | ( n1074 & n1091 ) | ( n1075 & n1091 ) ;
  assign n1099 = n1097 & n1098 ;
  assign n1100 = n1094 & ~n1099 ;
  assign n1101 = ( x40 & x41 ) | ( x40 & x42 ) | ( x41 & x42 ) ;
  assign n1102 = ( x37 & x38 ) | ( x37 & x39 ) | ( x38 & x39 ) ;
  assign n1103 = n1101 & ~n1102 ;
  assign n1104 = ~n1101 & n1102 ;
  assign n1105 = n1103 | n1104 ;
  assign n1106 = ~x37 & x38 ;
  assign n1107 = x37 & ~x38 ;
  assign n1108 = n1106 | n1107 ;
  assign n1109 = ~x39 & n1108 ;
  assign n1110 = x39 & ~n1108 ;
  assign n1111 = n1109 | n1110 ;
  assign n1112 = ~x40 & x41 ;
  assign n1113 = x40 & ~x41 ;
  assign n1114 = n1112 | n1113 ;
  assign n1115 = ~x42 & n1114 ;
  assign n1116 = x42 & ~n1114 ;
  assign n1117 = n1115 | n1116 ;
  assign n1118 = n1111 & n1117 ;
  assign n1119 = n1105 & ~n1118 ;
  assign n1120 = ~n1105 & n1118 ;
  assign n1121 = n1119 | n1120 ;
  assign n1122 = ( n1101 & n1102 ) | ( n1101 & n1118 ) | ( n1102 & n1118 ) ;
  assign n1123 = n1121 & n1122 ;
  assign n1124 = n1111 & ~n1117 ;
  assign n1125 = ~n1111 & n1117 ;
  assign n1126 = n1124 | n1125 ;
  assign n1127 = n1097 & n1126 ;
  assign n1128 = ~n1123 & n1127 ;
  assign n1129 = n1122 & n1126 ;
  assign n1130 = n1121 & ~n1129 ;
  assign n1131 = n1094 & n1098 ;
  assign n1132 = ~n1130 & n1131 ;
  assign n1133 = ( n1128 & n1130 ) | ( n1128 & ~n1132 ) | ( n1130 & ~n1132 ) ;
  assign n1134 = n1100 & n1133 ;
  assign n1135 = n1129 | n1131 ;
  assign n1136 = n1121 & n1127 ;
  assign n1137 = ~n1123 & n1136 ;
  assign n1138 = ~n1135 & n1137 ;
  assign n1139 = ~n1097 & n1098 ;
  assign n1140 = ( ~n1094 & n1098 ) | ( ~n1094 & n1139 ) | ( n1098 & n1139 ) ;
  assign n1141 = n1122 & ~n1126 ;
  assign n1142 = ( ~n1121 & n1122 ) | ( ~n1121 & n1141 ) | ( n1122 & n1141 ) ;
  assign n1143 = ( n1138 & n1140 ) | ( n1138 & n1142 ) | ( n1140 & n1142 ) ;
  assign n1144 = n1140 | n1142 ;
  assign n1145 = ( n1134 & n1143 ) | ( n1134 & n1144 ) | ( n1143 & n1144 ) ;
  assign n1146 = n1073 & n1145 ;
  assign n1147 = n1073 | n1145 ;
  assign n1148 = n1146 | n1147 ;
  assign n1149 = ~n1140 & n1142 ;
  assign n1150 = n1140 & ~n1142 ;
  assign n1151 = n1149 | n1150 ;
  assign n1152 = n1138 | n1151 ;
  assign n1153 = n1134 | n1152 ;
  assign n1154 = ~n1068 & n1070 ;
  assign n1155 = n1068 & ~n1070 ;
  assign n1156 = n1154 | n1155 ;
  assign n1157 = n1066 | n1156 ;
  assign n1158 = n1062 | n1157 ;
  assign n1159 = n1153 & n1158 ;
  assign n1160 = n1138 & n1151 ;
  assign n1161 = ( n1134 & n1151 ) | ( n1134 & n1160 ) | ( n1151 & n1160 ) ;
  assign n1162 = n1066 & n1156 ;
  assign n1163 = ( n1062 & n1156 ) | ( n1062 & n1162 ) | ( n1156 & n1162 ) ;
  assign n1164 = n1161 | n1163 ;
  assign n1165 = n1159 & ~n1164 ;
  assign n1166 = n1028 & n1066 ;
  assign n1167 = ( n1028 & ~n1061 ) | ( n1028 & n1166 ) | ( ~n1061 & n1166 ) ;
  assign n1168 = ~n1050 & n1054 ;
  assign n1169 = ( ~n1049 & n1054 ) | ( ~n1049 & n1168 ) | ( n1054 & n1168 ) ;
  assign n1170 = n1025 & ~n1026 ;
  assign n1171 = ( ~n1022 & n1025 ) | ( ~n1022 & n1170 ) | ( n1025 & n1170 ) ;
  assign n1172 = ~n1169 & n1171 ;
  assign n1173 = n1169 & ~n1171 ;
  assign n1174 = n1172 | n1173 ;
  assign n1175 = ~n1122 & n1126 ;
  assign n1176 = ( ~n1121 & n1126 ) | ( ~n1121 & n1175 ) | ( n1126 & n1175 ) ;
  assign n1177 = n1097 & ~n1098 ;
  assign n1178 = ( ~n1094 & n1097 ) | ( ~n1094 & n1177 ) | ( n1097 & n1177 ) ;
  assign n1179 = ~n1176 & n1178 ;
  assign n1180 = n1176 & ~n1178 ;
  assign n1181 = n1179 | n1180 ;
  assign n1182 = n1174 & n1181 ;
  assign n1183 = ( n1028 & n1058 ) | ( n1028 & ~n1059 ) | ( n1058 & ~n1059 ) ;
  assign n1184 = n1028 & n1058 ;
  assign n1185 = ( n1056 & n1183 ) | ( n1056 & n1184 ) | ( n1183 & n1184 ) ;
  assign n1186 = n1061 & ~n1185 ;
  assign n1187 = n1182 | n1186 ;
  assign n1188 = n1167 | n1187 ;
  assign n1189 = n1100 & ~n1138 ;
  assign n1190 = ( n1100 & n1130 ) | ( n1100 & n1131 ) | ( n1130 & n1131 ) ;
  assign n1191 = n1100 | n1130 ;
  assign n1192 = ( ~n1128 & n1190 ) | ( ~n1128 & n1191 ) | ( n1190 & n1191 ) ;
  assign n1193 = n1130 | n1131 ;
  assign n1194 = n1128 & ~n1193 ;
  assign n1195 = ( ~n1130 & n1192 ) | ( ~n1130 & n1194 ) | ( n1192 & n1194 ) ;
  assign n1196 = ( ~n1189 & n1192 ) | ( ~n1189 & n1195 ) | ( n1192 & n1195 ) ;
  assign n1197 = n1188 & n1196 ;
  assign n1198 = n1182 & n1186 ;
  assign n1199 = ( n1167 & n1182 ) | ( n1167 & n1198 ) | ( n1182 & n1198 ) ;
  assign n1200 = n1197 | n1199 ;
  assign n1201 = n1153 & ~n1161 ;
  assign n1202 = n1158 & ~n1163 ;
  assign n1203 = n1201 | n1202 ;
  assign n1204 = n1165 | n1203 ;
  assign n1205 = ( n1165 & n1200 ) | ( n1165 & n1204 ) | ( n1200 & n1204 ) ;
  assign n1206 = ( n1146 & n1148 ) | ( n1146 & n1205 ) | ( n1148 & n1205 ) ;
  assign n1207 = ~x67 & x68 ;
  assign n1208 = x67 & ~x68 ;
  assign n1209 = n1207 | n1208 ;
  assign n1210 = ~x69 & n1209 ;
  assign n1211 = x69 & ~n1209 ;
  assign n1212 = n1210 | n1211 ;
  assign n1213 = ~x70 & x71 ;
  assign n1214 = x70 & ~x71 ;
  assign n1215 = n1213 | n1214 ;
  assign n1216 = ~x72 & n1215 ;
  assign n1217 = x72 & ~n1215 ;
  assign n1218 = n1216 | n1217 ;
  assign n1219 = n1212 & n1218 ;
  assign n1220 = ( x70 & x71 ) | ( x70 & x72 ) | ( x71 & x72 ) ;
  assign n1221 = ( x67 & x68 ) | ( x67 & x69 ) | ( x68 & x69 ) ;
  assign n1222 = ~n1220 & n1221 ;
  assign n1223 = n1220 & ~n1221 ;
  assign n1224 = n1222 | n1223 ;
  assign n1225 = ~n1219 & n1224 ;
  assign n1226 = n1219 & ~n1224 ;
  assign n1227 = n1225 | n1226 ;
  assign n1228 = n1212 & ~n1218 ;
  assign n1229 = ~n1212 & n1218 ;
  assign n1230 = n1228 | n1229 ;
  assign n1231 = ( n1219 & n1220 ) | ( n1219 & n1221 ) | ( n1220 & n1221 ) ;
  assign n1232 = n1230 & n1231 ;
  assign n1233 = n1227 & ~n1232 ;
  assign n1234 = ( x76 & x77 ) | ( x76 & x78 ) | ( x77 & x78 ) ;
  assign n1235 = ( x73 & x74 ) | ( x73 & x75 ) | ( x74 & x75 ) ;
  assign n1236 = n1234 & ~n1235 ;
  assign n1237 = ~n1234 & n1235 ;
  assign n1238 = n1236 | n1237 ;
  assign n1239 = x73 & ~x74 ;
  assign n1240 = ~x73 & x74 ;
  assign n1241 = n1239 | n1240 ;
  assign n1242 = ~x75 & n1241 ;
  assign n1243 = x75 & ~n1241 ;
  assign n1244 = n1242 | n1243 ;
  assign n1245 = x76 & ~x77 ;
  assign n1246 = ~x76 & x77 ;
  assign n1247 = n1245 | n1246 ;
  assign n1248 = ~x78 & n1247 ;
  assign n1249 = x78 & ~n1247 ;
  assign n1250 = n1248 | n1249 ;
  assign n1251 = n1244 & n1250 ;
  assign n1252 = n1238 & ~n1251 ;
  assign n1253 = ~n1238 & n1251 ;
  assign n1254 = n1252 | n1253 ;
  assign n1255 = ( n1234 & n1235 ) | ( n1234 & n1251 ) | ( n1235 & n1251 ) ;
  assign n1256 = n1254 & n1255 ;
  assign n1257 = n1244 & ~n1250 ;
  assign n1258 = ~n1244 & n1250 ;
  assign n1259 = n1257 | n1258 ;
  assign n1260 = n1230 & n1259 ;
  assign n1261 = ~n1256 & n1260 ;
  assign n1262 = n1255 & n1259 ;
  assign n1263 = n1254 & ~n1262 ;
  assign n1264 = n1227 & n1231 ;
  assign n1265 = ~n1263 & n1264 ;
  assign n1266 = ( n1261 & n1263 ) | ( n1261 & ~n1265 ) | ( n1263 & ~n1265 ) ;
  assign n1267 = n1233 & n1266 ;
  assign n1268 = n1262 | n1264 ;
  assign n1269 = n1254 & n1260 ;
  assign n1270 = ~n1256 & n1269 ;
  assign n1271 = ~n1268 & n1270 ;
  assign n1272 = ~n1230 & n1231 ;
  assign n1273 = ( ~n1227 & n1231 ) | ( ~n1227 & n1272 ) | ( n1231 & n1272 ) ;
  assign n1274 = n1255 & ~n1259 ;
  assign n1275 = ( ~n1254 & n1255 ) | ( ~n1254 & n1274 ) | ( n1255 & n1274 ) ;
  assign n1276 = ( n1271 & n1273 ) | ( n1271 & n1275 ) | ( n1273 & n1275 ) ;
  assign n1277 = n1273 | n1275 ;
  assign n1278 = ( n1267 & n1276 ) | ( n1267 & n1277 ) | ( n1276 & n1277 ) ;
  assign n1279 = ~x55 & x56 ;
  assign n1280 = x55 & ~x56 ;
  assign n1281 = n1279 | n1280 ;
  assign n1282 = ~x57 & n1281 ;
  assign n1283 = x57 & ~n1281 ;
  assign n1284 = n1282 | n1283 ;
  assign n1285 = ~x58 & x59 ;
  assign n1286 = x58 & ~x59 ;
  assign n1287 = n1285 | n1286 ;
  assign n1288 = ~x60 & n1287 ;
  assign n1289 = x60 & ~n1287 ;
  assign n1290 = n1288 | n1289 ;
  assign n1291 = n1284 & n1290 ;
  assign n1292 = ( x58 & x59 ) | ( x58 & x60 ) | ( x59 & x60 ) ;
  assign n1293 = ( x55 & x56 ) | ( x55 & x57 ) | ( x56 & x57 ) ;
  assign n1294 = ~n1292 & n1293 ;
  assign n1295 = n1292 & ~n1293 ;
  assign n1296 = n1294 | n1295 ;
  assign n1297 = ~n1291 & n1296 ;
  assign n1298 = n1291 & ~n1296 ;
  assign n1299 = n1297 | n1298 ;
  assign n1300 = n1284 & ~n1290 ;
  assign n1301 = ~n1284 & n1290 ;
  assign n1302 = n1300 | n1301 ;
  assign n1303 = ( n1291 & n1292 ) | ( n1291 & n1293 ) | ( n1292 & n1293 ) ;
  assign n1304 = n1302 & n1303 ;
  assign n1305 = n1299 & ~n1304 ;
  assign n1306 = ( x64 & x65 ) | ( x64 & x66 ) | ( x65 & x66 ) ;
  assign n1307 = ( x61 & x62 ) | ( x61 & x63 ) | ( x62 & x63 ) ;
  assign n1308 = n1306 & ~n1307 ;
  assign n1309 = ~n1306 & n1307 ;
  assign n1310 = n1308 | n1309 ;
  assign n1311 = x61 & ~x62 ;
  assign n1312 = ~x61 & x62 ;
  assign n1313 = n1311 | n1312 ;
  assign n1314 = ~x63 & n1313 ;
  assign n1315 = x63 & ~n1313 ;
  assign n1316 = n1314 | n1315 ;
  assign n1317 = x64 & ~x65 ;
  assign n1318 = ~x64 & x65 ;
  assign n1319 = n1317 | n1318 ;
  assign n1320 = ~x66 & n1319 ;
  assign n1321 = x66 & ~n1319 ;
  assign n1322 = n1320 | n1321 ;
  assign n1323 = n1316 & n1322 ;
  assign n1324 = n1310 & ~n1323 ;
  assign n1325 = ~n1310 & n1323 ;
  assign n1326 = n1324 | n1325 ;
  assign n1327 = ( n1306 & n1307 ) | ( n1306 & n1323 ) | ( n1307 & n1323 ) ;
  assign n1328 = n1326 & n1327 ;
  assign n1329 = n1316 & ~n1322 ;
  assign n1330 = ~n1316 & n1322 ;
  assign n1331 = n1329 | n1330 ;
  assign n1332 = n1302 & n1331 ;
  assign n1333 = ~n1328 & n1332 ;
  assign n1334 = n1327 & n1331 ;
  assign n1335 = n1326 & ~n1334 ;
  assign n1336 = n1299 & n1303 ;
  assign n1337 = ~n1335 & n1336 ;
  assign n1338 = ( n1333 & n1335 ) | ( n1333 & ~n1337 ) | ( n1335 & ~n1337 ) ;
  assign n1339 = n1305 & n1338 ;
  assign n1340 = n1334 | n1336 ;
  assign n1341 = n1326 & n1332 ;
  assign n1342 = ~n1328 & n1341 ;
  assign n1343 = ~n1340 & n1342 ;
  assign n1344 = ~n1302 & n1303 ;
  assign n1345 = ( ~n1299 & n1303 ) | ( ~n1299 & n1344 ) | ( n1303 & n1344 ) ;
  assign n1346 = n1327 & ~n1331 ;
  assign n1347 = ( ~n1326 & n1327 ) | ( ~n1326 & n1346 ) | ( n1327 & n1346 ) ;
  assign n1348 = ( n1343 & n1345 ) | ( n1343 & n1347 ) | ( n1345 & n1347 ) ;
  assign n1349 = n1345 | n1347 ;
  assign n1350 = ( n1339 & n1348 ) | ( n1339 & n1349 ) | ( n1348 & n1349 ) ;
  assign n1351 = n1278 & n1350 ;
  assign n1352 = ~n1345 & n1347 ;
  assign n1353 = n1345 & ~n1347 ;
  assign n1354 = n1352 | n1353 ;
  assign n1355 = n1343 | n1354 ;
  assign n1356 = n1339 | n1355 ;
  assign n1357 = ~n1273 & n1275 ;
  assign n1358 = n1273 & ~n1275 ;
  assign n1359 = n1357 | n1358 ;
  assign n1360 = n1271 | n1359 ;
  assign n1361 = n1267 | n1360 ;
  assign n1362 = n1356 & n1361 ;
  assign n1363 = n1343 & n1354 ;
  assign n1364 = ( n1339 & n1354 ) | ( n1339 & n1363 ) | ( n1354 & n1363 ) ;
  assign n1365 = n1271 & n1359 ;
  assign n1366 = ( n1267 & n1359 ) | ( n1267 & n1365 ) | ( n1359 & n1365 ) ;
  assign n1367 = n1364 | n1366 ;
  assign n1368 = n1362 & ~n1367 ;
  assign n1369 = n1233 & n1271 ;
  assign n1370 = ( n1233 & ~n1266 ) | ( n1233 & n1369 ) | ( ~n1266 & n1369 ) ;
  assign n1371 = ~n1255 & n1259 ;
  assign n1372 = ( ~n1254 & n1259 ) | ( ~n1254 & n1371 ) | ( n1259 & n1371 ) ;
  assign n1373 = n1230 & ~n1231 ;
  assign n1374 = ( ~n1227 & n1230 ) | ( ~n1227 & n1373 ) | ( n1230 & n1373 ) ;
  assign n1375 = ~n1372 & n1374 ;
  assign n1376 = n1372 & ~n1374 ;
  assign n1377 = n1375 | n1376 ;
  assign n1378 = ~n1327 & n1331 ;
  assign n1379 = ( ~n1326 & n1331 ) | ( ~n1326 & n1378 ) | ( n1331 & n1378 ) ;
  assign n1380 = n1302 & ~n1303 ;
  assign n1381 = ( ~n1299 & n1302 ) | ( ~n1299 & n1380 ) | ( n1302 & n1380 ) ;
  assign n1382 = ~n1379 & n1381 ;
  assign n1383 = n1379 & ~n1381 ;
  assign n1384 = n1382 | n1383 ;
  assign n1385 = n1377 & n1384 ;
  assign n1386 = ( n1233 & n1263 ) | ( n1233 & ~n1264 ) | ( n1263 & ~n1264 ) ;
  assign n1387 = n1233 & n1263 ;
  assign n1388 = ( n1261 & n1386 ) | ( n1261 & n1387 ) | ( n1386 & n1387 ) ;
  assign n1389 = n1266 & ~n1388 ;
  assign n1390 = n1385 | n1389 ;
  assign n1391 = n1370 | n1390 ;
  assign n1392 = n1305 & ~n1343 ;
  assign n1393 = ( n1305 & n1335 ) | ( n1305 & n1336 ) | ( n1335 & n1336 ) ;
  assign n1394 = n1305 | n1335 ;
  assign n1395 = ( ~n1333 & n1393 ) | ( ~n1333 & n1394 ) | ( n1393 & n1394 ) ;
  assign n1396 = n1335 | n1336 ;
  assign n1397 = n1333 & ~n1396 ;
  assign n1398 = ( ~n1335 & n1395 ) | ( ~n1335 & n1397 ) | ( n1395 & n1397 ) ;
  assign n1399 = ( ~n1392 & n1395 ) | ( ~n1392 & n1398 ) | ( n1395 & n1398 ) ;
  assign n1400 = n1391 & n1399 ;
  assign n1401 = n1385 & n1389 ;
  assign n1402 = ( n1370 & n1385 ) | ( n1370 & n1401 ) | ( n1385 & n1401 ) ;
  assign n1403 = n1400 | n1402 ;
  assign n1404 = n1356 & ~n1364 ;
  assign n1405 = n1361 & ~n1366 ;
  assign n1406 = n1404 | n1405 ;
  assign n1407 = n1368 | n1406 ;
  assign n1408 = ( n1368 & n1403 ) | ( n1368 & n1407 ) | ( n1403 & n1407 ) ;
  assign n1409 = n1278 | n1350 ;
  assign n1410 = n1351 | n1409 ;
  assign n1411 = ( n1351 & n1408 ) | ( n1351 & n1410 ) | ( n1408 & n1410 ) ;
  assign n1412 = n1206 & n1411 ;
  assign n1413 = n1408 & n1409 ;
  assign n1414 = n1145 | n1351 ;
  assign n1415 = n1073 | n1351 ;
  assign n1416 = ( n1205 & n1414 ) | ( n1205 & n1415 ) | ( n1414 & n1415 ) ;
  assign n1417 = n1413 | n1416 ;
  assign n1418 = n1403 & n1406 ;
  assign n1419 = ~n1278 & n1350 ;
  assign n1420 = n1278 & ~n1350 ;
  assign n1421 = n1419 | n1420 ;
  assign n1422 = n1368 | n1421 ;
  assign n1423 = n1418 | n1422 ;
  assign n1424 = n1408 & n1421 ;
  assign n1425 = n1423 & ~n1424 ;
  assign n1426 = n1200 & n1203 ;
  assign n1427 = ~n1073 & n1145 ;
  assign n1428 = n1073 & ~n1145 ;
  assign n1429 = n1427 | n1428 ;
  assign n1430 = n1165 | n1429 ;
  assign n1431 = n1426 | n1430 ;
  assign n1432 = n1205 & n1429 ;
  assign n1433 = n1431 & ~n1432 ;
  assign n1434 = n1425 | n1433 ;
  assign n1435 = n1391 & ~n1402 ;
  assign n1436 = n1399 & ~n1435 ;
  assign n1437 = n1377 & ~n1384 ;
  assign n1438 = ~n1377 & n1384 ;
  assign n1439 = n1437 | n1438 ;
  assign n1440 = n1174 & ~n1181 ;
  assign n1441 = ~n1174 & n1181 ;
  assign n1442 = n1440 | n1441 ;
  assign n1443 = n1439 & n1442 ;
  assign n1444 = ~n1385 & n1391 ;
  assign n1445 = n1391 & ~n1399 ;
  assign n1446 = n1370 | n1389 ;
  assign n1447 = n1399 | n1446 ;
  assign n1448 = ( n1444 & n1445 ) | ( n1444 & ~n1447 ) | ( n1445 & ~n1447 ) ;
  assign n1449 = n1443 | n1448 ;
  assign n1450 = n1436 | n1449 ;
  assign n1451 = n1167 | n1186 ;
  assign n1452 = ( n1182 & n1196 ) | ( n1182 & ~n1451 ) | ( n1196 & ~n1451 ) ;
  assign n1453 = ( ~n1196 & n1451 ) | ( ~n1196 & n1452 ) | ( n1451 & n1452 ) ;
  assign n1454 = ( ~n1182 & n1452 ) | ( ~n1182 & n1453 ) | ( n1452 & n1453 ) ;
  assign n1455 = n1450 & n1454 ;
  assign n1456 = n1436 | n1448 ;
  assign n1457 = n1443 & n1456 ;
  assign n1458 = ( n1199 & ~n1201 ) | ( n1199 & n1202 ) | ( ~n1201 & n1202 ) ;
  assign n1459 = n1201 & ~n1202 ;
  assign n1460 = ( n1197 & n1458 ) | ( n1197 & ~n1459 ) | ( n1458 & ~n1459 ) ;
  assign n1461 = ( ~n1200 & n1201 ) | ( ~n1200 & n1460 ) | ( n1201 & n1460 ) ;
  assign n1462 = ( ~n1202 & n1460 ) | ( ~n1202 & n1461 ) | ( n1460 & n1461 ) ;
  assign n1463 = ( n1402 & ~n1404 ) | ( n1402 & n1405 ) | ( ~n1404 & n1405 ) ;
  assign n1464 = n1404 & ~n1405 ;
  assign n1465 = ( n1400 & n1463 ) | ( n1400 & ~n1464 ) | ( n1463 & ~n1464 ) ;
  assign n1466 = ( ~n1403 & n1404 ) | ( ~n1403 & n1465 ) | ( n1404 & n1465 ) ;
  assign n1467 = ( ~n1405 & n1465 ) | ( ~n1405 & n1466 ) | ( n1465 & n1466 ) ;
  assign n1468 = ( n1457 & n1462 ) | ( n1457 & n1467 ) | ( n1462 & n1467 ) ;
  assign n1469 = n1462 | n1467 ;
  assign n1470 = ( n1455 & n1468 ) | ( n1455 & n1469 ) | ( n1468 & n1469 ) ;
  assign n1471 = n1434 & n1470 ;
  assign n1472 = n1423 & n1431 ;
  assign n1473 = n1424 | n1432 ;
  assign n1474 = n1472 & ~n1473 ;
  assign n1475 = n1417 & n1474 ;
  assign n1476 = ( n1417 & n1471 ) | ( n1417 & n1475 ) | ( n1471 & n1475 ) ;
  assign n1477 = n1412 | n1476 ;
  assign n1853 = n1477 & n1852 ;
  assign n1854 = n1477 & ~n1853 ;
  assign n1855 = ( n1852 & ~n1853 ) | ( n1852 & n1854 ) | ( ~n1853 & n1854 ) ;
  assign n1856 = n1411 & ~n1412 ;
  assign n1857 = ( n1206 & ~n1412 ) | ( n1206 & n1856 ) | ( ~n1412 & n1856 ) ;
  assign n1858 = n1474 | n1857 ;
  assign n1859 = n1471 | n1858 ;
  assign n1860 = ~n1843 & n1847 ;
  assign n1861 = ( n1590 & n1800 ) | ( n1590 & n1838 ) | ( n1800 & n1838 ) ;
  assign n1862 = n1860 | n1861 ;
  assign n1863 = n1859 & n1862 ;
  assign n1864 = n1471 | n1474 ;
  assign n1865 = n1857 & n1864 ;
  assign n1866 = n1849 & n1860 ;
  assign n1867 = ( n1839 & n1860 ) | ( n1839 & n1866 ) | ( n1860 & n1866 ) ;
  assign n1868 = n1865 | n1867 ;
  assign n1869 = n1863 & ~n1868 ;
  assign n1870 = n1862 & ~n1867 ;
  assign n1871 = n1859 & ~n1865 ;
  assign n1872 = n1870 | n1871 ;
  assign n1873 = n1801 & ~n1849 ;
  assign n1874 = n1838 & n1873 ;
  assign n1875 = n1838 | n1873 ;
  assign n1876 = ~n1874 & n1875 ;
  assign n1877 = n1439 & ~n1442 ;
  assign n1878 = ~n1439 & n1442 ;
  assign n1879 = n1877 | n1878 ;
  assign n1880 = n1804 | n1807 ;
  assign n1881 = n1804 & ~n1807 ;
  assign n1882 = ( ~n1804 & n1880 ) | ( ~n1804 & n1881 ) | ( n1880 & n1881 ) ;
  assign n1883 = n1879 & n1882 ;
  assign n1884 = ~n1450 & n1454 ;
  assign n1885 = ( n1454 & n1457 ) | ( n1454 & n1884 ) | ( n1457 & n1884 ) ;
  assign n1886 = ~n1443 & n1456 ;
  assign n1887 = n1443 & ~n1448 ;
  assign n1888 = ~n1436 & n1887 ;
  assign n1889 = ~n1454 & n1888 ;
  assign n1890 = ( ~n1454 & n1886 ) | ( ~n1454 & n1889 ) | ( n1886 & n1889 ) ;
  assign n1891 = n1885 | n1890 ;
  assign n1892 = n1883 & n1891 ;
  assign n1893 = ~n1808 & n1816 ;
  assign n1894 = n1808 & ~n1815 ;
  assign n1895 = n1810 | n1821 ;
  assign n1896 = n1894 & ~n1895 ;
  assign n1897 = ( ~n1821 & n1893 ) | ( ~n1821 & n1896 ) | ( n1893 & n1896 ) ;
  assign n1898 = ~n1817 & n1823 ;
  assign n1899 = ( n1821 & n1897 ) | ( n1821 & ~n1898 ) | ( n1897 & ~n1898 ) ;
  assign n1900 = n1883 & n1899 ;
  assign n1901 = ( n1891 & n1899 ) | ( n1891 & n1900 ) | ( n1899 & n1900 ) ;
  assign n1902 = n1892 | n1901 ;
  assign n1903 = ( n1824 & n1830 ) | ( n1824 & ~n1837 ) | ( n1830 & ~n1837 ) ;
  assign n1904 = ( ~n1824 & n1837 ) | ( ~n1824 & n1903 ) | ( n1837 & n1903 ) ;
  assign n1905 = ( ~n1830 & n1903 ) | ( ~n1830 & n1904 ) | ( n1903 & n1904 ) ;
  assign n1907 = ( n1457 & ~n1462 ) | ( n1457 & n1467 ) | ( ~n1462 & n1467 ) ;
  assign n1908 = n1462 & ~n1467 ;
  assign n1909 = ( n1455 & n1907 ) | ( n1455 & ~n1908 ) | ( n1907 & ~n1908 ) ;
  assign n1906 = n1455 | n1457 ;
  assign n1910 = ( n1462 & ~n1906 ) | ( n1462 & n1909 ) | ( ~n1906 & n1909 ) ;
  assign n1911 = ( ~n1467 & n1909 ) | ( ~n1467 & n1910 ) | ( n1909 & n1910 ) ;
  assign n1912 = ( n1902 & n1905 ) | ( n1902 & n1911 ) | ( n1905 & n1911 ) ;
  assign n1913 = ( ~n1425 & n1433 ) | ( ~n1425 & n1470 ) | ( n1433 & n1470 ) ;
  assign n1914 = ( n1425 & ~n1470 ) | ( n1425 & n1913 ) | ( ~n1470 & n1913 ) ;
  assign n1915 = ( ~n1433 & n1913 ) | ( ~n1433 & n1914 ) | ( n1913 & n1914 ) ;
  assign n1916 = ( n1876 & n1912 ) | ( n1876 & n1915 ) | ( n1912 & n1915 ) ;
  assign n1917 = n1872 & n1916 ;
  assign n1918 = n1869 | n1917 ;
  assign n1919 = n1855 & n1918 ;
  assign n1920 = n1855 | n1869 ;
  assign n1921 = ~x979 & x980 ;
  assign n1922 = x979 & ~x980 ;
  assign n1923 = n1921 | n1922 ;
  assign n1924 = ~x981 & n1923 ;
  assign n1925 = x981 & ~n1923 ;
  assign n1926 = n1924 | n1925 ;
  assign n1927 = ~x982 & x983 ;
  assign n1928 = x982 & ~x983 ;
  assign n1929 = n1927 | n1928 ;
  assign n1930 = ~x984 & n1929 ;
  assign n1931 = x984 & ~n1929 ;
  assign n1932 = n1930 | n1931 ;
  assign n1933 = n1926 & n1932 ;
  assign n1934 = ( x982 & x983 ) | ( x982 & x984 ) | ( x983 & x984 ) ;
  assign n1935 = ( x979 & x980 ) | ( x979 & x981 ) | ( x980 & x981 ) ;
  assign n1936 = ~n1934 & n1935 ;
  assign n1937 = n1934 & ~n1935 ;
  assign n1938 = n1936 | n1937 ;
  assign n1939 = ~n1933 & n1938 ;
  assign n1940 = n1933 & ~n1938 ;
  assign n1941 = n1939 | n1940 ;
  assign n1942 = n1926 & ~n1932 ;
  assign n1943 = ~n1926 & n1932 ;
  assign n1944 = n1942 | n1943 ;
  assign n1945 = ( n1933 & n1934 ) | ( n1933 & n1935 ) | ( n1934 & n1935 ) ;
  assign n1946 = n1944 & n1945 ;
  assign n1947 = n1941 & ~n1946 ;
  assign n1948 = n1941 & n1945 ;
  assign n1949 = x985 & ~x986 ;
  assign n1950 = ~x985 & x986 ;
  assign n1951 = n1949 | n1950 ;
  assign n1952 = ~x987 & n1951 ;
  assign n1953 = x987 & ~n1951 ;
  assign n1954 = n1952 | n1953 ;
  assign n1955 = x988 & ~x989 ;
  assign n1956 = ~x988 & x989 ;
  assign n1957 = n1955 | n1956 ;
  assign n1958 = ~x990 & n1957 ;
  assign n1959 = x990 & ~n1957 ;
  assign n1960 = n1958 | n1959 ;
  assign n1961 = n1954 & ~n1960 ;
  assign n1962 = ~n1954 & n1960 ;
  assign n1963 = n1961 | n1962 ;
  assign n1964 = ( x988 & x989 ) | ( x988 & x990 ) | ( x989 & x990 ) ;
  assign n1965 = ( x985 & x986 ) | ( x985 & x987 ) | ( x986 & x987 ) ;
  assign n1966 = n1954 & n1960 ;
  assign n1967 = ( n1964 & n1965 ) | ( n1964 & n1966 ) | ( n1965 & n1966 ) ;
  assign n1968 = n1963 & n1967 ;
  assign n1969 = n1948 | n1968 ;
  assign n1970 = n1964 & ~n1965 ;
  assign n1971 = ~n1964 & n1965 ;
  assign n1972 = n1970 | n1971 ;
  assign n1973 = ~n1966 & n1972 ;
  assign n1974 = n1966 & ~n1972 ;
  assign n1975 = n1973 | n1974 ;
  assign n1976 = n1967 & n1975 ;
  assign n1977 = n1944 & n1963 ;
  assign n1978 = n1975 & n1977 ;
  assign n1979 = ~n1976 & n1978 ;
  assign n1980 = ~n1969 & n1979 ;
  assign n1981 = n1947 & n1980 ;
  assign n1982 = ~n1976 & n1977 ;
  assign n1983 = ~n1968 & n1975 ;
  assign n1984 = n1948 & ~n1983 ;
  assign n1985 = ( n1982 & n1983 ) | ( n1982 & ~n1984 ) | ( n1983 & ~n1984 ) ;
  assign n1986 = ( n1947 & n1981 ) | ( n1947 & ~n1985 ) | ( n1981 & ~n1985 ) ;
  assign n1987 = n1963 & ~n1967 ;
  assign n1988 = ( n1963 & ~n1975 ) | ( n1963 & n1987 ) | ( ~n1975 & n1987 ) ;
  assign n1989 = n1944 & ~n1945 ;
  assign n1990 = ( ~n1941 & n1944 ) | ( ~n1941 & n1989 ) | ( n1944 & n1989 ) ;
  assign n1991 = ~n1988 & n1990 ;
  assign n1992 = n1988 & ~n1990 ;
  assign n1993 = n1991 | n1992 ;
  assign n1994 = ( x976 & x977 ) | ( x976 & x978 ) | ( x977 & x978 ) ;
  assign n1995 = ( x973 & x974 ) | ( x973 & x975 ) | ( x974 & x975 ) ;
  assign n1996 = n1994 & ~n1995 ;
  assign n1997 = ~n1994 & n1995 ;
  assign n1998 = n1996 | n1997 ;
  assign n1999 = x973 & ~x974 ;
  assign n2000 = ~x973 & x974 ;
  assign n2001 = n1999 | n2000 ;
  assign n2002 = ~x975 & n2001 ;
  assign n2003 = x975 & ~n2001 ;
  assign n2004 = n2002 | n2003 ;
  assign n2005 = x976 & ~x977 ;
  assign n2006 = ~x976 & x977 ;
  assign n2007 = n2005 | n2006 ;
  assign n2008 = ~x978 & n2007 ;
  assign n2009 = x978 & ~n2007 ;
  assign n2010 = n2008 | n2009 ;
  assign n2011 = n2004 & n2010 ;
  assign n2012 = n1998 & ~n2011 ;
  assign n2013 = ~n1998 & n2011 ;
  assign n2014 = n2012 | n2013 ;
  assign n2015 = n2004 & ~n2010 ;
  assign n2016 = ~n2004 & n2010 ;
  assign n2017 = n2015 | n2016 ;
  assign n2018 = ( n1994 & n1995 ) | ( n1994 & n2011 ) | ( n1995 & n2011 ) ;
  assign n2019 = n2017 & ~n2018 ;
  assign n2020 = ( ~n2014 & n2017 ) | ( ~n2014 & n2019 ) | ( n2017 & n2019 ) ;
  assign n2021 = ~x967 & x968 ;
  assign n2022 = x967 & ~x968 ;
  assign n2023 = n2021 | n2022 ;
  assign n2024 = ~x969 & n2023 ;
  assign n2025 = x969 & ~n2023 ;
  assign n2026 = n2024 | n2025 ;
  assign n2027 = ~x970 & x971 ;
  assign n2028 = x970 & ~x971 ;
  assign n2029 = n2027 | n2028 ;
  assign n2030 = ~x972 & n2029 ;
  assign n2031 = x972 & ~n2029 ;
  assign n2032 = n2030 | n2031 ;
  assign n2033 = n2026 & n2032 ;
  assign n2034 = ( x970 & x971 ) | ( x970 & x972 ) | ( x971 & x972 ) ;
  assign n2035 = ( x967 & x968 ) | ( x967 & x969 ) | ( x968 & x969 ) ;
  assign n2036 = ~n2034 & n2035 ;
  assign n2037 = n2034 & ~n2035 ;
  assign n2038 = n2036 | n2037 ;
  assign n2039 = ~n2033 & n2038 ;
  assign n2040 = n2033 & ~n2038 ;
  assign n2041 = n2039 | n2040 ;
  assign n2042 = n2026 & ~n2032 ;
  assign n2043 = ~n2026 & n2032 ;
  assign n2044 = n2042 | n2043 ;
  assign n2045 = ( n2033 & n2034 ) | ( n2033 & n2035 ) | ( n2034 & n2035 ) ;
  assign n2046 = n2044 & ~n2045 ;
  assign n2047 = ( ~n2041 & n2044 ) | ( ~n2041 & n2046 ) | ( n2044 & n2046 ) ;
  assign n2048 = ~n2020 & n2047 ;
  assign n2049 = n2020 & ~n2047 ;
  assign n2050 = n2048 | n2049 ;
  assign n2051 = n1993 & n2050 ;
  assign n2052 = ( n1947 & ~n1948 ) | ( n1947 & n1983 ) | ( ~n1948 & n1983 ) ;
  assign n2053 = n1947 & n1983 ;
  assign n2054 = ( n1982 & n2052 ) | ( n1982 & n2053 ) | ( n2052 & n2053 ) ;
  assign n2055 = n1985 & ~n2054 ;
  assign n2056 = n2051 | n2055 ;
  assign n2057 = n1986 | n2056 ;
  assign n2058 = n2041 & n2045 ;
  assign n2059 = n2017 & n2018 ;
  assign n2060 = n2058 | n2059 ;
  assign n2061 = n2014 & n2018 ;
  assign n2062 = n2017 & n2044 ;
  assign n2063 = n2014 & n2062 ;
  assign n2064 = ~n2061 & n2063 ;
  assign n2065 = ~n2060 & n2064 ;
  assign n2066 = n2044 & n2045 ;
  assign n2067 = n2041 & ~n2066 ;
  assign n2068 = ~n2065 & n2067 ;
  assign n2069 = ~n2061 & n2062 ;
  assign n2070 = n2014 & ~n2059 ;
  assign n2071 = ( n2058 & n2067 ) | ( n2058 & n2070 ) | ( n2067 & n2070 ) ;
  assign n2072 = n2067 | n2070 ;
  assign n2073 = ( ~n2069 & n2071 ) | ( ~n2069 & n2072 ) | ( n2071 & n2072 ) ;
  assign n2074 = n2058 | n2070 ;
  assign n2075 = n2069 & ~n2074 ;
  assign n2076 = ( ~n2070 & n2073 ) | ( ~n2070 & n2075 ) | ( n2073 & n2075 ) ;
  assign n2077 = ( ~n2068 & n2073 ) | ( ~n2068 & n2076 ) | ( n2073 & n2076 ) ;
  assign n2078 = n2057 & n2077 ;
  assign n2079 = n2051 & n2055 ;
  assign n2080 = ( n1986 & n2051 ) | ( n1986 & n2079 ) | ( n2051 & n2079 ) ;
  assign n2081 = n2078 | n2080 ;
  assign n2082 = n2058 & ~n2070 ;
  assign n2083 = ( n2069 & n2070 ) | ( n2069 & ~n2082 ) | ( n2070 & ~n2082 ) ;
  assign n2084 = n2067 & n2083 ;
  assign n2085 = ~n2044 & n2045 ;
  assign n2086 = ( ~n2041 & n2045 ) | ( ~n2041 & n2085 ) | ( n2045 & n2085 ) ;
  assign n2087 = ~n2017 & n2018 ;
  assign n2088 = ( ~n2014 & n2018 ) | ( ~n2014 & n2087 ) | ( n2018 & n2087 ) ;
  assign n2089 = ~n2086 & n2088 ;
  assign n2090 = n2086 & ~n2088 ;
  assign n2091 = n2089 | n2090 ;
  assign n2092 = n2065 | n2091 ;
  assign n2093 = n2084 | n2092 ;
  assign n2094 = n2065 & n2091 ;
  assign n2095 = ( n2084 & n2091 ) | ( n2084 & n2094 ) | ( n2091 & n2094 ) ;
  assign n2096 = n2093 & ~n2095 ;
  assign n2097 = n1947 & n1985 ;
  assign n2098 = ~n1944 & n1945 ;
  assign n2099 = ( ~n1941 & n1945 ) | ( ~n1941 & n2098 ) | ( n1945 & n2098 ) ;
  assign n2100 = ~n1963 & n1967 ;
  assign n2101 = ( n1967 & ~n1975 ) | ( n1967 & n2100 ) | ( ~n1975 & n2100 ) ;
  assign n2102 = ~n2099 & n2101 ;
  assign n2103 = n2099 & ~n2101 ;
  assign n2104 = n2102 | n2103 ;
  assign n2105 = n1980 | n2104 ;
  assign n2106 = n2097 | n2105 ;
  assign n2107 = n1980 & n2104 ;
  assign n2108 = ( n2097 & n2104 ) | ( n2097 & n2107 ) | ( n2104 & n2107 ) ;
  assign n2109 = n2106 & ~n2108 ;
  assign n2110 = n2096 | n2109 ;
  assign n2111 = n2081 & n2110 ;
  assign n2112 = n2093 & n2106 ;
  assign n2113 = n2095 | n2108 ;
  assign n2114 = n2112 & ~n2113 ;
  assign n2115 = ( n1980 & n2099 ) | ( n1980 & n2101 ) | ( n2099 & n2101 ) ;
  assign n2116 = n2099 | n2101 ;
  assign n2117 = ( n2097 & n2115 ) | ( n2097 & n2116 ) | ( n2115 & n2116 ) ;
  assign n2118 = ( n2065 & n2086 ) | ( n2065 & n2088 ) | ( n2086 & n2088 ) ;
  assign n2119 = n2086 | n2088 ;
  assign n2120 = ( n2084 & n2118 ) | ( n2084 & n2119 ) | ( n2118 & n2119 ) ;
  assign n2121 = ~n2117 & n2120 ;
  assign n2122 = n2117 & ~n2120 ;
  assign n2123 = n2121 | n2122 ;
  assign n2124 = n2114 | n2123 ;
  assign n2125 = n2111 | n2124 ;
  assign n2126 = n2110 | n2114 ;
  assign n2127 = ( n2081 & n2114 ) | ( n2081 & n2126 ) | ( n2114 & n2126 ) ;
  assign n2128 = n2123 & n2127 ;
  assign n2129 = n2125 & ~n2128 ;
  assign n2130 = ( x958 & x959 ) | ( x958 & x960 ) | ( x959 & x960 ) ;
  assign n2131 = ( x955 & x956 ) | ( x955 & x957 ) | ( x956 & x957 ) ;
  assign n2132 = n2130 & ~n2131 ;
  assign n2133 = ~n2130 & n2131 ;
  assign n2134 = n2132 | n2133 ;
  assign n2135 = ~x955 & x956 ;
  assign n2136 = x955 & ~x956 ;
  assign n2137 = n2135 | n2136 ;
  assign n2138 = ~x957 & n2137 ;
  assign n2139 = x957 & ~n2137 ;
  assign n2140 = n2138 | n2139 ;
  assign n2141 = ~x958 & x959 ;
  assign n2142 = x958 & ~x959 ;
  assign n2143 = n2141 | n2142 ;
  assign n2144 = ~x960 & n2143 ;
  assign n2145 = x960 & ~n2143 ;
  assign n2146 = n2144 | n2145 ;
  assign n2147 = n2140 & n2146 ;
  assign n2148 = n2134 & ~n2147 ;
  assign n2149 = ~n2134 & n2147 ;
  assign n2150 = n2148 | n2149 ;
  assign n2151 = n2140 & ~n2146 ;
  assign n2152 = ~n2140 & n2146 ;
  assign n2153 = n2151 | n2152 ;
  assign n2154 = ( n2130 & n2131 ) | ( n2130 & n2147 ) | ( n2131 & n2147 ) ;
  assign n2155 = n2153 & n2154 ;
  assign n2156 = n2150 & ~n2155 ;
  assign n2157 = n2150 & n2154 ;
  assign n2158 = ~x961 & x962 ;
  assign n2159 = x961 & ~x962 ;
  assign n2160 = n2158 | n2159 ;
  assign n2161 = ~x963 & n2160 ;
  assign n2162 = x963 & ~n2160 ;
  assign n2163 = n2161 | n2162 ;
  assign n2164 = ~x964 & x965 ;
  assign n2165 = x964 & ~x965 ;
  assign n2166 = n2164 | n2165 ;
  assign n2167 = ~x966 & n2166 ;
  assign n2168 = x966 & ~n2166 ;
  assign n2169 = n2167 | n2168 ;
  assign n2170 = n2163 & ~n2169 ;
  assign n2171 = ~n2163 & n2169 ;
  assign n2172 = n2170 | n2171 ;
  assign n2173 = ( x964 & x965 ) | ( x964 & x966 ) | ( x965 & x966 ) ;
  assign n2174 = ( x961 & x962 ) | ( x961 & x963 ) | ( x962 & x963 ) ;
  assign n2175 = n2163 & n2169 ;
  assign n2176 = ( n2173 & n2174 ) | ( n2173 & n2175 ) | ( n2174 & n2175 ) ;
  assign n2177 = n2172 & n2176 ;
  assign n2178 = n2157 | n2177 ;
  assign n2179 = n2173 & ~n2174 ;
  assign n2180 = ~n2173 & n2174 ;
  assign n2181 = n2179 | n2180 ;
  assign n2182 = ~n2175 & n2181 ;
  assign n2183 = n2175 & ~n2181 ;
  assign n2184 = n2182 | n2183 ;
  assign n2185 = n2176 & n2184 ;
  assign n2186 = n2153 & n2172 ;
  assign n2187 = n2184 & n2186 ;
  assign n2188 = ~n2185 & n2187 ;
  assign n2189 = ~n2178 & n2188 ;
  assign n2190 = n2156 & n2189 ;
  assign n2191 = ~n2185 & n2186 ;
  assign n2192 = ~n2177 & n2184 ;
  assign n2193 = n2157 & ~n2192 ;
  assign n2194 = ( n2191 & n2192 ) | ( n2191 & ~n2193 ) | ( n2192 & ~n2193 ) ;
  assign n2195 = ( n2156 & n2190 ) | ( n2156 & ~n2194 ) | ( n2190 & ~n2194 ) ;
  assign n2196 = n2172 & ~n2176 ;
  assign n2197 = ( n2172 & ~n2184 ) | ( n2172 & n2196 ) | ( ~n2184 & n2196 ) ;
  assign n2198 = n2153 & ~n2154 ;
  assign n2199 = ( ~n2150 & n2153 ) | ( ~n2150 & n2198 ) | ( n2153 & n2198 ) ;
  assign n2200 = ~n2197 & n2199 ;
  assign n2201 = n2197 & ~n2199 ;
  assign n2202 = n2200 | n2201 ;
  assign n2203 = ( x952 & x953 ) | ( x952 & x954 ) | ( x953 & x954 ) ;
  assign n2204 = ( x949 & x950 ) | ( x949 & x951 ) | ( x950 & x951 ) ;
  assign n2205 = n2203 & ~n2204 ;
  assign n2206 = ~n2203 & n2204 ;
  assign n2207 = n2205 | n2206 ;
  assign n2208 = ~x949 & x950 ;
  assign n2209 = x949 & ~x950 ;
  assign n2210 = n2208 | n2209 ;
  assign n2211 = ~x951 & n2210 ;
  assign n2212 = x951 & ~n2210 ;
  assign n2213 = n2211 | n2212 ;
  assign n2214 = ~x952 & x953 ;
  assign n2215 = x952 & ~x953 ;
  assign n2216 = n2214 | n2215 ;
  assign n2217 = ~x954 & n2216 ;
  assign n2218 = x954 & ~n2216 ;
  assign n2219 = n2217 | n2218 ;
  assign n2220 = n2213 & n2219 ;
  assign n2221 = n2207 & ~n2220 ;
  assign n2222 = ~n2207 & n2220 ;
  assign n2223 = n2221 | n2222 ;
  assign n2224 = n2213 & ~n2219 ;
  assign n2225 = ~n2213 & n2219 ;
  assign n2226 = n2224 | n2225 ;
  assign n2227 = ( n2203 & n2204 ) | ( n2203 & n2220 ) | ( n2204 & n2220 ) ;
  assign n2228 = n2226 & ~n2227 ;
  assign n2229 = ( ~n2223 & n2226 ) | ( ~n2223 & n2228 ) | ( n2226 & n2228 ) ;
  assign n2230 = ~x943 & x944 ;
  assign n2231 = x943 & ~x944 ;
  assign n2232 = n2230 | n2231 ;
  assign n2233 = ~x945 & n2232 ;
  assign n2234 = x945 & ~n2232 ;
  assign n2235 = n2233 | n2234 ;
  assign n2236 = ~x946 & x947 ;
  assign n2237 = x946 & ~x947 ;
  assign n2238 = n2236 | n2237 ;
  assign n2239 = ~x948 & n2238 ;
  assign n2240 = x948 & ~n2238 ;
  assign n2241 = n2239 | n2240 ;
  assign n2242 = n2235 & ~n2241 ;
  assign n2243 = ~n2235 & n2241 ;
  assign n2244 = n2242 | n2243 ;
  assign n2245 = ( x946 & x947 ) | ( x946 & x948 ) | ( x947 & x948 ) ;
  assign n2246 = ( x943 & x944 ) | ( x943 & x945 ) | ( x944 & x945 ) ;
  assign n2247 = n2245 & ~n2246 ;
  assign n2248 = ~n2245 & n2246 ;
  assign n2249 = n2247 | n2248 ;
  assign n2250 = n2235 & n2241 ;
  assign n2251 = n2249 & ~n2250 ;
  assign n2252 = ~n2249 & n2250 ;
  assign n2253 = n2251 | n2252 ;
  assign n2254 = ( n2245 & n2246 ) | ( n2245 & n2250 ) | ( n2246 & n2250 ) ;
  assign n2255 = n2244 & ~n2254 ;
  assign n2256 = ( n2244 & ~n2253 ) | ( n2244 & n2255 ) | ( ~n2253 & n2255 ) ;
  assign n2257 = ~n2229 & n2256 ;
  assign n2258 = n2229 & ~n2256 ;
  assign n2259 = n2257 | n2258 ;
  assign n2260 = n2202 & n2259 ;
  assign n2261 = ( n2156 & ~n2157 ) | ( n2156 & n2192 ) | ( ~n2157 & n2192 ) ;
  assign n2262 = n2156 & n2192 ;
  assign n2263 = ( n2191 & n2261 ) | ( n2191 & n2262 ) | ( n2261 & n2262 ) ;
  assign n2264 = n2194 & ~n2263 ;
  assign n2265 = n2260 | n2264 ;
  assign n2266 = n2195 | n2265 ;
  assign n2267 = n2253 & n2254 ;
  assign n2268 = n2226 & n2227 ;
  assign n2269 = n2267 | n2268 ;
  assign n2270 = n2223 & n2227 ;
  assign n2271 = n2226 & n2244 ;
  assign n2272 = n2223 & n2271 ;
  assign n2273 = ~n2270 & n2272 ;
  assign n2274 = ~n2269 & n2273 ;
  assign n2275 = n2244 & n2254 ;
  assign n2276 = n2253 & ~n2275 ;
  assign n2277 = ~n2274 & n2276 ;
  assign n2278 = ~n2270 & n2271 ;
  assign n2279 = n2223 & ~n2268 ;
  assign n2280 = ( n2267 & n2276 ) | ( n2267 & n2279 ) | ( n2276 & n2279 ) ;
  assign n2281 = n2276 | n2279 ;
  assign n2282 = ( ~n2278 & n2280 ) | ( ~n2278 & n2281 ) | ( n2280 & n2281 ) ;
  assign n2283 = n2267 | n2279 ;
  assign n2284 = n2278 & ~n2283 ;
  assign n2285 = ( ~n2279 & n2282 ) | ( ~n2279 & n2284 ) | ( n2282 & n2284 ) ;
  assign n2286 = ( ~n2277 & n2282 ) | ( ~n2277 & n2285 ) | ( n2282 & n2285 ) ;
  assign n2287 = n2266 & n2286 ;
  assign n2288 = n2260 & n2264 ;
  assign n2289 = ( n2195 & n2260 ) | ( n2195 & n2288 ) | ( n2260 & n2288 ) ;
  assign n2290 = n2287 | n2289 ;
  assign n2291 = n2267 & ~n2279 ;
  assign n2292 = ( n2278 & n2279 ) | ( n2278 & ~n2291 ) | ( n2279 & ~n2291 ) ;
  assign n2293 = n2276 & n2292 ;
  assign n2294 = ~n2244 & n2254 ;
  assign n2295 = ( ~n2253 & n2254 ) | ( ~n2253 & n2294 ) | ( n2254 & n2294 ) ;
  assign n2296 = ~n2226 & n2227 ;
  assign n2297 = ( ~n2223 & n2227 ) | ( ~n2223 & n2296 ) | ( n2227 & n2296 ) ;
  assign n2298 = ~n2295 & n2297 ;
  assign n2299 = n2295 & ~n2297 ;
  assign n2300 = n2298 | n2299 ;
  assign n2301 = n2274 | n2300 ;
  assign n2302 = n2293 | n2301 ;
  assign n2303 = n2274 & n2300 ;
  assign n2304 = ( n2293 & n2300 ) | ( n2293 & n2303 ) | ( n2300 & n2303 ) ;
  assign n2305 = n2302 & ~n2304 ;
  assign n2306 = n2156 & n2194 ;
  assign n2307 = ~n2153 & n2154 ;
  assign n2308 = ( ~n2150 & n2154 ) | ( ~n2150 & n2307 ) | ( n2154 & n2307 ) ;
  assign n2309 = ~n2172 & n2176 ;
  assign n2310 = ( n2176 & ~n2184 ) | ( n2176 & n2309 ) | ( ~n2184 & n2309 ) ;
  assign n2311 = ~n2308 & n2310 ;
  assign n2312 = n2308 & ~n2310 ;
  assign n2313 = n2311 | n2312 ;
  assign n2314 = n2189 | n2313 ;
  assign n2315 = n2306 | n2314 ;
  assign n2316 = n2189 & n2313 ;
  assign n2317 = ( n2306 & n2313 ) | ( n2306 & n2316 ) | ( n2313 & n2316 ) ;
  assign n2318 = n2315 & ~n2317 ;
  assign n2319 = n2305 | n2318 ;
  assign n2320 = n2290 & n2319 ;
  assign n2321 = n2302 & n2315 ;
  assign n2322 = n2304 | n2317 ;
  assign n2323 = n2321 & ~n2322 ;
  assign n2324 = ( n2189 & n2308 ) | ( n2189 & n2310 ) | ( n2308 & n2310 ) ;
  assign n2325 = n2308 | n2310 ;
  assign n2326 = ( n2306 & n2324 ) | ( n2306 & n2325 ) | ( n2324 & n2325 ) ;
  assign n2327 = ( n2274 & n2295 ) | ( n2274 & n2297 ) | ( n2295 & n2297 ) ;
  assign n2328 = n2295 | n2297 ;
  assign n2329 = ( n2293 & n2327 ) | ( n2293 & n2328 ) | ( n2327 & n2328 ) ;
  assign n2330 = ~n2326 & n2329 ;
  assign n2331 = n2326 & ~n2329 ;
  assign n2332 = n2330 | n2331 ;
  assign n2333 = n2323 | n2332 ;
  assign n2334 = n2320 | n2333 ;
  assign n2335 = n2319 | n2323 ;
  assign n2336 = ( n2290 & n2323 ) | ( n2290 & n2335 ) | ( n2323 & n2335 ) ;
  assign n2337 = n2332 & n2336 ;
  assign n2338 = n2334 & ~n2337 ;
  assign n2339 = n2129 | n2338 ;
  assign n2340 = n2057 & ~n2080 ;
  assign n2341 = n2077 & ~n2340 ;
  assign n2342 = n1993 & ~n2050 ;
  assign n2343 = ~n1993 & n2050 ;
  assign n2344 = n2342 | n2343 ;
  assign n2345 = n2202 & ~n2259 ;
  assign n2346 = ~n2202 & n2259 ;
  assign n2347 = n2345 | n2346 ;
  assign n2348 = n2344 & n2347 ;
  assign n2349 = ~n2051 & n2057 ;
  assign n2350 = n2057 & ~n2077 ;
  assign n2351 = n1986 | n2055 ;
  assign n2352 = n2077 | n2351 ;
  assign n2353 = ( n2349 & n2350 ) | ( n2349 & ~n2352 ) | ( n2350 & ~n2352 ) ;
  assign n2354 = n2348 | n2353 ;
  assign n2355 = n2341 | n2354 ;
  assign n2356 = n2195 | n2264 ;
  assign n2357 = ( n2260 & n2286 ) | ( n2260 & ~n2356 ) | ( n2286 & ~n2356 ) ;
  assign n2358 = ( ~n2286 & n2356 ) | ( ~n2286 & n2357 ) | ( n2356 & n2357 ) ;
  assign n2359 = ( ~n2260 & n2357 ) | ( ~n2260 & n2358 ) | ( n2357 & n2358 ) ;
  assign n2360 = n2355 & n2359 ;
  assign n2361 = n2341 | n2353 ;
  assign n2362 = n2348 & n2361 ;
  assign n2363 = ( n2289 & ~n2305 ) | ( n2289 & n2318 ) | ( ~n2305 & n2318 ) ;
  assign n2364 = n2305 & ~n2318 ;
  assign n2365 = ( n2287 & n2363 ) | ( n2287 & ~n2364 ) | ( n2363 & ~n2364 ) ;
  assign n2366 = ( ~n2290 & n2305 ) | ( ~n2290 & n2365 ) | ( n2305 & n2365 ) ;
  assign n2367 = ( ~n2318 & n2365 ) | ( ~n2318 & n2366 ) | ( n2365 & n2366 ) ;
  assign n2368 = ( n2080 & ~n2096 ) | ( n2080 & n2109 ) | ( ~n2096 & n2109 ) ;
  assign n2369 = n2096 & ~n2109 ;
  assign n2370 = ( n2078 & n2368 ) | ( n2078 & ~n2369 ) | ( n2368 & ~n2369 ) ;
  assign n2371 = ( ~n2081 & n2096 ) | ( ~n2081 & n2370 ) | ( n2096 & n2370 ) ;
  assign n2372 = ( ~n2109 & n2370 ) | ( ~n2109 & n2371 ) | ( n2370 & n2371 ) ;
  assign n2373 = ( n2362 & n2367 ) | ( n2362 & n2372 ) | ( n2367 & n2372 ) ;
  assign n2374 = n2367 | n2372 ;
  assign n2375 = ( n2360 & n2373 ) | ( n2360 & n2374 ) | ( n2373 & n2374 ) ;
  assign n2376 = n2339 & n2375 ;
  assign n2377 = n2326 & n2329 ;
  assign n2378 = n2326 | n2329 ;
  assign n2379 = n2377 | n2378 ;
  assign n2380 = ( n2336 & n2377 ) | ( n2336 & n2379 ) | ( n2377 & n2379 ) ;
  assign n2381 = n2117 & n2120 ;
  assign n2382 = n2117 | n2120 ;
  assign n2383 = n2381 | n2382 ;
  assign n2384 = ( n2127 & n2381 ) | ( n2127 & n2383 ) | ( n2381 & n2383 ) ;
  assign n2385 = n2380 & n2384 ;
  assign n2386 = n2127 & n2382 ;
  assign n2387 = n2329 | n2381 ;
  assign n2388 = n2326 | n2381 ;
  assign n2389 = ( n2336 & n2387 ) | ( n2336 & n2388 ) | ( n2387 & n2388 ) ;
  assign n2390 = n2386 | n2389 ;
  assign n2391 = n2385 | n2390 ;
  assign n2392 = n2125 & n2334 ;
  assign n2393 = n2128 | n2337 ;
  assign n2394 = n2392 & ~n2393 ;
  assign n2395 = ( n2385 & n2391 ) | ( n2385 & n2394 ) | ( n2391 & n2394 ) ;
  assign n2396 = n2385 | n2391 ;
  assign n2397 = ( n2376 & n2395 ) | ( n2376 & n2396 ) | ( n2395 & n2396 ) ;
  assign n2398 = n1917 & n2397 ;
  assign n2399 = ( n1920 & n2397 ) | ( n1920 & n2398 ) | ( n2397 & n2398 ) ;
  assign n2400 = ~n1919 & n2399 ;
  assign n2401 = n1917 | n1920 ;
  assign n2402 = ~n1919 & n2401 ;
  assign n2403 = n2397 | n2402 ;
  assign n2404 = n2400 | n2403 ;
  assign n2405 = ~n1870 & n1871 ;
  assign n2406 = n1870 & ~n1871 ;
  assign n2407 = n2405 | n2406 ;
  assign n2408 = n1916 | n2407 ;
  assign n2409 = n2376 | n2394 ;
  assign n2410 = n2384 & ~n2385 ;
  assign n2411 = ( n2380 & ~n2385 ) | ( n2380 & n2410 ) | ( ~n2385 & n2410 ) ;
  assign n2412 = n2409 & n2411 ;
  assign n2413 = n2394 | n2411 ;
  assign n2414 = n2376 | n2413 ;
  assign n2415 = ~n2412 & n2414 ;
  assign n2416 = ~n1916 & n2415 ;
  assign n2417 = ( ~n2407 & n2415 ) | ( ~n2407 & n2416 ) | ( n2415 & n2416 ) ;
  assign n2418 = n2408 & n2417 ;
  assign n2419 = n1916 & n2407 ;
  assign n2420 = n2408 & ~n2419 ;
  assign n2421 = n2415 | n2420 ;
  assign n2422 = n1876 & n1915 ;
  assign n2423 = n1915 & ~n2422 ;
  assign n2424 = n1912 & ~n2422 ;
  assign n2425 = n1876 & n1912 ;
  assign n2426 = ( n2423 & n2424 ) | ( n2423 & n2425 ) | ( n2424 & n2425 ) ;
  assign n2427 = ~n1912 & n2422 ;
  assign n2428 = n1876 | n1912 ;
  assign n2429 = ( n2423 & ~n2427 ) | ( n2423 & n2428 ) | ( ~n2427 & n2428 ) ;
  assign n2430 = ~n2426 & n2429 ;
  assign n2431 = ( ~n2129 & n2338 ) | ( ~n2129 & n2375 ) | ( n2338 & n2375 ) ;
  assign n2432 = ( n2129 & ~n2375 ) | ( n2129 & n2431 ) | ( ~n2375 & n2431 ) ;
  assign n2433 = ( ~n2338 & n2431 ) | ( ~n2338 & n2432 ) | ( n2431 & n2432 ) ;
  assign n2434 = n1879 & ~n1882 ;
  assign n2435 = ~n1879 & n1882 ;
  assign n2436 = n2434 | n2435 ;
  assign n2437 = n2344 & ~n2347 ;
  assign n2438 = ~n2344 & n2347 ;
  assign n2439 = n2437 | n2438 ;
  assign n2440 = n2436 & n2439 ;
  assign n2441 = n1883 | n1891 ;
  assign n2442 = ~n1892 & n2441 ;
  assign n2443 = n1899 & ~n2442 ;
  assign n2444 = ~n1883 & n1891 ;
  assign n2445 = n1883 & ~n1891 ;
  assign n2446 = n2444 | n2445 ;
  assign n2447 = ~n1899 & n2446 ;
  assign n2448 = n2443 | n2447 ;
  assign n2449 = n2440 & n2448 ;
  assign n2450 = n1899 & ~n2440 ;
  assign n2451 = ( n2440 & n2446 ) | ( n2440 & ~n2450 ) | ( n2446 & ~n2450 ) ;
  assign n2452 = n2443 | n2451 ;
  assign n2453 = ~n2348 & n2361 ;
  assign n2454 = n2348 & ~n2353 ;
  assign n2455 = ~n2341 & n2454 ;
  assign n2456 = ~n2359 & n2455 ;
  assign n2457 = ( ~n2359 & n2453 ) | ( ~n2359 & n2456 ) | ( n2453 & n2456 ) ;
  assign n2458 = n2360 & ~n2362 ;
  assign n2459 = ( n2359 & n2457 ) | ( n2359 & ~n2458 ) | ( n2457 & ~n2458 ) ;
  assign n2460 = n2452 & n2459 ;
  assign n2461 = n2449 | n2460 ;
  assign n2463 = ( n2362 & ~n2367 ) | ( n2362 & n2372 ) | ( ~n2367 & n2372 ) ;
  assign n2464 = n2367 & ~n2372 ;
  assign n2465 = ( n2360 & n2463 ) | ( n2360 & ~n2464 ) | ( n2463 & ~n2464 ) ;
  assign n2462 = n2360 | n2362 ;
  assign n2466 = ( n2367 & ~n2462 ) | ( n2367 & n2465 ) | ( ~n2462 & n2465 ) ;
  assign n2467 = ( ~n2372 & n2465 ) | ( ~n2372 & n2466 ) | ( n2465 & n2466 ) ;
  assign n2468 = ~n1905 & n1911 ;
  assign n2469 = n1905 & ~n1911 ;
  assign n2470 = n2468 | n2469 ;
  assign n2471 = ~n1902 & n2470 ;
  assign n2472 = ( n1902 & ~n2470 ) | ( n1902 & n2471 ) | ( ~n2470 & n2471 ) ;
  assign n2473 = n2471 | n2472 ;
  assign n2474 = ( n2461 & n2467 ) | ( n2461 & n2473 ) | ( n2467 & n2473 ) ;
  assign n2475 = ( n2430 & n2433 ) | ( n2430 & n2474 ) | ( n2433 & n2474 ) ;
  assign n2476 = n2421 & n2475 ;
  assign n2477 = n2418 | n2476 ;
  assign n2478 = ( n2400 & n2404 ) | ( n2400 & n2477 ) | ( n2404 & n2477 ) ;
  assign n2479 = n1839 | n1849 ;
  assign n2480 = n1412 | n1843 ;
  assign n2481 = n1847 | n2480 ;
  assign n2482 = ( n2479 & n2480 ) | ( n2479 & n2481 ) | ( n2480 & n2481 ) ;
  assign n2483 = n1476 | n2482 ;
  assign n2484 = n1853 | n2483 ;
  assign n2485 = ( n1853 & n1869 ) | ( n1853 & n2484 ) | ( n1869 & n2484 ) ;
  assign n2486 = n1853 | n2484 ;
  assign n2487 = ( n1917 & n2485 ) | ( n1917 & n2486 ) | ( n2485 & n2486 ) ;
  assign n2488 = n2478 & ~n2487 ;
  assign n2492 = ( x886 & x887 ) | ( x886 & x888 ) | ( x887 & x888 ) ;
  assign n2493 = ( x883 & x884 ) | ( x883 & x885 ) | ( x884 & x885 ) ;
  assign n2494 = n2492 & ~n2493 ;
  assign n2495 = ~n2492 & n2493 ;
  assign n2496 = n2494 | n2495 ;
  assign n2497 = ~x883 & x884 ;
  assign n2498 = x883 & ~x884 ;
  assign n2499 = n2497 | n2498 ;
  assign n2500 = ~x885 & n2499 ;
  assign n2501 = x885 & ~n2499 ;
  assign n2502 = n2500 | n2501 ;
  assign n2503 = ~x886 & x887 ;
  assign n2504 = x886 & ~x887 ;
  assign n2505 = n2503 | n2504 ;
  assign n2506 = ~x888 & n2505 ;
  assign n2507 = x888 & ~n2505 ;
  assign n2508 = n2506 | n2507 ;
  assign n2509 = n2502 & n2508 ;
  assign n2510 = n2496 & ~n2509 ;
  assign n2511 = ~n2496 & n2509 ;
  assign n2512 = n2510 | n2511 ;
  assign n2513 = n2502 & ~n2508 ;
  assign n2514 = ~n2502 & n2508 ;
  assign n2515 = n2513 | n2514 ;
  assign n2516 = ( n2492 & n2493 ) | ( n2492 & n2509 ) | ( n2493 & n2509 ) ;
  assign n2517 = n2515 & n2516 ;
  assign n2518 = n2512 & ~n2517 ;
  assign n2519 = n2512 & n2516 ;
  assign n2520 = ~x889 & x890 ;
  assign n2521 = x889 & ~x890 ;
  assign n2522 = n2520 | n2521 ;
  assign n2523 = ~x891 & n2522 ;
  assign n2524 = x891 & ~n2522 ;
  assign n2525 = n2523 | n2524 ;
  assign n2526 = ~x892 & x893 ;
  assign n2527 = x892 & ~x893 ;
  assign n2528 = n2526 | n2527 ;
  assign n2529 = ~x894 & n2528 ;
  assign n2530 = x894 & ~n2528 ;
  assign n2531 = n2529 | n2530 ;
  assign n2532 = n2525 & ~n2531 ;
  assign n2533 = ~n2525 & n2531 ;
  assign n2534 = n2532 | n2533 ;
  assign n2535 = ( x892 & x893 ) | ( x892 & x894 ) | ( x893 & x894 ) ;
  assign n2536 = ( x889 & x890 ) | ( x889 & x891 ) | ( x890 & x891 ) ;
  assign n2537 = n2525 & n2531 ;
  assign n2538 = ( n2535 & n2536 ) | ( n2535 & n2537 ) | ( n2536 & n2537 ) ;
  assign n2539 = n2534 & n2538 ;
  assign n2540 = n2519 | n2539 ;
  assign n2541 = n2535 & ~n2536 ;
  assign n2542 = ~n2535 & n2536 ;
  assign n2543 = n2541 | n2542 ;
  assign n2544 = ~n2537 & n2543 ;
  assign n2545 = n2537 & ~n2543 ;
  assign n2546 = n2544 | n2545 ;
  assign n2547 = n2538 & n2546 ;
  assign n2548 = n2515 & n2534 ;
  assign n2549 = n2546 & n2548 ;
  assign n2550 = ~n2547 & n2549 ;
  assign n2551 = ~n2540 & n2550 ;
  assign n2552 = n2518 & n2551 ;
  assign n2553 = ~n2547 & n2548 ;
  assign n2554 = ~n2539 & n2546 ;
  assign n2555 = n2519 & ~n2554 ;
  assign n2556 = ( n2553 & n2554 ) | ( n2553 & ~n2555 ) | ( n2554 & ~n2555 ) ;
  assign n2557 = ( n2518 & n2552 ) | ( n2518 & ~n2556 ) | ( n2552 & ~n2556 ) ;
  assign n2558 = n2534 & ~n2538 ;
  assign n2559 = ( n2534 & ~n2546 ) | ( n2534 & n2558 ) | ( ~n2546 & n2558 ) ;
  assign n2560 = n2515 & ~n2516 ;
  assign n2561 = ( ~n2512 & n2515 ) | ( ~n2512 & n2560 ) | ( n2515 & n2560 ) ;
  assign n2562 = ~n2559 & n2561 ;
  assign n2563 = n2559 & ~n2561 ;
  assign n2564 = n2562 | n2563 ;
  assign n2565 = ( x880 & x881 ) | ( x880 & x882 ) | ( x881 & x882 ) ;
  assign n2566 = ( x877 & x878 ) | ( x877 & x879 ) | ( x878 & x879 ) ;
  assign n2567 = n2565 & ~n2566 ;
  assign n2568 = ~n2565 & n2566 ;
  assign n2569 = n2567 | n2568 ;
  assign n2570 = ~x877 & x878 ;
  assign n2571 = x877 & ~x878 ;
  assign n2572 = n2570 | n2571 ;
  assign n2573 = ~x879 & n2572 ;
  assign n2574 = x879 & ~n2572 ;
  assign n2575 = n2573 | n2574 ;
  assign n2576 = ~x880 & x881 ;
  assign n2577 = x880 & ~x881 ;
  assign n2578 = n2576 | n2577 ;
  assign n2579 = ~x882 & n2578 ;
  assign n2580 = x882 & ~n2578 ;
  assign n2581 = n2579 | n2580 ;
  assign n2582 = n2575 & n2581 ;
  assign n2583 = n2569 & ~n2582 ;
  assign n2584 = ~n2569 & n2582 ;
  assign n2585 = n2583 | n2584 ;
  assign n2586 = n2575 & ~n2581 ;
  assign n2587 = ~n2575 & n2581 ;
  assign n2588 = n2586 | n2587 ;
  assign n2589 = ( n2565 & n2566 ) | ( n2565 & n2582 ) | ( n2566 & n2582 ) ;
  assign n2590 = n2588 & ~n2589 ;
  assign n2591 = ( ~n2585 & n2588 ) | ( ~n2585 & n2590 ) | ( n2588 & n2590 ) ;
  assign n2592 = ~x871 & x872 ;
  assign n2593 = x871 & ~x872 ;
  assign n2594 = n2592 | n2593 ;
  assign n2595 = ~x873 & n2594 ;
  assign n2596 = x873 & ~n2594 ;
  assign n2597 = n2595 | n2596 ;
  assign n2598 = ~x874 & x875 ;
  assign n2599 = x874 & ~x875 ;
  assign n2600 = n2598 | n2599 ;
  assign n2601 = ~x876 & n2600 ;
  assign n2602 = x876 & ~n2600 ;
  assign n2603 = n2601 | n2602 ;
  assign n2604 = n2597 & ~n2603 ;
  assign n2605 = ~n2597 & n2603 ;
  assign n2606 = n2604 | n2605 ;
  assign n2607 = ( x874 & x875 ) | ( x874 & x876 ) | ( x875 & x876 ) ;
  assign n2608 = ( x871 & x872 ) | ( x871 & x873 ) | ( x872 & x873 ) ;
  assign n2609 = n2607 & ~n2608 ;
  assign n2610 = ~n2607 & n2608 ;
  assign n2611 = n2609 | n2610 ;
  assign n2612 = n2597 & n2603 ;
  assign n2613 = n2611 & ~n2612 ;
  assign n2614 = ~n2611 & n2612 ;
  assign n2615 = n2613 | n2614 ;
  assign n2616 = ( n2607 & n2608 ) | ( n2607 & n2612 ) | ( n2608 & n2612 ) ;
  assign n2617 = n2606 & ~n2616 ;
  assign n2618 = ( n2606 & ~n2615 ) | ( n2606 & n2617 ) | ( ~n2615 & n2617 ) ;
  assign n2619 = ~n2591 & n2618 ;
  assign n2620 = n2591 & ~n2618 ;
  assign n2621 = n2619 | n2620 ;
  assign n2622 = n2564 & n2621 ;
  assign n2623 = ( n2518 & ~n2519 ) | ( n2518 & n2554 ) | ( ~n2519 & n2554 ) ;
  assign n2624 = n2518 & n2554 ;
  assign n2625 = ( n2553 & n2623 ) | ( n2553 & n2624 ) | ( n2623 & n2624 ) ;
  assign n2626 = n2556 & ~n2625 ;
  assign n2627 = n2622 | n2626 ;
  assign n2628 = n2557 | n2627 ;
  assign n2629 = n2615 & n2616 ;
  assign n2630 = n2588 & n2589 ;
  assign n2631 = n2629 | n2630 ;
  assign n2632 = n2585 & n2589 ;
  assign n2633 = n2588 & n2606 ;
  assign n2634 = n2585 & n2633 ;
  assign n2635 = ~n2632 & n2634 ;
  assign n2636 = ~n2631 & n2635 ;
  assign n2637 = n2606 & n2616 ;
  assign n2638 = n2615 & ~n2637 ;
  assign n2639 = ~n2636 & n2638 ;
  assign n2640 = ~n2632 & n2633 ;
  assign n2641 = n2585 & ~n2630 ;
  assign n2642 = ( n2629 & n2638 ) | ( n2629 & n2641 ) | ( n2638 & n2641 ) ;
  assign n2643 = n2638 | n2641 ;
  assign n2644 = ( ~n2640 & n2642 ) | ( ~n2640 & n2643 ) | ( n2642 & n2643 ) ;
  assign n2645 = n2629 | n2641 ;
  assign n2646 = n2640 & ~n2645 ;
  assign n2647 = ( ~n2641 & n2644 ) | ( ~n2641 & n2646 ) | ( n2644 & n2646 ) ;
  assign n2648 = ( ~n2639 & n2644 ) | ( ~n2639 & n2647 ) | ( n2644 & n2647 ) ;
  assign n2649 = n2628 & n2648 ;
  assign n2650 = n2622 & n2626 ;
  assign n2651 = ( n2557 & n2622 ) | ( n2557 & n2650 ) | ( n2622 & n2650 ) ;
  assign n2652 = n2649 | n2651 ;
  assign n2653 = n2629 & ~n2641 ;
  assign n2654 = ( n2640 & n2641 ) | ( n2640 & ~n2653 ) | ( n2641 & ~n2653 ) ;
  assign n2655 = n2638 & n2654 ;
  assign n2656 = ~n2606 & n2616 ;
  assign n2657 = ( ~n2615 & n2616 ) | ( ~n2615 & n2656 ) | ( n2616 & n2656 ) ;
  assign n2658 = ~n2588 & n2589 ;
  assign n2659 = ( ~n2585 & n2589 ) | ( ~n2585 & n2658 ) | ( n2589 & n2658 ) ;
  assign n2660 = ~n2657 & n2659 ;
  assign n2661 = n2657 & ~n2659 ;
  assign n2662 = n2660 | n2661 ;
  assign n2663 = n2636 | n2662 ;
  assign n2664 = n2655 | n2663 ;
  assign n2665 = n2636 & n2662 ;
  assign n2666 = ( n2655 & n2662 ) | ( n2655 & n2665 ) | ( n2662 & n2665 ) ;
  assign n2667 = n2664 & ~n2666 ;
  assign n2668 = n2518 & n2556 ;
  assign n2669 = ~n2515 & n2516 ;
  assign n2670 = ( ~n2512 & n2516 ) | ( ~n2512 & n2669 ) | ( n2516 & n2669 ) ;
  assign n2671 = ~n2534 & n2538 ;
  assign n2672 = ( n2538 & ~n2546 ) | ( n2538 & n2671 ) | ( ~n2546 & n2671 ) ;
  assign n2673 = ~n2670 & n2672 ;
  assign n2674 = n2670 & ~n2672 ;
  assign n2675 = n2673 | n2674 ;
  assign n2676 = n2551 | n2675 ;
  assign n2677 = n2668 | n2676 ;
  assign n2678 = n2551 & n2675 ;
  assign n2679 = ( n2668 & n2675 ) | ( n2668 & n2678 ) | ( n2675 & n2678 ) ;
  assign n2680 = n2677 & ~n2679 ;
  assign n2681 = n2667 | n2680 ;
  assign n2682 = n2652 & n2681 ;
  assign n2683 = n2664 & n2677 ;
  assign n2684 = n2666 | n2679 ;
  assign n2685 = n2683 & ~n2684 ;
  assign n2686 = ( n2551 & n2670 ) | ( n2551 & n2672 ) | ( n2670 & n2672 ) ;
  assign n2687 = n2670 | n2672 ;
  assign n2688 = ( n2668 & n2686 ) | ( n2668 & n2687 ) | ( n2686 & n2687 ) ;
  assign n2689 = ( n2636 & n2657 ) | ( n2636 & n2659 ) | ( n2657 & n2659 ) ;
  assign n2690 = n2657 | n2659 ;
  assign n2691 = ( n2655 & n2689 ) | ( n2655 & n2690 ) | ( n2689 & n2690 ) ;
  assign n2692 = ~n2688 & n2691 ;
  assign n2693 = n2688 & ~n2691 ;
  assign n2694 = n2692 | n2693 ;
  assign n2695 = n2685 | n2694 ;
  assign n2696 = n2682 | n2695 ;
  assign n2697 = n2681 | n2685 ;
  assign n2698 = ( n2652 & n2685 ) | ( n2652 & n2697 ) | ( n2685 & n2697 ) ;
  assign n2699 = n2694 & n2698 ;
  assign n2700 = n2696 & ~n2699 ;
  assign n2701 = ( x862 & x863 ) | ( x862 & x864 ) | ( x863 & x864 ) ;
  assign n2702 = ( x859 & x860 ) | ( x859 & x861 ) | ( x860 & x861 ) ;
  assign n2703 = n2701 & ~n2702 ;
  assign n2704 = ~n2701 & n2702 ;
  assign n2705 = n2703 | n2704 ;
  assign n2706 = ~x859 & x860 ;
  assign n2707 = x859 & ~x860 ;
  assign n2708 = n2706 | n2707 ;
  assign n2709 = ~x861 & n2708 ;
  assign n2710 = x861 & ~n2708 ;
  assign n2711 = n2709 | n2710 ;
  assign n2712 = ~x862 & x863 ;
  assign n2713 = x862 & ~x863 ;
  assign n2714 = n2712 | n2713 ;
  assign n2715 = ~x864 & n2714 ;
  assign n2716 = x864 & ~n2714 ;
  assign n2717 = n2715 | n2716 ;
  assign n2718 = n2711 & n2717 ;
  assign n2719 = n2705 & ~n2718 ;
  assign n2720 = ~n2705 & n2718 ;
  assign n2721 = n2719 | n2720 ;
  assign n2722 = n2711 & ~n2717 ;
  assign n2723 = ~n2711 & n2717 ;
  assign n2724 = n2722 | n2723 ;
  assign n2725 = ( n2701 & n2702 ) | ( n2701 & n2718 ) | ( n2702 & n2718 ) ;
  assign n2726 = n2724 & n2725 ;
  assign n2727 = n2721 & ~n2726 ;
  assign n2728 = n2721 & n2725 ;
  assign n2729 = ~x865 & x866 ;
  assign n2730 = x865 & ~x866 ;
  assign n2731 = n2729 | n2730 ;
  assign n2732 = ~x867 & n2731 ;
  assign n2733 = x867 & ~n2731 ;
  assign n2734 = n2732 | n2733 ;
  assign n2735 = ~x868 & x869 ;
  assign n2736 = x868 & ~x869 ;
  assign n2737 = n2735 | n2736 ;
  assign n2738 = ~x870 & n2737 ;
  assign n2739 = x870 & ~n2737 ;
  assign n2740 = n2738 | n2739 ;
  assign n2741 = n2734 & ~n2740 ;
  assign n2742 = ~n2734 & n2740 ;
  assign n2743 = n2741 | n2742 ;
  assign n2744 = ( x868 & x869 ) | ( x868 & x870 ) | ( x869 & x870 ) ;
  assign n2745 = ( x865 & x866 ) | ( x865 & x867 ) | ( x866 & x867 ) ;
  assign n2746 = n2734 & n2740 ;
  assign n2747 = ( n2744 & n2745 ) | ( n2744 & n2746 ) | ( n2745 & n2746 ) ;
  assign n2748 = n2743 & n2747 ;
  assign n2749 = n2728 | n2748 ;
  assign n2750 = n2744 & ~n2745 ;
  assign n2751 = ~n2744 & n2745 ;
  assign n2752 = n2750 | n2751 ;
  assign n2753 = ~n2746 & n2752 ;
  assign n2754 = n2746 & ~n2752 ;
  assign n2755 = n2753 | n2754 ;
  assign n2756 = n2747 & n2755 ;
  assign n2757 = n2724 & n2743 ;
  assign n2758 = n2755 & n2757 ;
  assign n2759 = ~n2756 & n2758 ;
  assign n2760 = ~n2749 & n2759 ;
  assign n2761 = n2727 & n2760 ;
  assign n2762 = ~n2756 & n2757 ;
  assign n2763 = ~n2748 & n2755 ;
  assign n2764 = n2728 & ~n2763 ;
  assign n2765 = ( n2762 & n2763 ) | ( n2762 & ~n2764 ) | ( n2763 & ~n2764 ) ;
  assign n2766 = ( n2727 & n2761 ) | ( n2727 & ~n2765 ) | ( n2761 & ~n2765 ) ;
  assign n2767 = n2743 & ~n2747 ;
  assign n2768 = ( n2743 & ~n2755 ) | ( n2743 & n2767 ) | ( ~n2755 & n2767 ) ;
  assign n2769 = n2724 & ~n2725 ;
  assign n2770 = ( ~n2721 & n2724 ) | ( ~n2721 & n2769 ) | ( n2724 & n2769 ) ;
  assign n2771 = ~n2768 & n2770 ;
  assign n2772 = n2768 & ~n2770 ;
  assign n2773 = n2771 | n2772 ;
  assign n2774 = ( x856 & x857 ) | ( x856 & x858 ) | ( x857 & x858 ) ;
  assign n2775 = ( x853 & x854 ) | ( x853 & x855 ) | ( x854 & x855 ) ;
  assign n2776 = n2774 & ~n2775 ;
  assign n2777 = ~n2774 & n2775 ;
  assign n2778 = n2776 | n2777 ;
  assign n2779 = ~x853 & x854 ;
  assign n2780 = x853 & ~x854 ;
  assign n2781 = n2779 | n2780 ;
  assign n2782 = ~x855 & n2781 ;
  assign n2783 = x855 & ~n2781 ;
  assign n2784 = n2782 | n2783 ;
  assign n2785 = ~x856 & x857 ;
  assign n2786 = x856 & ~x857 ;
  assign n2787 = n2785 | n2786 ;
  assign n2788 = ~x858 & n2787 ;
  assign n2789 = x858 & ~n2787 ;
  assign n2790 = n2788 | n2789 ;
  assign n2791 = n2784 & n2790 ;
  assign n2792 = n2778 & ~n2791 ;
  assign n2793 = ~n2778 & n2791 ;
  assign n2794 = n2792 | n2793 ;
  assign n2795 = n2784 & ~n2790 ;
  assign n2796 = ~n2784 & n2790 ;
  assign n2797 = n2795 | n2796 ;
  assign n2798 = ( n2774 & n2775 ) | ( n2774 & n2791 ) | ( n2775 & n2791 ) ;
  assign n2799 = n2797 & ~n2798 ;
  assign n2800 = ( ~n2794 & n2797 ) | ( ~n2794 & n2799 ) | ( n2797 & n2799 ) ;
  assign n2801 = ~x847 & x848 ;
  assign n2802 = x847 & ~x848 ;
  assign n2803 = n2801 | n2802 ;
  assign n2804 = ~x849 & n2803 ;
  assign n2805 = x849 & ~n2803 ;
  assign n2806 = n2804 | n2805 ;
  assign n2807 = ~x850 & x851 ;
  assign n2808 = x850 & ~x851 ;
  assign n2809 = n2807 | n2808 ;
  assign n2810 = ~x852 & n2809 ;
  assign n2811 = x852 & ~n2809 ;
  assign n2812 = n2810 | n2811 ;
  assign n2813 = n2806 & ~n2812 ;
  assign n2814 = ~n2806 & n2812 ;
  assign n2815 = n2813 | n2814 ;
  assign n2816 = ( x850 & x851 ) | ( x850 & x852 ) | ( x851 & x852 ) ;
  assign n2817 = ( x847 & x848 ) | ( x847 & x849 ) | ( x848 & x849 ) ;
  assign n2818 = n2816 & ~n2817 ;
  assign n2819 = ~n2816 & n2817 ;
  assign n2820 = n2818 | n2819 ;
  assign n2821 = n2806 & n2812 ;
  assign n2822 = n2820 & ~n2821 ;
  assign n2823 = ~n2820 & n2821 ;
  assign n2824 = n2822 | n2823 ;
  assign n2825 = ( n2816 & n2817 ) | ( n2816 & n2821 ) | ( n2817 & n2821 ) ;
  assign n2826 = n2815 & ~n2825 ;
  assign n2827 = ( n2815 & ~n2824 ) | ( n2815 & n2826 ) | ( ~n2824 & n2826 ) ;
  assign n2828 = ~n2800 & n2827 ;
  assign n2829 = n2800 & ~n2827 ;
  assign n2830 = n2828 | n2829 ;
  assign n2831 = n2773 & n2830 ;
  assign n2832 = ( n2727 & ~n2728 ) | ( n2727 & n2763 ) | ( ~n2728 & n2763 ) ;
  assign n2833 = n2727 & n2763 ;
  assign n2834 = ( n2762 & n2832 ) | ( n2762 & n2833 ) | ( n2832 & n2833 ) ;
  assign n2835 = n2765 & ~n2834 ;
  assign n2836 = n2831 | n2835 ;
  assign n2837 = n2766 | n2836 ;
  assign n2838 = n2824 & n2825 ;
  assign n2839 = n2797 & n2798 ;
  assign n2840 = n2838 | n2839 ;
  assign n2841 = n2794 & n2798 ;
  assign n2842 = n2797 & n2815 ;
  assign n2843 = n2794 & n2842 ;
  assign n2844 = ~n2841 & n2843 ;
  assign n2845 = ~n2840 & n2844 ;
  assign n2846 = n2815 & n2825 ;
  assign n2847 = n2824 & ~n2846 ;
  assign n2848 = ~n2845 & n2847 ;
  assign n2849 = ~n2841 & n2842 ;
  assign n2850 = n2794 & ~n2839 ;
  assign n2851 = ( n2838 & n2847 ) | ( n2838 & n2850 ) | ( n2847 & n2850 ) ;
  assign n2852 = n2847 | n2850 ;
  assign n2853 = ( ~n2849 & n2851 ) | ( ~n2849 & n2852 ) | ( n2851 & n2852 ) ;
  assign n2854 = n2838 | n2850 ;
  assign n2855 = n2849 & ~n2854 ;
  assign n2856 = ( ~n2850 & n2853 ) | ( ~n2850 & n2855 ) | ( n2853 & n2855 ) ;
  assign n2857 = ( ~n2848 & n2853 ) | ( ~n2848 & n2856 ) | ( n2853 & n2856 ) ;
  assign n2858 = n2837 & n2857 ;
  assign n2859 = n2831 & n2835 ;
  assign n2860 = ( n2766 & n2831 ) | ( n2766 & n2859 ) | ( n2831 & n2859 ) ;
  assign n2861 = n2858 | n2860 ;
  assign n2862 = n2838 & ~n2850 ;
  assign n2863 = ( n2849 & n2850 ) | ( n2849 & ~n2862 ) | ( n2850 & ~n2862 ) ;
  assign n2864 = n2847 & n2863 ;
  assign n2865 = ~n2815 & n2825 ;
  assign n2866 = ( ~n2824 & n2825 ) | ( ~n2824 & n2865 ) | ( n2825 & n2865 ) ;
  assign n2867 = ~n2797 & n2798 ;
  assign n2868 = ( ~n2794 & n2798 ) | ( ~n2794 & n2867 ) | ( n2798 & n2867 ) ;
  assign n2869 = ~n2866 & n2868 ;
  assign n2870 = n2866 & ~n2868 ;
  assign n2871 = n2869 | n2870 ;
  assign n2872 = n2845 | n2871 ;
  assign n2873 = n2864 | n2872 ;
  assign n2874 = n2845 & n2871 ;
  assign n2875 = ( n2864 & n2871 ) | ( n2864 & n2874 ) | ( n2871 & n2874 ) ;
  assign n2876 = n2873 & ~n2875 ;
  assign n2877 = n2727 & n2765 ;
  assign n2878 = ~n2724 & n2725 ;
  assign n2879 = ( ~n2721 & n2725 ) | ( ~n2721 & n2878 ) | ( n2725 & n2878 ) ;
  assign n2880 = ~n2743 & n2747 ;
  assign n2881 = ( n2747 & ~n2755 ) | ( n2747 & n2880 ) | ( ~n2755 & n2880 ) ;
  assign n2882 = ~n2879 & n2881 ;
  assign n2883 = n2879 & ~n2881 ;
  assign n2884 = n2882 | n2883 ;
  assign n2885 = n2760 | n2884 ;
  assign n2886 = n2877 | n2885 ;
  assign n2887 = n2760 & n2884 ;
  assign n2888 = ( n2877 & n2884 ) | ( n2877 & n2887 ) | ( n2884 & n2887 ) ;
  assign n2889 = n2886 & ~n2888 ;
  assign n2890 = n2876 | n2889 ;
  assign n2891 = n2861 & n2890 ;
  assign n2892 = n2873 & n2886 ;
  assign n2893 = n2875 | n2888 ;
  assign n2894 = n2892 & ~n2893 ;
  assign n2895 = ( n2760 & n2879 ) | ( n2760 & n2881 ) | ( n2879 & n2881 ) ;
  assign n2896 = n2879 | n2881 ;
  assign n2897 = ( n2877 & n2895 ) | ( n2877 & n2896 ) | ( n2895 & n2896 ) ;
  assign n2898 = ( n2845 & n2866 ) | ( n2845 & n2868 ) | ( n2866 & n2868 ) ;
  assign n2899 = n2866 | n2868 ;
  assign n2900 = ( n2864 & n2898 ) | ( n2864 & n2899 ) | ( n2898 & n2899 ) ;
  assign n2901 = ~n2897 & n2900 ;
  assign n2902 = n2897 & ~n2900 ;
  assign n2903 = n2901 | n2902 ;
  assign n2904 = n2894 | n2903 ;
  assign n2905 = n2891 | n2904 ;
  assign n2906 = n2890 | n2894 ;
  assign n2907 = ( n2861 & n2894 ) | ( n2861 & n2906 ) | ( n2894 & n2906 ) ;
  assign n2908 = n2903 & n2907 ;
  assign n2909 = n2905 & ~n2908 ;
  assign n2910 = n2700 | n2909 ;
  assign n2911 = n2628 & ~n2651 ;
  assign n2912 = n2648 & ~n2911 ;
  assign n2913 = n2564 & ~n2621 ;
  assign n2914 = ~n2564 & n2621 ;
  assign n2915 = n2913 | n2914 ;
  assign n2916 = n2773 & ~n2830 ;
  assign n2917 = ~n2773 & n2830 ;
  assign n2918 = n2916 | n2917 ;
  assign n2919 = n2915 & n2918 ;
  assign n2920 = ~n2622 & n2628 ;
  assign n2921 = n2628 & ~n2648 ;
  assign n2922 = n2557 | n2626 ;
  assign n2923 = n2648 | n2922 ;
  assign n2924 = ( n2920 & n2921 ) | ( n2920 & ~n2923 ) | ( n2921 & ~n2923 ) ;
  assign n2925 = n2919 | n2924 ;
  assign n2926 = n2912 | n2925 ;
  assign n2927 = n2766 | n2835 ;
  assign n2928 = ( n2831 & n2857 ) | ( n2831 & ~n2927 ) | ( n2857 & ~n2927 ) ;
  assign n2929 = ( ~n2857 & n2927 ) | ( ~n2857 & n2928 ) | ( n2927 & n2928 ) ;
  assign n2930 = ( ~n2831 & n2928 ) | ( ~n2831 & n2929 ) | ( n2928 & n2929 ) ;
  assign n2931 = n2926 & n2930 ;
  assign n2932 = n2912 | n2924 ;
  assign n2933 = n2919 & n2932 ;
  assign n2934 = ( n2860 & ~n2876 ) | ( n2860 & n2889 ) | ( ~n2876 & n2889 ) ;
  assign n2935 = n2876 & ~n2889 ;
  assign n2936 = ( n2858 & n2934 ) | ( n2858 & ~n2935 ) | ( n2934 & ~n2935 ) ;
  assign n2937 = ( ~n2861 & n2876 ) | ( ~n2861 & n2936 ) | ( n2876 & n2936 ) ;
  assign n2938 = ( ~n2889 & n2936 ) | ( ~n2889 & n2937 ) | ( n2936 & n2937 ) ;
  assign n2939 = ( n2651 & ~n2667 ) | ( n2651 & n2680 ) | ( ~n2667 & n2680 ) ;
  assign n2940 = n2667 & ~n2680 ;
  assign n2941 = ( n2649 & n2939 ) | ( n2649 & ~n2940 ) | ( n2939 & ~n2940 ) ;
  assign n2942 = ( ~n2652 & n2667 ) | ( ~n2652 & n2941 ) | ( n2667 & n2941 ) ;
  assign n2943 = ( ~n2680 & n2941 ) | ( ~n2680 & n2942 ) | ( n2941 & n2942 ) ;
  assign n2944 = ( n2933 & n2938 ) | ( n2933 & n2943 ) | ( n2938 & n2943 ) ;
  assign n2945 = n2938 | n2943 ;
  assign n2946 = ( n2931 & n2944 ) | ( n2931 & n2945 ) | ( n2944 & n2945 ) ;
  assign n2947 = n2910 & n2946 ;
  assign n2948 = n2696 & n2905 ;
  assign n2949 = n2699 | n2908 ;
  assign n2950 = n2948 & ~n2949 ;
  assign n2951 = n2897 & n2900 ;
  assign n2952 = n2897 | n2900 ;
  assign n2953 = n2951 | n2952 ;
  assign n2954 = ( n2907 & n2951 ) | ( n2907 & n2953 ) | ( n2951 & n2953 ) ;
  assign n2955 = n2688 & n2691 ;
  assign n2956 = n2688 | n2691 ;
  assign n2957 = n2955 | n2956 ;
  assign n2958 = ( n2698 & n2955 ) | ( n2698 & n2957 ) | ( n2955 & n2957 ) ;
  assign n2959 = n2954 & n2958 ;
  assign n2960 = n2958 & ~n2959 ;
  assign n2961 = ( n2954 & ~n2959 ) | ( n2954 & n2960 ) | ( ~n2959 & n2960 ) ;
  assign n2962 = n2950 | n2961 ;
  assign n2963 = n2947 | n2962 ;
  assign n2964 = n2947 | n2950 ;
  assign n2965 = n2961 & n2964 ;
  assign n2966 = n2963 & ~n2965 ;
  assign n2967 = ( x934 & x935 ) | ( x934 & x936 ) | ( x935 & x936 ) ;
  assign n2968 = ( x931 & x932 ) | ( x931 & x933 ) | ( x932 & x933 ) ;
  assign n2969 = n2967 & ~n2968 ;
  assign n2970 = ~n2967 & n2968 ;
  assign n2971 = n2969 | n2970 ;
  assign n2972 = ~x931 & x932 ;
  assign n2973 = x931 & ~x932 ;
  assign n2974 = n2972 | n2973 ;
  assign n2975 = ~x933 & n2974 ;
  assign n2976 = x933 & ~n2974 ;
  assign n2977 = n2975 | n2976 ;
  assign n2978 = ~x934 & x935 ;
  assign n2979 = x934 & ~x935 ;
  assign n2980 = n2978 | n2979 ;
  assign n2981 = ~x936 & n2980 ;
  assign n2982 = x936 & ~n2980 ;
  assign n2983 = n2981 | n2982 ;
  assign n2984 = n2977 & n2983 ;
  assign n2985 = n2971 & ~n2984 ;
  assign n2986 = ~n2971 & n2984 ;
  assign n2987 = n2985 | n2986 ;
  assign n2988 = n2977 & ~n2983 ;
  assign n2989 = ~n2977 & n2983 ;
  assign n2990 = n2988 | n2989 ;
  assign n2991 = ( n2967 & n2968 ) | ( n2967 & n2984 ) | ( n2968 & n2984 ) ;
  assign n2992 = n2990 & n2991 ;
  assign n2993 = n2987 & ~n2992 ;
  assign n2994 = n2987 & n2991 ;
  assign n2995 = ~x937 & x938 ;
  assign n2996 = x937 & ~x938 ;
  assign n2997 = n2995 | n2996 ;
  assign n2998 = ~x939 & n2997 ;
  assign n2999 = x939 & ~n2997 ;
  assign n3000 = n2998 | n2999 ;
  assign n3001 = ~x940 & x941 ;
  assign n3002 = x940 & ~x941 ;
  assign n3003 = n3001 | n3002 ;
  assign n3004 = ~x942 & n3003 ;
  assign n3005 = x942 & ~n3003 ;
  assign n3006 = n3004 | n3005 ;
  assign n3007 = n3000 & ~n3006 ;
  assign n3008 = ~n3000 & n3006 ;
  assign n3009 = n3007 | n3008 ;
  assign n3010 = ( x940 & x941 ) | ( x940 & x942 ) | ( x941 & x942 ) ;
  assign n3011 = ( x937 & x938 ) | ( x937 & x939 ) | ( x938 & x939 ) ;
  assign n3012 = n3000 & n3006 ;
  assign n3013 = ( n3010 & n3011 ) | ( n3010 & n3012 ) | ( n3011 & n3012 ) ;
  assign n3014 = n3009 & n3013 ;
  assign n3015 = n2994 | n3014 ;
  assign n3016 = n3010 & ~n3011 ;
  assign n3017 = ~n3010 & n3011 ;
  assign n3018 = n3016 | n3017 ;
  assign n3019 = ~n3012 & n3018 ;
  assign n3020 = n3012 & ~n3018 ;
  assign n3021 = n3019 | n3020 ;
  assign n3022 = n3013 & n3021 ;
  assign n3023 = n2990 & n3009 ;
  assign n3024 = n3021 & n3023 ;
  assign n3025 = ~n3022 & n3024 ;
  assign n3026 = ~n3015 & n3025 ;
  assign n3027 = n2993 & n3026 ;
  assign n3028 = ~n3022 & n3023 ;
  assign n3029 = ~n3014 & n3021 ;
  assign n3030 = n2994 & ~n3029 ;
  assign n3031 = ( n3028 & n3029 ) | ( n3028 & ~n3030 ) | ( n3029 & ~n3030 ) ;
  assign n3032 = ( n2993 & n3027 ) | ( n2993 & ~n3031 ) | ( n3027 & ~n3031 ) ;
  assign n3033 = n3009 & ~n3013 ;
  assign n3034 = ( n3009 & ~n3021 ) | ( n3009 & n3033 ) | ( ~n3021 & n3033 ) ;
  assign n3035 = n2990 & ~n2991 ;
  assign n3036 = ( ~n2987 & n2990 ) | ( ~n2987 & n3035 ) | ( n2990 & n3035 ) ;
  assign n3037 = ~n3034 & n3036 ;
  assign n3038 = n3034 & ~n3036 ;
  assign n3039 = n3037 | n3038 ;
  assign n3040 = ( x928 & x929 ) | ( x928 & x930 ) | ( x929 & x930 ) ;
  assign n3041 = ( x925 & x926 ) | ( x925 & x927 ) | ( x926 & x927 ) ;
  assign n3042 = n3040 & ~n3041 ;
  assign n3043 = ~n3040 & n3041 ;
  assign n3044 = n3042 | n3043 ;
  assign n3045 = ~x925 & x926 ;
  assign n3046 = x925 & ~x926 ;
  assign n3047 = n3045 | n3046 ;
  assign n3048 = ~x927 & n3047 ;
  assign n3049 = x927 & ~n3047 ;
  assign n3050 = n3048 | n3049 ;
  assign n3051 = ~x928 & x929 ;
  assign n3052 = x928 & ~x929 ;
  assign n3053 = n3051 | n3052 ;
  assign n3054 = ~x930 & n3053 ;
  assign n3055 = x930 & ~n3053 ;
  assign n3056 = n3054 | n3055 ;
  assign n3057 = n3050 & n3056 ;
  assign n3058 = n3044 & ~n3057 ;
  assign n3059 = ~n3044 & n3057 ;
  assign n3060 = n3058 | n3059 ;
  assign n3061 = n3050 & ~n3056 ;
  assign n3062 = ~n3050 & n3056 ;
  assign n3063 = n3061 | n3062 ;
  assign n3064 = ( n3040 & n3041 ) | ( n3040 & n3057 ) | ( n3041 & n3057 ) ;
  assign n3065 = n3063 & ~n3064 ;
  assign n3066 = ( ~n3060 & n3063 ) | ( ~n3060 & n3065 ) | ( n3063 & n3065 ) ;
  assign n3067 = ~x919 & x920 ;
  assign n3068 = x919 & ~x920 ;
  assign n3069 = n3067 | n3068 ;
  assign n3070 = ~x921 & n3069 ;
  assign n3071 = x921 & ~n3069 ;
  assign n3072 = n3070 | n3071 ;
  assign n3073 = ~x922 & x923 ;
  assign n3074 = x922 & ~x923 ;
  assign n3075 = n3073 | n3074 ;
  assign n3076 = ~x924 & n3075 ;
  assign n3077 = x924 & ~n3075 ;
  assign n3078 = n3076 | n3077 ;
  assign n3079 = n3072 & ~n3078 ;
  assign n3080 = ~n3072 & n3078 ;
  assign n3081 = n3079 | n3080 ;
  assign n3082 = ( x922 & x923 ) | ( x922 & x924 ) | ( x923 & x924 ) ;
  assign n3083 = ( x919 & x920 ) | ( x919 & x921 ) | ( x920 & x921 ) ;
  assign n3084 = n3082 & ~n3083 ;
  assign n3085 = ~n3082 & n3083 ;
  assign n3086 = n3084 | n3085 ;
  assign n3087 = n3072 & n3078 ;
  assign n3088 = n3086 & ~n3087 ;
  assign n3089 = ~n3086 & n3087 ;
  assign n3090 = n3088 | n3089 ;
  assign n3091 = ( n3082 & n3083 ) | ( n3082 & n3087 ) | ( n3083 & n3087 ) ;
  assign n3092 = n3081 & ~n3091 ;
  assign n3093 = ( n3081 & ~n3090 ) | ( n3081 & n3092 ) | ( ~n3090 & n3092 ) ;
  assign n3094 = ~n3066 & n3093 ;
  assign n3095 = n3066 & ~n3093 ;
  assign n3096 = n3094 | n3095 ;
  assign n3097 = n3039 & n3096 ;
  assign n3098 = ( n2993 & ~n2994 ) | ( n2993 & n3029 ) | ( ~n2994 & n3029 ) ;
  assign n3099 = n2993 & n3029 ;
  assign n3100 = ( n3028 & n3098 ) | ( n3028 & n3099 ) | ( n3098 & n3099 ) ;
  assign n3101 = n3031 & ~n3100 ;
  assign n3102 = n3097 | n3101 ;
  assign n3103 = n3032 | n3102 ;
  assign n3104 = n3090 & n3091 ;
  assign n3105 = n3063 & n3064 ;
  assign n3106 = n3104 | n3105 ;
  assign n3107 = n3060 & n3064 ;
  assign n3108 = n3063 & n3081 ;
  assign n3109 = n3060 & n3108 ;
  assign n3110 = ~n3107 & n3109 ;
  assign n3111 = ~n3106 & n3110 ;
  assign n3112 = n3081 & n3091 ;
  assign n3113 = n3090 & ~n3112 ;
  assign n3114 = ~n3111 & n3113 ;
  assign n3115 = ~n3107 & n3108 ;
  assign n3116 = n3060 & ~n3105 ;
  assign n3117 = ( n3104 & n3113 ) | ( n3104 & n3116 ) | ( n3113 & n3116 ) ;
  assign n3118 = n3113 | n3116 ;
  assign n3119 = ( ~n3115 & n3117 ) | ( ~n3115 & n3118 ) | ( n3117 & n3118 ) ;
  assign n3120 = n3104 | n3116 ;
  assign n3121 = n3115 & ~n3120 ;
  assign n3122 = ( ~n3116 & n3119 ) | ( ~n3116 & n3121 ) | ( n3119 & n3121 ) ;
  assign n3123 = ( ~n3114 & n3119 ) | ( ~n3114 & n3122 ) | ( n3119 & n3122 ) ;
  assign n3124 = n3103 & n3123 ;
  assign n3125 = n3097 & n3101 ;
  assign n3126 = ( n3032 & n3097 ) | ( n3032 & n3125 ) | ( n3097 & n3125 ) ;
  assign n3127 = n3124 | n3126 ;
  assign n3128 = n3104 & ~n3116 ;
  assign n3129 = ( n3115 & n3116 ) | ( n3115 & ~n3128 ) | ( n3116 & ~n3128 ) ;
  assign n3130 = n3113 & n3129 ;
  assign n3131 = ~n3081 & n3091 ;
  assign n3132 = ( ~n3090 & n3091 ) | ( ~n3090 & n3131 ) | ( n3091 & n3131 ) ;
  assign n3133 = ~n3063 & n3064 ;
  assign n3134 = ( ~n3060 & n3064 ) | ( ~n3060 & n3133 ) | ( n3064 & n3133 ) ;
  assign n3135 = ~n3132 & n3134 ;
  assign n3136 = n3132 & ~n3134 ;
  assign n3137 = n3135 | n3136 ;
  assign n3138 = n3111 | n3137 ;
  assign n3139 = n3130 | n3138 ;
  assign n3140 = n3111 & n3137 ;
  assign n3141 = ( n3130 & n3137 ) | ( n3130 & n3140 ) | ( n3137 & n3140 ) ;
  assign n3142 = n3139 & ~n3141 ;
  assign n3143 = n2993 & n3031 ;
  assign n3144 = ~n2990 & n2991 ;
  assign n3145 = ( ~n2987 & n2991 ) | ( ~n2987 & n3144 ) | ( n2991 & n3144 ) ;
  assign n3146 = ~n3009 & n3013 ;
  assign n3147 = ( n3013 & ~n3021 ) | ( n3013 & n3146 ) | ( ~n3021 & n3146 ) ;
  assign n3148 = ~n3145 & n3147 ;
  assign n3149 = n3145 & ~n3147 ;
  assign n3150 = n3148 | n3149 ;
  assign n3151 = n3026 | n3150 ;
  assign n3152 = n3143 | n3151 ;
  assign n3153 = n3026 & n3150 ;
  assign n3154 = ( n3143 & n3150 ) | ( n3143 & n3153 ) | ( n3150 & n3153 ) ;
  assign n3155 = n3152 & ~n3154 ;
  assign n3156 = n3142 | n3155 ;
  assign n3157 = n3127 & n3156 ;
  assign n3158 = n3139 & n3152 ;
  assign n3159 = n3141 | n3154 ;
  assign n3160 = n3158 & ~n3159 ;
  assign n3161 = ( n3026 & n3145 ) | ( n3026 & n3147 ) | ( n3145 & n3147 ) ;
  assign n3162 = n3145 | n3147 ;
  assign n3163 = ( n3143 & n3161 ) | ( n3143 & n3162 ) | ( n3161 & n3162 ) ;
  assign n3164 = ( n3111 & n3132 ) | ( n3111 & n3134 ) | ( n3132 & n3134 ) ;
  assign n3165 = n3132 | n3134 ;
  assign n3166 = ( n3130 & n3164 ) | ( n3130 & n3165 ) | ( n3164 & n3165 ) ;
  assign n3167 = ~n3163 & n3166 ;
  assign n3168 = n3163 & ~n3166 ;
  assign n3169 = n3167 | n3168 ;
  assign n3170 = n3160 | n3169 ;
  assign n3171 = n3157 | n3170 ;
  assign n3172 = n3156 | n3160 ;
  assign n3173 = ( n3127 & n3160 ) | ( n3127 & n3172 ) | ( n3160 & n3172 ) ;
  assign n3174 = n3169 & n3173 ;
  assign n3175 = n3171 & ~n3174 ;
  assign n3176 = ( x910 & x911 ) | ( x910 & x912 ) | ( x911 & x912 ) ;
  assign n3177 = ( x907 & x908 ) | ( x907 & x909 ) | ( x908 & x909 ) ;
  assign n3178 = n3176 & ~n3177 ;
  assign n3179 = ~n3176 & n3177 ;
  assign n3180 = n3178 | n3179 ;
  assign n3181 = ~x907 & x908 ;
  assign n3182 = x907 & ~x908 ;
  assign n3183 = n3181 | n3182 ;
  assign n3184 = ~x909 & n3183 ;
  assign n3185 = x909 & ~n3183 ;
  assign n3186 = n3184 | n3185 ;
  assign n3187 = ~x910 & x911 ;
  assign n3188 = x910 & ~x911 ;
  assign n3189 = n3187 | n3188 ;
  assign n3190 = ~x912 & n3189 ;
  assign n3191 = x912 & ~n3189 ;
  assign n3192 = n3190 | n3191 ;
  assign n3193 = n3186 & n3192 ;
  assign n3194 = n3180 & ~n3193 ;
  assign n3195 = ~n3180 & n3193 ;
  assign n3196 = n3194 | n3195 ;
  assign n3197 = n3186 & ~n3192 ;
  assign n3198 = ~n3186 & n3192 ;
  assign n3199 = n3197 | n3198 ;
  assign n3200 = ( n3176 & n3177 ) | ( n3176 & n3193 ) | ( n3177 & n3193 ) ;
  assign n3201 = n3199 & n3200 ;
  assign n3202 = n3196 & ~n3201 ;
  assign n3203 = n3196 & n3200 ;
  assign n3204 = ~x913 & x914 ;
  assign n3205 = x913 & ~x914 ;
  assign n3206 = n3204 | n3205 ;
  assign n3207 = ~x915 & n3206 ;
  assign n3208 = x915 & ~n3206 ;
  assign n3209 = n3207 | n3208 ;
  assign n3210 = ~x916 & x917 ;
  assign n3211 = x916 & ~x917 ;
  assign n3212 = n3210 | n3211 ;
  assign n3213 = ~x918 & n3212 ;
  assign n3214 = x918 & ~n3212 ;
  assign n3215 = n3213 | n3214 ;
  assign n3216 = n3209 & ~n3215 ;
  assign n3217 = ~n3209 & n3215 ;
  assign n3218 = n3216 | n3217 ;
  assign n3219 = ( x916 & x917 ) | ( x916 & x918 ) | ( x917 & x918 ) ;
  assign n3220 = ( x913 & x914 ) | ( x913 & x915 ) | ( x914 & x915 ) ;
  assign n3221 = n3209 & n3215 ;
  assign n3222 = ( n3219 & n3220 ) | ( n3219 & n3221 ) | ( n3220 & n3221 ) ;
  assign n3223 = n3218 & n3222 ;
  assign n3224 = n3203 | n3223 ;
  assign n3225 = n3219 & ~n3220 ;
  assign n3226 = ~n3219 & n3220 ;
  assign n3227 = n3225 | n3226 ;
  assign n3228 = ~n3221 & n3227 ;
  assign n3229 = n3221 & ~n3227 ;
  assign n3230 = n3228 | n3229 ;
  assign n3231 = n3222 & n3230 ;
  assign n3232 = n3199 & n3218 ;
  assign n3233 = n3230 & n3232 ;
  assign n3234 = ~n3231 & n3233 ;
  assign n3235 = ~n3224 & n3234 ;
  assign n3236 = n3202 & n3235 ;
  assign n3237 = ~n3231 & n3232 ;
  assign n3238 = ~n3223 & n3230 ;
  assign n3239 = n3203 & ~n3238 ;
  assign n3240 = ( n3237 & n3238 ) | ( n3237 & ~n3239 ) | ( n3238 & ~n3239 ) ;
  assign n3241 = ( n3202 & n3236 ) | ( n3202 & ~n3240 ) | ( n3236 & ~n3240 ) ;
  assign n3242 = n3218 & ~n3222 ;
  assign n3243 = ( n3218 & ~n3230 ) | ( n3218 & n3242 ) | ( ~n3230 & n3242 ) ;
  assign n3244 = n3199 & ~n3200 ;
  assign n3245 = ( ~n3196 & n3199 ) | ( ~n3196 & n3244 ) | ( n3199 & n3244 ) ;
  assign n3246 = ~n3243 & n3245 ;
  assign n3247 = n3243 & ~n3245 ;
  assign n3248 = n3246 | n3247 ;
  assign n3249 = ( x904 & x905 ) | ( x904 & x906 ) | ( x905 & x906 ) ;
  assign n3250 = ( x901 & x902 ) | ( x901 & x903 ) | ( x902 & x903 ) ;
  assign n3251 = n3249 & ~n3250 ;
  assign n3252 = ~n3249 & n3250 ;
  assign n3253 = n3251 | n3252 ;
  assign n3254 = ~x901 & x902 ;
  assign n3255 = x901 & ~x902 ;
  assign n3256 = n3254 | n3255 ;
  assign n3257 = ~x903 & n3256 ;
  assign n3258 = x903 & ~n3256 ;
  assign n3259 = n3257 | n3258 ;
  assign n3260 = ~x904 & x905 ;
  assign n3261 = x904 & ~x905 ;
  assign n3262 = n3260 | n3261 ;
  assign n3263 = ~x906 & n3262 ;
  assign n3264 = x906 & ~n3262 ;
  assign n3265 = n3263 | n3264 ;
  assign n3266 = n3259 & n3265 ;
  assign n3267 = n3253 & ~n3266 ;
  assign n3268 = ~n3253 & n3266 ;
  assign n3269 = n3267 | n3268 ;
  assign n3270 = n3259 & ~n3265 ;
  assign n3271 = ~n3259 & n3265 ;
  assign n3272 = n3270 | n3271 ;
  assign n3273 = ( n3249 & n3250 ) | ( n3249 & n3266 ) | ( n3250 & n3266 ) ;
  assign n3274 = n3272 & ~n3273 ;
  assign n3275 = ( ~n3269 & n3272 ) | ( ~n3269 & n3274 ) | ( n3272 & n3274 ) ;
  assign n3276 = ~x895 & x896 ;
  assign n3277 = x895 & ~x896 ;
  assign n3278 = n3276 | n3277 ;
  assign n3279 = ~x897 & n3278 ;
  assign n3280 = x897 & ~n3278 ;
  assign n3281 = n3279 | n3280 ;
  assign n3282 = ~x898 & x899 ;
  assign n3283 = x898 & ~x899 ;
  assign n3284 = n3282 | n3283 ;
  assign n3285 = ~x900 & n3284 ;
  assign n3286 = x900 & ~n3284 ;
  assign n3287 = n3285 | n3286 ;
  assign n3288 = n3281 & ~n3287 ;
  assign n3289 = ~n3281 & n3287 ;
  assign n3290 = n3288 | n3289 ;
  assign n3291 = ( x898 & x899 ) | ( x898 & x900 ) | ( x899 & x900 ) ;
  assign n3292 = ( x895 & x896 ) | ( x895 & x897 ) | ( x896 & x897 ) ;
  assign n3293 = n3291 & ~n3292 ;
  assign n3294 = ~n3291 & n3292 ;
  assign n3295 = n3293 | n3294 ;
  assign n3296 = n3281 & n3287 ;
  assign n3297 = n3295 & ~n3296 ;
  assign n3298 = ~n3295 & n3296 ;
  assign n3299 = n3297 | n3298 ;
  assign n3300 = ( n3291 & n3292 ) | ( n3291 & n3296 ) | ( n3292 & n3296 ) ;
  assign n3301 = n3290 & ~n3300 ;
  assign n3302 = ( n3290 & ~n3299 ) | ( n3290 & n3301 ) | ( ~n3299 & n3301 ) ;
  assign n3303 = ~n3275 & n3302 ;
  assign n3304 = n3275 & ~n3302 ;
  assign n3305 = n3303 | n3304 ;
  assign n3306 = n3248 & n3305 ;
  assign n3307 = ( n3202 & ~n3203 ) | ( n3202 & n3238 ) | ( ~n3203 & n3238 ) ;
  assign n3308 = n3202 & n3238 ;
  assign n3309 = ( n3237 & n3307 ) | ( n3237 & n3308 ) | ( n3307 & n3308 ) ;
  assign n3310 = n3240 & ~n3309 ;
  assign n3311 = n3306 | n3310 ;
  assign n3312 = n3241 | n3311 ;
  assign n3313 = n3299 & n3300 ;
  assign n3314 = n3272 & n3273 ;
  assign n3315 = n3313 | n3314 ;
  assign n3316 = n3269 & n3273 ;
  assign n3317 = n3272 & n3290 ;
  assign n3318 = n3269 & n3317 ;
  assign n3319 = ~n3316 & n3318 ;
  assign n3320 = ~n3315 & n3319 ;
  assign n3321 = n3290 & n3300 ;
  assign n3322 = n3299 & ~n3321 ;
  assign n3323 = ~n3320 & n3322 ;
  assign n3324 = ~n3316 & n3317 ;
  assign n3325 = n3269 & ~n3314 ;
  assign n3326 = ( n3313 & n3322 ) | ( n3313 & n3325 ) | ( n3322 & n3325 ) ;
  assign n3327 = n3322 | n3325 ;
  assign n3328 = ( ~n3324 & n3326 ) | ( ~n3324 & n3327 ) | ( n3326 & n3327 ) ;
  assign n3329 = n3313 | n3325 ;
  assign n3330 = n3324 & ~n3329 ;
  assign n3331 = ( ~n3325 & n3328 ) | ( ~n3325 & n3330 ) | ( n3328 & n3330 ) ;
  assign n3332 = ( ~n3323 & n3328 ) | ( ~n3323 & n3331 ) | ( n3328 & n3331 ) ;
  assign n3333 = n3312 & n3332 ;
  assign n3334 = n3306 & n3310 ;
  assign n3335 = ( n3241 & n3306 ) | ( n3241 & n3334 ) | ( n3306 & n3334 ) ;
  assign n3336 = n3333 | n3335 ;
  assign n3337 = n3313 & ~n3325 ;
  assign n3338 = ( n3324 & n3325 ) | ( n3324 & ~n3337 ) | ( n3325 & ~n3337 ) ;
  assign n3339 = n3322 & n3338 ;
  assign n3340 = ~n3290 & n3300 ;
  assign n3341 = ( ~n3299 & n3300 ) | ( ~n3299 & n3340 ) | ( n3300 & n3340 ) ;
  assign n3342 = ~n3272 & n3273 ;
  assign n3343 = ( ~n3269 & n3273 ) | ( ~n3269 & n3342 ) | ( n3273 & n3342 ) ;
  assign n3344 = ~n3341 & n3343 ;
  assign n3345 = n3341 & ~n3343 ;
  assign n3346 = n3344 | n3345 ;
  assign n3347 = n3320 | n3346 ;
  assign n3348 = n3339 | n3347 ;
  assign n3349 = n3320 & n3346 ;
  assign n3350 = ( n3339 & n3346 ) | ( n3339 & n3349 ) | ( n3346 & n3349 ) ;
  assign n3351 = n3348 & ~n3350 ;
  assign n3352 = n3202 & n3240 ;
  assign n3353 = ~n3199 & n3200 ;
  assign n3354 = ( ~n3196 & n3200 ) | ( ~n3196 & n3353 ) | ( n3200 & n3353 ) ;
  assign n3355 = ~n3218 & n3222 ;
  assign n3356 = ( n3222 & ~n3230 ) | ( n3222 & n3355 ) | ( ~n3230 & n3355 ) ;
  assign n3357 = ~n3354 & n3356 ;
  assign n3358 = n3354 & ~n3356 ;
  assign n3359 = n3357 | n3358 ;
  assign n3360 = n3235 | n3359 ;
  assign n3361 = n3352 | n3360 ;
  assign n3362 = n3235 & n3359 ;
  assign n3363 = ( n3352 & n3359 ) | ( n3352 & n3362 ) | ( n3359 & n3362 ) ;
  assign n3364 = n3361 & ~n3363 ;
  assign n3365 = n3351 | n3364 ;
  assign n3366 = n3336 & n3365 ;
  assign n3367 = n3348 & n3361 ;
  assign n3368 = n3350 | n3363 ;
  assign n3369 = n3367 & ~n3368 ;
  assign n3370 = ( n3235 & n3354 ) | ( n3235 & n3356 ) | ( n3354 & n3356 ) ;
  assign n3371 = n3354 | n3356 ;
  assign n3372 = ( n3352 & n3370 ) | ( n3352 & n3371 ) | ( n3370 & n3371 ) ;
  assign n3373 = ( n3320 & n3341 ) | ( n3320 & n3343 ) | ( n3341 & n3343 ) ;
  assign n3374 = n3341 | n3343 ;
  assign n3375 = ( n3339 & n3373 ) | ( n3339 & n3374 ) | ( n3373 & n3374 ) ;
  assign n3376 = ~n3372 & n3375 ;
  assign n3377 = n3372 & ~n3375 ;
  assign n3378 = n3376 | n3377 ;
  assign n3379 = n3369 | n3378 ;
  assign n3380 = n3366 | n3379 ;
  assign n3381 = n3365 | n3369 ;
  assign n3382 = ( n3336 & n3369 ) | ( n3336 & n3381 ) | ( n3369 & n3381 ) ;
  assign n3383 = n3378 & n3382 ;
  assign n3384 = n3380 & ~n3383 ;
  assign n3385 = n3175 | n3384 ;
  assign n3386 = n3103 & ~n3126 ;
  assign n3387 = n3123 & ~n3386 ;
  assign n3388 = n3039 & ~n3096 ;
  assign n3389 = ~n3039 & n3096 ;
  assign n3390 = n3388 | n3389 ;
  assign n3391 = n3248 & ~n3305 ;
  assign n3392 = ~n3248 & n3305 ;
  assign n3393 = n3391 | n3392 ;
  assign n3394 = n3390 & n3393 ;
  assign n3395 = ~n3097 & n3103 ;
  assign n3396 = n3103 & ~n3123 ;
  assign n3397 = n3032 | n3101 ;
  assign n3398 = n3123 | n3397 ;
  assign n3399 = ( n3395 & n3396 ) | ( n3395 & ~n3398 ) | ( n3396 & ~n3398 ) ;
  assign n3400 = n3394 | n3399 ;
  assign n3401 = n3387 | n3400 ;
  assign n3402 = n3241 | n3310 ;
  assign n3403 = ( n3306 & n3332 ) | ( n3306 & ~n3402 ) | ( n3332 & ~n3402 ) ;
  assign n3404 = ( ~n3332 & n3402 ) | ( ~n3332 & n3403 ) | ( n3402 & n3403 ) ;
  assign n3405 = ( ~n3306 & n3403 ) | ( ~n3306 & n3404 ) | ( n3403 & n3404 ) ;
  assign n3406 = n3401 & n3405 ;
  assign n3407 = n3387 | n3399 ;
  assign n3408 = n3394 & n3407 ;
  assign n3409 = ( n3335 & ~n3351 ) | ( n3335 & n3364 ) | ( ~n3351 & n3364 ) ;
  assign n3410 = n3351 & ~n3364 ;
  assign n3411 = ( n3333 & n3409 ) | ( n3333 & ~n3410 ) | ( n3409 & ~n3410 ) ;
  assign n3412 = ( ~n3336 & n3351 ) | ( ~n3336 & n3411 ) | ( n3351 & n3411 ) ;
  assign n3413 = ( ~n3364 & n3411 ) | ( ~n3364 & n3412 ) | ( n3411 & n3412 ) ;
  assign n3414 = ( n3126 & ~n3142 ) | ( n3126 & n3155 ) | ( ~n3142 & n3155 ) ;
  assign n3415 = n3142 & ~n3155 ;
  assign n3416 = ( n3124 & n3414 ) | ( n3124 & ~n3415 ) | ( n3414 & ~n3415 ) ;
  assign n3417 = ( ~n3127 & n3142 ) | ( ~n3127 & n3416 ) | ( n3142 & n3416 ) ;
  assign n3418 = ( ~n3155 & n3416 ) | ( ~n3155 & n3417 ) | ( n3416 & n3417 ) ;
  assign n3419 = ( n3408 & n3413 ) | ( n3408 & n3418 ) | ( n3413 & n3418 ) ;
  assign n3420 = n3413 | n3418 ;
  assign n3421 = ( n3406 & n3419 ) | ( n3406 & n3420 ) | ( n3419 & n3420 ) ;
  assign n3422 = n3385 & n3421 ;
  assign n3423 = n3171 & n3380 ;
  assign n3424 = n3174 | n3383 ;
  assign n3425 = n3423 & ~n3424 ;
  assign n3426 = n3372 & n3375 ;
  assign n3427 = n3372 | n3375 ;
  assign n3428 = n3426 | n3427 ;
  assign n3429 = ( n3382 & n3426 ) | ( n3382 & n3428 ) | ( n3426 & n3428 ) ;
  assign n3430 = n3163 & n3166 ;
  assign n3431 = n3163 | n3166 ;
  assign n3432 = n3430 | n3431 ;
  assign n3433 = ( n3173 & n3430 ) | ( n3173 & n3432 ) | ( n3430 & n3432 ) ;
  assign n3434 = n3429 & n3433 ;
  assign n3435 = n3433 & ~n3434 ;
  assign n3436 = ( n3429 & ~n3434 ) | ( n3429 & n3435 ) | ( ~n3434 & n3435 ) ;
  assign n3437 = n3425 | n3436 ;
  assign n3438 = n3422 | n3437 ;
  assign n3439 = n3422 | n3425 ;
  assign n3440 = n3436 & n3439 ;
  assign n3441 = n3438 & ~n3440 ;
  assign n3442 = n2966 | n3441 ;
  assign n3443 = n3390 & ~n3393 ;
  assign n3444 = ~n3390 & n3393 ;
  assign n3445 = n3443 | n3444 ;
  assign n3446 = n2915 & ~n2918 ;
  assign n3447 = ~n2915 & n2918 ;
  assign n3448 = n3446 | n3447 ;
  assign n3449 = n3445 & n3448 ;
  assign n3450 = ~n3401 & n3405 ;
  assign n3451 = ( n3405 & n3408 ) | ( n3405 & n3450 ) | ( n3408 & n3450 ) ;
  assign n3452 = ~n3394 & n3407 ;
  assign n3453 = n3394 & ~n3399 ;
  assign n3454 = ~n3387 & n3453 ;
  assign n3455 = ~n3405 & n3454 ;
  assign n3456 = ( ~n3405 & n3452 ) | ( ~n3405 & n3455 ) | ( n3452 & n3455 ) ;
  assign n3457 = n3451 | n3456 ;
  assign n3458 = n3449 & n3457 ;
  assign n3459 = n3449 | n3452 ;
  assign n3460 = n3405 & ~n3449 ;
  assign n3461 = ( n3455 & n3459 ) | ( n3455 & ~n3460 ) | ( n3459 & ~n3460 ) ;
  assign n3462 = n3451 | n3461 ;
  assign n3463 = ~n2919 & n2932 ;
  assign n3464 = n2919 & ~n2924 ;
  assign n3465 = ~n2912 & n3464 ;
  assign n3466 = ~n2930 & n3465 ;
  assign n3467 = ( ~n2930 & n3463 ) | ( ~n2930 & n3466 ) | ( n3463 & n3466 ) ;
  assign n3468 = n2931 & ~n2933 ;
  assign n3469 = ( n2930 & n3467 ) | ( n2930 & ~n3468 ) | ( n3467 & ~n3468 ) ;
  assign n3470 = n3462 & n3469 ;
  assign n3471 = n3458 | n3470 ;
  assign n3473 = ( n2933 & ~n2938 ) | ( n2933 & n2943 ) | ( ~n2938 & n2943 ) ;
  assign n3474 = n2938 & ~n2943 ;
  assign n3475 = ( n2931 & n3473 ) | ( n2931 & ~n3474 ) | ( n3473 & ~n3474 ) ;
  assign n3472 = n2931 | n2933 ;
  assign n3476 = ( n2938 & ~n3472 ) | ( n2938 & n3475 ) | ( ~n3472 & n3475 ) ;
  assign n3477 = ( ~n2943 & n3475 ) | ( ~n2943 & n3476 ) | ( n3475 & n3476 ) ;
  assign n3479 = ( n3408 & ~n3413 ) | ( n3408 & n3418 ) | ( ~n3413 & n3418 ) ;
  assign n3480 = n3413 & ~n3418 ;
  assign n3481 = ( n3406 & n3479 ) | ( n3406 & ~n3480 ) | ( n3479 & ~n3480 ) ;
  assign n3478 = n3406 | n3408 ;
  assign n3482 = ( n3413 & ~n3478 ) | ( n3413 & n3481 ) | ( ~n3478 & n3481 ) ;
  assign n3483 = ( ~n3418 & n3481 ) | ( ~n3418 & n3482 ) | ( n3481 & n3482 ) ;
  assign n3484 = ( n3471 & n3477 ) | ( n3471 & n3483 ) | ( n3477 & n3483 ) ;
  assign n3485 = ( ~n3175 & n3384 ) | ( ~n3175 & n3421 ) | ( n3384 & n3421 ) ;
  assign n3486 = ( n3175 & ~n3421 ) | ( n3175 & n3485 ) | ( ~n3421 & n3485 ) ;
  assign n3487 = ( ~n3384 & n3485 ) | ( ~n3384 & n3486 ) | ( n3485 & n3486 ) ;
  assign n3488 = ( ~n2700 & n2909 ) | ( ~n2700 & n2946 ) | ( n2909 & n2946 ) ;
  assign n3489 = ( n2700 & ~n2946 ) | ( n2700 & n3488 ) | ( ~n2946 & n3488 ) ;
  assign n3490 = ( ~n2909 & n3488 ) | ( ~n2909 & n3489 ) | ( n3488 & n3489 ) ;
  assign n3491 = ( n3484 & n3487 ) | ( n3484 & n3490 ) | ( n3487 & n3490 ) ;
  assign n3492 = n3442 & n3491 ;
  assign n3493 = n3173 & n3431 ;
  assign n3494 = n3375 | n3430 ;
  assign n3495 = n3372 | n3430 ;
  assign n3496 = ( n3382 & n3494 ) | ( n3382 & n3495 ) | ( n3494 & n3495 ) ;
  assign n3497 = n3493 | n3496 ;
  assign n3498 = n3425 & n3497 ;
  assign n3499 = ( n3422 & n3497 ) | ( n3422 & n3498 ) | ( n3497 & n3498 ) ;
  assign n3500 = n3434 | n3499 ;
  assign n3501 = n2698 & n2956 ;
  assign n3502 = n2900 | n2955 ;
  assign n3503 = n2897 | n2955 ;
  assign n3504 = ( n2907 & n3502 ) | ( n2907 & n3503 ) | ( n3502 & n3503 ) ;
  assign n3505 = n3501 | n3504 ;
  assign n3506 = n2959 | n3505 ;
  assign n3507 = ( n2950 & n2959 ) | ( n2950 & n3506 ) | ( n2959 & n3506 ) ;
  assign n3508 = n2959 | n3506 ;
  assign n3509 = ( n2947 & n3507 ) | ( n2947 & n3508 ) | ( n3507 & n3508 ) ;
  assign n3510 = n3500 & n3509 ;
  assign n3511 = n2959 | n3434 ;
  assign n3512 = n3505 | n3511 ;
  assign n3513 = ( n2964 & n3511 ) | ( n2964 & n3512 ) | ( n3511 & n3512 ) ;
  assign n3514 = n3499 | n3513 ;
  assign n3515 = n3510 | n3514 ;
  assign n3516 = n2963 & n3438 ;
  assign n3517 = n2965 | n3440 ;
  assign n3518 = n3516 & ~n3517 ;
  assign n3519 = ( n3510 & n3515 ) | ( n3510 & n3518 ) | ( n3515 & n3518 ) ;
  assign n3520 = n3510 | n3515 ;
  assign n3521 = ( n3492 & n3519 ) | ( n3492 & n3520 ) | ( n3519 & n3520 ) ;
  assign n2489 = ~n2400 & n2487 ;
  assign n2490 = ~n2403 & n2489 ;
  assign n2491 = ( ~n2477 & n2489 ) | ( ~n2477 & n2490 ) | ( n2489 & n2490 ) ;
  assign n3522 = n2491 & n3521 ;
  assign n3523 = ( n2488 & n3521 ) | ( n2488 & n3522 ) | ( n3521 & n3522 ) ;
  assign n3524 = n2491 | n3521 ;
  assign n3525 = n2488 | n3524 ;
  assign n3526 = ~n3523 & n3525 ;
  assign n3527 = n3492 | n3518 ;
  assign n3528 = n3500 & ~n3510 ;
  assign n3529 = ( n3509 & ~n3510 ) | ( n3509 & n3528 ) | ( ~n3510 & n3528 ) ;
  assign n3530 = n3527 & n3529 ;
  assign n3531 = n3518 | n3529 ;
  assign n3532 = n3492 | n3531 ;
  assign n3533 = ~n3530 & n3532 ;
  assign n3534 = n1917 & ~n2397 ;
  assign n3535 = ( n1920 & ~n2397 ) | ( n1920 & n3534 ) | ( ~n2397 & n3534 ) ;
  assign n3536 = ~n1919 & n3535 ;
  assign n3537 = n2397 & ~n2402 ;
  assign n3538 = n3536 | n3537 ;
  assign n3539 = n2477 & n3538 ;
  assign n3540 = ( n2418 & n2476 ) | ( n2418 & ~n3538 ) | ( n2476 & ~n3538 ) ;
  assign n3541 = n3538 | n3540 ;
  assign n3542 = ~n3539 & n3541 ;
  assign n3543 = ( n1916 & ~n2407 ) | ( n1916 & n2415 ) | ( ~n2407 & n2415 ) ;
  assign n3544 = ( ~n1916 & n2407 ) | ( ~n1916 & n3543 ) | ( n2407 & n3543 ) ;
  assign n3545 = ( ~n2415 & n3543 ) | ( ~n2415 & n3544 ) | ( n3543 & n3544 ) ;
  assign n3546 = n2475 | n3545 ;
  assign n3547 = n2475 & n3545 ;
  assign n3548 = n3546 & ~n3547 ;
  assign n3549 = ( ~n2966 & n3441 ) | ( ~n2966 & n3491 ) | ( n3441 & n3491 ) ;
  assign n3550 = ( n2966 & ~n3491 ) | ( n2966 & n3549 ) | ( ~n3491 & n3549 ) ;
  assign n3551 = ( ~n3441 & n3549 ) | ( ~n3441 & n3550 ) | ( n3549 & n3550 ) ;
  assign n3552 = ~n2430 & n2433 ;
  assign n3553 = n2426 | n2433 ;
  assign n3554 = n2429 & ~n3553 ;
  assign n3555 = n3552 | n3554 ;
  assign n3556 = n2474 | n3555 ;
  assign n3557 = n2474 & n3555 ;
  assign n3558 = n3556 & ~n3557 ;
  assign n3559 = ( n3484 & ~n3487 ) | ( n3484 & n3490 ) | ( ~n3487 & n3490 ) ;
  assign n3560 = ( ~n3484 & n3487 ) | ( ~n3484 & n3559 ) | ( n3487 & n3559 ) ;
  assign n3561 = ( ~n3490 & n3559 ) | ( ~n3490 & n3560 ) | ( n3559 & n3560 ) ;
  assign n3562 = n3558 | n3561 ;
  assign n3563 = n2436 & ~n2439 ;
  assign n3564 = ~n2434 & n2439 ;
  assign n3565 = ~n2435 & n3564 ;
  assign n3566 = n3563 | n3565 ;
  assign n3567 = n3445 & ~n3448 ;
  assign n3568 = ~n3445 & n3448 ;
  assign n3569 = n3567 | n3568 ;
  assign n3570 = n3566 & n3569 ;
  assign n3571 = ~n2452 & n2459 ;
  assign n3572 = ( n2449 & n2459 ) | ( n2449 & n3571 ) | ( n2459 & n3571 ) ;
  assign n3573 = ~n2440 & n2448 ;
  assign n3574 = n1899 & n2440 ;
  assign n3575 = ( n2440 & ~n2446 ) | ( n2440 & n3574 ) | ( ~n2446 & n3574 ) ;
  assign n3576 = ~n2443 & n3575 ;
  assign n3577 = ~n2459 & n3576 ;
  assign n3578 = ( ~n2459 & n3573 ) | ( ~n2459 & n3577 ) | ( n3573 & n3577 ) ;
  assign n3579 = n3572 | n3578 ;
  assign n3580 = n3570 & n3579 ;
  assign n3581 = n3570 | n3578 ;
  assign n3582 = ( n3449 & ~n3457 ) | ( n3449 & n3469 ) | ( ~n3457 & n3469 ) ;
  assign n3583 = ( ~n3449 & n3457 ) | ( ~n3449 & n3582 ) | ( n3457 & n3582 ) ;
  assign n3584 = ( ~n3469 & n3582 ) | ( ~n3469 & n3583 ) | ( n3582 & n3583 ) ;
  assign n3585 = n3572 & n3584 ;
  assign n3586 = ( n3581 & n3584 ) | ( n3581 & n3585 ) | ( n3584 & n3585 ) ;
  assign n3587 = n3580 | n3586 ;
  assign n3588 = n1902 | n2470 ;
  assign n3589 = n1902 & n2470 ;
  assign n3590 = n3588 & ~n3589 ;
  assign n3591 = n2467 & ~n3590 ;
  assign n3592 = n1902 | n2467 ;
  assign n3593 = ( n2467 & n2470 ) | ( n2467 & n3592 ) | ( n2470 & n3592 ) ;
  assign n3594 = n3588 & ~n3593 ;
  assign n3595 = n2461 | n3594 ;
  assign n3596 = n3591 | n3595 ;
  assign n3597 = n2461 & n3594 ;
  assign n3598 = ( n2461 & n3591 ) | ( n2461 & n3597 ) | ( n3591 & n3597 ) ;
  assign n3599 = n3596 & ~n3598 ;
  assign n3600 = ( n3471 & ~n3477 ) | ( n3471 & n3483 ) | ( ~n3477 & n3483 ) ;
  assign n3601 = ( ~n3471 & n3477 ) | ( ~n3471 & n3600 ) | ( n3477 & n3600 ) ;
  assign n3602 = ( ~n3483 & n3600 ) | ( ~n3483 & n3601 ) | ( n3600 & n3601 ) ;
  assign n3603 = ( n3587 & n3599 ) | ( n3587 & n3602 ) | ( n3599 & n3602 ) ;
  assign n3604 = ( n2474 & n3555 ) | ( n2474 & ~n3561 ) | ( n3555 & ~n3561 ) ;
  assign n3605 = ( n3556 & n3603 ) | ( n3556 & ~n3604 ) | ( n3603 & ~n3604 ) ;
  assign n3606 = n3556 & ~n3604 ;
  assign n3607 = ( n3562 & n3605 ) | ( n3562 & n3606 ) | ( n3605 & n3606 ) ;
  assign n3608 = ( n3548 & n3551 ) | ( n3548 & n3607 ) | ( n3551 & n3607 ) ;
  assign n3609 = ( n3533 & n3542 ) | ( n3533 & n3608 ) | ( n3542 & n3608 ) ;
  assign n3610 = n3526 & n3609 ;
  assign n3611 = n3526 | n3609 ;
  assign n3612 = ~n3610 & n3611 ;
  assign n3613 = ~x403 & x404 ;
  assign n3614 = x403 & ~x404 ;
  assign n3615 = n3613 | n3614 ;
  assign n3616 = ~x405 & n3615 ;
  assign n3617 = x405 & ~n3615 ;
  assign n3618 = n3616 | n3617 ;
  assign n3619 = ~x406 & x407 ;
  assign n3620 = x406 & ~x407 ;
  assign n3621 = n3619 | n3620 ;
  assign n3622 = ~x408 & n3621 ;
  assign n3623 = x408 & ~n3621 ;
  assign n3624 = n3622 | n3623 ;
  assign n3625 = n3618 & n3624 ;
  assign n3626 = ( x406 & x407 ) | ( x406 & x408 ) | ( x407 & x408 ) ;
  assign n3627 = ( x403 & x404 ) | ( x403 & x405 ) | ( x404 & x405 ) ;
  assign n3628 = ~n3626 & n3627 ;
  assign n3629 = n3626 & ~n3627 ;
  assign n3630 = n3628 | n3629 ;
  assign n3631 = ~n3625 & n3630 ;
  assign n3632 = n3625 & ~n3630 ;
  assign n3633 = n3631 | n3632 ;
  assign n3634 = n3618 & ~n3624 ;
  assign n3635 = ~n3618 & n3624 ;
  assign n3636 = n3634 | n3635 ;
  assign n3637 = ( n3625 & n3626 ) | ( n3625 & n3627 ) | ( n3626 & n3627 ) ;
  assign n3638 = n3636 & n3637 ;
  assign n3639 = n3633 & ~n3638 ;
  assign n3640 = n3633 & n3637 ;
  assign n3641 = x409 & ~x410 ;
  assign n3642 = ~x409 & x410 ;
  assign n3643 = n3641 | n3642 ;
  assign n3644 = ~x411 & n3643 ;
  assign n3645 = x411 & ~n3643 ;
  assign n3646 = n3644 | n3645 ;
  assign n3647 = x412 & ~x413 ;
  assign n3648 = ~x412 & x413 ;
  assign n3649 = n3647 | n3648 ;
  assign n3650 = ~x414 & n3649 ;
  assign n3651 = x414 & ~n3649 ;
  assign n3652 = n3650 | n3651 ;
  assign n3653 = n3646 & ~n3652 ;
  assign n3654 = ~n3646 & n3652 ;
  assign n3655 = n3653 | n3654 ;
  assign n3656 = ( x412 & x413 ) | ( x412 & x414 ) | ( x413 & x414 ) ;
  assign n3657 = ( x409 & x410 ) | ( x409 & x411 ) | ( x410 & x411 ) ;
  assign n3658 = n3646 & n3652 ;
  assign n3659 = ( n3656 & n3657 ) | ( n3656 & n3658 ) | ( n3657 & n3658 ) ;
  assign n3660 = n3655 & n3659 ;
  assign n3661 = n3640 | n3660 ;
  assign n3662 = n3656 & ~n3657 ;
  assign n3663 = ~n3656 & n3657 ;
  assign n3664 = n3662 | n3663 ;
  assign n3665 = ~n3658 & n3664 ;
  assign n3666 = n3658 & ~n3664 ;
  assign n3667 = n3665 | n3666 ;
  assign n3668 = n3659 & n3667 ;
  assign n3669 = n3636 & n3655 ;
  assign n3670 = n3667 & n3669 ;
  assign n3671 = ~n3668 & n3670 ;
  assign n3672 = ~n3661 & n3671 ;
  assign n3673 = n3639 & n3672 ;
  assign n3674 = ~n3668 & n3669 ;
  assign n3675 = ~n3660 & n3667 ;
  assign n3676 = n3640 & ~n3675 ;
  assign n3677 = ( n3674 & n3675 ) | ( n3674 & ~n3676 ) | ( n3675 & ~n3676 ) ;
  assign n3678 = ( n3639 & n3673 ) | ( n3639 & ~n3677 ) | ( n3673 & ~n3677 ) ;
  assign n3679 = n3655 & ~n3659 ;
  assign n3680 = ( n3655 & ~n3667 ) | ( n3655 & n3679 ) | ( ~n3667 & n3679 ) ;
  assign n3681 = n3636 & ~n3637 ;
  assign n3682 = ( ~n3633 & n3636 ) | ( ~n3633 & n3681 ) | ( n3636 & n3681 ) ;
  assign n3683 = ~n3680 & n3682 ;
  assign n3684 = n3680 & ~n3682 ;
  assign n3685 = n3683 | n3684 ;
  assign n3686 = ( x400 & x401 ) | ( x400 & x402 ) | ( x401 & x402 ) ;
  assign n3687 = ( x397 & x398 ) | ( x397 & x399 ) | ( x398 & x399 ) ;
  assign n3688 = n3686 & ~n3687 ;
  assign n3689 = ~n3686 & n3687 ;
  assign n3690 = n3688 | n3689 ;
  assign n3691 = x397 & ~x398 ;
  assign n3692 = ~x397 & x398 ;
  assign n3693 = n3691 | n3692 ;
  assign n3694 = ~x399 & n3693 ;
  assign n3695 = x399 & ~n3693 ;
  assign n3696 = n3694 | n3695 ;
  assign n3697 = x400 & ~x401 ;
  assign n3698 = ~x400 & x401 ;
  assign n3699 = n3697 | n3698 ;
  assign n3700 = ~x402 & n3699 ;
  assign n3701 = x402 & ~n3699 ;
  assign n3702 = n3700 | n3701 ;
  assign n3703 = n3696 & n3702 ;
  assign n3704 = n3690 & ~n3703 ;
  assign n3705 = ~n3690 & n3703 ;
  assign n3706 = n3704 | n3705 ;
  assign n3707 = n3696 & ~n3702 ;
  assign n3708 = ~n3696 & n3702 ;
  assign n3709 = n3707 | n3708 ;
  assign n3710 = ( n3686 & n3687 ) | ( n3686 & n3703 ) | ( n3687 & n3703 ) ;
  assign n3711 = n3709 & ~n3710 ;
  assign n3712 = ( ~n3706 & n3709 ) | ( ~n3706 & n3711 ) | ( n3709 & n3711 ) ;
  assign n3713 = ~x391 & x392 ;
  assign n3714 = x391 & ~x392 ;
  assign n3715 = n3713 | n3714 ;
  assign n3716 = ~x393 & n3715 ;
  assign n3717 = x393 & ~n3715 ;
  assign n3718 = n3716 | n3717 ;
  assign n3719 = ~x394 & x395 ;
  assign n3720 = x394 & ~x395 ;
  assign n3721 = n3719 | n3720 ;
  assign n3722 = ~x396 & n3721 ;
  assign n3723 = x396 & ~n3721 ;
  assign n3724 = n3722 | n3723 ;
  assign n3725 = n3718 & n3724 ;
  assign n3726 = ( x394 & x395 ) | ( x394 & x396 ) | ( x395 & x396 ) ;
  assign n3727 = ( x391 & x392 ) | ( x391 & x393 ) | ( x392 & x393 ) ;
  assign n3728 = ~n3726 & n3727 ;
  assign n3729 = n3726 & ~n3727 ;
  assign n3730 = n3728 | n3729 ;
  assign n3731 = ~n3725 & n3730 ;
  assign n3732 = n3725 & ~n3730 ;
  assign n3733 = n3731 | n3732 ;
  assign n3734 = n3718 & ~n3724 ;
  assign n3735 = ~n3718 & n3724 ;
  assign n3736 = n3734 | n3735 ;
  assign n3737 = ( n3725 & n3726 ) | ( n3725 & n3727 ) | ( n3726 & n3727 ) ;
  assign n3738 = n3736 & ~n3737 ;
  assign n3739 = ( ~n3733 & n3736 ) | ( ~n3733 & n3738 ) | ( n3736 & n3738 ) ;
  assign n3740 = ~n3712 & n3739 ;
  assign n3741 = n3712 & ~n3739 ;
  assign n3742 = n3740 | n3741 ;
  assign n3743 = n3685 & n3742 ;
  assign n3744 = ( n3639 & ~n3640 ) | ( n3639 & n3675 ) | ( ~n3640 & n3675 ) ;
  assign n3745 = n3639 & n3675 ;
  assign n3746 = ( n3674 & n3744 ) | ( n3674 & n3745 ) | ( n3744 & n3745 ) ;
  assign n3747 = n3677 & ~n3746 ;
  assign n3748 = n3743 | n3747 ;
  assign n3749 = n3678 | n3748 ;
  assign n3750 = n3733 & n3737 ;
  assign n3751 = n3709 & n3710 ;
  assign n3752 = n3750 | n3751 ;
  assign n3753 = n3706 & n3710 ;
  assign n3754 = n3709 & n3736 ;
  assign n3755 = n3706 & n3754 ;
  assign n3756 = ~n3753 & n3755 ;
  assign n3757 = ~n3752 & n3756 ;
  assign n3758 = n3736 & n3737 ;
  assign n3759 = n3733 & ~n3758 ;
  assign n3760 = ~n3757 & n3759 ;
  assign n3761 = ~n3753 & n3754 ;
  assign n3762 = n3706 & ~n3751 ;
  assign n3763 = ( n3750 & n3759 ) | ( n3750 & n3762 ) | ( n3759 & n3762 ) ;
  assign n3764 = n3759 | n3762 ;
  assign n3765 = ( ~n3761 & n3763 ) | ( ~n3761 & n3764 ) | ( n3763 & n3764 ) ;
  assign n3766 = n3750 | n3762 ;
  assign n3767 = n3761 & ~n3766 ;
  assign n3768 = ( ~n3762 & n3765 ) | ( ~n3762 & n3767 ) | ( n3765 & n3767 ) ;
  assign n3769 = ( ~n3760 & n3765 ) | ( ~n3760 & n3768 ) | ( n3765 & n3768 ) ;
  assign n3770 = n3749 & n3769 ;
  assign n3771 = n3743 & n3747 ;
  assign n3772 = ( n3678 & n3743 ) | ( n3678 & n3771 ) | ( n3743 & n3771 ) ;
  assign n3773 = n3770 | n3772 ;
  assign n3774 = n3750 & ~n3762 ;
  assign n3775 = ( n3761 & n3762 ) | ( n3761 & ~n3774 ) | ( n3762 & ~n3774 ) ;
  assign n3776 = n3759 & n3775 ;
  assign n3777 = ~n3736 & n3737 ;
  assign n3778 = ( ~n3733 & n3737 ) | ( ~n3733 & n3777 ) | ( n3737 & n3777 ) ;
  assign n3779 = ~n3709 & n3710 ;
  assign n3780 = ( ~n3706 & n3710 ) | ( ~n3706 & n3779 ) | ( n3710 & n3779 ) ;
  assign n3781 = ~n3778 & n3780 ;
  assign n3782 = n3778 & ~n3780 ;
  assign n3783 = n3781 | n3782 ;
  assign n3784 = n3757 | n3783 ;
  assign n3785 = n3776 | n3784 ;
  assign n3786 = n3757 & n3783 ;
  assign n3787 = ( n3776 & n3783 ) | ( n3776 & n3786 ) | ( n3783 & n3786 ) ;
  assign n3788 = n3785 & ~n3787 ;
  assign n3789 = n3639 & n3677 ;
  assign n3790 = ~n3636 & n3637 ;
  assign n3791 = ( ~n3633 & n3637 ) | ( ~n3633 & n3790 ) | ( n3637 & n3790 ) ;
  assign n3792 = ~n3655 & n3659 ;
  assign n3793 = ( n3659 & ~n3667 ) | ( n3659 & n3792 ) | ( ~n3667 & n3792 ) ;
  assign n3794 = ~n3791 & n3793 ;
  assign n3795 = n3791 & ~n3793 ;
  assign n3796 = n3794 | n3795 ;
  assign n3797 = n3672 | n3796 ;
  assign n3798 = n3789 | n3797 ;
  assign n3799 = n3672 & n3796 ;
  assign n3800 = ( n3789 & n3796 ) | ( n3789 & n3799 ) | ( n3796 & n3799 ) ;
  assign n3801 = n3798 & ~n3800 ;
  assign n3802 = n3788 | n3801 ;
  assign n3803 = n3773 & n3802 ;
  assign n3804 = n3785 & n3798 ;
  assign n3805 = n3787 | n3800 ;
  assign n3806 = n3804 & ~n3805 ;
  assign n3807 = ( n3672 & n3791 ) | ( n3672 & n3793 ) | ( n3791 & n3793 ) ;
  assign n3808 = n3791 | n3793 ;
  assign n3809 = ( n3789 & n3807 ) | ( n3789 & n3808 ) | ( n3807 & n3808 ) ;
  assign n3810 = ( n3757 & n3778 ) | ( n3757 & n3780 ) | ( n3778 & n3780 ) ;
  assign n3811 = n3778 | n3780 ;
  assign n3812 = ( n3776 & n3810 ) | ( n3776 & n3811 ) | ( n3810 & n3811 ) ;
  assign n3813 = ~n3809 & n3812 ;
  assign n3814 = n3809 & ~n3812 ;
  assign n3815 = n3813 | n3814 ;
  assign n3816 = n3806 | n3815 ;
  assign n3817 = n3803 | n3816 ;
  assign n3818 = n3802 | n3806 ;
  assign n3819 = ( n3773 & n3806 ) | ( n3773 & n3818 ) | ( n3806 & n3818 ) ;
  assign n3820 = n3815 & n3819 ;
  assign n3821 = n3817 & ~n3820 ;
  assign n3822 = ( x382 & x383 ) | ( x382 & x384 ) | ( x383 & x384 ) ;
  assign n3823 = ( x379 & x380 ) | ( x379 & x381 ) | ( x380 & x381 ) ;
  assign n3824 = n3822 & ~n3823 ;
  assign n3825 = ~n3822 & n3823 ;
  assign n3826 = n3824 | n3825 ;
  assign n3827 = ~x379 & x380 ;
  assign n3828 = x379 & ~x380 ;
  assign n3829 = n3827 | n3828 ;
  assign n3830 = ~x381 & n3829 ;
  assign n3831 = x381 & ~n3829 ;
  assign n3832 = n3830 | n3831 ;
  assign n3833 = ~x382 & x383 ;
  assign n3834 = x382 & ~x383 ;
  assign n3835 = n3833 | n3834 ;
  assign n3836 = ~x384 & n3835 ;
  assign n3837 = x384 & ~n3835 ;
  assign n3838 = n3836 | n3837 ;
  assign n3839 = n3832 & n3838 ;
  assign n3840 = n3826 & ~n3839 ;
  assign n3841 = ~n3826 & n3839 ;
  assign n3842 = n3840 | n3841 ;
  assign n3843 = n3832 & ~n3838 ;
  assign n3844 = ~n3832 & n3838 ;
  assign n3845 = n3843 | n3844 ;
  assign n3846 = ( n3822 & n3823 ) | ( n3822 & n3839 ) | ( n3823 & n3839 ) ;
  assign n3847 = n3845 & n3846 ;
  assign n3848 = n3842 & ~n3847 ;
  assign n3849 = n3842 & n3846 ;
  assign n3850 = ~x385 & x386 ;
  assign n3851 = x385 & ~x386 ;
  assign n3852 = n3850 | n3851 ;
  assign n3853 = ~x387 & n3852 ;
  assign n3854 = x387 & ~n3852 ;
  assign n3855 = n3853 | n3854 ;
  assign n3856 = ~x388 & x389 ;
  assign n3857 = x388 & ~x389 ;
  assign n3858 = n3856 | n3857 ;
  assign n3859 = ~x390 & n3858 ;
  assign n3860 = x390 & ~n3858 ;
  assign n3861 = n3859 | n3860 ;
  assign n3862 = n3855 & ~n3861 ;
  assign n3863 = ~n3855 & n3861 ;
  assign n3864 = n3862 | n3863 ;
  assign n3865 = ( x388 & x389 ) | ( x388 & x390 ) | ( x389 & x390 ) ;
  assign n3866 = ( x385 & x386 ) | ( x385 & x387 ) | ( x386 & x387 ) ;
  assign n3867 = n3855 & n3861 ;
  assign n3868 = ( n3865 & n3866 ) | ( n3865 & n3867 ) | ( n3866 & n3867 ) ;
  assign n3869 = n3864 & n3868 ;
  assign n3870 = n3849 | n3869 ;
  assign n3871 = n3865 & ~n3866 ;
  assign n3872 = ~n3865 & n3866 ;
  assign n3873 = n3871 | n3872 ;
  assign n3874 = ~n3867 & n3873 ;
  assign n3875 = n3867 & ~n3873 ;
  assign n3876 = n3874 | n3875 ;
  assign n3877 = n3868 & n3876 ;
  assign n3878 = n3845 & n3864 ;
  assign n3879 = n3876 & n3878 ;
  assign n3880 = ~n3877 & n3879 ;
  assign n3881 = ~n3870 & n3880 ;
  assign n3882 = n3848 & n3881 ;
  assign n3883 = ~n3877 & n3878 ;
  assign n3884 = ~n3869 & n3876 ;
  assign n3885 = n3849 & ~n3884 ;
  assign n3886 = ( n3883 & n3884 ) | ( n3883 & ~n3885 ) | ( n3884 & ~n3885 ) ;
  assign n3887 = ( n3848 & n3882 ) | ( n3848 & ~n3886 ) | ( n3882 & ~n3886 ) ;
  assign n3888 = n3864 & ~n3868 ;
  assign n3889 = ( n3864 & ~n3876 ) | ( n3864 & n3888 ) | ( ~n3876 & n3888 ) ;
  assign n3890 = n3845 & ~n3846 ;
  assign n3891 = ( ~n3842 & n3845 ) | ( ~n3842 & n3890 ) | ( n3845 & n3890 ) ;
  assign n3892 = ~n3889 & n3891 ;
  assign n3893 = n3889 & ~n3891 ;
  assign n3894 = n3892 | n3893 ;
  assign n3895 = ( x376 & x377 ) | ( x376 & x378 ) | ( x377 & x378 ) ;
  assign n3896 = ( x373 & x374 ) | ( x373 & x375 ) | ( x374 & x375 ) ;
  assign n3897 = n3895 & ~n3896 ;
  assign n3898 = ~n3895 & n3896 ;
  assign n3899 = n3897 | n3898 ;
  assign n3900 = ~x373 & x374 ;
  assign n3901 = x373 & ~x374 ;
  assign n3902 = n3900 | n3901 ;
  assign n3903 = ~x375 & n3902 ;
  assign n3904 = x375 & ~n3902 ;
  assign n3905 = n3903 | n3904 ;
  assign n3906 = ~x376 & x377 ;
  assign n3907 = x376 & ~x377 ;
  assign n3908 = n3906 | n3907 ;
  assign n3909 = ~x378 & n3908 ;
  assign n3910 = x378 & ~n3908 ;
  assign n3911 = n3909 | n3910 ;
  assign n3912 = n3905 & n3911 ;
  assign n3913 = n3899 & ~n3912 ;
  assign n3914 = ~n3899 & n3912 ;
  assign n3915 = n3913 | n3914 ;
  assign n3916 = n3905 & ~n3911 ;
  assign n3917 = ~n3905 & n3911 ;
  assign n3918 = n3916 | n3917 ;
  assign n3919 = ( n3895 & n3896 ) | ( n3895 & n3912 ) | ( n3896 & n3912 ) ;
  assign n3920 = n3918 & ~n3919 ;
  assign n3921 = ( ~n3915 & n3918 ) | ( ~n3915 & n3920 ) | ( n3918 & n3920 ) ;
  assign n3922 = ~x367 & x368 ;
  assign n3923 = x367 & ~x368 ;
  assign n3924 = n3922 | n3923 ;
  assign n3925 = ~x369 & n3924 ;
  assign n3926 = x369 & ~n3924 ;
  assign n3927 = n3925 | n3926 ;
  assign n3928 = ~x370 & x371 ;
  assign n3929 = x370 & ~x371 ;
  assign n3930 = n3928 | n3929 ;
  assign n3931 = ~x372 & n3930 ;
  assign n3932 = x372 & ~n3930 ;
  assign n3933 = n3931 | n3932 ;
  assign n3934 = n3927 & ~n3933 ;
  assign n3935 = ~n3927 & n3933 ;
  assign n3936 = n3934 | n3935 ;
  assign n3937 = ( x370 & x371 ) | ( x370 & x372 ) | ( x371 & x372 ) ;
  assign n3938 = ( x367 & x368 ) | ( x367 & x369 ) | ( x368 & x369 ) ;
  assign n3939 = n3937 & ~n3938 ;
  assign n3940 = ~n3937 & n3938 ;
  assign n3941 = n3939 | n3940 ;
  assign n3942 = n3927 & n3933 ;
  assign n3943 = n3941 & ~n3942 ;
  assign n3944 = ~n3941 & n3942 ;
  assign n3945 = n3943 | n3944 ;
  assign n3946 = ( n3937 & n3938 ) | ( n3937 & n3942 ) | ( n3938 & n3942 ) ;
  assign n3947 = n3936 & ~n3946 ;
  assign n3948 = ( n3936 & ~n3945 ) | ( n3936 & n3947 ) | ( ~n3945 & n3947 ) ;
  assign n3949 = ~n3921 & n3948 ;
  assign n3950 = n3921 & ~n3948 ;
  assign n3951 = n3949 | n3950 ;
  assign n3952 = n3894 & n3951 ;
  assign n3953 = ( n3848 & ~n3849 ) | ( n3848 & n3884 ) | ( ~n3849 & n3884 ) ;
  assign n3954 = n3848 & n3884 ;
  assign n3955 = ( n3883 & n3953 ) | ( n3883 & n3954 ) | ( n3953 & n3954 ) ;
  assign n3956 = n3886 & ~n3955 ;
  assign n3957 = n3952 | n3956 ;
  assign n3958 = n3887 | n3957 ;
  assign n3959 = n3945 & n3946 ;
  assign n3960 = n3918 & n3919 ;
  assign n3961 = n3959 | n3960 ;
  assign n3962 = n3915 & n3919 ;
  assign n3963 = n3918 & n3936 ;
  assign n3964 = n3915 & n3963 ;
  assign n3965 = ~n3962 & n3964 ;
  assign n3966 = ~n3961 & n3965 ;
  assign n3967 = n3936 & n3946 ;
  assign n3968 = n3945 & ~n3967 ;
  assign n3969 = ~n3966 & n3968 ;
  assign n3970 = ~n3962 & n3963 ;
  assign n3971 = n3915 & ~n3960 ;
  assign n3972 = ( n3959 & n3968 ) | ( n3959 & n3971 ) | ( n3968 & n3971 ) ;
  assign n3973 = n3968 | n3971 ;
  assign n3974 = ( ~n3970 & n3972 ) | ( ~n3970 & n3973 ) | ( n3972 & n3973 ) ;
  assign n3975 = n3959 | n3971 ;
  assign n3976 = n3970 & ~n3975 ;
  assign n3977 = ( ~n3971 & n3974 ) | ( ~n3971 & n3976 ) | ( n3974 & n3976 ) ;
  assign n3978 = ( ~n3969 & n3974 ) | ( ~n3969 & n3977 ) | ( n3974 & n3977 ) ;
  assign n3979 = n3958 & n3978 ;
  assign n3980 = n3952 & n3956 ;
  assign n3981 = ( n3887 & n3952 ) | ( n3887 & n3980 ) | ( n3952 & n3980 ) ;
  assign n3982 = n3979 | n3981 ;
  assign n3983 = n3959 & ~n3971 ;
  assign n3984 = ( n3970 & n3971 ) | ( n3970 & ~n3983 ) | ( n3971 & ~n3983 ) ;
  assign n3985 = n3968 & n3984 ;
  assign n3986 = ~n3936 & n3946 ;
  assign n3987 = ( ~n3945 & n3946 ) | ( ~n3945 & n3986 ) | ( n3946 & n3986 ) ;
  assign n3988 = ~n3918 & n3919 ;
  assign n3989 = ( ~n3915 & n3919 ) | ( ~n3915 & n3988 ) | ( n3919 & n3988 ) ;
  assign n3990 = ~n3987 & n3989 ;
  assign n3991 = n3987 & ~n3989 ;
  assign n3992 = n3990 | n3991 ;
  assign n3993 = n3966 | n3992 ;
  assign n3994 = n3985 | n3993 ;
  assign n3995 = n3966 & n3992 ;
  assign n3996 = ( n3985 & n3992 ) | ( n3985 & n3995 ) | ( n3992 & n3995 ) ;
  assign n3997 = n3994 & ~n3996 ;
  assign n3998 = n3848 & n3886 ;
  assign n3999 = ~n3845 & n3846 ;
  assign n4000 = ( ~n3842 & n3846 ) | ( ~n3842 & n3999 ) | ( n3846 & n3999 ) ;
  assign n4001 = ~n3864 & n3868 ;
  assign n4002 = ( n3868 & ~n3876 ) | ( n3868 & n4001 ) | ( ~n3876 & n4001 ) ;
  assign n4003 = ~n4000 & n4002 ;
  assign n4004 = n4000 & ~n4002 ;
  assign n4005 = n4003 | n4004 ;
  assign n4006 = n3881 | n4005 ;
  assign n4007 = n3998 | n4006 ;
  assign n4008 = n3881 & n4005 ;
  assign n4009 = ( n3998 & n4005 ) | ( n3998 & n4008 ) | ( n4005 & n4008 ) ;
  assign n4010 = n4007 & ~n4009 ;
  assign n4011 = n3997 | n4010 ;
  assign n4012 = n3982 & n4011 ;
  assign n4013 = n3994 & n4007 ;
  assign n4014 = n3996 | n4009 ;
  assign n4015 = n4013 & ~n4014 ;
  assign n4016 = ( n3881 & n4000 ) | ( n3881 & n4002 ) | ( n4000 & n4002 ) ;
  assign n4017 = n4000 | n4002 ;
  assign n4018 = ( n3998 & n4016 ) | ( n3998 & n4017 ) | ( n4016 & n4017 ) ;
  assign n4019 = ( n3966 & n3987 ) | ( n3966 & n3989 ) | ( n3987 & n3989 ) ;
  assign n4020 = n3987 | n3989 ;
  assign n4021 = ( n3985 & n4019 ) | ( n3985 & n4020 ) | ( n4019 & n4020 ) ;
  assign n4022 = ~n4018 & n4021 ;
  assign n4023 = n4018 & ~n4021 ;
  assign n4024 = n4022 | n4023 ;
  assign n4025 = n4015 | n4024 ;
  assign n4026 = n4012 | n4025 ;
  assign n4027 = n4011 | n4015 ;
  assign n4028 = ( n3982 & n4015 ) | ( n3982 & n4027 ) | ( n4015 & n4027 ) ;
  assign n4029 = n4024 & n4028 ;
  assign n4030 = n4026 & ~n4029 ;
  assign n4031 = n3821 | n4030 ;
  assign n4032 = n3749 & ~n3772 ;
  assign n4033 = n3769 & ~n4032 ;
  assign n4034 = n3685 & ~n3742 ;
  assign n4035 = ~n3685 & n3742 ;
  assign n4036 = n4034 | n4035 ;
  assign n4037 = n3894 & ~n3951 ;
  assign n4038 = ~n3894 & n3951 ;
  assign n4039 = n4037 | n4038 ;
  assign n4040 = n4036 & n4039 ;
  assign n4041 = ~n3743 & n3749 ;
  assign n4042 = n3749 & ~n3769 ;
  assign n4043 = n3678 | n3747 ;
  assign n4044 = n3769 | n4043 ;
  assign n4045 = ( n4041 & n4042 ) | ( n4041 & ~n4044 ) | ( n4042 & ~n4044 ) ;
  assign n4046 = n4040 | n4045 ;
  assign n4047 = n4033 | n4046 ;
  assign n4048 = n3887 | n3956 ;
  assign n4049 = ( n3952 & n3978 ) | ( n3952 & ~n4048 ) | ( n3978 & ~n4048 ) ;
  assign n4050 = ( ~n3978 & n4048 ) | ( ~n3978 & n4049 ) | ( n4048 & n4049 ) ;
  assign n4051 = ( ~n3952 & n4049 ) | ( ~n3952 & n4050 ) | ( n4049 & n4050 ) ;
  assign n4052 = n4047 & n4051 ;
  assign n4053 = n4033 | n4045 ;
  assign n4054 = n4040 & n4053 ;
  assign n4055 = ( n3981 & ~n3997 ) | ( n3981 & n4010 ) | ( ~n3997 & n4010 ) ;
  assign n4056 = n3997 & ~n4010 ;
  assign n4057 = ( n3979 & n4055 ) | ( n3979 & ~n4056 ) | ( n4055 & ~n4056 ) ;
  assign n4058 = ( ~n3982 & n3997 ) | ( ~n3982 & n4057 ) | ( n3997 & n4057 ) ;
  assign n4059 = ( ~n4010 & n4057 ) | ( ~n4010 & n4058 ) | ( n4057 & n4058 ) ;
  assign n4060 = ( n3772 & ~n3788 ) | ( n3772 & n3801 ) | ( ~n3788 & n3801 ) ;
  assign n4061 = n3788 & ~n3801 ;
  assign n4062 = ( n3770 & n4060 ) | ( n3770 & ~n4061 ) | ( n4060 & ~n4061 ) ;
  assign n4063 = ( ~n3773 & n3788 ) | ( ~n3773 & n4062 ) | ( n3788 & n4062 ) ;
  assign n4064 = ( ~n3801 & n4062 ) | ( ~n3801 & n4063 ) | ( n4062 & n4063 ) ;
  assign n4065 = ( n4054 & n4059 ) | ( n4054 & n4064 ) | ( n4059 & n4064 ) ;
  assign n4066 = n4059 | n4064 ;
  assign n4067 = ( n4052 & n4065 ) | ( n4052 & n4066 ) | ( n4065 & n4066 ) ;
  assign n4068 = n4031 & n4067 ;
  assign n4069 = n3817 & n4026 ;
  assign n4070 = n3820 | n4029 ;
  assign n4071 = n4069 & ~n4070 ;
  assign n4072 = n4018 & n4021 ;
  assign n4073 = n4018 | n4021 ;
  assign n4074 = n4072 | n4073 ;
  assign n4075 = ( n4028 & n4072 ) | ( n4028 & n4074 ) | ( n4072 & n4074 ) ;
  assign n4076 = n3809 & n3812 ;
  assign n4077 = n3809 | n3812 ;
  assign n4078 = n4076 | n4077 ;
  assign n4079 = ( n3819 & n4076 ) | ( n3819 & n4078 ) | ( n4076 & n4078 ) ;
  assign n4080 = n4075 & n4079 ;
  assign n4081 = n4079 & ~n4080 ;
  assign n4082 = ( n4075 & ~n4080 ) | ( n4075 & n4081 ) | ( ~n4080 & n4081 ) ;
  assign n4083 = n4071 | n4082 ;
  assign n4084 = n4068 | n4083 ;
  assign n4085 = n4068 | n4071 ;
  assign n4086 = n4082 & n4085 ;
  assign n4087 = n4084 & ~n4086 ;
  assign n4088 = ~x451 & x452 ;
  assign n4089 = x451 & ~x452 ;
  assign n4090 = n4088 | n4089 ;
  assign n4091 = ~x453 & n4090 ;
  assign n4092 = x453 & ~n4090 ;
  assign n4093 = n4091 | n4092 ;
  assign n4094 = ~x454 & x455 ;
  assign n4095 = x454 & ~x455 ;
  assign n4096 = n4094 | n4095 ;
  assign n4097 = ~x456 & n4096 ;
  assign n4098 = x456 & ~n4096 ;
  assign n4099 = n4097 | n4098 ;
  assign n4100 = n4093 & n4099 ;
  assign n4101 = ( x454 & x455 ) | ( x454 & x456 ) | ( x455 & x456 ) ;
  assign n4102 = ( x451 & x452 ) | ( x451 & x453 ) | ( x452 & x453 ) ;
  assign n4103 = ~n4101 & n4102 ;
  assign n4104 = n4101 & ~n4102 ;
  assign n4105 = n4103 | n4104 ;
  assign n4106 = ~n4100 & n4105 ;
  assign n4107 = n4100 & ~n4105 ;
  assign n4108 = n4106 | n4107 ;
  assign n4109 = n4093 & ~n4099 ;
  assign n4110 = ~n4093 & n4099 ;
  assign n4111 = n4109 | n4110 ;
  assign n4112 = ( n4100 & n4101 ) | ( n4100 & n4102 ) | ( n4101 & n4102 ) ;
  assign n4113 = n4111 & n4112 ;
  assign n4114 = n4108 & ~n4113 ;
  assign n4115 = n4108 & n4112 ;
  assign n4116 = x457 & ~x458 ;
  assign n4117 = ~x457 & x458 ;
  assign n4118 = n4116 | n4117 ;
  assign n4119 = ~x459 & n4118 ;
  assign n4120 = x459 & ~n4118 ;
  assign n4121 = n4119 | n4120 ;
  assign n4122 = x460 & ~x461 ;
  assign n4123 = ~x460 & x461 ;
  assign n4124 = n4122 | n4123 ;
  assign n4125 = ~x462 & n4124 ;
  assign n4126 = x462 & ~n4124 ;
  assign n4127 = n4125 | n4126 ;
  assign n4128 = n4121 & ~n4127 ;
  assign n4129 = ~n4121 & n4127 ;
  assign n4130 = n4128 | n4129 ;
  assign n4131 = ( x460 & x461 ) | ( x460 & x462 ) | ( x461 & x462 ) ;
  assign n4132 = ( x457 & x458 ) | ( x457 & x459 ) | ( x458 & x459 ) ;
  assign n4133 = n4121 & n4127 ;
  assign n4134 = ( n4131 & n4132 ) | ( n4131 & n4133 ) | ( n4132 & n4133 ) ;
  assign n4135 = n4130 & n4134 ;
  assign n4136 = n4115 | n4135 ;
  assign n4137 = n4131 & ~n4132 ;
  assign n4138 = ~n4131 & n4132 ;
  assign n4139 = n4137 | n4138 ;
  assign n4140 = ~n4133 & n4139 ;
  assign n4141 = n4133 & ~n4139 ;
  assign n4142 = n4140 | n4141 ;
  assign n4143 = n4134 & n4142 ;
  assign n4144 = n4111 & n4130 ;
  assign n4145 = n4142 & n4144 ;
  assign n4146 = ~n4143 & n4145 ;
  assign n4147 = ~n4136 & n4146 ;
  assign n4148 = n4114 & n4147 ;
  assign n4149 = ~n4143 & n4144 ;
  assign n4150 = ~n4135 & n4142 ;
  assign n4151 = n4115 & ~n4150 ;
  assign n4152 = ( n4149 & n4150 ) | ( n4149 & ~n4151 ) | ( n4150 & ~n4151 ) ;
  assign n4153 = ( n4114 & n4148 ) | ( n4114 & ~n4152 ) | ( n4148 & ~n4152 ) ;
  assign n4154 = n4130 & ~n4134 ;
  assign n4155 = ( n4130 & ~n4142 ) | ( n4130 & n4154 ) | ( ~n4142 & n4154 ) ;
  assign n4156 = n4111 & ~n4112 ;
  assign n4157 = ( ~n4108 & n4111 ) | ( ~n4108 & n4156 ) | ( n4111 & n4156 ) ;
  assign n4158 = ~n4155 & n4157 ;
  assign n4159 = n4155 & ~n4157 ;
  assign n4160 = n4158 | n4159 ;
  assign n4161 = ( x448 & x449 ) | ( x448 & x450 ) | ( x449 & x450 ) ;
  assign n4162 = ( x445 & x446 ) | ( x445 & x447 ) | ( x446 & x447 ) ;
  assign n4163 = n4161 & ~n4162 ;
  assign n4164 = ~n4161 & n4162 ;
  assign n4165 = n4163 | n4164 ;
  assign n4166 = x445 & ~x446 ;
  assign n4167 = ~x445 & x446 ;
  assign n4168 = n4166 | n4167 ;
  assign n4169 = ~x447 & n4168 ;
  assign n4170 = x447 & ~n4168 ;
  assign n4171 = n4169 | n4170 ;
  assign n4172 = x448 & ~x449 ;
  assign n4173 = ~x448 & x449 ;
  assign n4174 = n4172 | n4173 ;
  assign n4175 = ~x450 & n4174 ;
  assign n4176 = x450 & ~n4174 ;
  assign n4177 = n4175 | n4176 ;
  assign n4178 = n4171 & n4177 ;
  assign n4179 = n4165 & ~n4178 ;
  assign n4180 = ~n4165 & n4178 ;
  assign n4181 = n4179 | n4180 ;
  assign n4182 = n4171 & ~n4177 ;
  assign n4183 = ~n4171 & n4177 ;
  assign n4184 = n4182 | n4183 ;
  assign n4185 = ( n4161 & n4162 ) | ( n4161 & n4178 ) | ( n4162 & n4178 ) ;
  assign n4186 = n4184 & ~n4185 ;
  assign n4187 = ( ~n4181 & n4184 ) | ( ~n4181 & n4186 ) | ( n4184 & n4186 ) ;
  assign n4188 = ~x439 & x440 ;
  assign n4189 = x439 & ~x440 ;
  assign n4190 = n4188 | n4189 ;
  assign n4191 = ~x441 & n4190 ;
  assign n4192 = x441 & ~n4190 ;
  assign n4193 = n4191 | n4192 ;
  assign n4194 = ~x442 & x443 ;
  assign n4195 = x442 & ~x443 ;
  assign n4196 = n4194 | n4195 ;
  assign n4197 = ~x444 & n4196 ;
  assign n4198 = x444 & ~n4196 ;
  assign n4199 = n4197 | n4198 ;
  assign n4200 = n4193 & n4199 ;
  assign n4201 = ( x442 & x443 ) | ( x442 & x444 ) | ( x443 & x444 ) ;
  assign n4202 = ( x439 & x440 ) | ( x439 & x441 ) | ( x440 & x441 ) ;
  assign n4203 = ~n4201 & n4202 ;
  assign n4204 = n4201 & ~n4202 ;
  assign n4205 = n4203 | n4204 ;
  assign n4206 = ~n4200 & n4205 ;
  assign n4207 = n4200 & ~n4205 ;
  assign n4208 = n4206 | n4207 ;
  assign n4209 = n4193 & ~n4199 ;
  assign n4210 = ~n4193 & n4199 ;
  assign n4211 = n4209 | n4210 ;
  assign n4212 = ( n4200 & n4201 ) | ( n4200 & n4202 ) | ( n4201 & n4202 ) ;
  assign n4213 = n4211 & ~n4212 ;
  assign n4214 = ( ~n4208 & n4211 ) | ( ~n4208 & n4213 ) | ( n4211 & n4213 ) ;
  assign n4215 = ~n4187 & n4214 ;
  assign n4216 = n4187 & ~n4214 ;
  assign n4217 = n4215 | n4216 ;
  assign n4218 = n4160 & n4217 ;
  assign n4219 = ( n4114 & ~n4115 ) | ( n4114 & n4150 ) | ( ~n4115 & n4150 ) ;
  assign n4220 = n4114 & n4150 ;
  assign n4221 = ( n4149 & n4219 ) | ( n4149 & n4220 ) | ( n4219 & n4220 ) ;
  assign n4222 = n4152 & ~n4221 ;
  assign n4223 = n4218 | n4222 ;
  assign n4224 = n4153 | n4223 ;
  assign n4225 = n4208 & n4212 ;
  assign n4226 = n4184 & n4185 ;
  assign n4227 = n4225 | n4226 ;
  assign n4228 = n4181 & n4185 ;
  assign n4229 = n4184 & n4211 ;
  assign n4230 = n4181 & n4229 ;
  assign n4231 = ~n4228 & n4230 ;
  assign n4232 = ~n4227 & n4231 ;
  assign n4233 = n4211 & n4212 ;
  assign n4234 = n4208 & ~n4233 ;
  assign n4235 = ~n4232 & n4234 ;
  assign n4236 = ~n4228 & n4229 ;
  assign n4237 = n4181 & ~n4226 ;
  assign n4238 = ( n4225 & n4234 ) | ( n4225 & n4237 ) | ( n4234 & n4237 ) ;
  assign n4239 = n4234 | n4237 ;
  assign n4240 = ( ~n4236 & n4238 ) | ( ~n4236 & n4239 ) | ( n4238 & n4239 ) ;
  assign n4241 = n4225 | n4237 ;
  assign n4242 = n4236 & ~n4241 ;
  assign n4243 = ( ~n4237 & n4240 ) | ( ~n4237 & n4242 ) | ( n4240 & n4242 ) ;
  assign n4244 = ( ~n4235 & n4240 ) | ( ~n4235 & n4243 ) | ( n4240 & n4243 ) ;
  assign n4245 = n4224 & n4244 ;
  assign n4246 = n4218 & n4222 ;
  assign n4247 = ( n4153 & n4218 ) | ( n4153 & n4246 ) | ( n4218 & n4246 ) ;
  assign n4248 = n4245 | n4247 ;
  assign n4249 = n4225 & ~n4237 ;
  assign n4250 = ( n4236 & n4237 ) | ( n4236 & ~n4249 ) | ( n4237 & ~n4249 ) ;
  assign n4251 = n4234 & n4250 ;
  assign n4252 = ~n4211 & n4212 ;
  assign n4253 = ( ~n4208 & n4212 ) | ( ~n4208 & n4252 ) | ( n4212 & n4252 ) ;
  assign n4254 = ~n4184 & n4185 ;
  assign n4255 = ( ~n4181 & n4185 ) | ( ~n4181 & n4254 ) | ( n4185 & n4254 ) ;
  assign n4256 = ~n4253 & n4255 ;
  assign n4257 = n4253 & ~n4255 ;
  assign n4258 = n4256 | n4257 ;
  assign n4259 = n4232 | n4258 ;
  assign n4260 = n4251 | n4259 ;
  assign n4261 = n4232 & n4258 ;
  assign n4262 = ( n4251 & n4258 ) | ( n4251 & n4261 ) | ( n4258 & n4261 ) ;
  assign n4263 = n4260 & ~n4262 ;
  assign n4264 = n4114 & n4152 ;
  assign n4265 = ~n4111 & n4112 ;
  assign n4266 = ( ~n4108 & n4112 ) | ( ~n4108 & n4265 ) | ( n4112 & n4265 ) ;
  assign n4267 = ~n4130 & n4134 ;
  assign n4268 = ( n4134 & ~n4142 ) | ( n4134 & n4267 ) | ( ~n4142 & n4267 ) ;
  assign n4269 = ~n4266 & n4268 ;
  assign n4270 = n4266 & ~n4268 ;
  assign n4271 = n4269 | n4270 ;
  assign n4272 = n4147 | n4271 ;
  assign n4273 = n4264 | n4272 ;
  assign n4274 = n4147 & n4271 ;
  assign n4275 = ( n4264 & n4271 ) | ( n4264 & n4274 ) | ( n4271 & n4274 ) ;
  assign n4276 = n4273 & ~n4275 ;
  assign n4277 = n4263 | n4276 ;
  assign n4278 = n4248 & n4277 ;
  assign n4279 = n4260 & n4273 ;
  assign n4280 = n4262 | n4275 ;
  assign n4281 = n4279 & ~n4280 ;
  assign n4282 = ( n4147 & n4266 ) | ( n4147 & n4268 ) | ( n4266 & n4268 ) ;
  assign n4283 = n4266 | n4268 ;
  assign n4284 = ( n4264 & n4282 ) | ( n4264 & n4283 ) | ( n4282 & n4283 ) ;
  assign n4285 = ( n4232 & n4253 ) | ( n4232 & n4255 ) | ( n4253 & n4255 ) ;
  assign n4286 = n4253 | n4255 ;
  assign n4287 = ( n4251 & n4285 ) | ( n4251 & n4286 ) | ( n4285 & n4286 ) ;
  assign n4288 = ~n4284 & n4287 ;
  assign n4289 = n4284 & ~n4287 ;
  assign n4290 = n4288 | n4289 ;
  assign n4291 = n4281 | n4290 ;
  assign n4292 = n4278 | n4291 ;
  assign n4293 = n4277 | n4281 ;
  assign n4294 = ( n4248 & n4281 ) | ( n4248 & n4293 ) | ( n4281 & n4293 ) ;
  assign n4295 = n4290 & n4294 ;
  assign n4296 = n4292 & ~n4295 ;
  assign n4297 = ~x427 & x428 ;
  assign n4298 = x427 & ~x428 ;
  assign n4299 = n4297 | n4298 ;
  assign n4300 = ~x429 & n4299 ;
  assign n4301 = x429 & ~n4299 ;
  assign n4302 = n4300 | n4301 ;
  assign n4303 = ~x430 & x431 ;
  assign n4304 = x430 & ~x431 ;
  assign n4305 = n4303 | n4304 ;
  assign n4306 = ~x432 & n4305 ;
  assign n4307 = x432 & ~n4305 ;
  assign n4308 = n4306 | n4307 ;
  assign n4309 = n4302 & n4308 ;
  assign n4310 = ( x430 & x431 ) | ( x430 & x432 ) | ( x431 & x432 ) ;
  assign n4311 = ( x427 & x428 ) | ( x427 & x429 ) | ( x428 & x429 ) ;
  assign n4312 = ~n4310 & n4311 ;
  assign n4313 = n4310 & ~n4311 ;
  assign n4314 = n4312 | n4313 ;
  assign n4315 = ~n4309 & n4314 ;
  assign n4316 = n4309 & ~n4314 ;
  assign n4317 = n4315 | n4316 ;
  assign n4318 = n4302 & ~n4308 ;
  assign n4319 = ~n4302 & n4308 ;
  assign n4320 = n4318 | n4319 ;
  assign n4321 = ( n4309 & n4310 ) | ( n4309 & n4311 ) | ( n4310 & n4311 ) ;
  assign n4322 = n4320 & n4321 ;
  assign n4323 = n4317 & ~n4322 ;
  assign n4324 = n4317 & n4321 ;
  assign n4325 = x433 & ~x434 ;
  assign n4326 = ~x433 & x434 ;
  assign n4327 = n4325 | n4326 ;
  assign n4328 = ~x435 & n4327 ;
  assign n4329 = x435 & ~n4327 ;
  assign n4330 = n4328 | n4329 ;
  assign n4331 = x436 & ~x437 ;
  assign n4332 = ~x436 & x437 ;
  assign n4333 = n4331 | n4332 ;
  assign n4334 = ~x438 & n4333 ;
  assign n4335 = x438 & ~n4333 ;
  assign n4336 = n4334 | n4335 ;
  assign n4337 = n4330 & ~n4336 ;
  assign n4338 = ~n4330 & n4336 ;
  assign n4339 = n4337 | n4338 ;
  assign n4340 = ( x436 & x437 ) | ( x436 & x438 ) | ( x437 & x438 ) ;
  assign n4341 = ( x433 & x434 ) | ( x433 & x435 ) | ( x434 & x435 ) ;
  assign n4342 = n4330 & n4336 ;
  assign n4343 = ( n4340 & n4341 ) | ( n4340 & n4342 ) | ( n4341 & n4342 ) ;
  assign n4344 = n4339 & n4343 ;
  assign n4345 = n4324 | n4344 ;
  assign n4346 = n4340 & ~n4341 ;
  assign n4347 = ~n4340 & n4341 ;
  assign n4348 = n4346 | n4347 ;
  assign n4349 = ~n4342 & n4348 ;
  assign n4350 = n4342 & ~n4348 ;
  assign n4351 = n4349 | n4350 ;
  assign n4352 = n4343 & n4351 ;
  assign n4353 = n4320 & n4339 ;
  assign n4354 = n4351 & n4353 ;
  assign n4355 = ~n4352 & n4354 ;
  assign n4356 = ~n4345 & n4355 ;
  assign n4357 = n4323 & n4356 ;
  assign n4358 = ~n4352 & n4353 ;
  assign n4359 = ~n4344 & n4351 ;
  assign n4360 = n4324 & ~n4359 ;
  assign n4361 = ( n4358 & n4359 ) | ( n4358 & ~n4360 ) | ( n4359 & ~n4360 ) ;
  assign n4362 = ( n4323 & n4357 ) | ( n4323 & ~n4361 ) | ( n4357 & ~n4361 ) ;
  assign n4363 = n4339 & ~n4343 ;
  assign n4364 = ( n4339 & ~n4351 ) | ( n4339 & n4363 ) | ( ~n4351 & n4363 ) ;
  assign n4365 = n4320 & ~n4321 ;
  assign n4366 = ( ~n4317 & n4320 ) | ( ~n4317 & n4365 ) | ( n4320 & n4365 ) ;
  assign n4367 = ~n4364 & n4366 ;
  assign n4368 = n4364 & ~n4366 ;
  assign n4369 = n4367 | n4368 ;
  assign n4370 = ( x424 & x425 ) | ( x424 & x426 ) | ( x425 & x426 ) ;
  assign n4371 = ( x421 & x422 ) | ( x421 & x423 ) | ( x422 & x423 ) ;
  assign n4372 = n4370 & ~n4371 ;
  assign n4373 = ~n4370 & n4371 ;
  assign n4374 = n4372 | n4373 ;
  assign n4375 = ~x421 & x422 ;
  assign n4376 = x421 & ~x422 ;
  assign n4377 = n4375 | n4376 ;
  assign n4378 = ~x423 & n4377 ;
  assign n4379 = x423 & ~n4377 ;
  assign n4380 = n4378 | n4379 ;
  assign n4381 = ~x424 & x425 ;
  assign n4382 = x424 & ~x425 ;
  assign n4383 = n4381 | n4382 ;
  assign n4384 = ~x426 & n4383 ;
  assign n4385 = x426 & ~n4383 ;
  assign n4386 = n4384 | n4385 ;
  assign n4387 = n4380 & n4386 ;
  assign n4388 = n4374 & ~n4387 ;
  assign n4389 = ~n4374 & n4387 ;
  assign n4390 = n4388 | n4389 ;
  assign n4391 = n4380 & ~n4386 ;
  assign n4392 = ~n4380 & n4386 ;
  assign n4393 = n4391 | n4392 ;
  assign n4394 = ( n4370 & n4371 ) | ( n4370 & n4387 ) | ( n4371 & n4387 ) ;
  assign n4395 = n4393 & ~n4394 ;
  assign n4396 = ( ~n4390 & n4393 ) | ( ~n4390 & n4395 ) | ( n4393 & n4395 ) ;
  assign n4397 = ~x415 & x416 ;
  assign n4398 = x415 & ~x416 ;
  assign n4399 = n4397 | n4398 ;
  assign n4400 = ~x417 & n4399 ;
  assign n4401 = x417 & ~n4399 ;
  assign n4402 = n4400 | n4401 ;
  assign n4403 = ~x418 & x419 ;
  assign n4404 = x418 & ~x419 ;
  assign n4405 = n4403 | n4404 ;
  assign n4406 = ~x420 & n4405 ;
  assign n4407 = x420 & ~n4405 ;
  assign n4408 = n4406 | n4407 ;
  assign n4409 = n4402 & ~n4408 ;
  assign n4410 = ~n4402 & n4408 ;
  assign n4411 = n4409 | n4410 ;
  assign n4412 = ( x418 & x419 ) | ( x418 & x420 ) | ( x419 & x420 ) ;
  assign n4413 = ( x415 & x416 ) | ( x415 & x417 ) | ( x416 & x417 ) ;
  assign n4414 = n4412 & ~n4413 ;
  assign n4415 = ~n4412 & n4413 ;
  assign n4416 = n4414 | n4415 ;
  assign n4417 = n4402 & n4408 ;
  assign n4418 = n4416 & ~n4417 ;
  assign n4419 = ~n4416 & n4417 ;
  assign n4420 = n4418 | n4419 ;
  assign n4421 = ( n4412 & n4413 ) | ( n4412 & n4417 ) | ( n4413 & n4417 ) ;
  assign n4422 = n4411 & ~n4421 ;
  assign n4423 = ( n4411 & ~n4420 ) | ( n4411 & n4422 ) | ( ~n4420 & n4422 ) ;
  assign n4424 = ~n4396 & n4423 ;
  assign n4425 = n4396 & ~n4423 ;
  assign n4426 = n4424 | n4425 ;
  assign n4427 = n4369 & n4426 ;
  assign n4428 = ( n4323 & ~n4324 ) | ( n4323 & n4359 ) | ( ~n4324 & n4359 ) ;
  assign n4429 = n4323 & n4359 ;
  assign n4430 = ( n4358 & n4428 ) | ( n4358 & n4429 ) | ( n4428 & n4429 ) ;
  assign n4431 = n4361 & ~n4430 ;
  assign n4432 = n4427 | n4431 ;
  assign n4433 = n4362 | n4432 ;
  assign n4434 = n4420 & n4421 ;
  assign n4435 = n4393 & n4394 ;
  assign n4436 = n4434 | n4435 ;
  assign n4437 = n4390 & n4394 ;
  assign n4438 = n4393 & n4411 ;
  assign n4439 = n4390 & n4438 ;
  assign n4440 = ~n4437 & n4439 ;
  assign n4441 = ~n4436 & n4440 ;
  assign n4442 = n4411 & n4421 ;
  assign n4443 = n4420 & ~n4442 ;
  assign n4444 = ~n4441 & n4443 ;
  assign n4445 = ~n4437 & n4438 ;
  assign n4446 = n4390 & ~n4435 ;
  assign n4447 = ( n4434 & n4443 ) | ( n4434 & n4446 ) | ( n4443 & n4446 ) ;
  assign n4448 = n4443 | n4446 ;
  assign n4449 = ( ~n4445 & n4447 ) | ( ~n4445 & n4448 ) | ( n4447 & n4448 ) ;
  assign n4450 = n4434 | n4446 ;
  assign n4451 = n4445 & ~n4450 ;
  assign n4452 = ( ~n4446 & n4449 ) | ( ~n4446 & n4451 ) | ( n4449 & n4451 ) ;
  assign n4453 = ( ~n4444 & n4449 ) | ( ~n4444 & n4452 ) | ( n4449 & n4452 ) ;
  assign n4454 = n4433 & n4453 ;
  assign n4455 = n4427 & n4431 ;
  assign n4456 = ( n4362 & n4427 ) | ( n4362 & n4455 ) | ( n4427 & n4455 ) ;
  assign n4457 = n4454 | n4456 ;
  assign n4458 = n4434 & ~n4446 ;
  assign n4459 = ( n4445 & n4446 ) | ( n4445 & ~n4458 ) | ( n4446 & ~n4458 ) ;
  assign n4460 = n4443 & n4459 ;
  assign n4461 = ~n4411 & n4421 ;
  assign n4462 = ( ~n4420 & n4421 ) | ( ~n4420 & n4461 ) | ( n4421 & n4461 ) ;
  assign n4463 = ~n4393 & n4394 ;
  assign n4464 = ( ~n4390 & n4394 ) | ( ~n4390 & n4463 ) | ( n4394 & n4463 ) ;
  assign n4465 = ~n4462 & n4464 ;
  assign n4466 = n4462 & ~n4464 ;
  assign n4467 = n4465 | n4466 ;
  assign n4468 = n4441 | n4467 ;
  assign n4469 = n4460 | n4468 ;
  assign n4470 = n4441 & n4467 ;
  assign n4471 = ( n4460 & n4467 ) | ( n4460 & n4470 ) | ( n4467 & n4470 ) ;
  assign n4472 = n4469 & ~n4471 ;
  assign n4473 = n4323 & n4361 ;
  assign n4474 = ~n4320 & n4321 ;
  assign n4475 = ( ~n4317 & n4321 ) | ( ~n4317 & n4474 ) | ( n4321 & n4474 ) ;
  assign n4476 = ~n4339 & n4343 ;
  assign n4477 = ( n4343 & ~n4351 ) | ( n4343 & n4476 ) | ( ~n4351 & n4476 ) ;
  assign n4478 = ~n4475 & n4477 ;
  assign n4479 = n4475 & ~n4477 ;
  assign n4480 = n4478 | n4479 ;
  assign n4481 = n4356 | n4480 ;
  assign n4482 = n4473 | n4481 ;
  assign n4483 = n4356 & n4480 ;
  assign n4484 = ( n4473 & n4480 ) | ( n4473 & n4483 ) | ( n4480 & n4483 ) ;
  assign n4485 = n4482 & ~n4484 ;
  assign n4486 = n4472 | n4485 ;
  assign n4487 = n4457 & n4486 ;
  assign n4488 = n4469 & n4482 ;
  assign n4489 = n4471 | n4484 ;
  assign n4490 = n4488 & ~n4489 ;
  assign n4491 = ( n4356 & n4475 ) | ( n4356 & n4477 ) | ( n4475 & n4477 ) ;
  assign n4492 = n4475 | n4477 ;
  assign n4493 = ( n4473 & n4491 ) | ( n4473 & n4492 ) | ( n4491 & n4492 ) ;
  assign n4494 = ( n4441 & n4462 ) | ( n4441 & n4464 ) | ( n4462 & n4464 ) ;
  assign n4495 = n4462 | n4464 ;
  assign n4496 = ( n4460 & n4494 ) | ( n4460 & n4495 ) | ( n4494 & n4495 ) ;
  assign n4497 = ~n4493 & n4496 ;
  assign n4498 = n4493 & ~n4496 ;
  assign n4499 = n4497 | n4498 ;
  assign n4500 = n4490 | n4499 ;
  assign n4501 = n4487 | n4500 ;
  assign n4502 = n4486 | n4490 ;
  assign n4503 = ( n4457 & n4490 ) | ( n4457 & n4502 ) | ( n4490 & n4502 ) ;
  assign n4504 = n4499 & n4503 ;
  assign n4505 = n4501 & ~n4504 ;
  assign n4506 = n4296 | n4505 ;
  assign n4507 = n4224 & ~n4247 ;
  assign n4508 = n4244 & ~n4507 ;
  assign n4509 = n4160 & ~n4217 ;
  assign n4510 = ~n4160 & n4217 ;
  assign n4511 = n4509 | n4510 ;
  assign n4512 = n4369 & ~n4426 ;
  assign n4513 = ~n4369 & n4426 ;
  assign n4514 = n4512 | n4513 ;
  assign n4515 = n4511 & n4514 ;
  assign n4516 = ~n4218 & n4224 ;
  assign n4517 = n4224 & ~n4244 ;
  assign n4518 = n4153 | n4222 ;
  assign n4519 = n4244 | n4518 ;
  assign n4520 = ( n4516 & n4517 ) | ( n4516 & ~n4519 ) | ( n4517 & ~n4519 ) ;
  assign n4521 = n4515 | n4520 ;
  assign n4522 = n4508 | n4521 ;
  assign n4523 = n4362 | n4431 ;
  assign n4524 = ( n4427 & n4453 ) | ( n4427 & ~n4523 ) | ( n4453 & ~n4523 ) ;
  assign n4525 = ( ~n4453 & n4523 ) | ( ~n4453 & n4524 ) | ( n4523 & n4524 ) ;
  assign n4526 = ( ~n4427 & n4524 ) | ( ~n4427 & n4525 ) | ( n4524 & n4525 ) ;
  assign n4527 = n4522 & n4526 ;
  assign n4528 = n4508 | n4520 ;
  assign n4529 = n4515 & n4528 ;
  assign n4530 = ( n4456 & ~n4472 ) | ( n4456 & n4485 ) | ( ~n4472 & n4485 ) ;
  assign n4531 = n4472 & ~n4485 ;
  assign n4532 = ( n4454 & n4530 ) | ( n4454 & ~n4531 ) | ( n4530 & ~n4531 ) ;
  assign n4533 = ( ~n4457 & n4472 ) | ( ~n4457 & n4532 ) | ( n4472 & n4532 ) ;
  assign n4534 = ( ~n4485 & n4532 ) | ( ~n4485 & n4533 ) | ( n4532 & n4533 ) ;
  assign n4535 = ( n4247 & ~n4263 ) | ( n4247 & n4276 ) | ( ~n4263 & n4276 ) ;
  assign n4536 = n4263 & ~n4276 ;
  assign n4537 = ( n4245 & n4535 ) | ( n4245 & ~n4536 ) | ( n4535 & ~n4536 ) ;
  assign n4538 = ( ~n4248 & n4263 ) | ( ~n4248 & n4537 ) | ( n4263 & n4537 ) ;
  assign n4539 = ( ~n4276 & n4537 ) | ( ~n4276 & n4538 ) | ( n4537 & n4538 ) ;
  assign n4540 = ( n4529 & n4534 ) | ( n4529 & n4539 ) | ( n4534 & n4539 ) ;
  assign n4541 = n4534 | n4539 ;
  assign n4542 = ( n4527 & n4540 ) | ( n4527 & n4541 ) | ( n4540 & n4541 ) ;
  assign n4543 = n4506 & n4542 ;
  assign n4544 = n4292 & n4501 ;
  assign n4545 = n4295 | n4504 ;
  assign n4546 = n4544 & ~n4545 ;
  assign n4547 = n4493 & n4496 ;
  assign n4548 = n4493 | n4496 ;
  assign n4549 = n4547 | n4548 ;
  assign n4550 = ( n4503 & n4547 ) | ( n4503 & n4549 ) | ( n4547 & n4549 ) ;
  assign n4551 = n4284 & n4287 ;
  assign n4552 = n4284 | n4287 ;
  assign n4553 = n4551 | n4552 ;
  assign n4554 = ( n4294 & n4551 ) | ( n4294 & n4553 ) | ( n4551 & n4553 ) ;
  assign n4555 = n4550 & n4554 ;
  assign n4556 = n4554 & ~n4555 ;
  assign n4557 = ( n4550 & ~n4555 ) | ( n4550 & n4556 ) | ( ~n4555 & n4556 ) ;
  assign n4558 = n4546 | n4557 ;
  assign n4559 = n4543 | n4558 ;
  assign n4560 = n4543 | n4546 ;
  assign n4561 = n4557 & n4560 ;
  assign n4562 = n4559 & ~n4561 ;
  assign n4563 = n4087 | n4562 ;
  assign n4564 = ( ~n4296 & n4505 ) | ( ~n4296 & n4542 ) | ( n4505 & n4542 ) ;
  assign n4565 = ( n4296 & ~n4542 ) | ( n4296 & n4564 ) | ( ~n4542 & n4564 ) ;
  assign n4566 = ( ~n4505 & n4564 ) | ( ~n4505 & n4565 ) | ( n4564 & n4565 ) ;
  assign n4567 = ( ~n3821 & n4030 ) | ( ~n3821 & n4067 ) | ( n4030 & n4067 ) ;
  assign n4568 = ( n3821 & ~n4067 ) | ( n3821 & n4567 ) | ( ~n4067 & n4567 ) ;
  assign n4569 = ( ~n4030 & n4567 ) | ( ~n4030 & n4568 ) | ( n4567 & n4568 ) ;
  assign n4570 = ~n4040 & n4053 ;
  assign n4571 = n4040 & ~n4045 ;
  assign n4572 = ~n4033 & n4571 ;
  assign n4573 = ~n4051 & n4572 ;
  assign n4574 = ( ~n4051 & n4570 ) | ( ~n4051 & n4573 ) | ( n4570 & n4573 ) ;
  assign n4575 = n4052 & ~n4054 ;
  assign n4576 = ( n4051 & n4574 ) | ( n4051 & ~n4575 ) | ( n4574 & ~n4575 ) ;
  assign n4577 = n4511 & ~n4514 ;
  assign n4578 = ~n4511 & n4514 ;
  assign n4579 = n4577 | n4578 ;
  assign n4580 = n4036 & ~n4039 ;
  assign n4581 = ~n4036 & n4039 ;
  assign n4582 = n4580 | n4581 ;
  assign n4583 = n4579 & n4582 ;
  assign n4584 = ~n4522 & n4526 ;
  assign n4585 = ( n4526 & n4529 ) | ( n4526 & n4584 ) | ( n4529 & n4584 ) ;
  assign n4586 = ~n4515 & n4528 ;
  assign n4587 = n4515 & ~n4520 ;
  assign n4588 = ~n4508 & n4587 ;
  assign n4589 = ~n4526 & n4588 ;
  assign n4590 = ( ~n4526 & n4586 ) | ( ~n4526 & n4589 ) | ( n4586 & n4589 ) ;
  assign n4591 = n4585 | n4590 ;
  assign n4592 = n4583 | n4591 ;
  assign n4593 = n4576 & n4592 ;
  assign n4594 = n4583 & n4591 ;
  assign n4596 = ( n4054 & ~n4059 ) | ( n4054 & n4064 ) | ( ~n4059 & n4064 ) ;
  assign n4597 = n4059 & ~n4064 ;
  assign n4598 = ( n4052 & n4596 ) | ( n4052 & ~n4597 ) | ( n4596 & ~n4597 ) ;
  assign n4595 = n4052 | n4054 ;
  assign n4599 = ( n4059 & ~n4595 ) | ( n4059 & n4598 ) | ( ~n4595 & n4598 ) ;
  assign n4600 = ( ~n4064 & n4598 ) | ( ~n4064 & n4599 ) | ( n4598 & n4599 ) ;
  assign n4602 = ( n4529 & ~n4534 ) | ( n4529 & n4539 ) | ( ~n4534 & n4539 ) ;
  assign n4603 = n4534 & ~n4539 ;
  assign n4604 = ( n4527 & n4602 ) | ( n4527 & ~n4603 ) | ( n4602 & ~n4603 ) ;
  assign n4601 = n4527 | n4529 ;
  assign n4605 = ( n4534 & ~n4601 ) | ( n4534 & n4604 ) | ( ~n4601 & n4604 ) ;
  assign n4606 = ( ~n4539 & n4604 ) | ( ~n4539 & n4605 ) | ( n4604 & n4605 ) ;
  assign n4607 = ( n4594 & n4600 ) | ( n4594 & n4606 ) | ( n4600 & n4606 ) ;
  assign n4608 = n4600 | n4606 ;
  assign n4609 = ( n4593 & n4607 ) | ( n4593 & n4608 ) | ( n4607 & n4608 ) ;
  assign n4610 = ( n4566 & n4569 ) | ( n4566 & n4609 ) | ( n4569 & n4609 ) ;
  assign n4611 = n4563 & n4610 ;
  assign n4612 = n4084 & n4559 ;
  assign n4613 = n4086 | n4561 ;
  assign n4614 = n4612 & ~n4613 ;
  assign n4623 = n3819 & n4077 ;
  assign n4624 = n4021 | n4076 ;
  assign n4625 = n4018 | n4076 ;
  assign n4626 = ( n4028 & n4624 ) | ( n4028 & n4625 ) | ( n4624 & n4625 ) ;
  assign n4627 = n4623 | n4626 ;
  assign n4628 = n4080 | n4627 ;
  assign n4629 = ( n4071 & n4080 ) | ( n4071 & n4628 ) | ( n4080 & n4628 ) ;
  assign n4630 = n4080 | n4628 ;
  assign n4631 = ( n4068 & n4629 ) | ( n4068 & n4630 ) | ( n4629 & n4630 ) ;
  assign n4615 = n4294 & n4552 ;
  assign n4616 = n4496 | n4551 ;
  assign n4617 = n4493 | n4551 ;
  assign n4618 = ( n4503 & n4616 ) | ( n4503 & n4617 ) | ( n4616 & n4617 ) ;
  assign n4619 = n4615 | n4618 ;
  assign n4620 = n4546 & n4619 ;
  assign n4621 = ( n4543 & n4619 ) | ( n4543 & n4620 ) | ( n4619 & n4620 ) ;
  assign n4622 = n4555 | n4621 ;
  assign n4632 = n4622 & n4631 ;
  assign n4633 = n4622 & ~n4632 ;
  assign n4634 = ( n4631 & ~n4632 ) | ( n4631 & n4633 ) | ( ~n4632 & n4633 ) ;
  assign n4635 = n4614 | n4634 ;
  assign n4636 = n4611 | n4635 ;
  assign n4637 = n4611 | n4614 ;
  assign n4638 = n4634 & n4637 ;
  assign n4639 = n4636 & ~n4638 ;
  assign n4640 = ( x310 & x311 ) | ( x310 & x312 ) | ( x311 & x312 ) ;
  assign n4641 = ( x307 & x308 ) | ( x307 & x309 ) | ( x308 & x309 ) ;
  assign n4642 = n4640 & ~n4641 ;
  assign n4643 = ~n4640 & n4641 ;
  assign n4644 = n4642 | n4643 ;
  assign n4645 = ~x307 & x308 ;
  assign n4646 = x307 & ~x308 ;
  assign n4647 = n4645 | n4646 ;
  assign n4648 = ~x309 & n4647 ;
  assign n4649 = x309 & ~n4647 ;
  assign n4650 = n4648 | n4649 ;
  assign n4651 = ~x310 & x311 ;
  assign n4652 = x310 & ~x311 ;
  assign n4653 = n4651 | n4652 ;
  assign n4654 = ~x312 & n4653 ;
  assign n4655 = x312 & ~n4653 ;
  assign n4656 = n4654 | n4655 ;
  assign n4657 = n4650 & n4656 ;
  assign n4658 = n4644 & ~n4657 ;
  assign n4659 = ~n4644 & n4657 ;
  assign n4660 = n4658 | n4659 ;
  assign n4661 = n4650 & ~n4656 ;
  assign n4662 = ~n4650 & n4656 ;
  assign n4663 = n4661 | n4662 ;
  assign n4664 = ( n4640 & n4641 ) | ( n4640 & n4657 ) | ( n4641 & n4657 ) ;
  assign n4665 = n4663 & n4664 ;
  assign n4666 = n4660 & ~n4665 ;
  assign n4667 = n4660 & n4664 ;
  assign n4668 = ~x313 & x314 ;
  assign n4669 = x313 & ~x314 ;
  assign n4670 = n4668 | n4669 ;
  assign n4671 = ~x315 & n4670 ;
  assign n4672 = x315 & ~n4670 ;
  assign n4673 = n4671 | n4672 ;
  assign n4674 = ~x316 & x317 ;
  assign n4675 = x316 & ~x317 ;
  assign n4676 = n4674 | n4675 ;
  assign n4677 = ~x318 & n4676 ;
  assign n4678 = x318 & ~n4676 ;
  assign n4679 = n4677 | n4678 ;
  assign n4680 = n4673 & ~n4679 ;
  assign n4681 = ~n4673 & n4679 ;
  assign n4682 = n4680 | n4681 ;
  assign n4683 = ( x316 & x317 ) | ( x316 & x318 ) | ( x317 & x318 ) ;
  assign n4684 = ( x313 & x314 ) | ( x313 & x315 ) | ( x314 & x315 ) ;
  assign n4685 = n4673 & n4679 ;
  assign n4686 = ( n4683 & n4684 ) | ( n4683 & n4685 ) | ( n4684 & n4685 ) ;
  assign n4687 = n4682 & n4686 ;
  assign n4688 = n4667 | n4687 ;
  assign n4689 = n4683 & ~n4684 ;
  assign n4690 = ~n4683 & n4684 ;
  assign n4691 = n4689 | n4690 ;
  assign n4692 = ~n4685 & n4691 ;
  assign n4693 = n4685 & ~n4691 ;
  assign n4694 = n4692 | n4693 ;
  assign n4695 = n4686 & n4694 ;
  assign n4696 = n4663 & n4682 ;
  assign n4697 = n4694 & n4696 ;
  assign n4698 = ~n4695 & n4697 ;
  assign n4699 = ~n4688 & n4698 ;
  assign n4700 = n4666 & n4699 ;
  assign n4701 = ~n4695 & n4696 ;
  assign n4702 = ~n4687 & n4694 ;
  assign n4703 = n4667 & ~n4702 ;
  assign n4704 = ( n4701 & n4702 ) | ( n4701 & ~n4703 ) | ( n4702 & ~n4703 ) ;
  assign n4705 = ( n4666 & n4700 ) | ( n4666 & ~n4704 ) | ( n4700 & ~n4704 ) ;
  assign n4706 = n4682 & ~n4686 ;
  assign n4707 = ( n4682 & ~n4694 ) | ( n4682 & n4706 ) | ( ~n4694 & n4706 ) ;
  assign n4708 = n4663 & ~n4664 ;
  assign n4709 = ( ~n4660 & n4663 ) | ( ~n4660 & n4708 ) | ( n4663 & n4708 ) ;
  assign n4710 = ~n4707 & n4709 ;
  assign n4711 = n4707 & ~n4709 ;
  assign n4712 = n4710 | n4711 ;
  assign n4713 = ( x304 & x305 ) | ( x304 & x306 ) | ( x305 & x306 ) ;
  assign n4714 = ( x301 & x302 ) | ( x301 & x303 ) | ( x302 & x303 ) ;
  assign n4715 = n4713 & ~n4714 ;
  assign n4716 = ~n4713 & n4714 ;
  assign n4717 = n4715 | n4716 ;
  assign n4718 = ~x301 & x302 ;
  assign n4719 = x301 & ~x302 ;
  assign n4720 = n4718 | n4719 ;
  assign n4721 = ~x303 & n4720 ;
  assign n4722 = x303 & ~n4720 ;
  assign n4723 = n4721 | n4722 ;
  assign n4724 = ~x304 & x305 ;
  assign n4725 = x304 & ~x305 ;
  assign n4726 = n4724 | n4725 ;
  assign n4727 = ~x306 & n4726 ;
  assign n4728 = x306 & ~n4726 ;
  assign n4729 = n4727 | n4728 ;
  assign n4730 = n4723 & n4729 ;
  assign n4731 = n4717 & ~n4730 ;
  assign n4732 = ~n4717 & n4730 ;
  assign n4733 = n4731 | n4732 ;
  assign n4734 = n4723 & ~n4729 ;
  assign n4735 = ~n4723 & n4729 ;
  assign n4736 = n4734 | n4735 ;
  assign n4737 = ( n4713 & n4714 ) | ( n4713 & n4730 ) | ( n4714 & n4730 ) ;
  assign n4738 = n4736 & ~n4737 ;
  assign n4739 = ( ~n4733 & n4736 ) | ( ~n4733 & n4738 ) | ( n4736 & n4738 ) ;
  assign n4740 = ~x295 & x296 ;
  assign n4741 = x295 & ~x296 ;
  assign n4742 = n4740 | n4741 ;
  assign n4743 = ~x297 & n4742 ;
  assign n4744 = x297 & ~n4742 ;
  assign n4745 = n4743 | n4744 ;
  assign n4746 = ~x298 & x299 ;
  assign n4747 = x298 & ~x299 ;
  assign n4748 = n4746 | n4747 ;
  assign n4749 = ~x300 & n4748 ;
  assign n4750 = x300 & ~n4748 ;
  assign n4751 = n4749 | n4750 ;
  assign n4752 = n4745 & ~n4751 ;
  assign n4753 = ~n4745 & n4751 ;
  assign n4754 = n4752 | n4753 ;
  assign n4755 = ( x298 & x299 ) | ( x298 & x300 ) | ( x299 & x300 ) ;
  assign n4756 = ( x295 & x296 ) | ( x295 & x297 ) | ( x296 & x297 ) ;
  assign n4757 = n4755 & ~n4756 ;
  assign n4758 = ~n4755 & n4756 ;
  assign n4759 = n4757 | n4758 ;
  assign n4760 = n4745 & n4751 ;
  assign n4761 = n4759 & ~n4760 ;
  assign n4762 = ~n4759 & n4760 ;
  assign n4763 = n4761 | n4762 ;
  assign n4764 = ( n4755 & n4756 ) | ( n4755 & n4760 ) | ( n4756 & n4760 ) ;
  assign n4765 = n4754 & ~n4764 ;
  assign n4766 = ( n4754 & ~n4763 ) | ( n4754 & n4765 ) | ( ~n4763 & n4765 ) ;
  assign n4767 = ~n4739 & n4766 ;
  assign n4768 = n4739 & ~n4766 ;
  assign n4769 = n4767 | n4768 ;
  assign n4770 = n4712 & n4769 ;
  assign n4771 = ( n4666 & ~n4667 ) | ( n4666 & n4702 ) | ( ~n4667 & n4702 ) ;
  assign n4772 = n4666 & n4702 ;
  assign n4773 = ( n4701 & n4771 ) | ( n4701 & n4772 ) | ( n4771 & n4772 ) ;
  assign n4774 = n4704 & ~n4773 ;
  assign n4775 = n4770 | n4774 ;
  assign n4776 = n4705 | n4775 ;
  assign n4777 = n4763 & n4764 ;
  assign n4778 = n4736 & n4737 ;
  assign n4779 = n4777 | n4778 ;
  assign n4780 = n4733 & n4737 ;
  assign n4781 = n4736 & n4754 ;
  assign n4782 = n4733 & n4781 ;
  assign n4783 = ~n4780 & n4782 ;
  assign n4784 = ~n4779 & n4783 ;
  assign n4785 = n4754 & n4764 ;
  assign n4786 = n4763 & ~n4785 ;
  assign n4787 = ~n4784 & n4786 ;
  assign n4788 = ~n4780 & n4781 ;
  assign n4789 = n4733 & ~n4778 ;
  assign n4790 = ( n4777 & n4786 ) | ( n4777 & n4789 ) | ( n4786 & n4789 ) ;
  assign n4791 = n4786 | n4789 ;
  assign n4792 = ( ~n4788 & n4790 ) | ( ~n4788 & n4791 ) | ( n4790 & n4791 ) ;
  assign n4793 = n4777 | n4789 ;
  assign n4794 = n4788 & ~n4793 ;
  assign n4795 = ( ~n4789 & n4792 ) | ( ~n4789 & n4794 ) | ( n4792 & n4794 ) ;
  assign n4796 = ( ~n4787 & n4792 ) | ( ~n4787 & n4795 ) | ( n4792 & n4795 ) ;
  assign n4797 = n4776 & n4796 ;
  assign n4798 = n4770 & n4774 ;
  assign n4799 = ( n4705 & n4770 ) | ( n4705 & n4798 ) | ( n4770 & n4798 ) ;
  assign n4800 = n4797 | n4799 ;
  assign n4801 = n4777 & ~n4789 ;
  assign n4802 = ( n4788 & n4789 ) | ( n4788 & ~n4801 ) | ( n4789 & ~n4801 ) ;
  assign n4803 = n4786 & n4802 ;
  assign n4804 = ~n4754 & n4764 ;
  assign n4805 = ( ~n4763 & n4764 ) | ( ~n4763 & n4804 ) | ( n4764 & n4804 ) ;
  assign n4806 = ~n4736 & n4737 ;
  assign n4807 = ( ~n4733 & n4737 ) | ( ~n4733 & n4806 ) | ( n4737 & n4806 ) ;
  assign n4808 = ~n4805 & n4807 ;
  assign n4809 = n4805 & ~n4807 ;
  assign n4810 = n4808 | n4809 ;
  assign n4811 = n4784 | n4810 ;
  assign n4812 = n4803 | n4811 ;
  assign n4813 = n4784 & n4810 ;
  assign n4814 = ( n4803 & n4810 ) | ( n4803 & n4813 ) | ( n4810 & n4813 ) ;
  assign n4815 = n4812 & ~n4814 ;
  assign n4816 = n4666 & n4704 ;
  assign n4817 = ~n4663 & n4664 ;
  assign n4818 = ( ~n4660 & n4664 ) | ( ~n4660 & n4817 ) | ( n4664 & n4817 ) ;
  assign n4819 = ~n4682 & n4686 ;
  assign n4820 = ( n4686 & ~n4694 ) | ( n4686 & n4819 ) | ( ~n4694 & n4819 ) ;
  assign n4821 = ~n4818 & n4820 ;
  assign n4822 = n4818 & ~n4820 ;
  assign n4823 = n4821 | n4822 ;
  assign n4824 = n4699 | n4823 ;
  assign n4825 = n4816 | n4824 ;
  assign n4826 = n4699 & n4823 ;
  assign n4827 = ( n4816 & n4823 ) | ( n4816 & n4826 ) | ( n4823 & n4826 ) ;
  assign n4828 = n4825 & ~n4827 ;
  assign n4829 = n4815 | n4828 ;
  assign n4830 = n4800 & n4829 ;
  assign n4831 = n4812 & n4825 ;
  assign n4832 = n4814 | n4827 ;
  assign n4833 = n4831 & ~n4832 ;
  assign n4834 = ( n4699 & n4818 ) | ( n4699 & n4820 ) | ( n4818 & n4820 ) ;
  assign n4835 = n4818 | n4820 ;
  assign n4836 = ( n4816 & n4834 ) | ( n4816 & n4835 ) | ( n4834 & n4835 ) ;
  assign n4837 = ( n4784 & n4805 ) | ( n4784 & n4807 ) | ( n4805 & n4807 ) ;
  assign n4838 = n4805 | n4807 ;
  assign n4839 = ( n4803 & n4837 ) | ( n4803 & n4838 ) | ( n4837 & n4838 ) ;
  assign n4840 = ~n4836 & n4839 ;
  assign n4841 = n4836 & ~n4839 ;
  assign n4842 = n4840 | n4841 ;
  assign n4843 = n4833 | n4842 ;
  assign n4844 = n4830 | n4843 ;
  assign n4845 = n4829 | n4833 ;
  assign n4846 = ( n4800 & n4833 ) | ( n4800 & n4845 ) | ( n4833 & n4845 ) ;
  assign n4847 = n4842 & n4846 ;
  assign n4848 = n4844 & ~n4847 ;
  assign n4849 = ( x286 & x287 ) | ( x286 & x288 ) | ( x287 & x288 ) ;
  assign n4850 = ( x283 & x284 ) | ( x283 & x285 ) | ( x284 & x285 ) ;
  assign n4851 = n4849 & ~n4850 ;
  assign n4852 = ~n4849 & n4850 ;
  assign n4853 = n4851 | n4852 ;
  assign n4854 = ~x283 & x284 ;
  assign n4855 = x283 & ~x284 ;
  assign n4856 = n4854 | n4855 ;
  assign n4857 = ~x285 & n4856 ;
  assign n4858 = x285 & ~n4856 ;
  assign n4859 = n4857 | n4858 ;
  assign n4860 = ~x286 & x287 ;
  assign n4861 = x286 & ~x287 ;
  assign n4862 = n4860 | n4861 ;
  assign n4863 = ~x288 & n4862 ;
  assign n4864 = x288 & ~n4862 ;
  assign n4865 = n4863 | n4864 ;
  assign n4866 = n4859 & n4865 ;
  assign n4867 = n4853 & ~n4866 ;
  assign n4868 = ~n4853 & n4866 ;
  assign n4869 = n4867 | n4868 ;
  assign n4870 = n4859 & ~n4865 ;
  assign n4871 = ~n4859 & n4865 ;
  assign n4872 = n4870 | n4871 ;
  assign n4873 = ( n4849 & n4850 ) | ( n4849 & n4866 ) | ( n4850 & n4866 ) ;
  assign n4874 = n4872 & n4873 ;
  assign n4875 = n4869 & ~n4874 ;
  assign n4876 = n4869 & n4873 ;
  assign n4877 = ~x289 & x290 ;
  assign n4878 = x289 & ~x290 ;
  assign n4879 = n4877 | n4878 ;
  assign n4880 = ~x291 & n4879 ;
  assign n4881 = x291 & ~n4879 ;
  assign n4882 = n4880 | n4881 ;
  assign n4883 = ~x292 & x293 ;
  assign n4884 = x292 & ~x293 ;
  assign n4885 = n4883 | n4884 ;
  assign n4886 = ~x294 & n4885 ;
  assign n4887 = x294 & ~n4885 ;
  assign n4888 = n4886 | n4887 ;
  assign n4889 = n4882 & ~n4888 ;
  assign n4890 = ~n4882 & n4888 ;
  assign n4891 = n4889 | n4890 ;
  assign n4892 = ( x292 & x293 ) | ( x292 & x294 ) | ( x293 & x294 ) ;
  assign n4893 = ( x289 & x290 ) | ( x289 & x291 ) | ( x290 & x291 ) ;
  assign n4894 = n4882 & n4888 ;
  assign n4895 = ( n4892 & n4893 ) | ( n4892 & n4894 ) | ( n4893 & n4894 ) ;
  assign n4896 = n4891 & n4895 ;
  assign n4897 = n4876 | n4896 ;
  assign n4898 = n4892 & ~n4893 ;
  assign n4899 = ~n4892 & n4893 ;
  assign n4900 = n4898 | n4899 ;
  assign n4901 = ~n4894 & n4900 ;
  assign n4902 = n4894 & ~n4900 ;
  assign n4903 = n4901 | n4902 ;
  assign n4904 = n4895 & n4903 ;
  assign n4905 = n4872 & n4891 ;
  assign n4906 = n4903 & n4905 ;
  assign n4907 = ~n4904 & n4906 ;
  assign n4908 = ~n4897 & n4907 ;
  assign n4909 = n4875 & n4908 ;
  assign n4910 = ~n4904 & n4905 ;
  assign n4911 = ~n4896 & n4903 ;
  assign n4912 = n4876 & ~n4911 ;
  assign n4913 = ( n4910 & n4911 ) | ( n4910 & ~n4912 ) | ( n4911 & ~n4912 ) ;
  assign n4914 = ( n4875 & n4909 ) | ( n4875 & ~n4913 ) | ( n4909 & ~n4913 ) ;
  assign n4915 = n4891 & ~n4895 ;
  assign n4916 = ( n4891 & ~n4903 ) | ( n4891 & n4915 ) | ( ~n4903 & n4915 ) ;
  assign n4917 = n4872 & ~n4873 ;
  assign n4918 = ( ~n4869 & n4872 ) | ( ~n4869 & n4917 ) | ( n4872 & n4917 ) ;
  assign n4919 = ~n4916 & n4918 ;
  assign n4920 = n4916 & ~n4918 ;
  assign n4921 = n4919 | n4920 ;
  assign n4922 = ( x280 & x281 ) | ( x280 & x282 ) | ( x281 & x282 ) ;
  assign n4923 = ( x277 & x278 ) | ( x277 & x279 ) | ( x278 & x279 ) ;
  assign n4924 = n4922 & ~n4923 ;
  assign n4925 = ~n4922 & n4923 ;
  assign n4926 = n4924 | n4925 ;
  assign n4927 = ~x277 & x278 ;
  assign n4928 = x277 & ~x278 ;
  assign n4929 = n4927 | n4928 ;
  assign n4930 = ~x279 & n4929 ;
  assign n4931 = x279 & ~n4929 ;
  assign n4932 = n4930 | n4931 ;
  assign n4933 = ~x280 & x281 ;
  assign n4934 = x280 & ~x281 ;
  assign n4935 = n4933 | n4934 ;
  assign n4936 = ~x282 & n4935 ;
  assign n4937 = x282 & ~n4935 ;
  assign n4938 = n4936 | n4937 ;
  assign n4939 = n4932 & n4938 ;
  assign n4940 = n4926 & ~n4939 ;
  assign n4941 = ~n4926 & n4939 ;
  assign n4942 = n4940 | n4941 ;
  assign n4943 = n4932 & ~n4938 ;
  assign n4944 = ~n4932 & n4938 ;
  assign n4945 = n4943 | n4944 ;
  assign n4946 = ( n4922 & n4923 ) | ( n4922 & n4939 ) | ( n4923 & n4939 ) ;
  assign n4947 = n4945 & ~n4946 ;
  assign n4948 = ( ~n4942 & n4945 ) | ( ~n4942 & n4947 ) | ( n4945 & n4947 ) ;
  assign n4949 = ~x271 & x272 ;
  assign n4950 = x271 & ~x272 ;
  assign n4951 = n4949 | n4950 ;
  assign n4952 = ~x273 & n4951 ;
  assign n4953 = x273 & ~n4951 ;
  assign n4954 = n4952 | n4953 ;
  assign n4955 = ~x274 & x275 ;
  assign n4956 = x274 & ~x275 ;
  assign n4957 = n4955 | n4956 ;
  assign n4958 = ~x276 & n4957 ;
  assign n4959 = x276 & ~n4957 ;
  assign n4960 = n4958 | n4959 ;
  assign n4961 = n4954 & ~n4960 ;
  assign n4962 = ~n4954 & n4960 ;
  assign n4963 = n4961 | n4962 ;
  assign n4964 = ( x274 & x275 ) | ( x274 & x276 ) | ( x275 & x276 ) ;
  assign n4965 = ( x271 & x272 ) | ( x271 & x273 ) | ( x272 & x273 ) ;
  assign n4966 = n4964 & ~n4965 ;
  assign n4967 = ~n4964 & n4965 ;
  assign n4968 = n4966 | n4967 ;
  assign n4969 = n4954 & n4960 ;
  assign n4970 = n4968 & ~n4969 ;
  assign n4971 = ~n4968 & n4969 ;
  assign n4972 = n4970 | n4971 ;
  assign n4973 = ( n4964 & n4965 ) | ( n4964 & n4969 ) | ( n4965 & n4969 ) ;
  assign n4974 = n4963 & ~n4973 ;
  assign n4975 = ( n4963 & ~n4972 ) | ( n4963 & n4974 ) | ( ~n4972 & n4974 ) ;
  assign n4976 = ~n4948 & n4975 ;
  assign n4977 = n4948 & ~n4975 ;
  assign n4978 = n4976 | n4977 ;
  assign n4979 = n4921 & n4978 ;
  assign n4980 = ( n4875 & ~n4876 ) | ( n4875 & n4911 ) | ( ~n4876 & n4911 ) ;
  assign n4981 = n4875 & n4911 ;
  assign n4982 = ( n4910 & n4980 ) | ( n4910 & n4981 ) | ( n4980 & n4981 ) ;
  assign n4983 = n4913 & ~n4982 ;
  assign n4984 = n4979 | n4983 ;
  assign n4985 = n4914 | n4984 ;
  assign n4986 = n4972 & n4973 ;
  assign n4987 = n4945 & n4946 ;
  assign n4988 = n4986 | n4987 ;
  assign n4989 = n4942 & n4946 ;
  assign n4990 = n4945 & n4963 ;
  assign n4991 = n4942 & n4990 ;
  assign n4992 = ~n4989 & n4991 ;
  assign n4993 = ~n4988 & n4992 ;
  assign n4994 = n4963 & n4973 ;
  assign n4995 = n4972 & ~n4994 ;
  assign n4996 = ~n4993 & n4995 ;
  assign n4997 = ~n4989 & n4990 ;
  assign n4998 = n4942 & ~n4987 ;
  assign n4999 = ( n4986 & n4995 ) | ( n4986 & n4998 ) | ( n4995 & n4998 ) ;
  assign n5000 = n4995 | n4998 ;
  assign n5001 = ( ~n4997 & n4999 ) | ( ~n4997 & n5000 ) | ( n4999 & n5000 ) ;
  assign n5002 = n4986 | n4998 ;
  assign n5003 = n4997 & ~n5002 ;
  assign n5004 = ( ~n4998 & n5001 ) | ( ~n4998 & n5003 ) | ( n5001 & n5003 ) ;
  assign n5005 = ( ~n4996 & n5001 ) | ( ~n4996 & n5004 ) | ( n5001 & n5004 ) ;
  assign n5006 = n4985 & n5005 ;
  assign n5007 = n4979 & n4983 ;
  assign n5008 = ( n4914 & n4979 ) | ( n4914 & n5007 ) | ( n4979 & n5007 ) ;
  assign n5009 = n5006 | n5008 ;
  assign n5010 = n4986 & ~n4998 ;
  assign n5011 = ( n4997 & n4998 ) | ( n4997 & ~n5010 ) | ( n4998 & ~n5010 ) ;
  assign n5012 = n4995 & n5011 ;
  assign n5013 = ~n4963 & n4973 ;
  assign n5014 = ( ~n4972 & n4973 ) | ( ~n4972 & n5013 ) | ( n4973 & n5013 ) ;
  assign n5015 = ~n4945 & n4946 ;
  assign n5016 = ( ~n4942 & n4946 ) | ( ~n4942 & n5015 ) | ( n4946 & n5015 ) ;
  assign n5017 = ~n5014 & n5016 ;
  assign n5018 = n5014 & ~n5016 ;
  assign n5019 = n5017 | n5018 ;
  assign n5020 = n4993 | n5019 ;
  assign n5021 = n5012 | n5020 ;
  assign n5022 = n4993 & n5019 ;
  assign n5023 = ( n5012 & n5019 ) | ( n5012 & n5022 ) | ( n5019 & n5022 ) ;
  assign n5024 = n5021 & ~n5023 ;
  assign n5025 = n4875 & n4913 ;
  assign n5026 = ~n4872 & n4873 ;
  assign n5027 = ( ~n4869 & n4873 ) | ( ~n4869 & n5026 ) | ( n4873 & n5026 ) ;
  assign n5028 = ~n4891 & n4895 ;
  assign n5029 = ( n4895 & ~n4903 ) | ( n4895 & n5028 ) | ( ~n4903 & n5028 ) ;
  assign n5030 = ~n5027 & n5029 ;
  assign n5031 = n5027 & ~n5029 ;
  assign n5032 = n5030 | n5031 ;
  assign n5033 = n4908 | n5032 ;
  assign n5034 = n5025 | n5033 ;
  assign n5035 = n4908 & n5032 ;
  assign n5036 = ( n5025 & n5032 ) | ( n5025 & n5035 ) | ( n5032 & n5035 ) ;
  assign n5037 = n5034 & ~n5036 ;
  assign n5038 = n5024 | n5037 ;
  assign n5039 = n5009 & n5038 ;
  assign n5040 = n5021 & n5034 ;
  assign n5041 = n5023 | n5036 ;
  assign n5042 = n5040 & ~n5041 ;
  assign n5043 = ( n4908 & n5027 ) | ( n4908 & n5029 ) | ( n5027 & n5029 ) ;
  assign n5044 = n5027 | n5029 ;
  assign n5045 = ( n5025 & n5043 ) | ( n5025 & n5044 ) | ( n5043 & n5044 ) ;
  assign n5046 = ( n4993 & n5014 ) | ( n4993 & n5016 ) | ( n5014 & n5016 ) ;
  assign n5047 = n5014 | n5016 ;
  assign n5048 = ( n5012 & n5046 ) | ( n5012 & n5047 ) | ( n5046 & n5047 ) ;
  assign n5049 = ~n5045 & n5048 ;
  assign n5050 = n5045 & ~n5048 ;
  assign n5051 = n5049 | n5050 ;
  assign n5052 = n5042 | n5051 ;
  assign n5053 = n5039 | n5052 ;
  assign n5054 = n5038 | n5042 ;
  assign n5055 = ( n5009 & n5042 ) | ( n5009 & n5054 ) | ( n5042 & n5054 ) ;
  assign n5056 = n5051 & n5055 ;
  assign n5057 = n5053 & ~n5056 ;
  assign n5058 = n4848 | n5057 ;
  assign n5059 = n4776 & ~n4799 ;
  assign n5060 = n4796 & ~n5059 ;
  assign n5061 = n4712 & ~n4769 ;
  assign n5062 = ~n4712 & n4769 ;
  assign n5063 = n5061 | n5062 ;
  assign n5064 = n4921 & ~n4978 ;
  assign n5065 = ~n4921 & n4978 ;
  assign n5066 = n5064 | n5065 ;
  assign n5067 = n5063 & n5066 ;
  assign n5068 = ~n4770 & n4776 ;
  assign n5069 = n4776 & ~n4796 ;
  assign n5070 = n4705 | n4774 ;
  assign n5071 = n4796 | n5070 ;
  assign n5072 = ( n5068 & n5069 ) | ( n5068 & ~n5071 ) | ( n5069 & ~n5071 ) ;
  assign n5073 = n5067 | n5072 ;
  assign n5074 = n5060 | n5073 ;
  assign n5075 = n4914 | n4983 ;
  assign n5076 = ( n4979 & n5005 ) | ( n4979 & ~n5075 ) | ( n5005 & ~n5075 ) ;
  assign n5077 = ( ~n5005 & n5075 ) | ( ~n5005 & n5076 ) | ( n5075 & n5076 ) ;
  assign n5078 = ( ~n4979 & n5076 ) | ( ~n4979 & n5077 ) | ( n5076 & n5077 ) ;
  assign n5079 = n5074 & n5078 ;
  assign n5080 = n5060 | n5072 ;
  assign n5081 = n5067 & n5080 ;
  assign n5082 = ( n5008 & ~n5024 ) | ( n5008 & n5037 ) | ( ~n5024 & n5037 ) ;
  assign n5083 = n5024 & ~n5037 ;
  assign n5084 = ( n5006 & n5082 ) | ( n5006 & ~n5083 ) | ( n5082 & ~n5083 ) ;
  assign n5085 = ( ~n5009 & n5024 ) | ( ~n5009 & n5084 ) | ( n5024 & n5084 ) ;
  assign n5086 = ( ~n5037 & n5084 ) | ( ~n5037 & n5085 ) | ( n5084 & n5085 ) ;
  assign n5087 = ( n4799 & ~n4815 ) | ( n4799 & n4828 ) | ( ~n4815 & n4828 ) ;
  assign n5088 = n4815 & ~n4828 ;
  assign n5089 = ( n4797 & n5087 ) | ( n4797 & ~n5088 ) | ( n5087 & ~n5088 ) ;
  assign n5090 = ( ~n4800 & n4815 ) | ( ~n4800 & n5089 ) | ( n4815 & n5089 ) ;
  assign n5091 = ( ~n4828 & n5089 ) | ( ~n4828 & n5090 ) | ( n5089 & n5090 ) ;
  assign n5092 = ( n5081 & n5086 ) | ( n5081 & n5091 ) | ( n5086 & n5091 ) ;
  assign n5093 = n5086 | n5091 ;
  assign n5094 = ( n5079 & n5092 ) | ( n5079 & n5093 ) | ( n5092 & n5093 ) ;
  assign n5095 = n5058 & n5094 ;
  assign n5096 = n4844 & n5053 ;
  assign n5097 = n4847 | n5056 ;
  assign n5098 = n5096 & ~n5097 ;
  assign n5099 = n5045 & n5048 ;
  assign n5100 = n5045 | n5048 ;
  assign n5101 = n5099 | n5100 ;
  assign n5102 = ( n5055 & n5099 ) | ( n5055 & n5101 ) | ( n5099 & n5101 ) ;
  assign n5103 = n4836 & n4839 ;
  assign n5104 = n4836 | n4839 ;
  assign n5105 = n5103 | n5104 ;
  assign n5106 = ( n4846 & n5103 ) | ( n4846 & n5105 ) | ( n5103 & n5105 ) ;
  assign n5107 = n5102 & n5106 ;
  assign n5108 = n5106 & ~n5107 ;
  assign n5109 = ( n5102 & ~n5107 ) | ( n5102 & n5108 ) | ( ~n5107 & n5108 ) ;
  assign n5110 = n5098 | n5109 ;
  assign n5111 = n5095 | n5110 ;
  assign n5112 = n5095 | n5098 ;
  assign n5113 = n5109 & n5112 ;
  assign n5114 = n5111 & ~n5113 ;
  assign n5115 = ~x355 & x356 ;
  assign n5116 = x355 & ~x356 ;
  assign n5117 = n5115 | n5116 ;
  assign n5118 = ~x357 & n5117 ;
  assign n5119 = x357 & ~n5117 ;
  assign n5120 = n5118 | n5119 ;
  assign n5121 = ~x358 & x359 ;
  assign n5122 = x358 & ~x359 ;
  assign n5123 = n5121 | n5122 ;
  assign n5124 = ~x360 & n5123 ;
  assign n5125 = x360 & ~n5123 ;
  assign n5126 = n5124 | n5125 ;
  assign n5127 = n5120 & n5126 ;
  assign n5128 = ( x358 & x359 ) | ( x358 & x360 ) | ( x359 & x360 ) ;
  assign n5129 = ( x355 & x356 ) | ( x355 & x357 ) | ( x356 & x357 ) ;
  assign n5130 = ~n5128 & n5129 ;
  assign n5131 = n5128 & ~n5129 ;
  assign n5132 = n5130 | n5131 ;
  assign n5133 = ~n5127 & n5132 ;
  assign n5134 = n5127 & ~n5132 ;
  assign n5135 = n5133 | n5134 ;
  assign n5136 = n5120 & ~n5126 ;
  assign n5137 = ~n5120 & n5126 ;
  assign n5138 = n5136 | n5137 ;
  assign n5139 = ( n5127 & n5128 ) | ( n5127 & n5129 ) | ( n5128 & n5129 ) ;
  assign n5140 = n5138 & n5139 ;
  assign n5141 = n5135 & ~n5140 ;
  assign n5142 = n5135 & n5139 ;
  assign n5143 = x361 & ~x362 ;
  assign n5144 = ~x361 & x362 ;
  assign n5145 = n5143 | n5144 ;
  assign n5146 = ~x363 & n5145 ;
  assign n5147 = x363 & ~n5145 ;
  assign n5148 = n5146 | n5147 ;
  assign n5149 = x364 & ~x365 ;
  assign n5150 = ~x364 & x365 ;
  assign n5151 = n5149 | n5150 ;
  assign n5152 = ~x366 & n5151 ;
  assign n5153 = x366 & ~n5151 ;
  assign n5154 = n5152 | n5153 ;
  assign n5155 = n5148 & ~n5154 ;
  assign n5156 = ~n5148 & n5154 ;
  assign n5157 = n5155 | n5156 ;
  assign n5158 = ( x364 & x365 ) | ( x364 & x366 ) | ( x365 & x366 ) ;
  assign n5159 = ( x361 & x362 ) | ( x361 & x363 ) | ( x362 & x363 ) ;
  assign n5160 = n5148 & n5154 ;
  assign n5161 = ( n5158 & n5159 ) | ( n5158 & n5160 ) | ( n5159 & n5160 ) ;
  assign n5162 = n5157 & n5161 ;
  assign n5163 = n5142 | n5162 ;
  assign n5164 = n5158 & ~n5159 ;
  assign n5165 = ~n5158 & n5159 ;
  assign n5166 = n5164 | n5165 ;
  assign n5167 = ~n5160 & n5166 ;
  assign n5168 = n5160 & ~n5166 ;
  assign n5169 = n5167 | n5168 ;
  assign n5170 = n5161 & n5169 ;
  assign n5171 = n5138 & n5157 ;
  assign n5172 = n5169 & n5171 ;
  assign n5173 = ~n5170 & n5172 ;
  assign n5174 = ~n5163 & n5173 ;
  assign n5175 = n5141 & n5174 ;
  assign n5176 = ~n5170 & n5171 ;
  assign n5177 = ~n5162 & n5169 ;
  assign n5178 = n5142 & ~n5177 ;
  assign n5179 = ( n5176 & n5177 ) | ( n5176 & ~n5178 ) | ( n5177 & ~n5178 ) ;
  assign n5180 = ( n5141 & n5175 ) | ( n5141 & ~n5179 ) | ( n5175 & ~n5179 ) ;
  assign n5181 = n5157 & ~n5161 ;
  assign n5182 = ( n5157 & ~n5169 ) | ( n5157 & n5181 ) | ( ~n5169 & n5181 ) ;
  assign n5183 = n5138 & ~n5139 ;
  assign n5184 = ( ~n5135 & n5138 ) | ( ~n5135 & n5183 ) | ( n5138 & n5183 ) ;
  assign n5185 = ~n5182 & n5184 ;
  assign n5186 = n5182 & ~n5184 ;
  assign n5187 = n5185 | n5186 ;
  assign n5188 = ( x352 & x353 ) | ( x352 & x354 ) | ( x353 & x354 ) ;
  assign n5189 = ( x349 & x350 ) | ( x349 & x351 ) | ( x350 & x351 ) ;
  assign n5190 = n5188 & ~n5189 ;
  assign n5191 = ~n5188 & n5189 ;
  assign n5192 = n5190 | n5191 ;
  assign n5193 = x349 & ~x350 ;
  assign n5194 = ~x349 & x350 ;
  assign n5195 = n5193 | n5194 ;
  assign n5196 = ~x351 & n5195 ;
  assign n5197 = x351 & ~n5195 ;
  assign n5198 = n5196 | n5197 ;
  assign n5199 = x352 & ~x353 ;
  assign n5200 = ~x352 & x353 ;
  assign n5201 = n5199 | n5200 ;
  assign n5202 = ~x354 & n5201 ;
  assign n5203 = x354 & ~n5201 ;
  assign n5204 = n5202 | n5203 ;
  assign n5205 = n5198 & n5204 ;
  assign n5206 = n5192 & ~n5205 ;
  assign n5207 = ~n5192 & n5205 ;
  assign n5208 = n5206 | n5207 ;
  assign n5209 = n5198 & ~n5204 ;
  assign n5210 = ~n5198 & n5204 ;
  assign n5211 = n5209 | n5210 ;
  assign n5212 = ( n5188 & n5189 ) | ( n5188 & n5205 ) | ( n5189 & n5205 ) ;
  assign n5213 = n5211 & ~n5212 ;
  assign n5214 = ( ~n5208 & n5211 ) | ( ~n5208 & n5213 ) | ( n5211 & n5213 ) ;
  assign n5215 = ~x343 & x344 ;
  assign n5216 = x343 & ~x344 ;
  assign n5217 = n5215 | n5216 ;
  assign n5218 = ~x345 & n5217 ;
  assign n5219 = x345 & ~n5217 ;
  assign n5220 = n5218 | n5219 ;
  assign n5221 = ~x346 & x347 ;
  assign n5222 = x346 & ~x347 ;
  assign n5223 = n5221 | n5222 ;
  assign n5224 = ~x348 & n5223 ;
  assign n5225 = x348 & ~n5223 ;
  assign n5226 = n5224 | n5225 ;
  assign n5227 = n5220 & n5226 ;
  assign n5228 = ( x346 & x347 ) | ( x346 & x348 ) | ( x347 & x348 ) ;
  assign n5229 = ( x343 & x344 ) | ( x343 & x345 ) | ( x344 & x345 ) ;
  assign n5230 = ~n5228 & n5229 ;
  assign n5231 = n5228 & ~n5229 ;
  assign n5232 = n5230 | n5231 ;
  assign n5233 = ~n5227 & n5232 ;
  assign n5234 = n5227 & ~n5232 ;
  assign n5235 = n5233 | n5234 ;
  assign n5236 = n5220 & ~n5226 ;
  assign n5237 = ~n5220 & n5226 ;
  assign n5238 = n5236 | n5237 ;
  assign n5239 = ( n5227 & n5228 ) | ( n5227 & n5229 ) | ( n5228 & n5229 ) ;
  assign n5240 = n5238 & ~n5239 ;
  assign n5241 = ( ~n5235 & n5238 ) | ( ~n5235 & n5240 ) | ( n5238 & n5240 ) ;
  assign n5242 = ~n5214 & n5241 ;
  assign n5243 = n5214 & ~n5241 ;
  assign n5244 = n5242 | n5243 ;
  assign n5245 = n5187 & n5244 ;
  assign n5246 = ( n5141 & ~n5142 ) | ( n5141 & n5177 ) | ( ~n5142 & n5177 ) ;
  assign n5247 = n5141 & n5177 ;
  assign n5248 = ( n5176 & n5246 ) | ( n5176 & n5247 ) | ( n5246 & n5247 ) ;
  assign n5249 = n5179 & ~n5248 ;
  assign n5250 = n5245 | n5249 ;
  assign n5251 = n5180 | n5250 ;
  assign n5252 = n5235 & n5239 ;
  assign n5253 = n5211 & n5212 ;
  assign n5254 = n5252 | n5253 ;
  assign n5255 = n5208 & n5212 ;
  assign n5256 = n5211 & n5238 ;
  assign n5257 = n5208 & n5256 ;
  assign n5258 = ~n5255 & n5257 ;
  assign n5259 = ~n5254 & n5258 ;
  assign n5260 = n5238 & n5239 ;
  assign n5261 = n5235 & ~n5260 ;
  assign n5262 = ~n5259 & n5261 ;
  assign n5263 = ~n5255 & n5256 ;
  assign n5264 = n5208 & ~n5253 ;
  assign n5265 = ( n5252 & n5261 ) | ( n5252 & n5264 ) | ( n5261 & n5264 ) ;
  assign n5266 = n5261 | n5264 ;
  assign n5267 = ( ~n5263 & n5265 ) | ( ~n5263 & n5266 ) | ( n5265 & n5266 ) ;
  assign n5268 = n5252 | n5264 ;
  assign n5269 = n5263 & ~n5268 ;
  assign n5270 = ( ~n5264 & n5267 ) | ( ~n5264 & n5269 ) | ( n5267 & n5269 ) ;
  assign n5271 = ( ~n5262 & n5267 ) | ( ~n5262 & n5270 ) | ( n5267 & n5270 ) ;
  assign n5272 = n5251 & n5271 ;
  assign n5273 = n5245 & n5249 ;
  assign n5274 = ( n5180 & n5245 ) | ( n5180 & n5273 ) | ( n5245 & n5273 ) ;
  assign n5275 = n5272 | n5274 ;
  assign n5276 = n5252 & ~n5264 ;
  assign n5277 = ( n5263 & n5264 ) | ( n5263 & ~n5276 ) | ( n5264 & ~n5276 ) ;
  assign n5278 = n5261 & n5277 ;
  assign n5279 = ~n5238 & n5239 ;
  assign n5280 = ( ~n5235 & n5239 ) | ( ~n5235 & n5279 ) | ( n5239 & n5279 ) ;
  assign n5281 = ~n5211 & n5212 ;
  assign n5282 = ( ~n5208 & n5212 ) | ( ~n5208 & n5281 ) | ( n5212 & n5281 ) ;
  assign n5283 = ~n5280 & n5282 ;
  assign n5284 = n5280 & ~n5282 ;
  assign n5285 = n5283 | n5284 ;
  assign n5286 = n5259 | n5285 ;
  assign n5287 = n5278 | n5286 ;
  assign n5288 = n5259 & n5285 ;
  assign n5289 = ( n5278 & n5285 ) | ( n5278 & n5288 ) | ( n5285 & n5288 ) ;
  assign n5290 = n5287 & ~n5289 ;
  assign n5291 = n5141 & n5179 ;
  assign n5292 = ~n5138 & n5139 ;
  assign n5293 = ( ~n5135 & n5139 ) | ( ~n5135 & n5292 ) | ( n5139 & n5292 ) ;
  assign n5294 = ~n5157 & n5161 ;
  assign n5295 = ( n5161 & ~n5169 ) | ( n5161 & n5294 ) | ( ~n5169 & n5294 ) ;
  assign n5296 = ~n5293 & n5295 ;
  assign n5297 = n5293 & ~n5295 ;
  assign n5298 = n5296 | n5297 ;
  assign n5299 = n5174 | n5298 ;
  assign n5300 = n5291 | n5299 ;
  assign n5301 = n5174 & n5298 ;
  assign n5302 = ( n5291 & n5298 ) | ( n5291 & n5301 ) | ( n5298 & n5301 ) ;
  assign n5303 = n5300 & ~n5302 ;
  assign n5304 = n5290 | n5303 ;
  assign n5305 = n5275 & n5304 ;
  assign n5306 = n5287 & n5300 ;
  assign n5307 = n5289 | n5302 ;
  assign n5308 = n5306 & ~n5307 ;
  assign n5309 = ( n5174 & n5293 ) | ( n5174 & n5295 ) | ( n5293 & n5295 ) ;
  assign n5310 = n5293 | n5295 ;
  assign n5311 = ( n5291 & n5309 ) | ( n5291 & n5310 ) | ( n5309 & n5310 ) ;
  assign n5312 = ( n5259 & n5280 ) | ( n5259 & n5282 ) | ( n5280 & n5282 ) ;
  assign n5313 = n5280 | n5282 ;
  assign n5314 = ( n5278 & n5312 ) | ( n5278 & n5313 ) | ( n5312 & n5313 ) ;
  assign n5315 = ~n5311 & n5314 ;
  assign n5316 = n5311 & ~n5314 ;
  assign n5317 = n5315 | n5316 ;
  assign n5318 = n5308 | n5317 ;
  assign n5319 = n5305 | n5318 ;
  assign n5320 = n5304 | n5308 ;
  assign n5321 = ( n5275 & n5308 ) | ( n5275 & n5320 ) | ( n5308 & n5320 ) ;
  assign n5322 = n5317 & n5321 ;
  assign n5323 = n5319 & ~n5322 ;
  assign n5324 = ~x331 & x332 ;
  assign n5325 = x331 & ~x332 ;
  assign n5326 = n5324 | n5325 ;
  assign n5327 = ~x333 & n5326 ;
  assign n5328 = x333 & ~n5326 ;
  assign n5329 = n5327 | n5328 ;
  assign n5330 = ~x334 & x335 ;
  assign n5331 = x334 & ~x335 ;
  assign n5332 = n5330 | n5331 ;
  assign n5333 = ~x336 & n5332 ;
  assign n5334 = x336 & ~n5332 ;
  assign n5335 = n5333 | n5334 ;
  assign n5336 = n5329 & n5335 ;
  assign n5337 = ( x334 & x335 ) | ( x334 & x336 ) | ( x335 & x336 ) ;
  assign n5338 = ( x331 & x332 ) | ( x331 & x333 ) | ( x332 & x333 ) ;
  assign n5339 = ~n5337 & n5338 ;
  assign n5340 = n5337 & ~n5338 ;
  assign n5341 = n5339 | n5340 ;
  assign n5342 = ~n5336 & n5341 ;
  assign n5343 = n5336 & ~n5341 ;
  assign n5344 = n5342 | n5343 ;
  assign n5345 = n5329 & ~n5335 ;
  assign n5346 = ~n5329 & n5335 ;
  assign n5347 = n5345 | n5346 ;
  assign n5348 = ( n5336 & n5337 ) | ( n5336 & n5338 ) | ( n5337 & n5338 ) ;
  assign n5349 = n5347 & n5348 ;
  assign n5350 = n5344 & ~n5349 ;
  assign n5351 = n5344 & n5348 ;
  assign n5352 = x337 & ~x338 ;
  assign n5353 = ~x337 & x338 ;
  assign n5354 = n5352 | n5353 ;
  assign n5355 = ~x339 & n5354 ;
  assign n5356 = x339 & ~n5354 ;
  assign n5357 = n5355 | n5356 ;
  assign n5358 = x340 & ~x341 ;
  assign n5359 = ~x340 & x341 ;
  assign n5360 = n5358 | n5359 ;
  assign n5361 = ~x342 & n5360 ;
  assign n5362 = x342 & ~n5360 ;
  assign n5363 = n5361 | n5362 ;
  assign n5364 = n5357 & ~n5363 ;
  assign n5365 = ~n5357 & n5363 ;
  assign n5366 = n5364 | n5365 ;
  assign n5367 = ( x340 & x341 ) | ( x340 & x342 ) | ( x341 & x342 ) ;
  assign n5368 = ( x337 & x338 ) | ( x337 & x339 ) | ( x338 & x339 ) ;
  assign n5369 = n5357 & n5363 ;
  assign n5370 = ( n5367 & n5368 ) | ( n5367 & n5369 ) | ( n5368 & n5369 ) ;
  assign n5371 = n5366 & n5370 ;
  assign n5372 = n5351 | n5371 ;
  assign n5373 = n5367 & ~n5368 ;
  assign n5374 = ~n5367 & n5368 ;
  assign n5375 = n5373 | n5374 ;
  assign n5376 = ~n5369 & n5375 ;
  assign n5377 = n5369 & ~n5375 ;
  assign n5378 = n5376 | n5377 ;
  assign n5379 = n5370 & n5378 ;
  assign n5380 = n5347 & n5366 ;
  assign n5381 = n5378 & n5380 ;
  assign n5382 = ~n5379 & n5381 ;
  assign n5383 = ~n5372 & n5382 ;
  assign n5384 = n5350 & n5383 ;
  assign n5385 = ~n5379 & n5380 ;
  assign n5386 = ~n5371 & n5378 ;
  assign n5387 = n5351 & ~n5386 ;
  assign n5388 = ( n5385 & n5386 ) | ( n5385 & ~n5387 ) | ( n5386 & ~n5387 ) ;
  assign n5389 = ( n5350 & n5384 ) | ( n5350 & ~n5388 ) | ( n5384 & ~n5388 ) ;
  assign n5390 = n5366 & ~n5370 ;
  assign n5391 = ( n5366 & ~n5378 ) | ( n5366 & n5390 ) | ( ~n5378 & n5390 ) ;
  assign n5392 = n5347 & ~n5348 ;
  assign n5393 = ( ~n5344 & n5347 ) | ( ~n5344 & n5392 ) | ( n5347 & n5392 ) ;
  assign n5394 = ~n5391 & n5393 ;
  assign n5395 = n5391 & ~n5393 ;
  assign n5396 = n5394 | n5395 ;
  assign n5397 = ( x328 & x329 ) | ( x328 & x330 ) | ( x329 & x330 ) ;
  assign n5398 = ( x325 & x326 ) | ( x325 & x327 ) | ( x326 & x327 ) ;
  assign n5399 = n5397 & ~n5398 ;
  assign n5400 = ~n5397 & n5398 ;
  assign n5401 = n5399 | n5400 ;
  assign n5402 = ~x325 & x326 ;
  assign n5403 = x325 & ~x326 ;
  assign n5404 = n5402 | n5403 ;
  assign n5405 = ~x327 & n5404 ;
  assign n5406 = x327 & ~n5404 ;
  assign n5407 = n5405 | n5406 ;
  assign n5408 = ~x328 & x329 ;
  assign n5409 = x328 & ~x329 ;
  assign n5410 = n5408 | n5409 ;
  assign n5411 = ~x330 & n5410 ;
  assign n5412 = x330 & ~n5410 ;
  assign n5413 = n5411 | n5412 ;
  assign n5414 = n5407 & n5413 ;
  assign n5415 = n5401 & ~n5414 ;
  assign n5416 = ~n5401 & n5414 ;
  assign n5417 = n5415 | n5416 ;
  assign n5418 = n5407 & ~n5413 ;
  assign n5419 = ~n5407 & n5413 ;
  assign n5420 = n5418 | n5419 ;
  assign n5421 = ( n5397 & n5398 ) | ( n5397 & n5414 ) | ( n5398 & n5414 ) ;
  assign n5422 = n5420 & ~n5421 ;
  assign n5423 = ( ~n5417 & n5420 ) | ( ~n5417 & n5422 ) | ( n5420 & n5422 ) ;
  assign n5424 = ~x319 & x320 ;
  assign n5425 = x319 & ~x320 ;
  assign n5426 = n5424 | n5425 ;
  assign n5427 = ~x321 & n5426 ;
  assign n5428 = x321 & ~n5426 ;
  assign n5429 = n5427 | n5428 ;
  assign n5430 = ~x322 & x323 ;
  assign n5431 = x322 & ~x323 ;
  assign n5432 = n5430 | n5431 ;
  assign n5433 = ~x324 & n5432 ;
  assign n5434 = x324 & ~n5432 ;
  assign n5435 = n5433 | n5434 ;
  assign n5436 = n5429 & ~n5435 ;
  assign n5437 = ~n5429 & n5435 ;
  assign n5438 = n5436 | n5437 ;
  assign n5439 = ( x322 & x323 ) | ( x322 & x324 ) | ( x323 & x324 ) ;
  assign n5440 = ( x319 & x320 ) | ( x319 & x321 ) | ( x320 & x321 ) ;
  assign n5441 = n5439 & ~n5440 ;
  assign n5442 = ~n5439 & n5440 ;
  assign n5443 = n5441 | n5442 ;
  assign n5444 = n5429 & n5435 ;
  assign n5445 = n5443 & ~n5444 ;
  assign n5446 = ~n5443 & n5444 ;
  assign n5447 = n5445 | n5446 ;
  assign n5448 = ( n5439 & n5440 ) | ( n5439 & n5444 ) | ( n5440 & n5444 ) ;
  assign n5449 = n5438 & ~n5448 ;
  assign n5450 = ( n5438 & ~n5447 ) | ( n5438 & n5449 ) | ( ~n5447 & n5449 ) ;
  assign n5451 = ~n5423 & n5450 ;
  assign n5452 = n5423 & ~n5450 ;
  assign n5453 = n5451 | n5452 ;
  assign n5454 = n5396 & n5453 ;
  assign n5455 = ( n5350 & ~n5351 ) | ( n5350 & n5386 ) | ( ~n5351 & n5386 ) ;
  assign n5456 = n5350 & n5386 ;
  assign n5457 = ( n5385 & n5455 ) | ( n5385 & n5456 ) | ( n5455 & n5456 ) ;
  assign n5458 = n5388 & ~n5457 ;
  assign n5459 = n5454 | n5458 ;
  assign n5460 = n5389 | n5459 ;
  assign n5461 = n5447 & n5448 ;
  assign n5462 = n5420 & n5421 ;
  assign n5463 = n5461 | n5462 ;
  assign n5464 = n5417 & n5421 ;
  assign n5465 = n5420 & n5438 ;
  assign n5466 = n5417 & n5465 ;
  assign n5467 = ~n5464 & n5466 ;
  assign n5468 = ~n5463 & n5467 ;
  assign n5469 = n5438 & n5448 ;
  assign n5470 = n5447 & ~n5469 ;
  assign n5471 = ~n5468 & n5470 ;
  assign n5472 = ~n5464 & n5465 ;
  assign n5473 = n5417 & ~n5462 ;
  assign n5474 = ( n5461 & n5470 ) | ( n5461 & n5473 ) | ( n5470 & n5473 ) ;
  assign n5475 = n5470 | n5473 ;
  assign n5476 = ( ~n5472 & n5474 ) | ( ~n5472 & n5475 ) | ( n5474 & n5475 ) ;
  assign n5477 = n5461 | n5473 ;
  assign n5478 = n5472 & ~n5477 ;
  assign n5479 = ( ~n5473 & n5476 ) | ( ~n5473 & n5478 ) | ( n5476 & n5478 ) ;
  assign n5480 = ( ~n5471 & n5476 ) | ( ~n5471 & n5479 ) | ( n5476 & n5479 ) ;
  assign n5481 = n5460 & n5480 ;
  assign n5482 = n5454 & n5458 ;
  assign n5483 = ( n5389 & n5454 ) | ( n5389 & n5482 ) | ( n5454 & n5482 ) ;
  assign n5484 = n5481 | n5483 ;
  assign n5485 = n5461 & ~n5473 ;
  assign n5486 = ( n5472 & n5473 ) | ( n5472 & ~n5485 ) | ( n5473 & ~n5485 ) ;
  assign n5487 = n5470 & n5486 ;
  assign n5488 = ~n5438 & n5448 ;
  assign n5489 = ( ~n5447 & n5448 ) | ( ~n5447 & n5488 ) | ( n5448 & n5488 ) ;
  assign n5490 = ~n5420 & n5421 ;
  assign n5491 = ( ~n5417 & n5421 ) | ( ~n5417 & n5490 ) | ( n5421 & n5490 ) ;
  assign n5492 = ~n5489 & n5491 ;
  assign n5493 = n5489 & ~n5491 ;
  assign n5494 = n5492 | n5493 ;
  assign n5495 = n5468 | n5494 ;
  assign n5496 = n5487 | n5495 ;
  assign n5497 = n5468 & n5494 ;
  assign n5498 = ( n5487 & n5494 ) | ( n5487 & n5497 ) | ( n5494 & n5497 ) ;
  assign n5499 = n5496 & ~n5498 ;
  assign n5500 = n5350 & n5388 ;
  assign n5501 = ~n5347 & n5348 ;
  assign n5502 = ( ~n5344 & n5348 ) | ( ~n5344 & n5501 ) | ( n5348 & n5501 ) ;
  assign n5503 = ~n5366 & n5370 ;
  assign n5504 = ( n5370 & ~n5378 ) | ( n5370 & n5503 ) | ( ~n5378 & n5503 ) ;
  assign n5505 = ~n5502 & n5504 ;
  assign n5506 = n5502 & ~n5504 ;
  assign n5507 = n5505 | n5506 ;
  assign n5508 = n5383 | n5507 ;
  assign n5509 = n5500 | n5508 ;
  assign n5510 = n5383 & n5507 ;
  assign n5511 = ( n5500 & n5507 ) | ( n5500 & n5510 ) | ( n5507 & n5510 ) ;
  assign n5512 = n5509 & ~n5511 ;
  assign n5513 = n5499 | n5512 ;
  assign n5514 = n5484 & n5513 ;
  assign n5515 = n5496 & n5509 ;
  assign n5516 = n5498 | n5511 ;
  assign n5517 = n5515 & ~n5516 ;
  assign n5518 = ( n5383 & n5502 ) | ( n5383 & n5504 ) | ( n5502 & n5504 ) ;
  assign n5519 = n5502 | n5504 ;
  assign n5520 = ( n5500 & n5518 ) | ( n5500 & n5519 ) | ( n5518 & n5519 ) ;
  assign n5521 = ( n5468 & n5489 ) | ( n5468 & n5491 ) | ( n5489 & n5491 ) ;
  assign n5522 = n5489 | n5491 ;
  assign n5523 = ( n5487 & n5521 ) | ( n5487 & n5522 ) | ( n5521 & n5522 ) ;
  assign n5524 = ~n5520 & n5523 ;
  assign n5525 = n5520 & ~n5523 ;
  assign n5526 = n5524 | n5525 ;
  assign n5527 = n5517 | n5526 ;
  assign n5528 = n5514 | n5527 ;
  assign n5529 = n5513 | n5517 ;
  assign n5530 = ( n5484 & n5517 ) | ( n5484 & n5529 ) | ( n5517 & n5529 ) ;
  assign n5531 = n5526 & n5530 ;
  assign n5532 = n5528 & ~n5531 ;
  assign n5533 = n5323 | n5532 ;
  assign n5534 = n5251 & ~n5274 ;
  assign n5535 = n5271 & ~n5534 ;
  assign n5536 = n5187 & ~n5244 ;
  assign n5537 = ~n5187 & n5244 ;
  assign n5538 = n5536 | n5537 ;
  assign n5539 = n5396 & ~n5453 ;
  assign n5540 = ~n5396 & n5453 ;
  assign n5541 = n5539 | n5540 ;
  assign n5542 = n5538 & n5541 ;
  assign n5543 = ~n5245 & n5251 ;
  assign n5544 = n5251 & ~n5271 ;
  assign n5545 = n5180 | n5249 ;
  assign n5546 = n5271 | n5545 ;
  assign n5547 = ( n5543 & n5544 ) | ( n5543 & ~n5546 ) | ( n5544 & ~n5546 ) ;
  assign n5548 = n5542 | n5547 ;
  assign n5549 = n5535 | n5548 ;
  assign n5550 = n5389 | n5458 ;
  assign n5551 = ( n5454 & n5480 ) | ( n5454 & ~n5550 ) | ( n5480 & ~n5550 ) ;
  assign n5552 = ( ~n5480 & n5550 ) | ( ~n5480 & n5551 ) | ( n5550 & n5551 ) ;
  assign n5553 = ( ~n5454 & n5551 ) | ( ~n5454 & n5552 ) | ( n5551 & n5552 ) ;
  assign n5554 = n5549 & n5553 ;
  assign n5555 = n5535 | n5547 ;
  assign n5556 = n5542 & n5555 ;
  assign n5557 = ( n5483 & ~n5499 ) | ( n5483 & n5512 ) | ( ~n5499 & n5512 ) ;
  assign n5558 = n5499 & ~n5512 ;
  assign n5559 = ( n5481 & n5557 ) | ( n5481 & ~n5558 ) | ( n5557 & ~n5558 ) ;
  assign n5560 = ( ~n5484 & n5499 ) | ( ~n5484 & n5559 ) | ( n5499 & n5559 ) ;
  assign n5561 = ( ~n5512 & n5559 ) | ( ~n5512 & n5560 ) | ( n5559 & n5560 ) ;
  assign n5562 = ( n5274 & ~n5290 ) | ( n5274 & n5303 ) | ( ~n5290 & n5303 ) ;
  assign n5563 = n5290 & ~n5303 ;
  assign n5564 = ( n5272 & n5562 ) | ( n5272 & ~n5563 ) | ( n5562 & ~n5563 ) ;
  assign n5565 = ( ~n5275 & n5290 ) | ( ~n5275 & n5564 ) | ( n5290 & n5564 ) ;
  assign n5566 = ( ~n5303 & n5564 ) | ( ~n5303 & n5565 ) | ( n5564 & n5565 ) ;
  assign n5567 = ( n5556 & n5561 ) | ( n5556 & n5566 ) | ( n5561 & n5566 ) ;
  assign n5568 = n5561 | n5566 ;
  assign n5569 = ( n5554 & n5567 ) | ( n5554 & n5568 ) | ( n5567 & n5568 ) ;
  assign n5570 = n5533 & n5569 ;
  assign n5571 = n5319 & n5528 ;
  assign n5572 = n5322 | n5531 ;
  assign n5573 = n5571 & ~n5572 ;
  assign n5574 = n5520 & n5523 ;
  assign n5575 = n5520 | n5523 ;
  assign n5576 = n5574 | n5575 ;
  assign n5577 = ( n5530 & n5574 ) | ( n5530 & n5576 ) | ( n5574 & n5576 ) ;
  assign n5578 = n5311 & n5314 ;
  assign n5579 = n5311 | n5314 ;
  assign n5580 = n5578 | n5579 ;
  assign n5581 = ( n5321 & n5578 ) | ( n5321 & n5580 ) | ( n5578 & n5580 ) ;
  assign n5582 = n5577 & n5581 ;
  assign n5583 = n5581 & ~n5582 ;
  assign n5584 = ( n5577 & ~n5582 ) | ( n5577 & n5583 ) | ( ~n5582 & n5583 ) ;
  assign n5585 = n5573 | n5584 ;
  assign n5586 = n5570 | n5585 ;
  assign n5587 = n5570 | n5573 ;
  assign n5588 = n5584 & n5587 ;
  assign n5589 = n5586 & ~n5588 ;
  assign n5590 = n5114 | n5589 ;
  assign n5591 = n5538 & ~n5541 ;
  assign n5592 = ~n5538 & n5541 ;
  assign n5593 = n5591 | n5592 ;
  assign n5594 = n5063 & ~n5066 ;
  assign n5595 = ~n5063 & n5066 ;
  assign n5596 = n5594 | n5595 ;
  assign n5597 = n5593 & n5596 ;
  assign n5598 = ~n5549 & n5553 ;
  assign n5599 = ( n5553 & n5556 ) | ( n5553 & n5598 ) | ( n5556 & n5598 ) ;
  assign n5600 = ~n5542 & n5555 ;
  assign n5601 = n5542 & ~n5547 ;
  assign n5602 = ~n5535 & n5601 ;
  assign n5603 = ~n5553 & n5602 ;
  assign n5604 = ( ~n5553 & n5600 ) | ( ~n5553 & n5603 ) | ( n5600 & n5603 ) ;
  assign n5605 = n5599 | n5604 ;
  assign n5606 = n5597 & n5605 ;
  assign n5607 = n5597 | n5600 ;
  assign n5608 = n5553 & ~n5597 ;
  assign n5609 = ( n5603 & n5607 ) | ( n5603 & ~n5608 ) | ( n5607 & ~n5608 ) ;
  assign n5610 = n5599 | n5609 ;
  assign n5611 = ~n5067 & n5080 ;
  assign n5612 = n5067 & ~n5072 ;
  assign n5613 = ~n5060 & n5612 ;
  assign n5614 = ~n5078 & n5613 ;
  assign n5615 = ( ~n5078 & n5611 ) | ( ~n5078 & n5614 ) | ( n5611 & n5614 ) ;
  assign n5616 = n5079 & ~n5081 ;
  assign n5617 = ( n5078 & n5615 ) | ( n5078 & ~n5616 ) | ( n5615 & ~n5616 ) ;
  assign n5618 = n5610 & n5617 ;
  assign n5619 = n5606 | n5618 ;
  assign n5621 = ( n5081 & ~n5086 ) | ( n5081 & n5091 ) | ( ~n5086 & n5091 ) ;
  assign n5622 = n5086 & ~n5091 ;
  assign n5623 = ( n5079 & n5621 ) | ( n5079 & ~n5622 ) | ( n5621 & ~n5622 ) ;
  assign n5620 = n5079 | n5081 ;
  assign n5624 = ( n5086 & ~n5620 ) | ( n5086 & n5623 ) | ( ~n5620 & n5623 ) ;
  assign n5625 = ( ~n5091 & n5623 ) | ( ~n5091 & n5624 ) | ( n5623 & n5624 ) ;
  assign n5627 = ( n5556 & ~n5561 ) | ( n5556 & n5566 ) | ( ~n5561 & n5566 ) ;
  assign n5628 = n5561 & ~n5566 ;
  assign n5629 = ( n5554 & n5627 ) | ( n5554 & ~n5628 ) | ( n5627 & ~n5628 ) ;
  assign n5626 = n5554 | n5556 ;
  assign n5630 = ( n5561 & ~n5626 ) | ( n5561 & n5629 ) | ( ~n5626 & n5629 ) ;
  assign n5631 = ( ~n5566 & n5629 ) | ( ~n5566 & n5630 ) | ( n5629 & n5630 ) ;
  assign n5632 = ( n5619 & n5625 ) | ( n5619 & n5631 ) | ( n5625 & n5631 ) ;
  assign n5633 = ( ~n5323 & n5532 ) | ( ~n5323 & n5569 ) | ( n5532 & n5569 ) ;
  assign n5634 = ( n5323 & ~n5569 ) | ( n5323 & n5633 ) | ( ~n5569 & n5633 ) ;
  assign n5635 = ( ~n5532 & n5633 ) | ( ~n5532 & n5634 ) | ( n5633 & n5634 ) ;
  assign n5636 = ( ~n4848 & n5057 ) | ( ~n4848 & n5094 ) | ( n5057 & n5094 ) ;
  assign n5637 = ( n4848 & ~n5094 ) | ( n4848 & n5636 ) | ( ~n5094 & n5636 ) ;
  assign n5638 = ( ~n5057 & n5636 ) | ( ~n5057 & n5637 ) | ( n5636 & n5637 ) ;
  assign n5639 = ( n5632 & n5635 ) | ( n5632 & n5638 ) | ( n5635 & n5638 ) ;
  assign n5640 = n5590 & n5639 ;
  assign n5641 = n5111 & n5586 ;
  assign n5642 = n5113 | n5588 ;
  assign n5643 = n5641 & ~n5642 ;
  assign n5652 = n4846 & n5104 ;
  assign n5653 = n5048 | n5103 ;
  assign n5654 = n5045 | n5103 ;
  assign n5655 = ( n5055 & n5653 ) | ( n5055 & n5654 ) | ( n5653 & n5654 ) ;
  assign n5656 = n5652 | n5655 ;
  assign n5657 = n5107 | n5656 ;
  assign n5658 = ( n5098 & n5107 ) | ( n5098 & n5657 ) | ( n5107 & n5657 ) ;
  assign n5659 = n5107 | n5657 ;
  assign n5660 = ( n5095 & n5658 ) | ( n5095 & n5659 ) | ( n5658 & n5659 ) ;
  assign n5644 = n5321 & n5579 ;
  assign n5645 = n5523 | n5578 ;
  assign n5646 = n5520 | n5578 ;
  assign n5647 = ( n5530 & n5645 ) | ( n5530 & n5646 ) | ( n5645 & n5646 ) ;
  assign n5648 = n5644 | n5647 ;
  assign n5649 = n5573 & n5648 ;
  assign n5650 = ( n5570 & n5648 ) | ( n5570 & n5649 ) | ( n5648 & n5649 ) ;
  assign n5651 = n5582 | n5650 ;
  assign n5661 = n5651 & n5660 ;
  assign n5662 = n5651 & ~n5661 ;
  assign n5663 = ( n5660 & ~n5661 ) | ( n5660 & n5662 ) | ( ~n5661 & n5662 ) ;
  assign n5664 = n5643 | n5663 ;
  assign n5665 = n5640 | n5664 ;
  assign n5666 = n5640 | n5643 ;
  assign n5667 = n5663 & n5666 ;
  assign n5668 = n5665 & ~n5667 ;
  assign n5669 = n4639 | n5668 ;
  assign n5670 = ( ~n5114 & n5589 ) | ( ~n5114 & n5639 ) | ( n5589 & n5639 ) ;
  assign n5671 = ( n5114 & ~n5639 ) | ( n5114 & n5670 ) | ( ~n5639 & n5670 ) ;
  assign n5672 = ( ~n5589 & n5670 ) | ( ~n5589 & n5671 ) | ( n5670 & n5671 ) ;
  assign n5673 = ( ~n4087 & n4562 ) | ( ~n4087 & n4610 ) | ( n4562 & n4610 ) ;
  assign n5674 = ( n4087 & ~n4610 ) | ( n4087 & n5673 ) | ( ~n4610 & n5673 ) ;
  assign n5675 = ( ~n4562 & n5673 ) | ( ~n4562 & n5674 ) | ( n5673 & n5674 ) ;
  assign n5676 = n4579 & ~n4582 ;
  assign n5677 = ~n4579 & n4582 ;
  assign n5678 = n5676 | n5677 ;
  assign n5679 = n5593 & ~n5596 ;
  assign n5680 = ~n5593 & n5596 ;
  assign n5681 = n5679 | n5680 ;
  assign n5682 = n5678 & n5681 ;
  assign n5683 = n4592 & ~n4594 ;
  assign n5684 = n4576 & ~n5683 ;
  assign n5685 = ~n4583 & n4591 ;
  assign n5686 = n4583 & ~n4591 ;
  assign n5687 = n5685 | n5686 ;
  assign n5688 = ~n4576 & n5687 ;
  assign n5689 = n5684 | n5688 ;
  assign n5690 = n5682 & n5689 ;
  assign n5691 = n4576 & ~n5682 ;
  assign n5692 = ( n5682 & n5687 ) | ( n5682 & ~n5691 ) | ( n5687 & ~n5691 ) ;
  assign n5693 = n5684 | n5692 ;
  assign n5694 = ( n5597 & ~n5605 ) | ( n5597 & n5617 ) | ( ~n5605 & n5617 ) ;
  assign n5695 = ( ~n5597 & n5605 ) | ( ~n5597 & n5694 ) | ( n5605 & n5694 ) ;
  assign n5696 = ( ~n5617 & n5694 ) | ( ~n5617 & n5695 ) | ( n5694 & n5695 ) ;
  assign n5697 = n5693 & n5696 ;
  assign n5698 = n5690 | n5697 ;
  assign n5699 = ( n5619 & ~n5625 ) | ( n5619 & n5631 ) | ( ~n5625 & n5631 ) ;
  assign n5700 = ( ~n5619 & n5625 ) | ( ~n5619 & n5699 ) | ( n5625 & n5699 ) ;
  assign n5701 = ( ~n5631 & n5699 ) | ( ~n5631 & n5700 ) | ( n5699 & n5700 ) ;
  assign n5703 = ( n4594 & ~n4600 ) | ( n4594 & n4606 ) | ( ~n4600 & n4606 ) ;
  assign n5704 = n4600 & ~n4606 ;
  assign n5705 = ( n4593 & n5703 ) | ( n4593 & ~n5704 ) | ( n5703 & ~n5704 ) ;
  assign n5702 = n4593 | n4594 ;
  assign n5706 = ( n4600 & ~n5702 ) | ( n4600 & n5705 ) | ( ~n5702 & n5705 ) ;
  assign n5707 = ( ~n4606 & n5705 ) | ( ~n4606 & n5706 ) | ( n5705 & n5706 ) ;
  assign n5708 = ( n5698 & n5701 ) | ( n5698 & n5707 ) | ( n5701 & n5707 ) ;
  assign n5709 = ( ~n4566 & n4569 ) | ( ~n4566 & n4609 ) | ( n4569 & n4609 ) ;
  assign n5710 = ( n4566 & ~n4609 ) | ( n4566 & n5709 ) | ( ~n4609 & n5709 ) ;
  assign n5711 = ( ~n4569 & n5709 ) | ( ~n4569 & n5710 ) | ( n5709 & n5710 ) ;
  assign n5712 = ( n5632 & ~n5635 ) | ( n5632 & n5638 ) | ( ~n5635 & n5638 ) ;
  assign n5713 = ( ~n5632 & n5635 ) | ( ~n5632 & n5712 ) | ( n5635 & n5712 ) ;
  assign n5714 = ( ~n5638 & n5712 ) | ( ~n5638 & n5713 ) | ( n5712 & n5713 ) ;
  assign n5715 = ( n5708 & n5711 ) | ( n5708 & n5714 ) | ( n5711 & n5714 ) ;
  assign n5716 = ( n5672 & n5675 ) | ( n5672 & n5715 ) | ( n5675 & n5715 ) ;
  assign n5717 = n5669 & n5716 ;
  assign n5718 = n4636 & n5665 ;
  assign n5719 = n4638 | n5667 ;
  assign n5720 = n5718 & ~n5719 ;
  assign n5728 = n5107 | n5582 ;
  assign n5729 = n5656 | n5728 ;
  assign n5730 = ( n5112 & n5728 ) | ( n5112 & n5729 ) | ( n5728 & n5729 ) ;
  assign n5731 = n5650 | n5730 ;
  assign n5732 = n5661 | n5731 ;
  assign n5733 = ( n5643 & n5661 ) | ( n5643 & n5732 ) | ( n5661 & n5732 ) ;
  assign n5734 = n5661 | n5732 ;
  assign n5735 = ( n5640 & n5733 ) | ( n5640 & n5734 ) | ( n5733 & n5734 ) ;
  assign n5721 = n4080 | n4555 ;
  assign n5722 = n4627 | n5721 ;
  assign n5723 = ( n4085 & n5721 ) | ( n4085 & n5722 ) | ( n5721 & n5722 ) ;
  assign n5724 = n4621 | n5723 ;
  assign n5725 = n4614 & n5724 ;
  assign n5726 = ( n4611 & n5724 ) | ( n4611 & n5725 ) | ( n5724 & n5725 ) ;
  assign n5727 = n4632 | n5726 ;
  assign n5736 = n5727 & n5735 ;
  assign n5737 = n5727 & ~n5736 ;
  assign n5738 = ( n5735 & ~n5736 ) | ( n5735 & n5737 ) | ( ~n5736 & n5737 ) ;
  assign n5739 = n5720 | n5738 ;
  assign n5740 = n5717 | n5739 ;
  assign n5741 = n5717 | n5720 ;
  assign n5742 = n5738 & n5741 ;
  assign n5743 = n5740 & ~n5742 ;
  assign n5744 = ~x211 & x212 ;
  assign n5745 = x211 & ~x212 ;
  assign n5746 = n5744 | n5745 ;
  assign n5747 = ~x213 & n5746 ;
  assign n5748 = x213 & ~n5746 ;
  assign n5749 = n5747 | n5748 ;
  assign n5750 = ~x214 & x215 ;
  assign n5751 = x214 & ~x215 ;
  assign n5752 = n5750 | n5751 ;
  assign n5753 = ~x216 & n5752 ;
  assign n5754 = x216 & ~n5752 ;
  assign n5755 = n5753 | n5754 ;
  assign n5756 = n5749 & n5755 ;
  assign n5757 = ( x214 & x215 ) | ( x214 & x216 ) | ( x215 & x216 ) ;
  assign n5758 = ( x211 & x212 ) | ( x211 & x213 ) | ( x212 & x213 ) ;
  assign n5759 = ~n5757 & n5758 ;
  assign n5760 = n5757 & ~n5758 ;
  assign n5761 = n5759 | n5760 ;
  assign n5762 = ~n5756 & n5761 ;
  assign n5763 = n5756 & ~n5761 ;
  assign n5764 = n5762 | n5763 ;
  assign n5765 = n5749 & ~n5755 ;
  assign n5766 = ~n5749 & n5755 ;
  assign n5767 = n5765 | n5766 ;
  assign n5768 = ( n5756 & n5757 ) | ( n5756 & n5758 ) | ( n5757 & n5758 ) ;
  assign n5769 = n5767 & n5768 ;
  assign n5770 = n5764 & ~n5769 ;
  assign n5771 = n5764 & n5768 ;
  assign n5772 = x217 & ~x218 ;
  assign n5773 = ~x217 & x218 ;
  assign n5774 = n5772 | n5773 ;
  assign n5775 = ~x219 & n5774 ;
  assign n5776 = x219 & ~n5774 ;
  assign n5777 = n5775 | n5776 ;
  assign n5778 = x220 & ~x221 ;
  assign n5779 = ~x220 & x221 ;
  assign n5780 = n5778 | n5779 ;
  assign n5781 = ~x222 & n5780 ;
  assign n5782 = x222 & ~n5780 ;
  assign n5783 = n5781 | n5782 ;
  assign n5784 = n5777 & ~n5783 ;
  assign n5785 = ~n5777 & n5783 ;
  assign n5786 = n5784 | n5785 ;
  assign n5787 = ( x220 & x221 ) | ( x220 & x222 ) | ( x221 & x222 ) ;
  assign n5788 = ( x217 & x218 ) | ( x217 & x219 ) | ( x218 & x219 ) ;
  assign n5789 = n5777 & n5783 ;
  assign n5790 = ( n5787 & n5788 ) | ( n5787 & n5789 ) | ( n5788 & n5789 ) ;
  assign n5791 = n5786 & n5790 ;
  assign n5792 = n5771 | n5791 ;
  assign n5793 = n5787 & ~n5788 ;
  assign n5794 = ~n5787 & n5788 ;
  assign n5795 = n5793 | n5794 ;
  assign n5796 = ~n5789 & n5795 ;
  assign n5797 = n5789 & ~n5795 ;
  assign n5798 = n5796 | n5797 ;
  assign n5799 = n5790 & n5798 ;
  assign n5800 = n5767 & n5786 ;
  assign n5801 = n5798 & n5800 ;
  assign n5802 = ~n5799 & n5801 ;
  assign n5803 = ~n5792 & n5802 ;
  assign n5804 = n5770 & n5803 ;
  assign n5805 = ~n5799 & n5800 ;
  assign n5806 = ~n5791 & n5798 ;
  assign n5807 = n5771 & ~n5806 ;
  assign n5808 = ( n5805 & n5806 ) | ( n5805 & ~n5807 ) | ( n5806 & ~n5807 ) ;
  assign n5809 = ( n5770 & n5804 ) | ( n5770 & ~n5808 ) | ( n5804 & ~n5808 ) ;
  assign n5810 = n5786 & ~n5790 ;
  assign n5811 = ( n5786 & ~n5798 ) | ( n5786 & n5810 ) | ( ~n5798 & n5810 ) ;
  assign n5812 = n5767 & ~n5768 ;
  assign n5813 = ( ~n5764 & n5767 ) | ( ~n5764 & n5812 ) | ( n5767 & n5812 ) ;
  assign n5814 = ~n5811 & n5813 ;
  assign n5815 = n5811 & ~n5813 ;
  assign n5816 = n5814 | n5815 ;
  assign n5817 = ( x208 & x209 ) | ( x208 & x210 ) | ( x209 & x210 ) ;
  assign n5818 = ( x205 & x206 ) | ( x205 & x207 ) | ( x206 & x207 ) ;
  assign n5819 = n5817 & ~n5818 ;
  assign n5820 = ~n5817 & n5818 ;
  assign n5821 = n5819 | n5820 ;
  assign n5822 = x205 & ~x206 ;
  assign n5823 = ~x205 & x206 ;
  assign n5824 = n5822 | n5823 ;
  assign n5825 = ~x207 & n5824 ;
  assign n5826 = x207 & ~n5824 ;
  assign n5827 = n5825 | n5826 ;
  assign n5828 = x208 & ~x209 ;
  assign n5829 = ~x208 & x209 ;
  assign n5830 = n5828 | n5829 ;
  assign n5831 = ~x210 & n5830 ;
  assign n5832 = x210 & ~n5830 ;
  assign n5833 = n5831 | n5832 ;
  assign n5834 = n5827 & n5833 ;
  assign n5835 = n5821 & ~n5834 ;
  assign n5836 = ~n5821 & n5834 ;
  assign n5837 = n5835 | n5836 ;
  assign n5838 = n5827 & ~n5833 ;
  assign n5839 = ~n5827 & n5833 ;
  assign n5840 = n5838 | n5839 ;
  assign n5841 = ( n5817 & n5818 ) | ( n5817 & n5834 ) | ( n5818 & n5834 ) ;
  assign n5842 = n5840 & ~n5841 ;
  assign n5843 = ( ~n5837 & n5840 ) | ( ~n5837 & n5842 ) | ( n5840 & n5842 ) ;
  assign n5844 = ~x199 & x200 ;
  assign n5845 = x199 & ~x200 ;
  assign n5846 = n5844 | n5845 ;
  assign n5847 = ~x201 & n5846 ;
  assign n5848 = x201 & ~n5846 ;
  assign n5849 = n5847 | n5848 ;
  assign n5850 = ~x202 & x203 ;
  assign n5851 = x202 & ~x203 ;
  assign n5852 = n5850 | n5851 ;
  assign n5853 = ~x204 & n5852 ;
  assign n5854 = x204 & ~n5852 ;
  assign n5855 = n5853 | n5854 ;
  assign n5856 = n5849 & n5855 ;
  assign n5857 = ( x202 & x203 ) | ( x202 & x204 ) | ( x203 & x204 ) ;
  assign n5858 = ( x199 & x200 ) | ( x199 & x201 ) | ( x200 & x201 ) ;
  assign n5859 = ~n5857 & n5858 ;
  assign n5860 = n5857 & ~n5858 ;
  assign n5861 = n5859 | n5860 ;
  assign n5862 = ~n5856 & n5861 ;
  assign n5863 = n5856 & ~n5861 ;
  assign n5864 = n5862 | n5863 ;
  assign n5865 = n5849 & ~n5855 ;
  assign n5866 = ~n5849 & n5855 ;
  assign n5867 = n5865 | n5866 ;
  assign n5868 = ( n5856 & n5857 ) | ( n5856 & n5858 ) | ( n5857 & n5858 ) ;
  assign n5869 = n5867 & ~n5868 ;
  assign n5870 = ( ~n5864 & n5867 ) | ( ~n5864 & n5869 ) | ( n5867 & n5869 ) ;
  assign n5871 = ~n5843 & n5870 ;
  assign n5872 = n5843 & ~n5870 ;
  assign n5873 = n5871 | n5872 ;
  assign n5874 = n5816 & n5873 ;
  assign n5875 = ( n5770 & ~n5771 ) | ( n5770 & n5806 ) | ( ~n5771 & n5806 ) ;
  assign n5876 = n5770 & n5806 ;
  assign n5877 = ( n5805 & n5875 ) | ( n5805 & n5876 ) | ( n5875 & n5876 ) ;
  assign n5878 = n5808 & ~n5877 ;
  assign n5879 = n5874 | n5878 ;
  assign n5880 = n5809 | n5879 ;
  assign n5881 = n5864 & n5868 ;
  assign n5882 = n5840 & n5841 ;
  assign n5883 = n5881 | n5882 ;
  assign n5884 = n5837 & n5841 ;
  assign n5885 = n5840 & n5867 ;
  assign n5886 = n5837 & n5885 ;
  assign n5887 = ~n5884 & n5886 ;
  assign n5888 = ~n5883 & n5887 ;
  assign n5889 = n5867 & n5868 ;
  assign n5890 = n5864 & ~n5889 ;
  assign n5891 = ~n5888 & n5890 ;
  assign n5892 = ~n5884 & n5885 ;
  assign n5893 = n5837 & ~n5882 ;
  assign n5894 = ( n5881 & n5890 ) | ( n5881 & n5893 ) | ( n5890 & n5893 ) ;
  assign n5895 = n5890 | n5893 ;
  assign n5896 = ( ~n5892 & n5894 ) | ( ~n5892 & n5895 ) | ( n5894 & n5895 ) ;
  assign n5897 = n5881 | n5893 ;
  assign n5898 = n5892 & ~n5897 ;
  assign n5899 = ( ~n5893 & n5896 ) | ( ~n5893 & n5898 ) | ( n5896 & n5898 ) ;
  assign n5900 = ( ~n5891 & n5896 ) | ( ~n5891 & n5899 ) | ( n5896 & n5899 ) ;
  assign n5901 = n5880 & n5900 ;
  assign n5902 = n5874 & n5878 ;
  assign n5903 = ( n5809 & n5874 ) | ( n5809 & n5902 ) | ( n5874 & n5902 ) ;
  assign n5904 = n5901 | n5903 ;
  assign n5905 = n5881 & ~n5893 ;
  assign n5906 = ( n5892 & n5893 ) | ( n5892 & ~n5905 ) | ( n5893 & ~n5905 ) ;
  assign n5907 = n5890 & n5906 ;
  assign n5908 = ~n5867 & n5868 ;
  assign n5909 = ( ~n5864 & n5868 ) | ( ~n5864 & n5908 ) | ( n5868 & n5908 ) ;
  assign n5910 = ~n5840 & n5841 ;
  assign n5911 = ( ~n5837 & n5841 ) | ( ~n5837 & n5910 ) | ( n5841 & n5910 ) ;
  assign n5912 = ~n5909 & n5911 ;
  assign n5913 = n5909 & ~n5911 ;
  assign n5914 = n5912 | n5913 ;
  assign n5915 = n5888 | n5914 ;
  assign n5916 = n5907 | n5915 ;
  assign n5917 = n5888 & n5914 ;
  assign n5918 = ( n5907 & n5914 ) | ( n5907 & n5917 ) | ( n5914 & n5917 ) ;
  assign n5919 = n5916 & ~n5918 ;
  assign n5920 = n5770 & n5808 ;
  assign n5921 = ~n5767 & n5768 ;
  assign n5922 = ( ~n5764 & n5768 ) | ( ~n5764 & n5921 ) | ( n5768 & n5921 ) ;
  assign n5923 = ~n5786 & n5790 ;
  assign n5924 = ( n5790 & ~n5798 ) | ( n5790 & n5923 ) | ( ~n5798 & n5923 ) ;
  assign n5925 = ~n5922 & n5924 ;
  assign n5926 = n5922 & ~n5924 ;
  assign n5927 = n5925 | n5926 ;
  assign n5928 = n5803 | n5927 ;
  assign n5929 = n5920 | n5928 ;
  assign n5930 = n5803 & n5927 ;
  assign n5931 = ( n5920 & n5927 ) | ( n5920 & n5930 ) | ( n5927 & n5930 ) ;
  assign n5932 = n5929 & ~n5931 ;
  assign n5933 = n5919 | n5932 ;
  assign n5934 = n5904 & n5933 ;
  assign n5935 = n5916 & n5929 ;
  assign n5936 = n5918 | n5931 ;
  assign n5937 = n5935 & ~n5936 ;
  assign n5938 = ( n5803 & n5922 ) | ( n5803 & n5924 ) | ( n5922 & n5924 ) ;
  assign n5939 = n5922 | n5924 ;
  assign n5940 = ( n5920 & n5938 ) | ( n5920 & n5939 ) | ( n5938 & n5939 ) ;
  assign n5941 = ( n5888 & n5909 ) | ( n5888 & n5911 ) | ( n5909 & n5911 ) ;
  assign n5942 = n5909 | n5911 ;
  assign n5943 = ( n5907 & n5941 ) | ( n5907 & n5942 ) | ( n5941 & n5942 ) ;
  assign n5944 = ~n5940 & n5943 ;
  assign n5945 = n5940 & ~n5943 ;
  assign n5946 = n5944 | n5945 ;
  assign n5947 = n5937 | n5946 ;
  assign n5948 = n5934 | n5947 ;
  assign n5949 = n5933 | n5937 ;
  assign n5950 = ( n5904 & n5937 ) | ( n5904 & n5949 ) | ( n5937 & n5949 ) ;
  assign n5951 = n5946 & n5950 ;
  assign n5952 = n5948 & ~n5951 ;
  assign n5953 = ( x190 & x191 ) | ( x190 & x192 ) | ( x191 & x192 ) ;
  assign n5954 = ( x187 & x188 ) | ( x187 & x189 ) | ( x188 & x189 ) ;
  assign n5955 = n5953 & ~n5954 ;
  assign n5956 = ~n5953 & n5954 ;
  assign n5957 = n5955 | n5956 ;
  assign n5958 = ~x187 & x188 ;
  assign n5959 = x187 & ~x188 ;
  assign n5960 = n5958 | n5959 ;
  assign n5961 = ~x189 & n5960 ;
  assign n5962 = x189 & ~n5960 ;
  assign n5963 = n5961 | n5962 ;
  assign n5964 = ~x190 & x191 ;
  assign n5965 = x190 & ~x191 ;
  assign n5966 = n5964 | n5965 ;
  assign n5967 = ~x192 & n5966 ;
  assign n5968 = x192 & ~n5966 ;
  assign n5969 = n5967 | n5968 ;
  assign n5970 = n5963 & n5969 ;
  assign n5971 = n5957 & ~n5970 ;
  assign n5972 = ~n5957 & n5970 ;
  assign n5973 = n5971 | n5972 ;
  assign n5974 = n5963 & ~n5969 ;
  assign n5975 = ~n5963 & n5969 ;
  assign n5976 = n5974 | n5975 ;
  assign n5977 = ( n5953 & n5954 ) | ( n5953 & n5970 ) | ( n5954 & n5970 ) ;
  assign n5978 = n5976 & n5977 ;
  assign n5979 = n5973 & ~n5978 ;
  assign n5980 = n5973 & n5977 ;
  assign n5981 = ~x193 & x194 ;
  assign n5982 = x193 & ~x194 ;
  assign n5983 = n5981 | n5982 ;
  assign n5984 = ~x195 & n5983 ;
  assign n5985 = x195 & ~n5983 ;
  assign n5986 = n5984 | n5985 ;
  assign n5987 = ~x196 & x197 ;
  assign n5988 = x196 & ~x197 ;
  assign n5989 = n5987 | n5988 ;
  assign n5990 = ~x198 & n5989 ;
  assign n5991 = x198 & ~n5989 ;
  assign n5992 = n5990 | n5991 ;
  assign n5993 = n5986 & ~n5992 ;
  assign n5994 = ~n5986 & n5992 ;
  assign n5995 = n5993 | n5994 ;
  assign n5996 = ( x196 & x197 ) | ( x196 & x198 ) | ( x197 & x198 ) ;
  assign n5997 = ( x193 & x194 ) | ( x193 & x195 ) | ( x194 & x195 ) ;
  assign n5998 = n5986 & n5992 ;
  assign n5999 = ( n5996 & n5997 ) | ( n5996 & n5998 ) | ( n5997 & n5998 ) ;
  assign n6000 = n5995 & n5999 ;
  assign n6001 = n5980 | n6000 ;
  assign n6002 = n5996 & ~n5997 ;
  assign n6003 = ~n5996 & n5997 ;
  assign n6004 = n6002 | n6003 ;
  assign n6005 = ~n5998 & n6004 ;
  assign n6006 = n5998 & ~n6004 ;
  assign n6007 = n6005 | n6006 ;
  assign n6008 = n5999 & n6007 ;
  assign n6009 = n5976 & n5995 ;
  assign n6010 = n6007 & n6009 ;
  assign n6011 = ~n6008 & n6010 ;
  assign n6012 = ~n6001 & n6011 ;
  assign n6013 = n5979 & n6012 ;
  assign n6014 = ~n6008 & n6009 ;
  assign n6015 = ~n6000 & n6007 ;
  assign n6016 = n5980 & ~n6015 ;
  assign n6017 = ( n6014 & n6015 ) | ( n6014 & ~n6016 ) | ( n6015 & ~n6016 ) ;
  assign n6018 = ( n5979 & n6013 ) | ( n5979 & ~n6017 ) | ( n6013 & ~n6017 ) ;
  assign n6019 = n5995 & ~n5999 ;
  assign n6020 = ( n5995 & ~n6007 ) | ( n5995 & n6019 ) | ( ~n6007 & n6019 ) ;
  assign n6021 = n5976 & ~n5977 ;
  assign n6022 = ( ~n5973 & n5976 ) | ( ~n5973 & n6021 ) | ( n5976 & n6021 ) ;
  assign n6023 = ~n6020 & n6022 ;
  assign n6024 = n6020 & ~n6022 ;
  assign n6025 = n6023 | n6024 ;
  assign n6026 = ( x184 & x185 ) | ( x184 & x186 ) | ( x185 & x186 ) ;
  assign n6027 = ( x181 & x182 ) | ( x181 & x183 ) | ( x182 & x183 ) ;
  assign n6028 = n6026 & ~n6027 ;
  assign n6029 = ~n6026 & n6027 ;
  assign n6030 = n6028 | n6029 ;
  assign n6031 = ~x181 & x182 ;
  assign n6032 = x181 & ~x182 ;
  assign n6033 = n6031 | n6032 ;
  assign n6034 = ~x183 & n6033 ;
  assign n6035 = x183 & ~n6033 ;
  assign n6036 = n6034 | n6035 ;
  assign n6037 = ~x184 & x185 ;
  assign n6038 = x184 & ~x185 ;
  assign n6039 = n6037 | n6038 ;
  assign n6040 = ~x186 & n6039 ;
  assign n6041 = x186 & ~n6039 ;
  assign n6042 = n6040 | n6041 ;
  assign n6043 = n6036 & n6042 ;
  assign n6044 = n6030 & ~n6043 ;
  assign n6045 = ~n6030 & n6043 ;
  assign n6046 = n6044 | n6045 ;
  assign n6047 = n6036 & ~n6042 ;
  assign n6048 = ~n6036 & n6042 ;
  assign n6049 = n6047 | n6048 ;
  assign n6050 = ( n6026 & n6027 ) | ( n6026 & n6043 ) | ( n6027 & n6043 ) ;
  assign n6051 = n6049 & ~n6050 ;
  assign n6052 = ( ~n6046 & n6049 ) | ( ~n6046 & n6051 ) | ( n6049 & n6051 ) ;
  assign n6053 = ~x175 & x176 ;
  assign n6054 = x175 & ~x176 ;
  assign n6055 = n6053 | n6054 ;
  assign n6056 = ~x177 & n6055 ;
  assign n6057 = x177 & ~n6055 ;
  assign n6058 = n6056 | n6057 ;
  assign n6059 = ~x178 & x179 ;
  assign n6060 = x178 & ~x179 ;
  assign n6061 = n6059 | n6060 ;
  assign n6062 = ~x180 & n6061 ;
  assign n6063 = x180 & ~n6061 ;
  assign n6064 = n6062 | n6063 ;
  assign n6065 = n6058 & ~n6064 ;
  assign n6066 = ~n6058 & n6064 ;
  assign n6067 = n6065 | n6066 ;
  assign n6068 = ( x178 & x179 ) | ( x178 & x180 ) | ( x179 & x180 ) ;
  assign n6069 = ( x175 & x176 ) | ( x175 & x177 ) | ( x176 & x177 ) ;
  assign n6070 = n6068 & ~n6069 ;
  assign n6071 = ~n6068 & n6069 ;
  assign n6072 = n6070 | n6071 ;
  assign n6073 = n6058 & n6064 ;
  assign n6074 = n6072 & ~n6073 ;
  assign n6075 = ~n6072 & n6073 ;
  assign n6076 = n6074 | n6075 ;
  assign n6077 = ( n6068 & n6069 ) | ( n6068 & n6073 ) | ( n6069 & n6073 ) ;
  assign n6078 = n6067 & ~n6077 ;
  assign n6079 = ( n6067 & ~n6076 ) | ( n6067 & n6078 ) | ( ~n6076 & n6078 ) ;
  assign n6080 = ~n6052 & n6079 ;
  assign n6081 = n6052 & ~n6079 ;
  assign n6082 = n6080 | n6081 ;
  assign n6083 = n6025 & n6082 ;
  assign n6084 = ( n5979 & ~n5980 ) | ( n5979 & n6015 ) | ( ~n5980 & n6015 ) ;
  assign n6085 = n5979 & n6015 ;
  assign n6086 = ( n6014 & n6084 ) | ( n6014 & n6085 ) | ( n6084 & n6085 ) ;
  assign n6087 = n6017 & ~n6086 ;
  assign n6088 = n6083 | n6087 ;
  assign n6089 = n6018 | n6088 ;
  assign n6090 = n6076 & n6077 ;
  assign n6091 = n6049 & n6050 ;
  assign n6092 = n6090 | n6091 ;
  assign n6093 = n6046 & n6050 ;
  assign n6094 = n6049 & n6067 ;
  assign n6095 = n6046 & n6094 ;
  assign n6096 = ~n6093 & n6095 ;
  assign n6097 = ~n6092 & n6096 ;
  assign n6098 = n6067 & n6077 ;
  assign n6099 = n6076 & ~n6098 ;
  assign n6100 = ~n6097 & n6099 ;
  assign n6101 = ~n6093 & n6094 ;
  assign n6102 = n6046 & ~n6091 ;
  assign n6103 = ( n6090 & n6099 ) | ( n6090 & n6102 ) | ( n6099 & n6102 ) ;
  assign n6104 = n6099 | n6102 ;
  assign n6105 = ( ~n6101 & n6103 ) | ( ~n6101 & n6104 ) | ( n6103 & n6104 ) ;
  assign n6106 = n6090 | n6102 ;
  assign n6107 = n6101 & ~n6106 ;
  assign n6108 = ( ~n6102 & n6105 ) | ( ~n6102 & n6107 ) | ( n6105 & n6107 ) ;
  assign n6109 = ( ~n6100 & n6105 ) | ( ~n6100 & n6108 ) | ( n6105 & n6108 ) ;
  assign n6110 = n6089 & n6109 ;
  assign n6111 = n6083 & n6087 ;
  assign n6112 = ( n6018 & n6083 ) | ( n6018 & n6111 ) | ( n6083 & n6111 ) ;
  assign n6113 = n6110 | n6112 ;
  assign n6114 = n6090 & ~n6102 ;
  assign n6115 = ( n6101 & n6102 ) | ( n6101 & ~n6114 ) | ( n6102 & ~n6114 ) ;
  assign n6116 = n6099 & n6115 ;
  assign n6117 = ~n6067 & n6077 ;
  assign n6118 = ( ~n6076 & n6077 ) | ( ~n6076 & n6117 ) | ( n6077 & n6117 ) ;
  assign n6119 = ~n6049 & n6050 ;
  assign n6120 = ( ~n6046 & n6050 ) | ( ~n6046 & n6119 ) | ( n6050 & n6119 ) ;
  assign n6121 = ~n6118 & n6120 ;
  assign n6122 = n6118 & ~n6120 ;
  assign n6123 = n6121 | n6122 ;
  assign n6124 = n6097 | n6123 ;
  assign n6125 = n6116 | n6124 ;
  assign n6126 = n6097 & n6123 ;
  assign n6127 = ( n6116 & n6123 ) | ( n6116 & n6126 ) | ( n6123 & n6126 ) ;
  assign n6128 = n6125 & ~n6127 ;
  assign n6129 = n5979 & n6017 ;
  assign n6130 = ~n5976 & n5977 ;
  assign n6131 = ( ~n5973 & n5977 ) | ( ~n5973 & n6130 ) | ( n5977 & n6130 ) ;
  assign n6132 = ~n5995 & n5999 ;
  assign n6133 = ( n5999 & ~n6007 ) | ( n5999 & n6132 ) | ( ~n6007 & n6132 ) ;
  assign n6134 = ~n6131 & n6133 ;
  assign n6135 = n6131 & ~n6133 ;
  assign n6136 = n6134 | n6135 ;
  assign n6137 = n6012 | n6136 ;
  assign n6138 = n6129 | n6137 ;
  assign n6139 = n6012 & n6136 ;
  assign n6140 = ( n6129 & n6136 ) | ( n6129 & n6139 ) | ( n6136 & n6139 ) ;
  assign n6141 = n6138 & ~n6140 ;
  assign n6142 = n6128 | n6141 ;
  assign n6143 = n6113 & n6142 ;
  assign n6144 = n6125 & n6138 ;
  assign n6145 = n6127 | n6140 ;
  assign n6146 = n6144 & ~n6145 ;
  assign n6147 = ( n6012 & n6131 ) | ( n6012 & n6133 ) | ( n6131 & n6133 ) ;
  assign n6148 = n6131 | n6133 ;
  assign n6149 = ( n6129 & n6147 ) | ( n6129 & n6148 ) | ( n6147 & n6148 ) ;
  assign n6150 = ( n6097 & n6118 ) | ( n6097 & n6120 ) | ( n6118 & n6120 ) ;
  assign n6151 = n6118 | n6120 ;
  assign n6152 = ( n6116 & n6150 ) | ( n6116 & n6151 ) | ( n6150 & n6151 ) ;
  assign n6153 = ~n6149 & n6152 ;
  assign n6154 = n6149 & ~n6152 ;
  assign n6155 = n6153 | n6154 ;
  assign n6156 = n6146 | n6155 ;
  assign n6157 = n6143 | n6156 ;
  assign n6158 = n6142 | n6146 ;
  assign n6159 = ( n6113 & n6146 ) | ( n6113 & n6158 ) | ( n6146 & n6158 ) ;
  assign n6160 = n6155 & n6159 ;
  assign n6161 = n6157 & ~n6160 ;
  assign n6162 = n5952 | n6161 ;
  assign n6163 = n5880 & ~n5903 ;
  assign n6164 = n5900 & ~n6163 ;
  assign n6165 = n5816 & ~n5873 ;
  assign n6166 = ~n5816 & n5873 ;
  assign n6167 = n6165 | n6166 ;
  assign n6168 = n6025 & ~n6082 ;
  assign n6169 = ~n6025 & n6082 ;
  assign n6170 = n6168 | n6169 ;
  assign n6171 = n6167 & n6170 ;
  assign n6172 = ~n5874 & n5880 ;
  assign n6173 = n5880 & ~n5900 ;
  assign n6174 = n5809 | n5878 ;
  assign n6175 = n5900 | n6174 ;
  assign n6176 = ( n6172 & n6173 ) | ( n6172 & ~n6175 ) | ( n6173 & ~n6175 ) ;
  assign n6177 = n6171 | n6176 ;
  assign n6178 = n6164 | n6177 ;
  assign n6179 = n6018 | n6087 ;
  assign n6180 = ( n6083 & n6109 ) | ( n6083 & ~n6179 ) | ( n6109 & ~n6179 ) ;
  assign n6181 = ( ~n6109 & n6179 ) | ( ~n6109 & n6180 ) | ( n6179 & n6180 ) ;
  assign n6182 = ( ~n6083 & n6180 ) | ( ~n6083 & n6181 ) | ( n6180 & n6181 ) ;
  assign n6183 = n6178 & n6182 ;
  assign n6184 = n6164 | n6176 ;
  assign n6185 = n6171 & n6184 ;
  assign n6186 = ( n6112 & ~n6128 ) | ( n6112 & n6141 ) | ( ~n6128 & n6141 ) ;
  assign n6187 = n6128 & ~n6141 ;
  assign n6188 = ( n6110 & n6186 ) | ( n6110 & ~n6187 ) | ( n6186 & ~n6187 ) ;
  assign n6189 = ( ~n6113 & n6128 ) | ( ~n6113 & n6188 ) | ( n6128 & n6188 ) ;
  assign n6190 = ( ~n6141 & n6188 ) | ( ~n6141 & n6189 ) | ( n6188 & n6189 ) ;
  assign n6191 = ( n5903 & ~n5919 ) | ( n5903 & n5932 ) | ( ~n5919 & n5932 ) ;
  assign n6192 = n5919 & ~n5932 ;
  assign n6193 = ( n5901 & n6191 ) | ( n5901 & ~n6192 ) | ( n6191 & ~n6192 ) ;
  assign n6194 = ( ~n5904 & n5919 ) | ( ~n5904 & n6193 ) | ( n5919 & n6193 ) ;
  assign n6195 = ( ~n5932 & n6193 ) | ( ~n5932 & n6194 ) | ( n6193 & n6194 ) ;
  assign n6196 = ( n6185 & n6190 ) | ( n6185 & n6195 ) | ( n6190 & n6195 ) ;
  assign n6197 = n6190 | n6195 ;
  assign n6198 = ( n6183 & n6196 ) | ( n6183 & n6197 ) | ( n6196 & n6197 ) ;
  assign n6199 = n6162 & n6198 ;
  assign n6200 = n5948 & n6157 ;
  assign n6201 = n5951 | n6160 ;
  assign n6202 = n6200 & ~n6201 ;
  assign n6203 = n6149 & n6152 ;
  assign n6204 = n6149 | n6152 ;
  assign n6205 = n6203 | n6204 ;
  assign n6206 = ( n6159 & n6203 ) | ( n6159 & n6205 ) | ( n6203 & n6205 ) ;
  assign n6207 = n5940 & n5943 ;
  assign n6208 = n5940 | n5943 ;
  assign n6209 = n6207 | n6208 ;
  assign n6210 = ( n5950 & n6207 ) | ( n5950 & n6209 ) | ( n6207 & n6209 ) ;
  assign n6211 = n6206 & n6210 ;
  assign n6212 = n6210 & ~n6211 ;
  assign n6213 = ( n6206 & ~n6211 ) | ( n6206 & n6212 ) | ( ~n6211 & n6212 ) ;
  assign n6214 = n6202 | n6213 ;
  assign n6215 = n6199 | n6214 ;
  assign n6216 = n6199 | n6202 ;
  assign n6217 = n6213 & n6216 ;
  assign n6218 = n6215 & ~n6217 ;
  assign n6219 = ~x259 & x260 ;
  assign n6220 = x259 & ~x260 ;
  assign n6221 = n6219 | n6220 ;
  assign n6222 = ~x261 & n6221 ;
  assign n6223 = x261 & ~n6221 ;
  assign n6224 = n6222 | n6223 ;
  assign n6225 = ~x262 & x263 ;
  assign n6226 = x262 & ~x263 ;
  assign n6227 = n6225 | n6226 ;
  assign n6228 = ~x264 & n6227 ;
  assign n6229 = x264 & ~n6227 ;
  assign n6230 = n6228 | n6229 ;
  assign n6231 = n6224 & n6230 ;
  assign n6232 = ( x262 & x263 ) | ( x262 & x264 ) | ( x263 & x264 ) ;
  assign n6233 = ( x259 & x260 ) | ( x259 & x261 ) | ( x260 & x261 ) ;
  assign n6234 = ~n6232 & n6233 ;
  assign n6235 = n6232 & ~n6233 ;
  assign n6236 = n6234 | n6235 ;
  assign n6237 = ~n6231 & n6236 ;
  assign n6238 = n6231 & ~n6236 ;
  assign n6239 = n6237 | n6238 ;
  assign n6240 = n6224 & ~n6230 ;
  assign n6241 = ~n6224 & n6230 ;
  assign n6242 = n6240 | n6241 ;
  assign n6243 = ( n6231 & n6232 ) | ( n6231 & n6233 ) | ( n6232 & n6233 ) ;
  assign n6244 = n6242 & n6243 ;
  assign n6245 = n6239 & ~n6244 ;
  assign n6246 = n6239 & n6243 ;
  assign n6247 = x265 & ~x266 ;
  assign n6248 = ~x265 & x266 ;
  assign n6249 = n6247 | n6248 ;
  assign n6250 = ~x267 & n6249 ;
  assign n6251 = x267 & ~n6249 ;
  assign n6252 = n6250 | n6251 ;
  assign n6253 = x268 & ~x269 ;
  assign n6254 = ~x268 & x269 ;
  assign n6255 = n6253 | n6254 ;
  assign n6256 = ~x270 & n6255 ;
  assign n6257 = x270 & ~n6255 ;
  assign n6258 = n6256 | n6257 ;
  assign n6259 = n6252 & ~n6258 ;
  assign n6260 = ~n6252 & n6258 ;
  assign n6261 = n6259 | n6260 ;
  assign n6262 = ( x268 & x269 ) | ( x268 & x270 ) | ( x269 & x270 ) ;
  assign n6263 = ( x265 & x266 ) | ( x265 & x267 ) | ( x266 & x267 ) ;
  assign n6264 = n6252 & n6258 ;
  assign n6265 = ( n6262 & n6263 ) | ( n6262 & n6264 ) | ( n6263 & n6264 ) ;
  assign n6266 = n6261 & n6265 ;
  assign n6267 = n6246 | n6266 ;
  assign n6268 = n6262 & ~n6263 ;
  assign n6269 = ~n6262 & n6263 ;
  assign n6270 = n6268 | n6269 ;
  assign n6271 = ~n6264 & n6270 ;
  assign n6272 = n6264 & ~n6270 ;
  assign n6273 = n6271 | n6272 ;
  assign n6274 = n6265 & n6273 ;
  assign n6275 = n6242 & n6261 ;
  assign n6276 = n6273 & n6275 ;
  assign n6277 = ~n6274 & n6276 ;
  assign n6278 = ~n6267 & n6277 ;
  assign n6279 = n6245 & n6278 ;
  assign n6280 = ~n6274 & n6275 ;
  assign n6281 = ~n6266 & n6273 ;
  assign n6282 = n6246 & ~n6281 ;
  assign n6283 = ( n6280 & n6281 ) | ( n6280 & ~n6282 ) | ( n6281 & ~n6282 ) ;
  assign n6284 = ( n6245 & n6279 ) | ( n6245 & ~n6283 ) | ( n6279 & ~n6283 ) ;
  assign n6285 = n6261 & ~n6265 ;
  assign n6286 = ( n6261 & ~n6273 ) | ( n6261 & n6285 ) | ( ~n6273 & n6285 ) ;
  assign n6287 = n6242 & ~n6243 ;
  assign n6288 = ( ~n6239 & n6242 ) | ( ~n6239 & n6287 ) | ( n6242 & n6287 ) ;
  assign n6289 = ~n6286 & n6288 ;
  assign n6290 = n6286 & ~n6288 ;
  assign n6291 = n6289 | n6290 ;
  assign n6292 = ( x256 & x257 ) | ( x256 & x258 ) | ( x257 & x258 ) ;
  assign n6293 = ( x253 & x254 ) | ( x253 & x255 ) | ( x254 & x255 ) ;
  assign n6294 = n6292 & ~n6293 ;
  assign n6295 = ~n6292 & n6293 ;
  assign n6296 = n6294 | n6295 ;
  assign n6297 = x253 & ~x254 ;
  assign n6298 = ~x253 & x254 ;
  assign n6299 = n6297 | n6298 ;
  assign n6300 = ~x255 & n6299 ;
  assign n6301 = x255 & ~n6299 ;
  assign n6302 = n6300 | n6301 ;
  assign n6303 = x256 & ~x257 ;
  assign n6304 = ~x256 & x257 ;
  assign n6305 = n6303 | n6304 ;
  assign n6306 = ~x258 & n6305 ;
  assign n6307 = x258 & ~n6305 ;
  assign n6308 = n6306 | n6307 ;
  assign n6309 = n6302 & n6308 ;
  assign n6310 = n6296 & ~n6309 ;
  assign n6311 = ~n6296 & n6309 ;
  assign n6312 = n6310 | n6311 ;
  assign n6313 = n6302 & ~n6308 ;
  assign n6314 = ~n6302 & n6308 ;
  assign n6315 = n6313 | n6314 ;
  assign n6316 = ( n6292 & n6293 ) | ( n6292 & n6309 ) | ( n6293 & n6309 ) ;
  assign n6317 = n6315 & ~n6316 ;
  assign n6318 = ( ~n6312 & n6315 ) | ( ~n6312 & n6317 ) | ( n6315 & n6317 ) ;
  assign n6319 = ~x247 & x248 ;
  assign n6320 = x247 & ~x248 ;
  assign n6321 = n6319 | n6320 ;
  assign n6322 = ~x249 & n6321 ;
  assign n6323 = x249 & ~n6321 ;
  assign n6324 = n6322 | n6323 ;
  assign n6325 = ~x250 & x251 ;
  assign n6326 = x250 & ~x251 ;
  assign n6327 = n6325 | n6326 ;
  assign n6328 = ~x252 & n6327 ;
  assign n6329 = x252 & ~n6327 ;
  assign n6330 = n6328 | n6329 ;
  assign n6331 = n6324 & n6330 ;
  assign n6332 = ( x250 & x251 ) | ( x250 & x252 ) | ( x251 & x252 ) ;
  assign n6333 = ( x247 & x248 ) | ( x247 & x249 ) | ( x248 & x249 ) ;
  assign n6334 = ~n6332 & n6333 ;
  assign n6335 = n6332 & ~n6333 ;
  assign n6336 = n6334 | n6335 ;
  assign n6337 = ~n6331 & n6336 ;
  assign n6338 = n6331 & ~n6336 ;
  assign n6339 = n6337 | n6338 ;
  assign n6340 = n6324 & ~n6330 ;
  assign n6341 = ~n6324 & n6330 ;
  assign n6342 = n6340 | n6341 ;
  assign n6343 = ( n6331 & n6332 ) | ( n6331 & n6333 ) | ( n6332 & n6333 ) ;
  assign n6344 = n6342 & ~n6343 ;
  assign n6345 = ( ~n6339 & n6342 ) | ( ~n6339 & n6344 ) | ( n6342 & n6344 ) ;
  assign n6346 = ~n6318 & n6345 ;
  assign n6347 = n6318 & ~n6345 ;
  assign n6348 = n6346 | n6347 ;
  assign n6349 = n6291 & n6348 ;
  assign n6350 = ( n6245 & ~n6246 ) | ( n6245 & n6281 ) | ( ~n6246 & n6281 ) ;
  assign n6351 = n6245 & n6281 ;
  assign n6352 = ( n6280 & n6350 ) | ( n6280 & n6351 ) | ( n6350 & n6351 ) ;
  assign n6353 = n6283 & ~n6352 ;
  assign n6354 = n6349 | n6353 ;
  assign n6355 = n6284 | n6354 ;
  assign n6356 = n6339 & n6343 ;
  assign n6357 = n6315 & n6316 ;
  assign n6358 = n6356 | n6357 ;
  assign n6359 = n6312 & n6316 ;
  assign n6360 = n6315 & n6342 ;
  assign n6361 = n6312 & n6360 ;
  assign n6362 = ~n6359 & n6361 ;
  assign n6363 = ~n6358 & n6362 ;
  assign n6364 = n6342 & n6343 ;
  assign n6365 = n6339 & ~n6364 ;
  assign n6366 = ~n6363 & n6365 ;
  assign n6367 = ~n6359 & n6360 ;
  assign n6368 = n6312 & ~n6357 ;
  assign n6369 = ( n6356 & n6365 ) | ( n6356 & n6368 ) | ( n6365 & n6368 ) ;
  assign n6370 = n6365 | n6368 ;
  assign n6371 = ( ~n6367 & n6369 ) | ( ~n6367 & n6370 ) | ( n6369 & n6370 ) ;
  assign n6372 = n6356 | n6368 ;
  assign n6373 = n6367 & ~n6372 ;
  assign n6374 = ( ~n6368 & n6371 ) | ( ~n6368 & n6373 ) | ( n6371 & n6373 ) ;
  assign n6375 = ( ~n6366 & n6371 ) | ( ~n6366 & n6374 ) | ( n6371 & n6374 ) ;
  assign n6376 = n6355 & n6375 ;
  assign n6377 = n6349 & n6353 ;
  assign n6378 = ( n6284 & n6349 ) | ( n6284 & n6377 ) | ( n6349 & n6377 ) ;
  assign n6379 = n6376 | n6378 ;
  assign n6380 = n6356 & ~n6368 ;
  assign n6381 = ( n6367 & n6368 ) | ( n6367 & ~n6380 ) | ( n6368 & ~n6380 ) ;
  assign n6382 = n6365 & n6381 ;
  assign n6383 = ~n6342 & n6343 ;
  assign n6384 = ( ~n6339 & n6343 ) | ( ~n6339 & n6383 ) | ( n6343 & n6383 ) ;
  assign n6385 = ~n6315 & n6316 ;
  assign n6386 = ( ~n6312 & n6316 ) | ( ~n6312 & n6385 ) | ( n6316 & n6385 ) ;
  assign n6387 = ~n6384 & n6386 ;
  assign n6388 = n6384 & ~n6386 ;
  assign n6389 = n6387 | n6388 ;
  assign n6390 = n6363 | n6389 ;
  assign n6391 = n6382 | n6390 ;
  assign n6392 = n6363 & n6389 ;
  assign n6393 = ( n6382 & n6389 ) | ( n6382 & n6392 ) | ( n6389 & n6392 ) ;
  assign n6394 = n6391 & ~n6393 ;
  assign n6395 = n6245 & n6283 ;
  assign n6396 = ~n6242 & n6243 ;
  assign n6397 = ( ~n6239 & n6243 ) | ( ~n6239 & n6396 ) | ( n6243 & n6396 ) ;
  assign n6398 = ~n6261 & n6265 ;
  assign n6399 = ( n6265 & ~n6273 ) | ( n6265 & n6398 ) | ( ~n6273 & n6398 ) ;
  assign n6400 = ~n6397 & n6399 ;
  assign n6401 = n6397 & ~n6399 ;
  assign n6402 = n6400 | n6401 ;
  assign n6403 = n6278 | n6402 ;
  assign n6404 = n6395 | n6403 ;
  assign n6405 = n6278 & n6402 ;
  assign n6406 = ( n6395 & n6402 ) | ( n6395 & n6405 ) | ( n6402 & n6405 ) ;
  assign n6407 = n6404 & ~n6406 ;
  assign n6408 = n6394 | n6407 ;
  assign n6409 = n6379 & n6408 ;
  assign n6410 = n6391 & n6404 ;
  assign n6411 = n6393 | n6406 ;
  assign n6412 = n6410 & ~n6411 ;
  assign n6413 = ( n6278 & n6397 ) | ( n6278 & n6399 ) | ( n6397 & n6399 ) ;
  assign n6414 = n6397 | n6399 ;
  assign n6415 = ( n6395 & n6413 ) | ( n6395 & n6414 ) | ( n6413 & n6414 ) ;
  assign n6416 = ( n6363 & n6384 ) | ( n6363 & n6386 ) | ( n6384 & n6386 ) ;
  assign n6417 = n6384 | n6386 ;
  assign n6418 = ( n6382 & n6416 ) | ( n6382 & n6417 ) | ( n6416 & n6417 ) ;
  assign n6419 = ~n6415 & n6418 ;
  assign n6420 = n6415 & ~n6418 ;
  assign n6421 = n6419 | n6420 ;
  assign n6422 = n6412 | n6421 ;
  assign n6423 = n6409 | n6422 ;
  assign n6424 = n6408 | n6412 ;
  assign n6425 = ( n6379 & n6412 ) | ( n6379 & n6424 ) | ( n6412 & n6424 ) ;
  assign n6426 = n6421 & n6425 ;
  assign n6427 = n6423 & ~n6426 ;
  assign n6428 = ~x235 & x236 ;
  assign n6429 = x235 & ~x236 ;
  assign n6430 = n6428 | n6429 ;
  assign n6431 = ~x237 & n6430 ;
  assign n6432 = x237 & ~n6430 ;
  assign n6433 = n6431 | n6432 ;
  assign n6434 = ~x238 & x239 ;
  assign n6435 = x238 & ~x239 ;
  assign n6436 = n6434 | n6435 ;
  assign n6437 = ~x240 & n6436 ;
  assign n6438 = x240 & ~n6436 ;
  assign n6439 = n6437 | n6438 ;
  assign n6440 = n6433 & n6439 ;
  assign n6441 = ( x238 & x239 ) | ( x238 & x240 ) | ( x239 & x240 ) ;
  assign n6442 = ( x235 & x236 ) | ( x235 & x237 ) | ( x236 & x237 ) ;
  assign n6443 = ~n6441 & n6442 ;
  assign n6444 = n6441 & ~n6442 ;
  assign n6445 = n6443 | n6444 ;
  assign n6446 = ~n6440 & n6445 ;
  assign n6447 = n6440 & ~n6445 ;
  assign n6448 = n6446 | n6447 ;
  assign n6449 = n6433 & ~n6439 ;
  assign n6450 = ~n6433 & n6439 ;
  assign n6451 = n6449 | n6450 ;
  assign n6452 = ( n6440 & n6441 ) | ( n6440 & n6442 ) | ( n6441 & n6442 ) ;
  assign n6453 = n6451 & n6452 ;
  assign n6454 = n6448 & ~n6453 ;
  assign n6455 = n6448 & n6452 ;
  assign n6456 = x241 & ~x242 ;
  assign n6457 = ~x241 & x242 ;
  assign n6458 = n6456 | n6457 ;
  assign n6459 = ~x243 & n6458 ;
  assign n6460 = x243 & ~n6458 ;
  assign n6461 = n6459 | n6460 ;
  assign n6462 = x244 & ~x245 ;
  assign n6463 = ~x244 & x245 ;
  assign n6464 = n6462 | n6463 ;
  assign n6465 = ~x246 & n6464 ;
  assign n6466 = x246 & ~n6464 ;
  assign n6467 = n6465 | n6466 ;
  assign n6468 = n6461 & ~n6467 ;
  assign n6469 = ~n6461 & n6467 ;
  assign n6470 = n6468 | n6469 ;
  assign n6471 = ( x244 & x245 ) | ( x244 & x246 ) | ( x245 & x246 ) ;
  assign n6472 = ( x241 & x242 ) | ( x241 & x243 ) | ( x242 & x243 ) ;
  assign n6473 = n6461 & n6467 ;
  assign n6474 = ( n6471 & n6472 ) | ( n6471 & n6473 ) | ( n6472 & n6473 ) ;
  assign n6475 = n6470 & n6474 ;
  assign n6476 = n6455 | n6475 ;
  assign n6477 = n6471 & ~n6472 ;
  assign n6478 = ~n6471 & n6472 ;
  assign n6479 = n6477 | n6478 ;
  assign n6480 = ~n6473 & n6479 ;
  assign n6481 = n6473 & ~n6479 ;
  assign n6482 = n6480 | n6481 ;
  assign n6483 = n6474 & n6482 ;
  assign n6484 = n6451 & n6470 ;
  assign n6485 = n6482 & n6484 ;
  assign n6486 = ~n6483 & n6485 ;
  assign n6487 = ~n6476 & n6486 ;
  assign n6488 = n6454 & n6487 ;
  assign n6489 = ~n6483 & n6484 ;
  assign n6490 = ~n6475 & n6482 ;
  assign n6491 = n6455 & ~n6490 ;
  assign n6492 = ( n6489 & n6490 ) | ( n6489 & ~n6491 ) | ( n6490 & ~n6491 ) ;
  assign n6493 = ( n6454 & n6488 ) | ( n6454 & ~n6492 ) | ( n6488 & ~n6492 ) ;
  assign n6494 = n6470 & ~n6474 ;
  assign n6495 = ( n6470 & ~n6482 ) | ( n6470 & n6494 ) | ( ~n6482 & n6494 ) ;
  assign n6496 = n6451 & ~n6452 ;
  assign n6497 = ( ~n6448 & n6451 ) | ( ~n6448 & n6496 ) | ( n6451 & n6496 ) ;
  assign n6498 = ~n6495 & n6497 ;
  assign n6499 = n6495 & ~n6497 ;
  assign n6500 = n6498 | n6499 ;
  assign n6501 = ( x232 & x233 ) | ( x232 & x234 ) | ( x233 & x234 ) ;
  assign n6502 = ( x229 & x230 ) | ( x229 & x231 ) | ( x230 & x231 ) ;
  assign n6503 = n6501 & ~n6502 ;
  assign n6504 = ~n6501 & n6502 ;
  assign n6505 = n6503 | n6504 ;
  assign n6506 = ~x229 & x230 ;
  assign n6507 = x229 & ~x230 ;
  assign n6508 = n6506 | n6507 ;
  assign n6509 = ~x231 & n6508 ;
  assign n6510 = x231 & ~n6508 ;
  assign n6511 = n6509 | n6510 ;
  assign n6512 = ~x232 & x233 ;
  assign n6513 = x232 & ~x233 ;
  assign n6514 = n6512 | n6513 ;
  assign n6515 = ~x234 & n6514 ;
  assign n6516 = x234 & ~n6514 ;
  assign n6517 = n6515 | n6516 ;
  assign n6518 = n6511 & n6517 ;
  assign n6519 = n6505 & ~n6518 ;
  assign n6520 = ~n6505 & n6518 ;
  assign n6521 = n6519 | n6520 ;
  assign n6522 = n6511 & ~n6517 ;
  assign n6523 = ~n6511 & n6517 ;
  assign n6524 = n6522 | n6523 ;
  assign n6525 = ( n6501 & n6502 ) | ( n6501 & n6518 ) | ( n6502 & n6518 ) ;
  assign n6526 = n6524 & ~n6525 ;
  assign n6527 = ( ~n6521 & n6524 ) | ( ~n6521 & n6526 ) | ( n6524 & n6526 ) ;
  assign n6528 = ~x223 & x224 ;
  assign n6529 = x223 & ~x224 ;
  assign n6530 = n6528 | n6529 ;
  assign n6531 = ~x225 & n6530 ;
  assign n6532 = x225 & ~n6530 ;
  assign n6533 = n6531 | n6532 ;
  assign n6534 = ~x226 & x227 ;
  assign n6535 = x226 & ~x227 ;
  assign n6536 = n6534 | n6535 ;
  assign n6537 = ~x228 & n6536 ;
  assign n6538 = x228 & ~n6536 ;
  assign n6539 = n6537 | n6538 ;
  assign n6540 = n6533 & ~n6539 ;
  assign n6541 = ~n6533 & n6539 ;
  assign n6542 = n6540 | n6541 ;
  assign n6543 = ( x226 & x227 ) | ( x226 & x228 ) | ( x227 & x228 ) ;
  assign n6544 = ( x223 & x224 ) | ( x223 & x225 ) | ( x224 & x225 ) ;
  assign n6545 = n6543 & ~n6544 ;
  assign n6546 = ~n6543 & n6544 ;
  assign n6547 = n6545 | n6546 ;
  assign n6548 = n6533 & n6539 ;
  assign n6549 = n6547 & ~n6548 ;
  assign n6550 = ~n6547 & n6548 ;
  assign n6551 = n6549 | n6550 ;
  assign n6552 = ( n6543 & n6544 ) | ( n6543 & n6548 ) | ( n6544 & n6548 ) ;
  assign n6553 = n6542 & ~n6552 ;
  assign n6554 = ( n6542 & ~n6551 ) | ( n6542 & n6553 ) | ( ~n6551 & n6553 ) ;
  assign n6555 = ~n6527 & n6554 ;
  assign n6556 = n6527 & ~n6554 ;
  assign n6557 = n6555 | n6556 ;
  assign n6558 = n6500 & n6557 ;
  assign n6559 = ( n6454 & ~n6455 ) | ( n6454 & n6490 ) | ( ~n6455 & n6490 ) ;
  assign n6560 = n6454 & n6490 ;
  assign n6561 = ( n6489 & n6559 ) | ( n6489 & n6560 ) | ( n6559 & n6560 ) ;
  assign n6562 = n6492 & ~n6561 ;
  assign n6563 = n6558 | n6562 ;
  assign n6564 = n6493 | n6563 ;
  assign n6565 = n6551 & n6552 ;
  assign n6566 = n6524 & n6525 ;
  assign n6567 = n6565 | n6566 ;
  assign n6568 = n6521 & n6525 ;
  assign n6569 = n6524 & n6542 ;
  assign n6570 = n6521 & n6569 ;
  assign n6571 = ~n6568 & n6570 ;
  assign n6572 = ~n6567 & n6571 ;
  assign n6573 = n6542 & n6552 ;
  assign n6574 = n6551 & ~n6573 ;
  assign n6575 = ~n6572 & n6574 ;
  assign n6576 = ~n6568 & n6569 ;
  assign n6577 = n6521 & ~n6566 ;
  assign n6578 = ( n6565 & n6574 ) | ( n6565 & n6577 ) | ( n6574 & n6577 ) ;
  assign n6579 = n6574 | n6577 ;
  assign n6580 = ( ~n6576 & n6578 ) | ( ~n6576 & n6579 ) | ( n6578 & n6579 ) ;
  assign n6581 = n6565 | n6577 ;
  assign n6582 = n6576 & ~n6581 ;
  assign n6583 = ( ~n6577 & n6580 ) | ( ~n6577 & n6582 ) | ( n6580 & n6582 ) ;
  assign n6584 = ( ~n6575 & n6580 ) | ( ~n6575 & n6583 ) | ( n6580 & n6583 ) ;
  assign n6585 = n6564 & n6584 ;
  assign n6586 = n6558 & n6562 ;
  assign n6587 = ( n6493 & n6558 ) | ( n6493 & n6586 ) | ( n6558 & n6586 ) ;
  assign n6588 = n6585 | n6587 ;
  assign n6589 = n6565 & ~n6577 ;
  assign n6590 = ( n6576 & n6577 ) | ( n6576 & ~n6589 ) | ( n6577 & ~n6589 ) ;
  assign n6591 = n6574 & n6590 ;
  assign n6592 = ~n6542 & n6552 ;
  assign n6593 = ( ~n6551 & n6552 ) | ( ~n6551 & n6592 ) | ( n6552 & n6592 ) ;
  assign n6594 = ~n6524 & n6525 ;
  assign n6595 = ( ~n6521 & n6525 ) | ( ~n6521 & n6594 ) | ( n6525 & n6594 ) ;
  assign n6596 = ~n6593 & n6595 ;
  assign n6597 = n6593 & ~n6595 ;
  assign n6598 = n6596 | n6597 ;
  assign n6599 = n6572 | n6598 ;
  assign n6600 = n6591 | n6599 ;
  assign n6601 = n6572 & n6598 ;
  assign n6602 = ( n6591 & n6598 ) | ( n6591 & n6601 ) | ( n6598 & n6601 ) ;
  assign n6603 = n6600 & ~n6602 ;
  assign n6604 = n6454 & n6492 ;
  assign n6605 = ~n6451 & n6452 ;
  assign n6606 = ( ~n6448 & n6452 ) | ( ~n6448 & n6605 ) | ( n6452 & n6605 ) ;
  assign n6607 = ~n6470 & n6474 ;
  assign n6608 = ( n6474 & ~n6482 ) | ( n6474 & n6607 ) | ( ~n6482 & n6607 ) ;
  assign n6609 = ~n6606 & n6608 ;
  assign n6610 = n6606 & ~n6608 ;
  assign n6611 = n6609 | n6610 ;
  assign n6612 = n6487 | n6611 ;
  assign n6613 = n6604 | n6612 ;
  assign n6614 = n6487 & n6611 ;
  assign n6615 = ( n6604 & n6611 ) | ( n6604 & n6614 ) | ( n6611 & n6614 ) ;
  assign n6616 = n6613 & ~n6615 ;
  assign n6617 = n6603 | n6616 ;
  assign n6618 = n6588 & n6617 ;
  assign n6619 = n6600 & n6613 ;
  assign n6620 = n6602 | n6615 ;
  assign n6621 = n6619 & ~n6620 ;
  assign n6622 = ( n6487 & n6606 ) | ( n6487 & n6608 ) | ( n6606 & n6608 ) ;
  assign n6623 = n6606 | n6608 ;
  assign n6624 = ( n6604 & n6622 ) | ( n6604 & n6623 ) | ( n6622 & n6623 ) ;
  assign n6625 = ( n6572 & n6593 ) | ( n6572 & n6595 ) | ( n6593 & n6595 ) ;
  assign n6626 = n6593 | n6595 ;
  assign n6627 = ( n6591 & n6625 ) | ( n6591 & n6626 ) | ( n6625 & n6626 ) ;
  assign n6628 = ~n6624 & n6627 ;
  assign n6629 = n6624 & ~n6627 ;
  assign n6630 = n6628 | n6629 ;
  assign n6631 = n6621 | n6630 ;
  assign n6632 = n6618 | n6631 ;
  assign n6633 = n6617 | n6621 ;
  assign n6634 = ( n6588 & n6621 ) | ( n6588 & n6633 ) | ( n6621 & n6633 ) ;
  assign n6635 = n6630 & n6634 ;
  assign n6636 = n6632 & ~n6635 ;
  assign n6637 = n6427 | n6636 ;
  assign n6638 = n6355 & ~n6378 ;
  assign n6639 = n6375 & ~n6638 ;
  assign n6640 = n6291 & ~n6348 ;
  assign n6641 = ~n6291 & n6348 ;
  assign n6642 = n6640 | n6641 ;
  assign n6643 = n6500 & ~n6557 ;
  assign n6644 = ~n6500 & n6557 ;
  assign n6645 = n6643 | n6644 ;
  assign n6646 = n6642 & n6645 ;
  assign n6647 = ~n6349 & n6355 ;
  assign n6648 = n6355 & ~n6375 ;
  assign n6649 = n6284 | n6353 ;
  assign n6650 = n6375 | n6649 ;
  assign n6651 = ( n6647 & n6648 ) | ( n6647 & ~n6650 ) | ( n6648 & ~n6650 ) ;
  assign n6652 = n6646 | n6651 ;
  assign n6653 = n6639 | n6652 ;
  assign n6654 = n6493 | n6562 ;
  assign n6655 = ( n6558 & n6584 ) | ( n6558 & ~n6654 ) | ( n6584 & ~n6654 ) ;
  assign n6656 = ( ~n6584 & n6654 ) | ( ~n6584 & n6655 ) | ( n6654 & n6655 ) ;
  assign n6657 = ( ~n6558 & n6655 ) | ( ~n6558 & n6656 ) | ( n6655 & n6656 ) ;
  assign n6658 = n6653 & n6657 ;
  assign n6659 = n6639 | n6651 ;
  assign n6660 = n6646 & n6659 ;
  assign n6661 = ( n6587 & ~n6603 ) | ( n6587 & n6616 ) | ( ~n6603 & n6616 ) ;
  assign n6662 = n6603 & ~n6616 ;
  assign n6663 = ( n6585 & n6661 ) | ( n6585 & ~n6662 ) | ( n6661 & ~n6662 ) ;
  assign n6664 = ( ~n6588 & n6603 ) | ( ~n6588 & n6663 ) | ( n6603 & n6663 ) ;
  assign n6665 = ( ~n6616 & n6663 ) | ( ~n6616 & n6664 ) | ( n6663 & n6664 ) ;
  assign n6666 = ( n6378 & ~n6394 ) | ( n6378 & n6407 ) | ( ~n6394 & n6407 ) ;
  assign n6667 = n6394 & ~n6407 ;
  assign n6668 = ( n6376 & n6666 ) | ( n6376 & ~n6667 ) | ( n6666 & ~n6667 ) ;
  assign n6669 = ( ~n6379 & n6394 ) | ( ~n6379 & n6668 ) | ( n6394 & n6668 ) ;
  assign n6670 = ( ~n6407 & n6668 ) | ( ~n6407 & n6669 ) | ( n6668 & n6669 ) ;
  assign n6671 = ( n6660 & n6665 ) | ( n6660 & n6670 ) | ( n6665 & n6670 ) ;
  assign n6672 = n6665 | n6670 ;
  assign n6673 = ( n6658 & n6671 ) | ( n6658 & n6672 ) | ( n6671 & n6672 ) ;
  assign n6674 = n6637 & n6673 ;
  assign n6675 = n6423 & n6632 ;
  assign n6676 = n6426 | n6635 ;
  assign n6677 = n6675 & ~n6676 ;
  assign n6678 = n6624 & n6627 ;
  assign n6679 = n6624 | n6627 ;
  assign n6680 = n6678 | n6679 ;
  assign n6681 = ( n6634 & n6678 ) | ( n6634 & n6680 ) | ( n6678 & n6680 ) ;
  assign n6682 = n6415 & n6418 ;
  assign n6683 = n6415 | n6418 ;
  assign n6684 = n6682 | n6683 ;
  assign n6685 = ( n6425 & n6682 ) | ( n6425 & n6684 ) | ( n6682 & n6684 ) ;
  assign n6686 = n6681 & n6685 ;
  assign n6687 = n6685 & ~n6686 ;
  assign n6688 = ( n6681 & ~n6686 ) | ( n6681 & n6687 ) | ( ~n6686 & n6687 ) ;
  assign n6689 = n6677 | n6688 ;
  assign n6690 = n6674 | n6689 ;
  assign n6691 = n6674 | n6677 ;
  assign n6692 = n6688 & n6691 ;
  assign n6693 = n6690 & ~n6692 ;
  assign n6694 = n6218 | n6693 ;
  assign n6695 = ( ~n6427 & n6636 ) | ( ~n6427 & n6673 ) | ( n6636 & n6673 ) ;
  assign n6696 = ( n6427 & ~n6673 ) | ( n6427 & n6695 ) | ( ~n6673 & n6695 ) ;
  assign n6697 = ( ~n6636 & n6695 ) | ( ~n6636 & n6696 ) | ( n6695 & n6696 ) ;
  assign n6698 = ( ~n5952 & n6161 ) | ( ~n5952 & n6198 ) | ( n6161 & n6198 ) ;
  assign n6699 = ( n5952 & ~n6198 ) | ( n5952 & n6698 ) | ( ~n6198 & n6698 ) ;
  assign n6700 = ( ~n6161 & n6698 ) | ( ~n6161 & n6699 ) | ( n6698 & n6699 ) ;
  assign n6701 = ~n6171 & n6184 ;
  assign n6702 = n6171 & ~n6176 ;
  assign n6703 = ~n6164 & n6702 ;
  assign n6704 = ~n6182 & n6703 ;
  assign n6705 = ( ~n6182 & n6701 ) | ( ~n6182 & n6704 ) | ( n6701 & n6704 ) ;
  assign n6706 = n6183 & ~n6185 ;
  assign n6707 = ( n6182 & n6705 ) | ( n6182 & ~n6706 ) | ( n6705 & ~n6706 ) ;
  assign n6708 = n6642 & ~n6645 ;
  assign n6709 = ~n6642 & n6645 ;
  assign n6710 = n6708 | n6709 ;
  assign n6711 = n6167 & ~n6170 ;
  assign n6712 = ~n6167 & n6170 ;
  assign n6713 = n6711 | n6712 ;
  assign n6714 = n6710 & n6713 ;
  assign n6715 = ~n6653 & n6657 ;
  assign n6716 = ( n6657 & n6660 ) | ( n6657 & n6715 ) | ( n6660 & n6715 ) ;
  assign n6717 = ~n6646 & n6659 ;
  assign n6718 = n6646 & ~n6651 ;
  assign n6719 = ~n6639 & n6718 ;
  assign n6720 = ~n6657 & n6719 ;
  assign n6721 = ( ~n6657 & n6717 ) | ( ~n6657 & n6720 ) | ( n6717 & n6720 ) ;
  assign n6722 = n6716 | n6721 ;
  assign n6723 = n6714 | n6722 ;
  assign n6724 = n6707 & n6723 ;
  assign n6725 = n6714 & n6722 ;
  assign n6727 = ( n6185 & ~n6190 ) | ( n6185 & n6195 ) | ( ~n6190 & n6195 ) ;
  assign n6728 = n6190 & ~n6195 ;
  assign n6729 = ( n6183 & n6727 ) | ( n6183 & ~n6728 ) | ( n6727 & ~n6728 ) ;
  assign n6726 = n6183 | n6185 ;
  assign n6730 = ( n6190 & ~n6726 ) | ( n6190 & n6729 ) | ( ~n6726 & n6729 ) ;
  assign n6731 = ( ~n6195 & n6729 ) | ( ~n6195 & n6730 ) | ( n6729 & n6730 ) ;
  assign n6733 = ( n6660 & ~n6665 ) | ( n6660 & n6670 ) | ( ~n6665 & n6670 ) ;
  assign n6734 = n6665 & ~n6670 ;
  assign n6735 = ( n6658 & n6733 ) | ( n6658 & ~n6734 ) | ( n6733 & ~n6734 ) ;
  assign n6732 = n6658 | n6660 ;
  assign n6736 = ( n6665 & ~n6732 ) | ( n6665 & n6735 ) | ( ~n6732 & n6735 ) ;
  assign n6737 = ( ~n6670 & n6735 ) | ( ~n6670 & n6736 ) | ( n6735 & n6736 ) ;
  assign n6738 = ( n6725 & n6731 ) | ( n6725 & n6737 ) | ( n6731 & n6737 ) ;
  assign n6739 = n6731 | n6737 ;
  assign n6740 = ( n6724 & n6738 ) | ( n6724 & n6739 ) | ( n6738 & n6739 ) ;
  assign n6741 = ( n6697 & n6700 ) | ( n6697 & n6740 ) | ( n6700 & n6740 ) ;
  assign n6742 = n6694 & n6741 ;
  assign n6743 = n6215 & n6690 ;
  assign n6744 = n6217 | n6692 ;
  assign n6745 = n6743 & ~n6744 ;
  assign n6754 = n5950 & n6208 ;
  assign n6755 = n6152 | n6207 ;
  assign n6756 = n6149 | n6207 ;
  assign n6757 = ( n6159 & n6755 ) | ( n6159 & n6756 ) | ( n6755 & n6756 ) ;
  assign n6758 = n6754 | n6757 ;
  assign n6759 = n6211 | n6758 ;
  assign n6760 = ( n6202 & n6211 ) | ( n6202 & n6759 ) | ( n6211 & n6759 ) ;
  assign n6761 = n6211 | n6759 ;
  assign n6762 = ( n6199 & n6760 ) | ( n6199 & n6761 ) | ( n6760 & n6761 ) ;
  assign n6746 = n6425 & n6683 ;
  assign n6747 = n6627 | n6682 ;
  assign n6748 = n6624 | n6682 ;
  assign n6749 = ( n6634 & n6747 ) | ( n6634 & n6748 ) | ( n6747 & n6748 ) ;
  assign n6750 = n6746 | n6749 ;
  assign n6751 = n6677 & n6750 ;
  assign n6752 = ( n6674 & n6750 ) | ( n6674 & n6751 ) | ( n6750 & n6751 ) ;
  assign n6753 = n6686 | n6752 ;
  assign n6763 = n6753 & n6762 ;
  assign n6764 = n6753 & ~n6763 ;
  assign n6765 = ( n6762 & ~n6763 ) | ( n6762 & n6764 ) | ( ~n6763 & n6764 ) ;
  assign n6766 = n6745 | n6765 ;
  assign n6767 = n6742 | n6766 ;
  assign n6768 = n6742 | n6745 ;
  assign n6769 = n6765 & n6768 ;
  assign n6770 = n6767 & ~n6769 ;
  assign n6771 = ( x118 & x119 ) | ( x118 & x120 ) | ( x119 & x120 ) ;
  assign n6772 = ( x115 & x116 ) | ( x115 & x117 ) | ( x116 & x117 ) ;
  assign n6773 = n6771 & ~n6772 ;
  assign n6774 = ~n6771 & n6772 ;
  assign n6775 = n6773 | n6774 ;
  assign n6776 = ~x115 & x116 ;
  assign n6777 = x115 & ~x116 ;
  assign n6778 = n6776 | n6777 ;
  assign n6779 = ~x117 & n6778 ;
  assign n6780 = x117 & ~n6778 ;
  assign n6781 = n6779 | n6780 ;
  assign n6782 = ~x118 & x119 ;
  assign n6783 = x118 & ~x119 ;
  assign n6784 = n6782 | n6783 ;
  assign n6785 = ~x120 & n6784 ;
  assign n6786 = x120 & ~n6784 ;
  assign n6787 = n6785 | n6786 ;
  assign n6788 = n6781 & n6787 ;
  assign n6789 = n6775 & ~n6788 ;
  assign n6790 = ~n6775 & n6788 ;
  assign n6791 = n6789 | n6790 ;
  assign n6792 = n6781 & ~n6787 ;
  assign n6793 = ~n6781 & n6787 ;
  assign n6794 = n6792 | n6793 ;
  assign n6795 = ( n6771 & n6772 ) | ( n6771 & n6788 ) | ( n6772 & n6788 ) ;
  assign n6796 = n6794 & n6795 ;
  assign n6797 = n6791 & ~n6796 ;
  assign n6798 = n6791 & n6795 ;
  assign n6799 = ~x121 & x122 ;
  assign n6800 = x121 & ~x122 ;
  assign n6801 = n6799 | n6800 ;
  assign n6802 = ~x123 & n6801 ;
  assign n6803 = x123 & ~n6801 ;
  assign n6804 = n6802 | n6803 ;
  assign n6805 = ~x124 & x125 ;
  assign n6806 = x124 & ~x125 ;
  assign n6807 = n6805 | n6806 ;
  assign n6808 = ~x126 & n6807 ;
  assign n6809 = x126 & ~n6807 ;
  assign n6810 = n6808 | n6809 ;
  assign n6811 = n6804 & ~n6810 ;
  assign n6812 = ~n6804 & n6810 ;
  assign n6813 = n6811 | n6812 ;
  assign n6814 = ( x124 & x125 ) | ( x124 & x126 ) | ( x125 & x126 ) ;
  assign n6815 = ( x121 & x122 ) | ( x121 & x123 ) | ( x122 & x123 ) ;
  assign n6816 = n6804 & n6810 ;
  assign n6817 = ( n6814 & n6815 ) | ( n6814 & n6816 ) | ( n6815 & n6816 ) ;
  assign n6818 = n6813 & n6817 ;
  assign n6819 = n6798 | n6818 ;
  assign n6820 = n6814 & ~n6815 ;
  assign n6821 = ~n6814 & n6815 ;
  assign n6822 = n6820 | n6821 ;
  assign n6823 = ~n6816 & n6822 ;
  assign n6824 = n6816 & ~n6822 ;
  assign n6825 = n6823 | n6824 ;
  assign n6826 = n6817 & n6825 ;
  assign n6827 = n6794 & n6813 ;
  assign n6828 = n6825 & n6827 ;
  assign n6829 = ~n6826 & n6828 ;
  assign n6830 = ~n6819 & n6829 ;
  assign n6831 = n6797 & n6830 ;
  assign n6832 = ~n6826 & n6827 ;
  assign n6833 = ~n6818 & n6825 ;
  assign n6834 = n6798 & ~n6833 ;
  assign n6835 = ( n6832 & n6833 ) | ( n6832 & ~n6834 ) | ( n6833 & ~n6834 ) ;
  assign n6836 = ( n6797 & n6831 ) | ( n6797 & ~n6835 ) | ( n6831 & ~n6835 ) ;
  assign n6837 = n6813 & ~n6817 ;
  assign n6838 = ( n6813 & ~n6825 ) | ( n6813 & n6837 ) | ( ~n6825 & n6837 ) ;
  assign n6839 = n6794 & ~n6795 ;
  assign n6840 = ( ~n6791 & n6794 ) | ( ~n6791 & n6839 ) | ( n6794 & n6839 ) ;
  assign n6841 = ~n6838 & n6840 ;
  assign n6842 = n6838 & ~n6840 ;
  assign n6843 = n6841 | n6842 ;
  assign n6844 = ( x112 & x113 ) | ( x112 & x114 ) | ( x113 & x114 ) ;
  assign n6845 = ( x109 & x110 ) | ( x109 & x111 ) | ( x110 & x111 ) ;
  assign n6846 = n6844 & ~n6845 ;
  assign n6847 = ~n6844 & n6845 ;
  assign n6848 = n6846 | n6847 ;
  assign n6849 = ~x109 & x110 ;
  assign n6850 = x109 & ~x110 ;
  assign n6851 = n6849 | n6850 ;
  assign n6852 = ~x111 & n6851 ;
  assign n6853 = x111 & ~n6851 ;
  assign n6854 = n6852 | n6853 ;
  assign n6855 = ~x112 & x113 ;
  assign n6856 = x112 & ~x113 ;
  assign n6857 = n6855 | n6856 ;
  assign n6858 = ~x114 & n6857 ;
  assign n6859 = x114 & ~n6857 ;
  assign n6860 = n6858 | n6859 ;
  assign n6861 = n6854 & n6860 ;
  assign n6862 = n6848 & ~n6861 ;
  assign n6863 = ~n6848 & n6861 ;
  assign n6864 = n6862 | n6863 ;
  assign n6865 = n6854 & ~n6860 ;
  assign n6866 = ~n6854 & n6860 ;
  assign n6867 = n6865 | n6866 ;
  assign n6868 = ( n6844 & n6845 ) | ( n6844 & n6861 ) | ( n6845 & n6861 ) ;
  assign n6869 = n6867 & ~n6868 ;
  assign n6870 = ( ~n6864 & n6867 ) | ( ~n6864 & n6869 ) | ( n6867 & n6869 ) ;
  assign n6871 = ~x103 & x104 ;
  assign n6872 = x103 & ~x104 ;
  assign n6873 = n6871 | n6872 ;
  assign n6874 = ~x105 & n6873 ;
  assign n6875 = x105 & ~n6873 ;
  assign n6876 = n6874 | n6875 ;
  assign n6877 = ~x106 & x107 ;
  assign n6878 = x106 & ~x107 ;
  assign n6879 = n6877 | n6878 ;
  assign n6880 = ~x108 & n6879 ;
  assign n6881 = x108 & ~n6879 ;
  assign n6882 = n6880 | n6881 ;
  assign n6883 = n6876 & ~n6882 ;
  assign n6884 = ~n6876 & n6882 ;
  assign n6885 = n6883 | n6884 ;
  assign n6886 = ( x106 & x107 ) | ( x106 & x108 ) | ( x107 & x108 ) ;
  assign n6887 = ( x103 & x104 ) | ( x103 & x105 ) | ( x104 & x105 ) ;
  assign n6888 = n6886 & ~n6887 ;
  assign n6889 = ~n6886 & n6887 ;
  assign n6890 = n6888 | n6889 ;
  assign n6891 = n6876 & n6882 ;
  assign n6892 = n6890 & ~n6891 ;
  assign n6893 = ~n6890 & n6891 ;
  assign n6894 = n6892 | n6893 ;
  assign n6895 = ( n6886 & n6887 ) | ( n6886 & n6891 ) | ( n6887 & n6891 ) ;
  assign n6896 = n6885 & ~n6895 ;
  assign n6897 = ( n6885 & ~n6894 ) | ( n6885 & n6896 ) | ( ~n6894 & n6896 ) ;
  assign n6898 = ~n6870 & n6897 ;
  assign n6899 = n6870 & ~n6897 ;
  assign n6900 = n6898 | n6899 ;
  assign n6901 = n6843 & n6900 ;
  assign n6902 = ( n6797 & ~n6798 ) | ( n6797 & n6833 ) | ( ~n6798 & n6833 ) ;
  assign n6903 = n6797 & n6833 ;
  assign n6904 = ( n6832 & n6902 ) | ( n6832 & n6903 ) | ( n6902 & n6903 ) ;
  assign n6905 = n6835 & ~n6904 ;
  assign n6906 = n6901 | n6905 ;
  assign n6907 = n6836 | n6906 ;
  assign n6908 = n6894 & n6895 ;
  assign n6909 = n6867 & n6868 ;
  assign n6910 = n6908 | n6909 ;
  assign n6911 = n6864 & n6868 ;
  assign n6912 = n6867 & n6885 ;
  assign n6913 = n6864 & n6912 ;
  assign n6914 = ~n6911 & n6913 ;
  assign n6915 = ~n6910 & n6914 ;
  assign n6916 = n6885 & n6895 ;
  assign n6917 = n6894 & ~n6916 ;
  assign n6918 = ~n6915 & n6917 ;
  assign n6919 = ~n6911 & n6912 ;
  assign n6920 = n6864 & ~n6909 ;
  assign n6921 = ( n6908 & n6917 ) | ( n6908 & n6920 ) | ( n6917 & n6920 ) ;
  assign n6922 = n6917 | n6920 ;
  assign n6923 = ( ~n6919 & n6921 ) | ( ~n6919 & n6922 ) | ( n6921 & n6922 ) ;
  assign n6924 = n6908 | n6920 ;
  assign n6925 = n6919 & ~n6924 ;
  assign n6926 = ( ~n6920 & n6923 ) | ( ~n6920 & n6925 ) | ( n6923 & n6925 ) ;
  assign n6927 = ( ~n6918 & n6923 ) | ( ~n6918 & n6926 ) | ( n6923 & n6926 ) ;
  assign n6928 = n6907 & n6927 ;
  assign n6929 = n6901 & n6905 ;
  assign n6930 = ( n6836 & n6901 ) | ( n6836 & n6929 ) | ( n6901 & n6929 ) ;
  assign n6931 = n6928 | n6930 ;
  assign n6932 = n6908 & ~n6920 ;
  assign n6933 = ( n6919 & n6920 ) | ( n6919 & ~n6932 ) | ( n6920 & ~n6932 ) ;
  assign n6934 = n6917 & n6933 ;
  assign n6935 = ~n6885 & n6895 ;
  assign n6936 = ( ~n6894 & n6895 ) | ( ~n6894 & n6935 ) | ( n6895 & n6935 ) ;
  assign n6937 = ~n6867 & n6868 ;
  assign n6938 = ( ~n6864 & n6868 ) | ( ~n6864 & n6937 ) | ( n6868 & n6937 ) ;
  assign n6939 = ~n6936 & n6938 ;
  assign n6940 = n6936 & ~n6938 ;
  assign n6941 = n6939 | n6940 ;
  assign n6942 = n6915 | n6941 ;
  assign n6943 = n6934 | n6942 ;
  assign n6944 = n6915 & n6941 ;
  assign n6945 = ( n6934 & n6941 ) | ( n6934 & n6944 ) | ( n6941 & n6944 ) ;
  assign n6946 = n6943 & ~n6945 ;
  assign n6947 = n6797 & n6835 ;
  assign n6948 = ~n6794 & n6795 ;
  assign n6949 = ( ~n6791 & n6795 ) | ( ~n6791 & n6948 ) | ( n6795 & n6948 ) ;
  assign n6950 = ~n6813 & n6817 ;
  assign n6951 = ( n6817 & ~n6825 ) | ( n6817 & n6950 ) | ( ~n6825 & n6950 ) ;
  assign n6952 = ~n6949 & n6951 ;
  assign n6953 = n6949 & ~n6951 ;
  assign n6954 = n6952 | n6953 ;
  assign n6955 = n6830 | n6954 ;
  assign n6956 = n6947 | n6955 ;
  assign n6957 = n6830 & n6954 ;
  assign n6958 = ( n6947 & n6954 ) | ( n6947 & n6957 ) | ( n6954 & n6957 ) ;
  assign n6959 = n6956 & ~n6958 ;
  assign n6960 = n6946 | n6959 ;
  assign n6961 = n6931 & n6960 ;
  assign n6962 = n6943 & n6956 ;
  assign n6963 = n6945 | n6958 ;
  assign n6964 = n6962 & ~n6963 ;
  assign n6965 = ( n6830 & n6949 ) | ( n6830 & n6951 ) | ( n6949 & n6951 ) ;
  assign n6966 = n6949 | n6951 ;
  assign n6967 = ( n6947 & n6965 ) | ( n6947 & n6966 ) | ( n6965 & n6966 ) ;
  assign n6968 = ( n6915 & n6936 ) | ( n6915 & n6938 ) | ( n6936 & n6938 ) ;
  assign n6969 = n6936 | n6938 ;
  assign n6970 = ( n6934 & n6968 ) | ( n6934 & n6969 ) | ( n6968 & n6969 ) ;
  assign n6971 = ~n6967 & n6970 ;
  assign n6972 = n6967 & ~n6970 ;
  assign n6973 = n6971 | n6972 ;
  assign n6974 = n6964 | n6973 ;
  assign n6975 = n6961 | n6974 ;
  assign n6976 = n6960 | n6964 ;
  assign n6977 = ( n6931 & n6964 ) | ( n6931 & n6976 ) | ( n6964 & n6976 ) ;
  assign n6978 = n6973 & n6977 ;
  assign n6979 = n6975 & ~n6978 ;
  assign n6980 = ( x94 & x95 ) | ( x94 & x96 ) | ( x95 & x96 ) ;
  assign n6981 = ( x91 & x92 ) | ( x91 & x93 ) | ( x92 & x93 ) ;
  assign n6982 = n6980 & ~n6981 ;
  assign n6983 = ~n6980 & n6981 ;
  assign n6984 = n6982 | n6983 ;
  assign n6985 = ~x91 & x92 ;
  assign n6986 = x91 & ~x92 ;
  assign n6987 = n6985 | n6986 ;
  assign n6988 = ~x93 & n6987 ;
  assign n6989 = x93 & ~n6987 ;
  assign n6990 = n6988 | n6989 ;
  assign n6991 = ~x94 & x95 ;
  assign n6992 = x94 & ~x95 ;
  assign n6993 = n6991 | n6992 ;
  assign n6994 = ~x96 & n6993 ;
  assign n6995 = x96 & ~n6993 ;
  assign n6996 = n6994 | n6995 ;
  assign n6997 = n6990 & n6996 ;
  assign n6998 = n6984 & ~n6997 ;
  assign n6999 = ~n6984 & n6997 ;
  assign n7000 = n6998 | n6999 ;
  assign n7001 = n6990 & ~n6996 ;
  assign n7002 = ~n6990 & n6996 ;
  assign n7003 = n7001 | n7002 ;
  assign n7004 = ( n6980 & n6981 ) | ( n6980 & n6997 ) | ( n6981 & n6997 ) ;
  assign n7005 = n7003 & n7004 ;
  assign n7006 = n7000 & ~n7005 ;
  assign n7007 = n7000 & n7004 ;
  assign n7008 = ~x97 & x98 ;
  assign n7009 = x97 & ~x98 ;
  assign n7010 = n7008 | n7009 ;
  assign n7011 = ~x99 & n7010 ;
  assign n7012 = x99 & ~n7010 ;
  assign n7013 = n7011 | n7012 ;
  assign n7014 = ~x100 & x101 ;
  assign n7015 = x100 & ~x101 ;
  assign n7016 = n7014 | n7015 ;
  assign n7017 = ~x102 & n7016 ;
  assign n7018 = x102 & ~n7016 ;
  assign n7019 = n7017 | n7018 ;
  assign n7020 = n7013 & ~n7019 ;
  assign n7021 = ~n7013 & n7019 ;
  assign n7022 = n7020 | n7021 ;
  assign n7023 = ( x100 & x101 ) | ( x100 & x102 ) | ( x101 & x102 ) ;
  assign n7024 = ( x97 & x98 ) | ( x97 & x99 ) | ( x98 & x99 ) ;
  assign n7025 = n7013 & n7019 ;
  assign n7026 = ( n7023 & n7024 ) | ( n7023 & n7025 ) | ( n7024 & n7025 ) ;
  assign n7027 = n7022 & n7026 ;
  assign n7028 = n7007 | n7027 ;
  assign n7029 = n7023 & ~n7024 ;
  assign n7030 = ~n7023 & n7024 ;
  assign n7031 = n7029 | n7030 ;
  assign n7032 = ~n7025 & n7031 ;
  assign n7033 = n7025 & ~n7031 ;
  assign n7034 = n7032 | n7033 ;
  assign n7035 = n7026 & n7034 ;
  assign n7036 = n7003 & n7022 ;
  assign n7037 = n7034 & n7036 ;
  assign n7038 = ~n7035 & n7037 ;
  assign n7039 = ~n7028 & n7038 ;
  assign n7040 = n7006 & n7039 ;
  assign n7041 = ~n7035 & n7036 ;
  assign n7042 = ~n7027 & n7034 ;
  assign n7043 = n7007 & ~n7042 ;
  assign n7044 = ( n7041 & n7042 ) | ( n7041 & ~n7043 ) | ( n7042 & ~n7043 ) ;
  assign n7045 = ( n7006 & n7040 ) | ( n7006 & ~n7044 ) | ( n7040 & ~n7044 ) ;
  assign n7046 = n7022 & ~n7026 ;
  assign n7047 = ( n7022 & ~n7034 ) | ( n7022 & n7046 ) | ( ~n7034 & n7046 ) ;
  assign n7048 = n7003 & ~n7004 ;
  assign n7049 = ( ~n7000 & n7003 ) | ( ~n7000 & n7048 ) | ( n7003 & n7048 ) ;
  assign n7050 = ~n7047 & n7049 ;
  assign n7051 = n7047 & ~n7049 ;
  assign n7052 = n7050 | n7051 ;
  assign n7053 = ( x88 & x89 ) | ( x88 & x90 ) | ( x89 & x90 ) ;
  assign n7054 = ( x85 & x86 ) | ( x85 & x87 ) | ( x86 & x87 ) ;
  assign n7055 = n7053 & ~n7054 ;
  assign n7056 = ~n7053 & n7054 ;
  assign n7057 = n7055 | n7056 ;
  assign n7058 = ~x85 & x86 ;
  assign n7059 = x85 & ~x86 ;
  assign n7060 = n7058 | n7059 ;
  assign n7061 = ~x87 & n7060 ;
  assign n7062 = x87 & ~n7060 ;
  assign n7063 = n7061 | n7062 ;
  assign n7064 = ~x88 & x89 ;
  assign n7065 = x88 & ~x89 ;
  assign n7066 = n7064 | n7065 ;
  assign n7067 = ~x90 & n7066 ;
  assign n7068 = x90 & ~n7066 ;
  assign n7069 = n7067 | n7068 ;
  assign n7070 = n7063 & n7069 ;
  assign n7071 = n7057 & ~n7070 ;
  assign n7072 = ~n7057 & n7070 ;
  assign n7073 = n7071 | n7072 ;
  assign n7074 = n7063 & ~n7069 ;
  assign n7075 = ~n7063 & n7069 ;
  assign n7076 = n7074 | n7075 ;
  assign n7077 = ( n7053 & n7054 ) | ( n7053 & n7070 ) | ( n7054 & n7070 ) ;
  assign n7078 = n7076 & ~n7077 ;
  assign n7079 = ( ~n7073 & n7076 ) | ( ~n7073 & n7078 ) | ( n7076 & n7078 ) ;
  assign n7080 = ~x79 & x80 ;
  assign n7081 = x79 & ~x80 ;
  assign n7082 = n7080 | n7081 ;
  assign n7083 = ~x81 & n7082 ;
  assign n7084 = x81 & ~n7082 ;
  assign n7085 = n7083 | n7084 ;
  assign n7086 = ~x82 & x83 ;
  assign n7087 = x82 & ~x83 ;
  assign n7088 = n7086 | n7087 ;
  assign n7089 = ~x84 & n7088 ;
  assign n7090 = x84 & ~n7088 ;
  assign n7091 = n7089 | n7090 ;
  assign n7092 = n7085 & ~n7091 ;
  assign n7093 = ~n7085 & n7091 ;
  assign n7094 = n7092 | n7093 ;
  assign n7095 = ( x82 & x83 ) | ( x82 & x84 ) | ( x83 & x84 ) ;
  assign n7096 = ( x79 & x80 ) | ( x79 & x81 ) | ( x80 & x81 ) ;
  assign n7097 = n7095 & ~n7096 ;
  assign n7098 = ~n7095 & n7096 ;
  assign n7099 = n7097 | n7098 ;
  assign n7100 = n7085 & n7091 ;
  assign n7101 = n7099 & ~n7100 ;
  assign n7102 = ~n7099 & n7100 ;
  assign n7103 = n7101 | n7102 ;
  assign n7104 = ( n7095 & n7096 ) | ( n7095 & n7100 ) | ( n7096 & n7100 ) ;
  assign n7105 = n7094 & ~n7104 ;
  assign n7106 = ( n7094 & ~n7103 ) | ( n7094 & n7105 ) | ( ~n7103 & n7105 ) ;
  assign n7107 = ~n7079 & n7106 ;
  assign n7108 = n7079 & ~n7106 ;
  assign n7109 = n7107 | n7108 ;
  assign n7110 = n7052 & n7109 ;
  assign n7111 = ( n7006 & ~n7007 ) | ( n7006 & n7042 ) | ( ~n7007 & n7042 ) ;
  assign n7112 = n7006 & n7042 ;
  assign n7113 = ( n7041 & n7111 ) | ( n7041 & n7112 ) | ( n7111 & n7112 ) ;
  assign n7114 = n7044 & ~n7113 ;
  assign n7115 = n7110 | n7114 ;
  assign n7116 = n7045 | n7115 ;
  assign n7117 = n7103 & n7104 ;
  assign n7118 = n7076 & n7077 ;
  assign n7119 = n7117 | n7118 ;
  assign n7120 = n7073 & n7077 ;
  assign n7121 = n7076 & n7094 ;
  assign n7122 = n7073 & n7121 ;
  assign n7123 = ~n7120 & n7122 ;
  assign n7124 = ~n7119 & n7123 ;
  assign n7125 = n7094 & n7104 ;
  assign n7126 = n7103 & ~n7125 ;
  assign n7127 = ~n7124 & n7126 ;
  assign n7128 = ~n7120 & n7121 ;
  assign n7129 = n7073 & ~n7118 ;
  assign n7130 = ( n7117 & n7126 ) | ( n7117 & n7129 ) | ( n7126 & n7129 ) ;
  assign n7131 = n7126 | n7129 ;
  assign n7132 = ( ~n7128 & n7130 ) | ( ~n7128 & n7131 ) | ( n7130 & n7131 ) ;
  assign n7133 = n7117 | n7129 ;
  assign n7134 = n7128 & ~n7133 ;
  assign n7135 = ( ~n7129 & n7132 ) | ( ~n7129 & n7134 ) | ( n7132 & n7134 ) ;
  assign n7136 = ( ~n7127 & n7132 ) | ( ~n7127 & n7135 ) | ( n7132 & n7135 ) ;
  assign n7137 = n7116 & n7136 ;
  assign n7138 = n7110 & n7114 ;
  assign n7139 = ( n7045 & n7110 ) | ( n7045 & n7138 ) | ( n7110 & n7138 ) ;
  assign n7140 = n7137 | n7139 ;
  assign n7141 = n7117 & ~n7129 ;
  assign n7142 = ( n7128 & n7129 ) | ( n7128 & ~n7141 ) | ( n7129 & ~n7141 ) ;
  assign n7143 = n7126 & n7142 ;
  assign n7144 = ~n7094 & n7104 ;
  assign n7145 = ( ~n7103 & n7104 ) | ( ~n7103 & n7144 ) | ( n7104 & n7144 ) ;
  assign n7146 = ~n7076 & n7077 ;
  assign n7147 = ( ~n7073 & n7077 ) | ( ~n7073 & n7146 ) | ( n7077 & n7146 ) ;
  assign n7148 = ~n7145 & n7147 ;
  assign n7149 = n7145 & ~n7147 ;
  assign n7150 = n7148 | n7149 ;
  assign n7151 = n7124 | n7150 ;
  assign n7152 = n7143 | n7151 ;
  assign n7153 = n7124 & n7150 ;
  assign n7154 = ( n7143 & n7150 ) | ( n7143 & n7153 ) | ( n7150 & n7153 ) ;
  assign n7155 = n7152 & ~n7154 ;
  assign n7156 = n7006 & n7044 ;
  assign n7157 = ~n7003 & n7004 ;
  assign n7158 = ( ~n7000 & n7004 ) | ( ~n7000 & n7157 ) | ( n7004 & n7157 ) ;
  assign n7159 = ~n7022 & n7026 ;
  assign n7160 = ( n7026 & ~n7034 ) | ( n7026 & n7159 ) | ( ~n7034 & n7159 ) ;
  assign n7161 = ~n7158 & n7160 ;
  assign n7162 = n7158 & ~n7160 ;
  assign n7163 = n7161 | n7162 ;
  assign n7164 = n7039 | n7163 ;
  assign n7165 = n7156 | n7164 ;
  assign n7166 = n7039 & n7163 ;
  assign n7167 = ( n7156 & n7163 ) | ( n7156 & n7166 ) | ( n7163 & n7166 ) ;
  assign n7168 = n7165 & ~n7167 ;
  assign n7169 = n7155 | n7168 ;
  assign n7170 = n7140 & n7169 ;
  assign n7171 = n7152 & n7165 ;
  assign n7172 = n7154 | n7167 ;
  assign n7173 = n7171 & ~n7172 ;
  assign n7174 = ( n7039 & n7158 ) | ( n7039 & n7160 ) | ( n7158 & n7160 ) ;
  assign n7175 = n7158 | n7160 ;
  assign n7176 = ( n7156 & n7174 ) | ( n7156 & n7175 ) | ( n7174 & n7175 ) ;
  assign n7177 = ( n7124 & n7145 ) | ( n7124 & n7147 ) | ( n7145 & n7147 ) ;
  assign n7178 = n7145 | n7147 ;
  assign n7179 = ( n7143 & n7177 ) | ( n7143 & n7178 ) | ( n7177 & n7178 ) ;
  assign n7180 = ~n7176 & n7179 ;
  assign n7181 = n7176 & ~n7179 ;
  assign n7182 = n7180 | n7181 ;
  assign n7183 = n7173 | n7182 ;
  assign n7184 = n7170 | n7183 ;
  assign n7185 = n7169 | n7173 ;
  assign n7186 = ( n7140 & n7173 ) | ( n7140 & n7185 ) | ( n7173 & n7185 ) ;
  assign n7187 = n7182 & n7186 ;
  assign n7188 = n7184 & ~n7187 ;
  assign n7189 = n6979 | n7188 ;
  assign n7190 = n6907 & ~n6930 ;
  assign n7191 = n6927 & ~n7190 ;
  assign n7192 = n6843 & ~n6900 ;
  assign n7193 = ~n6843 & n6900 ;
  assign n7194 = n7192 | n7193 ;
  assign n7195 = n7052 & ~n7109 ;
  assign n7196 = ~n7052 & n7109 ;
  assign n7197 = n7195 | n7196 ;
  assign n7198 = n7194 & n7197 ;
  assign n7199 = ~n6901 & n6907 ;
  assign n7200 = n6907 & ~n6927 ;
  assign n7201 = n6836 | n6905 ;
  assign n7202 = n6927 | n7201 ;
  assign n7203 = ( n7199 & n7200 ) | ( n7199 & ~n7202 ) | ( n7200 & ~n7202 ) ;
  assign n7204 = n7198 | n7203 ;
  assign n7205 = n7191 | n7204 ;
  assign n7206 = n7045 | n7114 ;
  assign n7207 = ( n7110 & n7136 ) | ( n7110 & ~n7206 ) | ( n7136 & ~n7206 ) ;
  assign n7208 = ( ~n7136 & n7206 ) | ( ~n7136 & n7207 ) | ( n7206 & n7207 ) ;
  assign n7209 = ( ~n7110 & n7207 ) | ( ~n7110 & n7208 ) | ( n7207 & n7208 ) ;
  assign n7210 = n7205 & n7209 ;
  assign n7211 = n7191 | n7203 ;
  assign n7212 = n7198 & n7211 ;
  assign n7213 = ( n7139 & ~n7155 ) | ( n7139 & n7168 ) | ( ~n7155 & n7168 ) ;
  assign n7214 = n7155 & ~n7168 ;
  assign n7215 = ( n7137 & n7213 ) | ( n7137 & ~n7214 ) | ( n7213 & ~n7214 ) ;
  assign n7216 = ( ~n7140 & n7155 ) | ( ~n7140 & n7215 ) | ( n7155 & n7215 ) ;
  assign n7217 = ( ~n7168 & n7215 ) | ( ~n7168 & n7216 ) | ( n7215 & n7216 ) ;
  assign n7218 = ( n6930 & ~n6946 ) | ( n6930 & n6959 ) | ( ~n6946 & n6959 ) ;
  assign n7219 = n6946 & ~n6959 ;
  assign n7220 = ( n6928 & n7218 ) | ( n6928 & ~n7219 ) | ( n7218 & ~n7219 ) ;
  assign n7221 = ( ~n6931 & n6946 ) | ( ~n6931 & n7220 ) | ( n6946 & n7220 ) ;
  assign n7222 = ( ~n6959 & n7220 ) | ( ~n6959 & n7221 ) | ( n7220 & n7221 ) ;
  assign n7223 = ( n7212 & n7217 ) | ( n7212 & n7222 ) | ( n7217 & n7222 ) ;
  assign n7224 = n7217 | n7222 ;
  assign n7225 = ( n7210 & n7223 ) | ( n7210 & n7224 ) | ( n7223 & n7224 ) ;
  assign n7226 = n7189 & n7225 ;
  assign n7227 = n6975 & n7184 ;
  assign n7228 = n6978 | n7187 ;
  assign n7229 = n7227 & ~n7228 ;
  assign n7230 = n7176 & n7179 ;
  assign n7231 = n7176 | n7179 ;
  assign n7232 = n7230 | n7231 ;
  assign n7233 = ( n7186 & n7230 ) | ( n7186 & n7232 ) | ( n7230 & n7232 ) ;
  assign n7234 = n6967 & n6970 ;
  assign n7235 = n6967 | n6970 ;
  assign n7236 = n7234 | n7235 ;
  assign n7237 = ( n6977 & n7234 ) | ( n6977 & n7236 ) | ( n7234 & n7236 ) ;
  assign n7238 = n7233 & n7237 ;
  assign n7239 = n7237 & ~n7238 ;
  assign n7240 = ( n7233 & ~n7238 ) | ( n7233 & n7239 ) | ( ~n7238 & n7239 ) ;
  assign n7241 = n7229 | n7240 ;
  assign n7242 = n7226 | n7241 ;
  assign n7243 = n7226 | n7229 ;
  assign n7244 = n7240 & n7243 ;
  assign n7245 = n7242 & ~n7244 ;
  assign n7246 = ( x166 & x167 ) | ( x166 & x168 ) | ( x167 & x168 ) ;
  assign n7247 = ( x163 & x164 ) | ( x163 & x165 ) | ( x164 & x165 ) ;
  assign n7248 = n7246 & ~n7247 ;
  assign n7249 = ~n7246 & n7247 ;
  assign n7250 = n7248 | n7249 ;
  assign n7251 = ~x163 & x164 ;
  assign n7252 = x163 & ~x164 ;
  assign n7253 = n7251 | n7252 ;
  assign n7254 = ~x165 & n7253 ;
  assign n7255 = x165 & ~n7253 ;
  assign n7256 = n7254 | n7255 ;
  assign n7257 = ~x166 & x167 ;
  assign n7258 = x166 & ~x167 ;
  assign n7259 = n7257 | n7258 ;
  assign n7260 = ~x168 & n7259 ;
  assign n7261 = x168 & ~n7259 ;
  assign n7262 = n7260 | n7261 ;
  assign n7263 = n7256 & n7262 ;
  assign n7264 = n7250 & ~n7263 ;
  assign n7265 = ~n7250 & n7263 ;
  assign n7266 = n7264 | n7265 ;
  assign n7267 = n7256 & ~n7262 ;
  assign n7268 = ~n7256 & n7262 ;
  assign n7269 = n7267 | n7268 ;
  assign n7270 = ( n7246 & n7247 ) | ( n7246 & n7263 ) | ( n7247 & n7263 ) ;
  assign n7271 = n7269 & n7270 ;
  assign n7272 = n7266 & ~n7271 ;
  assign n7273 = n7266 & n7270 ;
  assign n7274 = ~x169 & x170 ;
  assign n7275 = x169 & ~x170 ;
  assign n7276 = n7274 | n7275 ;
  assign n7277 = ~x171 & n7276 ;
  assign n7278 = x171 & ~n7276 ;
  assign n7279 = n7277 | n7278 ;
  assign n7280 = ~x172 & x173 ;
  assign n7281 = x172 & ~x173 ;
  assign n7282 = n7280 | n7281 ;
  assign n7283 = ~x174 & n7282 ;
  assign n7284 = x174 & ~n7282 ;
  assign n7285 = n7283 | n7284 ;
  assign n7286 = n7279 & ~n7285 ;
  assign n7287 = ~n7279 & n7285 ;
  assign n7288 = n7286 | n7287 ;
  assign n7289 = ( x172 & x173 ) | ( x172 & x174 ) | ( x173 & x174 ) ;
  assign n7290 = ( x169 & x170 ) | ( x169 & x171 ) | ( x170 & x171 ) ;
  assign n7291 = n7279 & n7285 ;
  assign n7292 = ( n7289 & n7290 ) | ( n7289 & n7291 ) | ( n7290 & n7291 ) ;
  assign n7293 = n7288 & n7292 ;
  assign n7294 = n7273 | n7293 ;
  assign n7295 = n7289 & ~n7290 ;
  assign n7296 = ~n7289 & n7290 ;
  assign n7297 = n7295 | n7296 ;
  assign n7298 = ~n7291 & n7297 ;
  assign n7299 = n7291 & ~n7297 ;
  assign n7300 = n7298 | n7299 ;
  assign n7301 = n7292 & n7300 ;
  assign n7302 = n7269 & n7288 ;
  assign n7303 = n7300 & n7302 ;
  assign n7304 = ~n7301 & n7303 ;
  assign n7305 = ~n7294 & n7304 ;
  assign n7306 = n7272 & n7305 ;
  assign n7307 = ~n7301 & n7302 ;
  assign n7308 = ~n7293 & n7300 ;
  assign n7309 = n7273 & ~n7308 ;
  assign n7310 = ( n7307 & n7308 ) | ( n7307 & ~n7309 ) | ( n7308 & ~n7309 ) ;
  assign n7311 = ( n7272 & n7306 ) | ( n7272 & ~n7310 ) | ( n7306 & ~n7310 ) ;
  assign n7312 = n7288 & ~n7292 ;
  assign n7313 = ( n7288 & ~n7300 ) | ( n7288 & n7312 ) | ( ~n7300 & n7312 ) ;
  assign n7314 = n7269 & ~n7270 ;
  assign n7315 = ( ~n7266 & n7269 ) | ( ~n7266 & n7314 ) | ( n7269 & n7314 ) ;
  assign n7316 = ~n7313 & n7315 ;
  assign n7317 = n7313 & ~n7315 ;
  assign n7318 = n7316 | n7317 ;
  assign n7319 = ( x160 & x161 ) | ( x160 & x162 ) | ( x161 & x162 ) ;
  assign n7320 = ( x157 & x158 ) | ( x157 & x159 ) | ( x158 & x159 ) ;
  assign n7321 = n7319 & ~n7320 ;
  assign n7322 = ~n7319 & n7320 ;
  assign n7323 = n7321 | n7322 ;
  assign n7324 = ~x157 & x158 ;
  assign n7325 = x157 & ~x158 ;
  assign n7326 = n7324 | n7325 ;
  assign n7327 = ~x159 & n7326 ;
  assign n7328 = x159 & ~n7326 ;
  assign n7329 = n7327 | n7328 ;
  assign n7330 = ~x160 & x161 ;
  assign n7331 = x160 & ~x161 ;
  assign n7332 = n7330 | n7331 ;
  assign n7333 = ~x162 & n7332 ;
  assign n7334 = x162 & ~n7332 ;
  assign n7335 = n7333 | n7334 ;
  assign n7336 = n7329 & n7335 ;
  assign n7337 = n7323 & ~n7336 ;
  assign n7338 = ~n7323 & n7336 ;
  assign n7339 = n7337 | n7338 ;
  assign n7340 = n7329 & ~n7335 ;
  assign n7341 = ~n7329 & n7335 ;
  assign n7342 = n7340 | n7341 ;
  assign n7343 = ( n7319 & n7320 ) | ( n7319 & n7336 ) | ( n7320 & n7336 ) ;
  assign n7344 = n7342 & ~n7343 ;
  assign n7345 = ( ~n7339 & n7342 ) | ( ~n7339 & n7344 ) | ( n7342 & n7344 ) ;
  assign n7346 = ~x151 & x152 ;
  assign n7347 = x151 & ~x152 ;
  assign n7348 = n7346 | n7347 ;
  assign n7349 = ~x153 & n7348 ;
  assign n7350 = x153 & ~n7348 ;
  assign n7351 = n7349 | n7350 ;
  assign n7352 = ~x154 & x155 ;
  assign n7353 = x154 & ~x155 ;
  assign n7354 = n7352 | n7353 ;
  assign n7355 = ~x156 & n7354 ;
  assign n7356 = x156 & ~n7354 ;
  assign n7357 = n7355 | n7356 ;
  assign n7358 = n7351 & ~n7357 ;
  assign n7359 = ~n7351 & n7357 ;
  assign n7360 = n7358 | n7359 ;
  assign n7361 = ( x154 & x155 ) | ( x154 & x156 ) | ( x155 & x156 ) ;
  assign n7362 = ( x151 & x152 ) | ( x151 & x153 ) | ( x152 & x153 ) ;
  assign n7363 = n7361 & ~n7362 ;
  assign n7364 = ~n7361 & n7362 ;
  assign n7365 = n7363 | n7364 ;
  assign n7366 = n7351 & n7357 ;
  assign n7367 = n7365 & ~n7366 ;
  assign n7368 = ~n7365 & n7366 ;
  assign n7369 = n7367 | n7368 ;
  assign n7370 = ( n7361 & n7362 ) | ( n7361 & n7366 ) | ( n7362 & n7366 ) ;
  assign n7371 = n7360 & ~n7370 ;
  assign n7372 = ( n7360 & ~n7369 ) | ( n7360 & n7371 ) | ( ~n7369 & n7371 ) ;
  assign n7373 = ~n7345 & n7372 ;
  assign n7374 = n7345 & ~n7372 ;
  assign n7375 = n7373 | n7374 ;
  assign n7376 = n7318 & n7375 ;
  assign n7377 = ( n7272 & ~n7273 ) | ( n7272 & n7308 ) | ( ~n7273 & n7308 ) ;
  assign n7378 = n7272 & n7308 ;
  assign n7379 = ( n7307 & n7377 ) | ( n7307 & n7378 ) | ( n7377 & n7378 ) ;
  assign n7380 = n7310 & ~n7379 ;
  assign n7381 = n7376 | n7380 ;
  assign n7382 = n7311 | n7381 ;
  assign n7383 = n7369 & n7370 ;
  assign n7384 = n7342 & n7343 ;
  assign n7385 = n7383 | n7384 ;
  assign n7386 = n7339 & n7343 ;
  assign n7387 = n7342 & n7360 ;
  assign n7388 = n7339 & n7387 ;
  assign n7389 = ~n7386 & n7388 ;
  assign n7390 = ~n7385 & n7389 ;
  assign n7391 = n7360 & n7370 ;
  assign n7392 = n7369 & ~n7391 ;
  assign n7393 = ~n7390 & n7392 ;
  assign n7394 = ~n7386 & n7387 ;
  assign n7395 = n7339 & ~n7384 ;
  assign n7396 = ( n7383 & n7392 ) | ( n7383 & n7395 ) | ( n7392 & n7395 ) ;
  assign n7397 = n7392 | n7395 ;
  assign n7398 = ( ~n7394 & n7396 ) | ( ~n7394 & n7397 ) | ( n7396 & n7397 ) ;
  assign n7399 = n7383 | n7395 ;
  assign n7400 = n7394 & ~n7399 ;
  assign n7401 = ( ~n7395 & n7398 ) | ( ~n7395 & n7400 ) | ( n7398 & n7400 ) ;
  assign n7402 = ( ~n7393 & n7398 ) | ( ~n7393 & n7401 ) | ( n7398 & n7401 ) ;
  assign n7403 = n7382 & n7402 ;
  assign n7404 = n7376 & n7380 ;
  assign n7405 = ( n7311 & n7376 ) | ( n7311 & n7404 ) | ( n7376 & n7404 ) ;
  assign n7406 = n7403 | n7405 ;
  assign n7407 = n7383 & ~n7395 ;
  assign n7408 = ( n7394 & n7395 ) | ( n7394 & ~n7407 ) | ( n7395 & ~n7407 ) ;
  assign n7409 = n7392 & n7408 ;
  assign n7410 = ~n7360 & n7370 ;
  assign n7411 = ( ~n7369 & n7370 ) | ( ~n7369 & n7410 ) | ( n7370 & n7410 ) ;
  assign n7412 = ~n7342 & n7343 ;
  assign n7413 = ( ~n7339 & n7343 ) | ( ~n7339 & n7412 ) | ( n7343 & n7412 ) ;
  assign n7414 = ~n7411 & n7413 ;
  assign n7415 = n7411 & ~n7413 ;
  assign n7416 = n7414 | n7415 ;
  assign n7417 = n7390 | n7416 ;
  assign n7418 = n7409 | n7417 ;
  assign n7419 = n7390 & n7416 ;
  assign n7420 = ( n7409 & n7416 ) | ( n7409 & n7419 ) | ( n7416 & n7419 ) ;
  assign n7421 = n7418 & ~n7420 ;
  assign n7422 = n7272 & n7310 ;
  assign n7423 = ~n7269 & n7270 ;
  assign n7424 = ( ~n7266 & n7270 ) | ( ~n7266 & n7423 ) | ( n7270 & n7423 ) ;
  assign n7425 = ~n7288 & n7292 ;
  assign n7426 = ( n7292 & ~n7300 ) | ( n7292 & n7425 ) | ( ~n7300 & n7425 ) ;
  assign n7427 = ~n7424 & n7426 ;
  assign n7428 = n7424 & ~n7426 ;
  assign n7429 = n7427 | n7428 ;
  assign n7430 = n7305 | n7429 ;
  assign n7431 = n7422 | n7430 ;
  assign n7432 = n7305 & n7429 ;
  assign n7433 = ( n7422 & n7429 ) | ( n7422 & n7432 ) | ( n7429 & n7432 ) ;
  assign n7434 = n7431 & ~n7433 ;
  assign n7435 = n7421 | n7434 ;
  assign n7436 = n7406 & n7435 ;
  assign n7437 = n7418 & n7431 ;
  assign n7438 = n7420 | n7433 ;
  assign n7439 = n7437 & ~n7438 ;
  assign n7440 = ( n7305 & n7424 ) | ( n7305 & n7426 ) | ( n7424 & n7426 ) ;
  assign n7441 = n7424 | n7426 ;
  assign n7442 = ( n7422 & n7440 ) | ( n7422 & n7441 ) | ( n7440 & n7441 ) ;
  assign n7443 = ( n7390 & n7411 ) | ( n7390 & n7413 ) | ( n7411 & n7413 ) ;
  assign n7444 = n7411 | n7413 ;
  assign n7445 = ( n7409 & n7443 ) | ( n7409 & n7444 ) | ( n7443 & n7444 ) ;
  assign n7446 = ~n7442 & n7445 ;
  assign n7447 = n7442 & ~n7445 ;
  assign n7448 = n7446 | n7447 ;
  assign n7449 = n7439 | n7448 ;
  assign n7450 = n7436 | n7449 ;
  assign n7451 = n7435 | n7439 ;
  assign n7452 = ( n7406 & n7439 ) | ( n7406 & n7451 ) | ( n7439 & n7451 ) ;
  assign n7453 = n7448 & n7452 ;
  assign n7454 = n7450 & ~n7453 ;
  assign n7455 = ( x142 & x143 ) | ( x142 & x144 ) | ( x143 & x144 ) ;
  assign n7456 = ( x139 & x140 ) | ( x139 & x141 ) | ( x140 & x141 ) ;
  assign n7457 = n7455 & ~n7456 ;
  assign n7458 = ~n7455 & n7456 ;
  assign n7459 = n7457 | n7458 ;
  assign n7460 = ~x139 & x140 ;
  assign n7461 = x139 & ~x140 ;
  assign n7462 = n7460 | n7461 ;
  assign n7463 = ~x141 & n7462 ;
  assign n7464 = x141 & ~n7462 ;
  assign n7465 = n7463 | n7464 ;
  assign n7466 = ~x142 & x143 ;
  assign n7467 = x142 & ~x143 ;
  assign n7468 = n7466 | n7467 ;
  assign n7469 = ~x144 & n7468 ;
  assign n7470 = x144 & ~n7468 ;
  assign n7471 = n7469 | n7470 ;
  assign n7472 = n7465 & n7471 ;
  assign n7473 = n7459 & ~n7472 ;
  assign n7474 = ~n7459 & n7472 ;
  assign n7475 = n7473 | n7474 ;
  assign n7476 = n7465 & ~n7471 ;
  assign n7477 = ~n7465 & n7471 ;
  assign n7478 = n7476 | n7477 ;
  assign n7479 = ( n7455 & n7456 ) | ( n7455 & n7472 ) | ( n7456 & n7472 ) ;
  assign n7480 = n7478 & n7479 ;
  assign n7481 = n7475 & ~n7480 ;
  assign n7482 = n7475 & n7479 ;
  assign n7483 = ~x145 & x146 ;
  assign n7484 = x145 & ~x146 ;
  assign n7485 = n7483 | n7484 ;
  assign n7486 = ~x147 & n7485 ;
  assign n7487 = x147 & ~n7485 ;
  assign n7488 = n7486 | n7487 ;
  assign n7489 = ~x148 & x149 ;
  assign n7490 = x148 & ~x149 ;
  assign n7491 = n7489 | n7490 ;
  assign n7492 = ~x150 & n7491 ;
  assign n7493 = x150 & ~n7491 ;
  assign n7494 = n7492 | n7493 ;
  assign n7495 = n7488 & ~n7494 ;
  assign n7496 = ~n7488 & n7494 ;
  assign n7497 = n7495 | n7496 ;
  assign n7498 = ( x148 & x149 ) | ( x148 & x150 ) | ( x149 & x150 ) ;
  assign n7499 = ( x145 & x146 ) | ( x145 & x147 ) | ( x146 & x147 ) ;
  assign n7500 = n7488 & n7494 ;
  assign n7501 = ( n7498 & n7499 ) | ( n7498 & n7500 ) | ( n7499 & n7500 ) ;
  assign n7502 = n7497 & n7501 ;
  assign n7503 = n7482 | n7502 ;
  assign n7504 = n7498 & ~n7499 ;
  assign n7505 = ~n7498 & n7499 ;
  assign n7506 = n7504 | n7505 ;
  assign n7507 = ~n7500 & n7506 ;
  assign n7508 = n7500 & ~n7506 ;
  assign n7509 = n7507 | n7508 ;
  assign n7510 = n7501 & n7509 ;
  assign n7511 = n7478 & n7497 ;
  assign n7512 = n7509 & n7511 ;
  assign n7513 = ~n7510 & n7512 ;
  assign n7514 = ~n7503 & n7513 ;
  assign n7515 = n7481 & n7514 ;
  assign n7516 = ~n7510 & n7511 ;
  assign n7517 = ~n7502 & n7509 ;
  assign n7518 = n7482 & ~n7517 ;
  assign n7519 = ( n7516 & n7517 ) | ( n7516 & ~n7518 ) | ( n7517 & ~n7518 ) ;
  assign n7520 = ( n7481 & n7515 ) | ( n7481 & ~n7519 ) | ( n7515 & ~n7519 ) ;
  assign n7521 = n7497 & ~n7501 ;
  assign n7522 = ( n7497 & ~n7509 ) | ( n7497 & n7521 ) | ( ~n7509 & n7521 ) ;
  assign n7523 = n7478 & ~n7479 ;
  assign n7524 = ( ~n7475 & n7478 ) | ( ~n7475 & n7523 ) | ( n7478 & n7523 ) ;
  assign n7525 = ~n7522 & n7524 ;
  assign n7526 = n7522 & ~n7524 ;
  assign n7527 = n7525 | n7526 ;
  assign n7528 = ( x136 & x137 ) | ( x136 & x138 ) | ( x137 & x138 ) ;
  assign n7529 = ( x133 & x134 ) | ( x133 & x135 ) | ( x134 & x135 ) ;
  assign n7530 = n7528 & ~n7529 ;
  assign n7531 = ~n7528 & n7529 ;
  assign n7532 = n7530 | n7531 ;
  assign n7533 = ~x133 & x134 ;
  assign n7534 = x133 & ~x134 ;
  assign n7535 = n7533 | n7534 ;
  assign n7536 = ~x135 & n7535 ;
  assign n7537 = x135 & ~n7535 ;
  assign n7538 = n7536 | n7537 ;
  assign n7539 = ~x136 & x137 ;
  assign n7540 = x136 & ~x137 ;
  assign n7541 = n7539 | n7540 ;
  assign n7542 = ~x138 & n7541 ;
  assign n7543 = x138 & ~n7541 ;
  assign n7544 = n7542 | n7543 ;
  assign n7545 = n7538 & n7544 ;
  assign n7546 = n7532 & ~n7545 ;
  assign n7547 = ~n7532 & n7545 ;
  assign n7548 = n7546 | n7547 ;
  assign n7549 = n7538 & ~n7544 ;
  assign n7550 = ~n7538 & n7544 ;
  assign n7551 = n7549 | n7550 ;
  assign n7552 = ( n7528 & n7529 ) | ( n7528 & n7545 ) | ( n7529 & n7545 ) ;
  assign n7553 = n7551 & ~n7552 ;
  assign n7554 = ( ~n7548 & n7551 ) | ( ~n7548 & n7553 ) | ( n7551 & n7553 ) ;
  assign n7555 = ~x127 & x128 ;
  assign n7556 = x127 & ~x128 ;
  assign n7557 = n7555 | n7556 ;
  assign n7558 = ~x129 & n7557 ;
  assign n7559 = x129 & ~n7557 ;
  assign n7560 = n7558 | n7559 ;
  assign n7561 = ~x130 & x131 ;
  assign n7562 = x130 & ~x131 ;
  assign n7563 = n7561 | n7562 ;
  assign n7564 = ~x132 & n7563 ;
  assign n7565 = x132 & ~n7563 ;
  assign n7566 = n7564 | n7565 ;
  assign n7567 = n7560 & ~n7566 ;
  assign n7568 = ~n7560 & n7566 ;
  assign n7569 = n7567 | n7568 ;
  assign n7570 = ( x130 & x131 ) | ( x130 & x132 ) | ( x131 & x132 ) ;
  assign n7571 = ( x127 & x128 ) | ( x127 & x129 ) | ( x128 & x129 ) ;
  assign n7572 = n7570 & ~n7571 ;
  assign n7573 = ~n7570 & n7571 ;
  assign n7574 = n7572 | n7573 ;
  assign n7575 = n7560 & n7566 ;
  assign n7576 = n7574 & ~n7575 ;
  assign n7577 = ~n7574 & n7575 ;
  assign n7578 = n7576 | n7577 ;
  assign n7579 = ( n7570 & n7571 ) | ( n7570 & n7575 ) | ( n7571 & n7575 ) ;
  assign n7580 = n7569 & ~n7579 ;
  assign n7581 = ( n7569 & ~n7578 ) | ( n7569 & n7580 ) | ( ~n7578 & n7580 ) ;
  assign n7582 = ~n7554 & n7581 ;
  assign n7583 = n7554 & ~n7581 ;
  assign n7584 = n7582 | n7583 ;
  assign n7585 = n7527 & n7584 ;
  assign n7586 = ( n7481 & ~n7482 ) | ( n7481 & n7517 ) | ( ~n7482 & n7517 ) ;
  assign n7587 = n7481 & n7517 ;
  assign n7588 = ( n7516 & n7586 ) | ( n7516 & n7587 ) | ( n7586 & n7587 ) ;
  assign n7589 = n7519 & ~n7588 ;
  assign n7590 = n7585 | n7589 ;
  assign n7591 = n7520 | n7590 ;
  assign n7592 = n7578 & n7579 ;
  assign n7593 = n7551 & n7552 ;
  assign n7594 = n7592 | n7593 ;
  assign n7595 = n7548 & n7552 ;
  assign n7596 = n7551 & n7569 ;
  assign n7597 = n7548 & n7596 ;
  assign n7598 = ~n7595 & n7597 ;
  assign n7599 = ~n7594 & n7598 ;
  assign n7600 = n7569 & n7579 ;
  assign n7601 = n7578 & ~n7600 ;
  assign n7602 = ~n7599 & n7601 ;
  assign n7603 = ~n7595 & n7596 ;
  assign n7604 = n7548 & ~n7593 ;
  assign n7605 = ( n7592 & n7601 ) | ( n7592 & n7604 ) | ( n7601 & n7604 ) ;
  assign n7606 = n7601 | n7604 ;
  assign n7607 = ( ~n7603 & n7605 ) | ( ~n7603 & n7606 ) | ( n7605 & n7606 ) ;
  assign n7608 = n7592 | n7604 ;
  assign n7609 = n7603 & ~n7608 ;
  assign n7610 = ( ~n7604 & n7607 ) | ( ~n7604 & n7609 ) | ( n7607 & n7609 ) ;
  assign n7611 = ( ~n7602 & n7607 ) | ( ~n7602 & n7610 ) | ( n7607 & n7610 ) ;
  assign n7612 = n7591 & n7611 ;
  assign n7613 = n7585 & n7589 ;
  assign n7614 = ( n7520 & n7585 ) | ( n7520 & n7613 ) | ( n7585 & n7613 ) ;
  assign n7615 = n7612 | n7614 ;
  assign n7616 = n7592 & ~n7604 ;
  assign n7617 = ( n7603 & n7604 ) | ( n7603 & ~n7616 ) | ( n7604 & ~n7616 ) ;
  assign n7618 = n7601 & n7617 ;
  assign n7619 = ~n7569 & n7579 ;
  assign n7620 = ( ~n7578 & n7579 ) | ( ~n7578 & n7619 ) | ( n7579 & n7619 ) ;
  assign n7621 = ~n7551 & n7552 ;
  assign n7622 = ( ~n7548 & n7552 ) | ( ~n7548 & n7621 ) | ( n7552 & n7621 ) ;
  assign n7623 = ~n7620 & n7622 ;
  assign n7624 = n7620 & ~n7622 ;
  assign n7625 = n7623 | n7624 ;
  assign n7626 = n7599 | n7625 ;
  assign n7627 = n7618 | n7626 ;
  assign n7628 = n7599 & n7625 ;
  assign n7629 = ( n7618 & n7625 ) | ( n7618 & n7628 ) | ( n7625 & n7628 ) ;
  assign n7630 = n7627 & ~n7629 ;
  assign n7631 = n7481 & n7519 ;
  assign n7632 = ~n7478 & n7479 ;
  assign n7633 = ( ~n7475 & n7479 ) | ( ~n7475 & n7632 ) | ( n7479 & n7632 ) ;
  assign n7634 = ~n7497 & n7501 ;
  assign n7635 = ( n7501 & ~n7509 ) | ( n7501 & n7634 ) | ( ~n7509 & n7634 ) ;
  assign n7636 = ~n7633 & n7635 ;
  assign n7637 = n7633 & ~n7635 ;
  assign n7638 = n7636 | n7637 ;
  assign n7639 = n7514 | n7638 ;
  assign n7640 = n7631 | n7639 ;
  assign n7641 = n7514 & n7638 ;
  assign n7642 = ( n7631 & n7638 ) | ( n7631 & n7641 ) | ( n7638 & n7641 ) ;
  assign n7643 = n7640 & ~n7642 ;
  assign n7644 = n7630 | n7643 ;
  assign n7645 = n7615 & n7644 ;
  assign n7646 = n7627 & n7640 ;
  assign n7647 = n7629 | n7642 ;
  assign n7648 = n7646 & ~n7647 ;
  assign n7649 = ( n7514 & n7633 ) | ( n7514 & n7635 ) | ( n7633 & n7635 ) ;
  assign n7650 = n7633 | n7635 ;
  assign n7651 = ( n7631 & n7649 ) | ( n7631 & n7650 ) | ( n7649 & n7650 ) ;
  assign n7652 = ( n7599 & n7620 ) | ( n7599 & n7622 ) | ( n7620 & n7622 ) ;
  assign n7653 = n7620 | n7622 ;
  assign n7654 = ( n7618 & n7652 ) | ( n7618 & n7653 ) | ( n7652 & n7653 ) ;
  assign n7655 = ~n7651 & n7654 ;
  assign n7656 = n7651 & ~n7654 ;
  assign n7657 = n7655 | n7656 ;
  assign n7658 = n7648 | n7657 ;
  assign n7659 = n7645 | n7658 ;
  assign n7660 = n7644 | n7648 ;
  assign n7661 = ( n7615 & n7648 ) | ( n7615 & n7660 ) | ( n7648 & n7660 ) ;
  assign n7662 = n7657 & n7661 ;
  assign n7663 = n7659 & ~n7662 ;
  assign n7664 = n7454 | n7663 ;
  assign n7665 = n7382 & ~n7405 ;
  assign n7666 = n7402 & ~n7665 ;
  assign n7667 = n7318 & ~n7375 ;
  assign n7668 = ~n7318 & n7375 ;
  assign n7669 = n7667 | n7668 ;
  assign n7670 = n7527 & ~n7584 ;
  assign n7671 = ~n7527 & n7584 ;
  assign n7672 = n7670 | n7671 ;
  assign n7673 = n7669 & n7672 ;
  assign n7674 = ~n7376 & n7382 ;
  assign n7675 = n7382 & ~n7402 ;
  assign n7676 = n7311 | n7380 ;
  assign n7677 = n7402 | n7676 ;
  assign n7678 = ( n7674 & n7675 ) | ( n7674 & ~n7677 ) | ( n7675 & ~n7677 ) ;
  assign n7679 = n7673 | n7678 ;
  assign n7680 = n7666 | n7679 ;
  assign n7681 = n7520 | n7589 ;
  assign n7682 = ( n7585 & n7611 ) | ( n7585 & ~n7681 ) | ( n7611 & ~n7681 ) ;
  assign n7683 = ( ~n7611 & n7681 ) | ( ~n7611 & n7682 ) | ( n7681 & n7682 ) ;
  assign n7684 = ( ~n7585 & n7682 ) | ( ~n7585 & n7683 ) | ( n7682 & n7683 ) ;
  assign n7685 = n7680 & n7684 ;
  assign n7686 = n7666 | n7678 ;
  assign n7687 = n7673 & n7686 ;
  assign n7688 = ( n7614 & ~n7630 ) | ( n7614 & n7643 ) | ( ~n7630 & n7643 ) ;
  assign n7689 = n7630 & ~n7643 ;
  assign n7690 = ( n7612 & n7688 ) | ( n7612 & ~n7689 ) | ( n7688 & ~n7689 ) ;
  assign n7691 = ( ~n7615 & n7630 ) | ( ~n7615 & n7690 ) | ( n7630 & n7690 ) ;
  assign n7692 = ( ~n7643 & n7690 ) | ( ~n7643 & n7691 ) | ( n7690 & n7691 ) ;
  assign n7693 = ( n7405 & ~n7421 ) | ( n7405 & n7434 ) | ( ~n7421 & n7434 ) ;
  assign n7694 = n7421 & ~n7434 ;
  assign n7695 = ( n7403 & n7693 ) | ( n7403 & ~n7694 ) | ( n7693 & ~n7694 ) ;
  assign n7696 = ( ~n7406 & n7421 ) | ( ~n7406 & n7695 ) | ( n7421 & n7695 ) ;
  assign n7697 = ( ~n7434 & n7695 ) | ( ~n7434 & n7696 ) | ( n7695 & n7696 ) ;
  assign n7698 = ( n7687 & n7692 ) | ( n7687 & n7697 ) | ( n7692 & n7697 ) ;
  assign n7699 = n7692 | n7697 ;
  assign n7700 = ( n7685 & n7698 ) | ( n7685 & n7699 ) | ( n7698 & n7699 ) ;
  assign n7701 = n7664 & n7700 ;
  assign n7702 = n7450 & n7659 ;
  assign n7703 = n7453 | n7662 ;
  assign n7704 = n7702 & ~n7703 ;
  assign n7705 = n7651 & n7654 ;
  assign n7706 = n7651 | n7654 ;
  assign n7707 = n7705 | n7706 ;
  assign n7708 = ( n7661 & n7705 ) | ( n7661 & n7707 ) | ( n7705 & n7707 ) ;
  assign n7709 = n7442 & n7445 ;
  assign n7710 = n7442 | n7445 ;
  assign n7711 = n7709 | n7710 ;
  assign n7712 = ( n7452 & n7709 ) | ( n7452 & n7711 ) | ( n7709 & n7711 ) ;
  assign n7713 = n7708 & n7712 ;
  assign n7714 = n7712 & ~n7713 ;
  assign n7715 = ( n7708 & ~n7713 ) | ( n7708 & n7714 ) | ( ~n7713 & n7714 ) ;
  assign n7716 = n7704 | n7715 ;
  assign n7717 = n7701 | n7716 ;
  assign n7718 = n7701 | n7704 ;
  assign n7719 = n7715 & n7718 ;
  assign n7720 = n7717 & ~n7719 ;
  assign n7721 = n7245 | n7720 ;
  assign n7722 = n7669 & ~n7672 ;
  assign n7723 = ~n7669 & n7672 ;
  assign n7724 = n7722 | n7723 ;
  assign n7725 = n7194 & ~n7197 ;
  assign n7726 = ~n7194 & n7197 ;
  assign n7727 = n7725 | n7726 ;
  assign n7728 = n7724 & n7727 ;
  assign n7729 = ~n7680 & n7684 ;
  assign n7730 = ( n7684 & n7687 ) | ( n7684 & n7729 ) | ( n7687 & n7729 ) ;
  assign n7731 = ~n7673 & n7686 ;
  assign n7732 = n7673 & ~n7678 ;
  assign n7733 = ~n7666 & n7732 ;
  assign n7734 = ~n7684 & n7733 ;
  assign n7735 = ( ~n7684 & n7731 ) | ( ~n7684 & n7734 ) | ( n7731 & n7734 ) ;
  assign n7736 = n7730 | n7735 ;
  assign n7737 = n7728 & n7736 ;
  assign n7738 = n7728 | n7731 ;
  assign n7739 = n7684 & ~n7728 ;
  assign n7740 = ( n7734 & n7738 ) | ( n7734 & ~n7739 ) | ( n7738 & ~n7739 ) ;
  assign n7741 = n7730 | n7740 ;
  assign n7742 = ~n7198 & n7211 ;
  assign n7743 = n7198 & ~n7203 ;
  assign n7744 = ~n7191 & n7743 ;
  assign n7745 = ~n7209 & n7744 ;
  assign n7746 = ( ~n7209 & n7742 ) | ( ~n7209 & n7745 ) | ( n7742 & n7745 ) ;
  assign n7747 = n7210 & ~n7212 ;
  assign n7748 = ( n7209 & n7746 ) | ( n7209 & ~n7747 ) | ( n7746 & ~n7747 ) ;
  assign n7749 = n7741 & n7748 ;
  assign n7750 = n7737 | n7749 ;
  assign n7752 = ( n7212 & ~n7217 ) | ( n7212 & n7222 ) | ( ~n7217 & n7222 ) ;
  assign n7753 = n7217 & ~n7222 ;
  assign n7754 = ( n7210 & n7752 ) | ( n7210 & ~n7753 ) | ( n7752 & ~n7753 ) ;
  assign n7751 = n7210 | n7212 ;
  assign n7755 = ( n7217 & ~n7751 ) | ( n7217 & n7754 ) | ( ~n7751 & n7754 ) ;
  assign n7756 = ( ~n7222 & n7754 ) | ( ~n7222 & n7755 ) | ( n7754 & n7755 ) ;
  assign n7758 = ( n7687 & ~n7692 ) | ( n7687 & n7697 ) | ( ~n7692 & n7697 ) ;
  assign n7759 = n7692 & ~n7697 ;
  assign n7760 = ( n7685 & n7758 ) | ( n7685 & ~n7759 ) | ( n7758 & ~n7759 ) ;
  assign n7757 = n7685 | n7687 ;
  assign n7761 = ( n7692 & ~n7757 ) | ( n7692 & n7760 ) | ( ~n7757 & n7760 ) ;
  assign n7762 = ( ~n7697 & n7760 ) | ( ~n7697 & n7761 ) | ( n7760 & n7761 ) ;
  assign n7763 = ( n7750 & n7756 ) | ( n7750 & n7762 ) | ( n7756 & n7762 ) ;
  assign n7764 = ( ~n7454 & n7663 ) | ( ~n7454 & n7700 ) | ( n7663 & n7700 ) ;
  assign n7765 = ( n7454 & ~n7700 ) | ( n7454 & n7764 ) | ( ~n7700 & n7764 ) ;
  assign n7766 = ( ~n7663 & n7764 ) | ( ~n7663 & n7765 ) | ( n7764 & n7765 ) ;
  assign n7767 = ( ~n6979 & n7188 ) | ( ~n6979 & n7225 ) | ( n7188 & n7225 ) ;
  assign n7768 = ( n6979 & ~n7225 ) | ( n6979 & n7767 ) | ( ~n7225 & n7767 ) ;
  assign n7769 = ( ~n7188 & n7767 ) | ( ~n7188 & n7768 ) | ( n7767 & n7768 ) ;
  assign n7770 = ( n7763 & n7766 ) | ( n7763 & n7769 ) | ( n7766 & n7769 ) ;
  assign n7771 = n7721 & n7770 ;
  assign n7772 = n7242 & n7717 ;
  assign n7773 = n7244 | n7719 ;
  assign n7774 = n7772 & ~n7773 ;
  assign n7783 = n6977 & n7235 ;
  assign n7784 = n7179 | n7234 ;
  assign n7785 = n7176 | n7234 ;
  assign n7786 = ( n7186 & n7784 ) | ( n7186 & n7785 ) | ( n7784 & n7785 ) ;
  assign n7787 = n7783 | n7786 ;
  assign n7788 = n7238 | n7787 ;
  assign n7789 = ( n7229 & n7238 ) | ( n7229 & n7788 ) | ( n7238 & n7788 ) ;
  assign n7790 = n7238 | n7788 ;
  assign n7791 = ( n7226 & n7789 ) | ( n7226 & n7790 ) | ( n7789 & n7790 ) ;
  assign n7775 = n7452 & n7710 ;
  assign n7776 = n7654 | n7709 ;
  assign n7777 = n7651 | n7709 ;
  assign n7778 = ( n7661 & n7776 ) | ( n7661 & n7777 ) | ( n7776 & n7777 ) ;
  assign n7779 = n7775 | n7778 ;
  assign n7780 = n7704 & n7779 ;
  assign n7781 = ( n7701 & n7779 ) | ( n7701 & n7780 ) | ( n7779 & n7780 ) ;
  assign n7782 = n7713 | n7781 ;
  assign n7792 = n7782 & n7791 ;
  assign n7793 = n7782 & ~n7792 ;
  assign n7794 = ( n7791 & ~n7792 ) | ( n7791 & n7793 ) | ( ~n7792 & n7793 ) ;
  assign n7795 = n7774 | n7794 ;
  assign n7796 = n7771 | n7795 ;
  assign n7797 = n7771 | n7774 ;
  assign n7798 = n7794 & n7797 ;
  assign n7799 = n7796 & ~n7798 ;
  assign n7800 = n6770 | n7799 ;
  assign n7801 = ( ~n7245 & n7720 ) | ( ~n7245 & n7770 ) | ( n7720 & n7770 ) ;
  assign n7802 = ( n7245 & ~n7770 ) | ( n7245 & n7801 ) | ( ~n7770 & n7801 ) ;
  assign n7803 = ( ~n7720 & n7801 ) | ( ~n7720 & n7802 ) | ( n7801 & n7802 ) ;
  assign n7804 = ( ~n6218 & n6693 ) | ( ~n6218 & n6741 ) | ( n6693 & n6741 ) ;
  assign n7805 = ( n6218 & ~n6741 ) | ( n6218 & n7804 ) | ( ~n6741 & n7804 ) ;
  assign n7806 = ( ~n6693 & n7804 ) | ( ~n6693 & n7805 ) | ( n7804 & n7805 ) ;
  assign n7807 = n6710 & ~n6713 ;
  assign n7808 = ~n6710 & n6713 ;
  assign n7809 = n7807 | n7808 ;
  assign n7810 = n7724 & ~n7727 ;
  assign n7811 = ~n7724 & n7727 ;
  assign n7812 = n7810 | n7811 ;
  assign n7813 = n7809 & n7812 ;
  assign n7814 = n6723 & ~n6725 ;
  assign n7815 = n6707 & ~n7814 ;
  assign n7816 = ~n6714 & n6722 ;
  assign n7817 = n6714 & ~n6722 ;
  assign n7818 = n7816 | n7817 ;
  assign n7819 = ~n6707 & n7818 ;
  assign n7820 = n7815 | n7819 ;
  assign n7821 = n7813 & n7820 ;
  assign n7822 = n6707 & ~n7813 ;
  assign n7823 = ( n7813 & n7818 ) | ( n7813 & ~n7822 ) | ( n7818 & ~n7822 ) ;
  assign n7824 = n7815 | n7823 ;
  assign n7825 = ( n7728 & ~n7736 ) | ( n7728 & n7748 ) | ( ~n7736 & n7748 ) ;
  assign n7826 = ( ~n7728 & n7736 ) | ( ~n7728 & n7825 ) | ( n7736 & n7825 ) ;
  assign n7827 = ( ~n7748 & n7825 ) | ( ~n7748 & n7826 ) | ( n7825 & n7826 ) ;
  assign n7828 = n7824 & n7827 ;
  assign n7829 = n7821 | n7828 ;
  assign n7830 = ( n7750 & ~n7756 ) | ( n7750 & n7762 ) | ( ~n7756 & n7762 ) ;
  assign n7831 = ( ~n7750 & n7756 ) | ( ~n7750 & n7830 ) | ( n7756 & n7830 ) ;
  assign n7832 = ( ~n7762 & n7830 ) | ( ~n7762 & n7831 ) | ( n7830 & n7831 ) ;
  assign n7834 = ( n6725 & ~n6731 ) | ( n6725 & n6737 ) | ( ~n6731 & n6737 ) ;
  assign n7835 = n6731 & ~n6737 ;
  assign n7836 = ( n6724 & n7834 ) | ( n6724 & ~n7835 ) | ( n7834 & ~n7835 ) ;
  assign n7833 = n6724 | n6725 ;
  assign n7837 = ( n6731 & ~n7833 ) | ( n6731 & n7836 ) | ( ~n7833 & n7836 ) ;
  assign n7838 = ( ~n6737 & n7836 ) | ( ~n6737 & n7837 ) | ( n7836 & n7837 ) ;
  assign n7839 = ( n7829 & n7832 ) | ( n7829 & n7838 ) | ( n7832 & n7838 ) ;
  assign n7840 = ( ~n6697 & n6700 ) | ( ~n6697 & n6740 ) | ( n6700 & n6740 ) ;
  assign n7841 = ( n6697 & ~n6740 ) | ( n6697 & n7840 ) | ( ~n6740 & n7840 ) ;
  assign n7842 = ( ~n6700 & n7840 ) | ( ~n6700 & n7841 ) | ( n7840 & n7841 ) ;
  assign n7843 = ( n7763 & ~n7766 ) | ( n7763 & n7769 ) | ( ~n7766 & n7769 ) ;
  assign n7844 = ( ~n7763 & n7766 ) | ( ~n7763 & n7843 ) | ( n7766 & n7843 ) ;
  assign n7845 = ( ~n7769 & n7843 ) | ( ~n7769 & n7844 ) | ( n7843 & n7844 ) ;
  assign n7846 = ( n7839 & n7842 ) | ( n7839 & n7845 ) | ( n7842 & n7845 ) ;
  assign n7847 = ( n7803 & n7806 ) | ( n7803 & n7846 ) | ( n7806 & n7846 ) ;
  assign n7848 = n7800 & n7847 ;
  assign n7849 = n6767 & n7796 ;
  assign n7850 = n6769 | n7798 ;
  assign n7851 = n7849 & ~n7850 ;
  assign n7859 = n7238 | n7713 ;
  assign n7860 = n7787 | n7859 ;
  assign n7861 = ( n7243 & n7859 ) | ( n7243 & n7860 ) | ( n7859 & n7860 ) ;
  assign n7862 = n7781 | n7861 ;
  assign n7863 = n7792 | n7862 ;
  assign n7864 = ( n7774 & n7792 ) | ( n7774 & n7863 ) | ( n7792 & n7863 ) ;
  assign n7865 = n7792 | n7863 ;
  assign n7866 = ( n7771 & n7864 ) | ( n7771 & n7865 ) | ( n7864 & n7865 ) ;
  assign n7852 = n6211 | n6686 ;
  assign n7853 = n6758 | n7852 ;
  assign n7854 = ( n6216 & n7852 ) | ( n6216 & n7853 ) | ( n7852 & n7853 ) ;
  assign n7855 = n6752 | n7854 ;
  assign n7856 = n6745 & n7855 ;
  assign n7857 = ( n6742 & n7855 ) | ( n6742 & n7856 ) | ( n7855 & n7856 ) ;
  assign n7858 = n6763 | n7857 ;
  assign n7867 = n7858 & n7866 ;
  assign n7868 = n7858 & ~n7867 ;
  assign n7869 = ( n7866 & ~n7867 ) | ( n7866 & n7868 ) | ( ~n7867 & n7868 ) ;
  assign n7870 = n7851 | n7869 ;
  assign n7871 = n7848 | n7870 ;
  assign n7872 = n7848 | n7851 ;
  assign n7873 = n7869 & n7872 ;
  assign n7874 = n7871 & ~n7873 ;
  assign n7875 = ( ~n4639 & n5668 ) | ( ~n4639 & n5716 ) | ( n5668 & n5716 ) ;
  assign n7876 = ( n4639 & ~n5716 ) | ( n4639 & n7875 ) | ( ~n5716 & n7875 ) ;
  assign n7877 = ( ~n5668 & n7875 ) | ( ~n5668 & n7876 ) | ( n7875 & n7876 ) ;
  assign n7878 = ( ~n6770 & n7799 ) | ( ~n6770 & n7847 ) | ( n7799 & n7847 ) ;
  assign n7879 = ( n6770 & ~n7847 ) | ( n6770 & n7878 ) | ( ~n7847 & n7878 ) ;
  assign n7880 = ( ~n7799 & n7878 ) | ( ~n7799 & n7879 ) | ( n7878 & n7879 ) ;
  assign n7881 = n5678 & ~n5681 ;
  assign n7882 = ~n5678 & n5681 ;
  assign n7883 = n7881 | n7882 ;
  assign n7884 = n7809 & ~n7812 ;
  assign n7885 = ~n7809 & n7812 ;
  assign n7886 = n7884 | n7885 ;
  assign n7887 = n7883 & n7886 ;
  assign n7888 = ~n5693 & n5696 ;
  assign n7889 = ( n5690 & n5696 ) | ( n5690 & n7888 ) | ( n5696 & n7888 ) ;
  assign n7890 = ~n5682 & n5689 ;
  assign n7891 = n4576 & n5682 ;
  assign n7892 = ( n5682 & ~n5687 ) | ( n5682 & n7891 ) | ( ~n5687 & n7891 ) ;
  assign n7893 = ~n5684 & n7892 ;
  assign n7894 = ~n5696 & n7893 ;
  assign n7895 = ( ~n5696 & n7890 ) | ( ~n5696 & n7894 ) | ( n7890 & n7894 ) ;
  assign n7896 = n7889 | n7895 ;
  assign n7897 = n7887 & n7896 ;
  assign n7898 = ~n7813 & n7820 ;
  assign n7899 = n6707 & n7813 ;
  assign n7900 = ( n7813 & ~n7818 ) | ( n7813 & n7899 ) | ( ~n7818 & n7899 ) ;
  assign n7901 = ~n7815 & n7900 ;
  assign n7902 = ~n7827 & n7901 ;
  assign n7903 = ( ~n7827 & n7898 ) | ( ~n7827 & n7902 ) | ( n7898 & n7902 ) ;
  assign n7904 = ~n7821 & n7828 ;
  assign n7905 = ( n7827 & n7903 ) | ( n7827 & ~n7904 ) | ( n7903 & ~n7904 ) ;
  assign n7906 = n7887 | n7896 ;
  assign n7907 = n7905 & n7906 ;
  assign n7908 = n7897 | n7907 ;
  assign n7909 = ( n7829 & ~n7832 ) | ( n7829 & n7838 ) | ( ~n7832 & n7838 ) ;
  assign n7910 = ( ~n7829 & n7832 ) | ( ~n7829 & n7909 ) | ( n7832 & n7909 ) ;
  assign n7911 = ( ~n7838 & n7909 ) | ( ~n7838 & n7910 ) | ( n7909 & n7910 ) ;
  assign n7912 = ( n5698 & ~n5701 ) | ( n5698 & n5707 ) | ( ~n5701 & n5707 ) ;
  assign n7913 = ( ~n5698 & n5701 ) | ( ~n5698 & n7912 ) | ( n5701 & n7912 ) ;
  assign n7914 = ( ~n5707 & n7912 ) | ( ~n5707 & n7913 ) | ( n7912 & n7913 ) ;
  assign n7915 = ( n7908 & n7911 ) | ( n7908 & n7914 ) | ( n7911 & n7914 ) ;
  assign n7916 = ( n7803 & ~n7806 ) | ( n7803 & n7846 ) | ( ~n7806 & n7846 ) ;
  assign n7917 = ( ~n7803 & n7806 ) | ( ~n7803 & n7846 ) | ( n7806 & n7846 ) ;
  assign n7918 = ( ~n7846 & n7916 ) | ( ~n7846 & n7917 ) | ( n7916 & n7917 ) ;
  assign n7919 = ( n5672 & ~n5675 ) | ( n5672 & n5715 ) | ( ~n5675 & n5715 ) ;
  assign n7920 = ( ~n5672 & n5675 ) | ( ~n5672 & n5715 ) | ( n5675 & n5715 ) ;
  assign n7921 = ( ~n5715 & n7919 ) | ( ~n5715 & n7920 ) | ( n7919 & n7920 ) ;
  assign n7922 = ( n7839 & ~n7842 ) | ( n7839 & n7845 ) | ( ~n7842 & n7845 ) ;
  assign n7923 = ( ~n7839 & n7842 ) | ( ~n7839 & n7922 ) | ( n7842 & n7922 ) ;
  assign n7924 = ( ~n7845 & n7922 ) | ( ~n7845 & n7923 ) | ( n7922 & n7923 ) ;
  assign n7925 = ( n7918 & n7921 ) | ( n7918 & n7924 ) | ( n7921 & n7924 ) ;
  assign n7926 = ( n5708 & ~n5711 ) | ( n5708 & n5714 ) | ( ~n5711 & n5714 ) ;
  assign n7927 = ( ~n5708 & n5711 ) | ( ~n5708 & n7926 ) | ( n5711 & n7926 ) ;
  assign n7928 = ( ~n5714 & n7926 ) | ( ~n5714 & n7927 ) | ( n7926 & n7927 ) ;
  assign n7929 = ( n7918 & n7921 ) | ( n7918 & n7928 ) | ( n7921 & n7928 ) ;
  assign n7930 = ( n7915 & n7925 ) | ( n7915 & n7929 ) | ( n7925 & n7929 ) ;
  assign n7931 = ( n7877 & n7880 ) | ( n7877 & n7930 ) | ( n7880 & n7930 ) ;
  assign n7932 = ( n5743 & ~n7874 ) | ( n5743 & n7931 ) | ( ~n7874 & n7931 ) ;
  assign n7933 = ( n7874 & ~n7931 ) | ( n7874 & n7932 ) | ( ~n7931 & n7932 ) ;
  assign n7934 = ( ~n5743 & n7932 ) | ( ~n5743 & n7933 ) | ( n7932 & n7933 ) ;
  assign n7935 = n3533 | n3539 ;
  assign n7936 = n3541 & ~n7935 ;
  assign n7937 = n3533 & n3539 ;
  assign n7938 = ( n3533 & ~n3541 ) | ( n3533 & n7937 ) | ( ~n3541 & n7937 ) ;
  assign n7939 = n7936 | n7938 ;
  assign n7940 = n3608 & n7939 ;
  assign n7941 = n3608 | n7939 ;
  assign n7942 = ~n7940 & n7941 ;
  assign n7943 = ( n7877 & ~n7880 ) | ( n7877 & n7930 ) | ( ~n7880 & n7930 ) ;
  assign n7944 = ( ~n7877 & n7880 ) | ( ~n7877 & n7943 ) | ( n7880 & n7943 ) ;
  assign n7945 = ( ~n7930 & n7943 ) | ( ~n7930 & n7944 ) | ( n7943 & n7944 ) ;
  assign n7946 = n3547 | n3551 ;
  assign n7947 = n3546 & ~n7946 ;
  assign n7948 = ~n3548 & n3551 ;
  assign n7949 = n7947 | n7948 ;
  assign n7950 = n3607 & n7949 ;
  assign n7951 = n3607 | n7949 ;
  assign n7952 = ~n7950 & n7951 ;
  assign n7953 = ~n3558 & n3561 ;
  assign n7954 = n2474 | n3561 ;
  assign n7955 = ( n3555 & n3561 ) | ( n3555 & n7954 ) | ( n3561 & n7954 ) ;
  assign n7956 = n3556 & ~n7955 ;
  assign n7957 = n3603 & n7956 ;
  assign n7958 = ( n3603 & n7953 ) | ( n3603 & n7957 ) | ( n7953 & n7957 ) ;
  assign n7959 = n3603 | n7956 ;
  assign n7960 = n7953 | n7959 ;
  assign n7961 = ~n7958 & n7960 ;
  assign n7962 = ~n3599 & n3602 ;
  assign n7963 = n3599 & ~n3602 ;
  assign n7964 = n7962 | n7963 ;
  assign n7965 = n3587 & n7964 ;
  assign n7966 = n3587 | n7964 ;
  assign n7967 = ~n7965 & n7966 ;
  assign n7968 = n7883 & ~n7886 ;
  assign n7969 = ~n7883 & n7886 ;
  assign n7970 = n7968 | n7969 ;
  assign n7971 = n3566 | n3569 ;
  assign n7972 = n3566 & ~n3569 ;
  assign n7973 = ( ~n3566 & n7971 ) | ( ~n3566 & n7972 ) | ( n7971 & n7972 ) ;
  assign n7974 = n7970 & n7973 ;
  assign n7975 = ~n7897 & n7906 ;
  assign n7976 = n7905 & ~n7975 ;
  assign n7977 = ~n7887 & n7896 ;
  assign n7978 = n7887 & ~n7896 ;
  assign n7979 = n7977 | n7978 ;
  assign n7980 = ~n7905 & n7979 ;
  assign n7981 = n7976 | n7980 ;
  assign n7982 = n7974 & n7981 ;
  assign n7983 = n7905 & ~n7974 ;
  assign n7984 = ( n7974 & n7979 ) | ( n7974 & ~n7983 ) | ( n7979 & ~n7983 ) ;
  assign n7985 = n7976 | n7984 ;
  assign n7986 = ( n3570 & ~n3579 ) | ( n3570 & n3584 ) | ( ~n3579 & n3584 ) ;
  assign n7987 = ( ~n3570 & n3579 ) | ( ~n3570 & n7986 ) | ( n3579 & n7986 ) ;
  assign n7988 = ( ~n3584 & n7986 ) | ( ~n3584 & n7987 ) | ( n7986 & n7987 ) ;
  assign n7989 = n7985 & n7988 ;
  assign n7990 = n7982 | n7989 ;
  assign n7991 = ( n7908 & ~n7911 ) | ( n7908 & n7914 ) | ( ~n7911 & n7914 ) ;
  assign n7992 = ( ~n7908 & n7911 ) | ( ~n7908 & n7991 ) | ( n7911 & n7991 ) ;
  assign n7993 = ( ~n7914 & n7991 ) | ( ~n7914 & n7992 ) | ( n7991 & n7992 ) ;
  assign n7994 = ( n7967 & n7990 ) | ( n7967 & n7993 ) | ( n7990 & n7993 ) ;
  assign n7995 = ( n7915 & n7924 ) | ( n7915 & ~n7928 ) | ( n7924 & ~n7928 ) ;
  assign n7996 = ( ~n7915 & n7928 ) | ( ~n7915 & n7995 ) | ( n7928 & n7995 ) ;
  assign n7997 = ( ~n7924 & n7995 ) | ( ~n7924 & n7996 ) | ( n7995 & n7996 ) ;
  assign n7998 = ( n7961 & n7994 ) | ( n7961 & n7997 ) | ( n7994 & n7997 ) ;
  assign n7999 = ( n7915 & n7924 ) | ( n7915 & n7928 ) | ( n7924 & n7928 ) ;
  assign n8000 = ( n7918 & ~n7921 ) | ( n7918 & n7924 ) | ( ~n7921 & n7924 ) ;
  assign n8001 = ( n7918 & ~n7921 ) | ( n7918 & n7928 ) | ( ~n7921 & n7928 ) ;
  assign n8002 = ( n7915 & n8000 ) | ( n7915 & n8001 ) | ( n8000 & n8001 ) ;
  assign n8003 = ( ~n7918 & n7921 ) | ( ~n7918 & n8002 ) | ( n7921 & n8002 ) ;
  assign n8004 = ( ~n7999 & n8002 ) | ( ~n7999 & n8003 ) | ( n8002 & n8003 ) ;
  assign n8005 = ( n7952 & n7998 ) | ( n7952 & n8004 ) | ( n7998 & n8004 ) ;
  assign n8006 = ( n7942 & n7945 ) | ( n7942 & n8005 ) | ( n7945 & n8005 ) ;
  assign n8007 = ( n3612 & n7934 ) | ( n3612 & n8006 ) | ( n7934 & n8006 ) ;
  assign n8008 = n5740 & n7871 ;
  assign n8009 = n5742 | n7873 ;
  assign n8010 = n8008 & ~n8009 ;
  assign n8011 = n5743 | n7874 ;
  assign n8012 = n7931 & n8011 ;
  assign n8013 = n8010 | n8012 ;
  assign n8021 = n6763 | n7792 ;
  assign n8022 = n7862 | n8021 ;
  assign n8023 = ( n7797 & n8021 ) | ( n7797 & n8022 ) | ( n8021 & n8022 ) ;
  assign n8024 = n7857 | n8023 ;
  assign n8025 = n7867 | n8024 ;
  assign n8026 = ( n7851 & n7867 ) | ( n7851 & n8025 ) | ( n7867 & n8025 ) ;
  assign n8027 = n7867 | n8025 ;
  assign n8028 = ( n7848 & n8026 ) | ( n7848 & n8027 ) | ( n8026 & n8027 ) ;
  assign n8014 = n4632 | n5661 ;
  assign n8015 = n5731 | n8014 ;
  assign n8016 = ( n5666 & n8014 ) | ( n5666 & n8015 ) | ( n8014 & n8015 ) ;
  assign n8017 = n5726 | n8016 ;
  assign n8018 = n5720 & n8017 ;
  assign n8019 = ( n5717 & n8017 ) | ( n5717 & n8018 ) | ( n8017 & n8018 ) ;
  assign n8020 = n5736 | n8019 ;
  assign n8029 = n8020 & n8028 ;
  assign n8030 = n8020 & ~n8029 ;
  assign n8031 = ( n8028 & ~n8029 ) | ( n8028 & n8030 ) | ( ~n8029 & n8030 ) ;
  assign n8032 = n8013 & n8031 ;
  assign n8033 = n2478 & n2487 ;
  assign n8034 = ( n3523 & n3610 ) | ( n3523 & n8033 ) | ( n3610 & n8033 ) ;
  assign n8035 = n3523 | n8033 ;
  assign n8036 = n3525 | n8035 ;
  assign n8037 = ( n3609 & n8035 ) | ( n3609 & n8036 ) | ( n8035 & n8036 ) ;
  assign n8038 = ~n8034 & n8037 ;
  assign n8039 = n8010 | n8031 ;
  assign n8040 = n8012 | n8039 ;
  assign n8041 = n8038 & n8040 ;
  assign n8042 = ~n8032 & n8041 ;
  assign n8043 = ~n8032 & n8040 ;
  assign n8044 = n8038 | n8043 ;
  assign n8045 = ~n8042 & n8044 ;
  assign n8046 = n8007 | n8045 ;
  assign n8047 = ( x598 & x599 ) | ( x598 & x600 ) | ( x599 & x600 ) ;
  assign n8048 = ( x595 & x596 ) | ( x595 & x597 ) | ( x596 & x597 ) ;
  assign n8049 = n8047 & ~n8048 ;
  assign n8050 = ~n8047 & n8048 ;
  assign n8051 = n8049 | n8050 ;
  assign n8052 = ~x595 & x596 ;
  assign n8053 = x595 & ~x596 ;
  assign n8054 = n8052 | n8053 ;
  assign n8055 = ~x597 & n8054 ;
  assign n8056 = x597 & ~n8054 ;
  assign n8057 = n8055 | n8056 ;
  assign n8058 = ~x598 & x599 ;
  assign n8059 = x598 & ~x599 ;
  assign n8060 = n8058 | n8059 ;
  assign n8061 = ~x600 & n8060 ;
  assign n8062 = x600 & ~n8060 ;
  assign n8063 = n8061 | n8062 ;
  assign n8064 = n8057 & n8063 ;
  assign n8065 = n8051 & ~n8064 ;
  assign n8066 = ~n8051 & n8064 ;
  assign n8067 = n8065 | n8066 ;
  assign n8068 = n8057 & ~n8063 ;
  assign n8069 = ~n8057 & n8063 ;
  assign n8070 = n8068 | n8069 ;
  assign n8071 = ( n8047 & n8048 ) | ( n8047 & n8064 ) | ( n8048 & n8064 ) ;
  assign n8072 = n8070 & n8071 ;
  assign n8073 = n8067 & ~n8072 ;
  assign n8074 = n8067 & n8071 ;
  assign n8075 = ~x601 & x602 ;
  assign n8076 = x601 & ~x602 ;
  assign n8077 = n8075 | n8076 ;
  assign n8078 = ~x603 & n8077 ;
  assign n8079 = x603 & ~n8077 ;
  assign n8080 = n8078 | n8079 ;
  assign n8081 = ~x604 & x605 ;
  assign n8082 = x604 & ~x605 ;
  assign n8083 = n8081 | n8082 ;
  assign n8084 = ~x606 & n8083 ;
  assign n8085 = x606 & ~n8083 ;
  assign n8086 = n8084 | n8085 ;
  assign n8087 = n8080 & ~n8086 ;
  assign n8088 = ~n8080 & n8086 ;
  assign n8089 = n8087 | n8088 ;
  assign n8090 = ( x604 & x605 ) | ( x604 & x606 ) | ( x605 & x606 ) ;
  assign n8091 = ( x601 & x602 ) | ( x601 & x603 ) | ( x602 & x603 ) ;
  assign n8092 = n8080 & n8086 ;
  assign n8093 = ( n8090 & n8091 ) | ( n8090 & n8092 ) | ( n8091 & n8092 ) ;
  assign n8094 = n8089 & n8093 ;
  assign n8095 = n8074 | n8094 ;
  assign n8096 = n8090 & ~n8091 ;
  assign n8097 = ~n8090 & n8091 ;
  assign n8098 = n8096 | n8097 ;
  assign n8099 = ~n8092 & n8098 ;
  assign n8100 = n8092 & ~n8098 ;
  assign n8101 = n8099 | n8100 ;
  assign n8102 = n8093 & n8101 ;
  assign n8103 = n8070 & n8089 ;
  assign n8104 = n8101 & n8103 ;
  assign n8105 = ~n8102 & n8104 ;
  assign n8106 = ~n8095 & n8105 ;
  assign n8107 = n8073 & n8106 ;
  assign n8108 = ~n8102 & n8103 ;
  assign n8109 = ~n8094 & n8101 ;
  assign n8110 = n8074 & ~n8109 ;
  assign n8111 = ( n8108 & n8109 ) | ( n8108 & ~n8110 ) | ( n8109 & ~n8110 ) ;
  assign n8112 = ( n8073 & n8107 ) | ( n8073 & ~n8111 ) | ( n8107 & ~n8111 ) ;
  assign n8113 = n8089 & ~n8093 ;
  assign n8114 = ( n8089 & ~n8101 ) | ( n8089 & n8113 ) | ( ~n8101 & n8113 ) ;
  assign n8115 = n8070 & ~n8071 ;
  assign n8116 = ( ~n8067 & n8070 ) | ( ~n8067 & n8115 ) | ( n8070 & n8115 ) ;
  assign n8117 = ~n8114 & n8116 ;
  assign n8118 = n8114 & ~n8116 ;
  assign n8119 = n8117 | n8118 ;
  assign n8120 = ( x592 & x593 ) | ( x592 & x594 ) | ( x593 & x594 ) ;
  assign n8121 = ( x589 & x590 ) | ( x589 & x591 ) | ( x590 & x591 ) ;
  assign n8122 = n8120 & ~n8121 ;
  assign n8123 = ~n8120 & n8121 ;
  assign n8124 = n8122 | n8123 ;
  assign n8125 = ~x589 & x590 ;
  assign n8126 = x589 & ~x590 ;
  assign n8127 = n8125 | n8126 ;
  assign n8128 = ~x591 & n8127 ;
  assign n8129 = x591 & ~n8127 ;
  assign n8130 = n8128 | n8129 ;
  assign n8131 = ~x592 & x593 ;
  assign n8132 = x592 & ~x593 ;
  assign n8133 = n8131 | n8132 ;
  assign n8134 = ~x594 & n8133 ;
  assign n8135 = x594 & ~n8133 ;
  assign n8136 = n8134 | n8135 ;
  assign n8137 = n8130 & n8136 ;
  assign n8138 = n8124 & ~n8137 ;
  assign n8139 = ~n8124 & n8137 ;
  assign n8140 = n8138 | n8139 ;
  assign n8141 = n8130 & ~n8136 ;
  assign n8142 = ~n8130 & n8136 ;
  assign n8143 = n8141 | n8142 ;
  assign n8144 = ( n8120 & n8121 ) | ( n8120 & n8137 ) | ( n8121 & n8137 ) ;
  assign n8145 = n8143 & ~n8144 ;
  assign n8146 = ( ~n8140 & n8143 ) | ( ~n8140 & n8145 ) | ( n8143 & n8145 ) ;
  assign n8147 = ~x583 & x584 ;
  assign n8148 = x583 & ~x584 ;
  assign n8149 = n8147 | n8148 ;
  assign n8150 = ~x585 & n8149 ;
  assign n8151 = x585 & ~n8149 ;
  assign n8152 = n8150 | n8151 ;
  assign n8153 = ~x586 & x587 ;
  assign n8154 = x586 & ~x587 ;
  assign n8155 = n8153 | n8154 ;
  assign n8156 = ~x588 & n8155 ;
  assign n8157 = x588 & ~n8155 ;
  assign n8158 = n8156 | n8157 ;
  assign n8159 = n8152 & ~n8158 ;
  assign n8160 = ~n8152 & n8158 ;
  assign n8161 = n8159 | n8160 ;
  assign n8162 = ( x586 & x587 ) | ( x586 & x588 ) | ( x587 & x588 ) ;
  assign n8163 = ( x583 & x584 ) | ( x583 & x585 ) | ( x584 & x585 ) ;
  assign n8164 = n8162 & ~n8163 ;
  assign n8165 = ~n8162 & n8163 ;
  assign n8166 = n8164 | n8165 ;
  assign n8167 = n8152 & n8158 ;
  assign n8168 = n8166 & ~n8167 ;
  assign n8169 = ~n8166 & n8167 ;
  assign n8170 = n8168 | n8169 ;
  assign n8171 = ( n8162 & n8163 ) | ( n8162 & n8167 ) | ( n8163 & n8167 ) ;
  assign n8172 = n8161 & ~n8171 ;
  assign n8173 = ( n8161 & ~n8170 ) | ( n8161 & n8172 ) | ( ~n8170 & n8172 ) ;
  assign n8174 = ~n8146 & n8173 ;
  assign n8175 = n8146 & ~n8173 ;
  assign n8176 = n8174 | n8175 ;
  assign n8177 = n8119 & n8176 ;
  assign n8178 = ( n8073 & ~n8074 ) | ( n8073 & n8109 ) | ( ~n8074 & n8109 ) ;
  assign n8179 = n8073 & n8109 ;
  assign n8180 = ( n8108 & n8178 ) | ( n8108 & n8179 ) | ( n8178 & n8179 ) ;
  assign n8181 = n8111 & ~n8180 ;
  assign n8182 = n8177 | n8181 ;
  assign n8183 = n8112 | n8182 ;
  assign n8184 = n8170 & n8171 ;
  assign n8185 = n8143 & n8144 ;
  assign n8186 = n8184 | n8185 ;
  assign n8187 = n8140 & n8144 ;
  assign n8188 = n8143 & n8161 ;
  assign n8189 = n8140 & n8188 ;
  assign n8190 = ~n8187 & n8189 ;
  assign n8191 = ~n8186 & n8190 ;
  assign n8192 = n8161 & n8171 ;
  assign n8193 = n8170 & ~n8192 ;
  assign n8194 = ~n8191 & n8193 ;
  assign n8195 = ~n8187 & n8188 ;
  assign n8196 = n8140 & ~n8185 ;
  assign n8197 = ( n8184 & n8193 ) | ( n8184 & n8196 ) | ( n8193 & n8196 ) ;
  assign n8198 = n8193 | n8196 ;
  assign n8199 = ( ~n8195 & n8197 ) | ( ~n8195 & n8198 ) | ( n8197 & n8198 ) ;
  assign n8200 = n8184 | n8196 ;
  assign n8201 = n8195 & ~n8200 ;
  assign n8202 = ( ~n8196 & n8199 ) | ( ~n8196 & n8201 ) | ( n8199 & n8201 ) ;
  assign n8203 = ( ~n8194 & n8199 ) | ( ~n8194 & n8202 ) | ( n8199 & n8202 ) ;
  assign n8204 = n8183 & n8203 ;
  assign n8205 = n8177 & n8181 ;
  assign n8206 = ( n8112 & n8177 ) | ( n8112 & n8205 ) | ( n8177 & n8205 ) ;
  assign n8207 = n8204 | n8206 ;
  assign n8208 = n8184 & ~n8196 ;
  assign n8209 = ( n8195 & n8196 ) | ( n8195 & ~n8208 ) | ( n8196 & ~n8208 ) ;
  assign n8210 = n8193 & n8209 ;
  assign n8211 = ~n8161 & n8171 ;
  assign n8212 = ( ~n8170 & n8171 ) | ( ~n8170 & n8211 ) | ( n8171 & n8211 ) ;
  assign n8213 = ~n8143 & n8144 ;
  assign n8214 = ( ~n8140 & n8144 ) | ( ~n8140 & n8213 ) | ( n8144 & n8213 ) ;
  assign n8215 = ~n8212 & n8214 ;
  assign n8216 = n8212 & ~n8214 ;
  assign n8217 = n8215 | n8216 ;
  assign n8218 = n8191 | n8217 ;
  assign n8219 = n8210 | n8218 ;
  assign n8220 = n8191 & n8217 ;
  assign n8221 = ( n8210 & n8217 ) | ( n8210 & n8220 ) | ( n8217 & n8220 ) ;
  assign n8222 = n8219 & ~n8221 ;
  assign n8223 = n8073 & n8111 ;
  assign n8224 = ~n8070 & n8071 ;
  assign n8225 = ( ~n8067 & n8071 ) | ( ~n8067 & n8224 ) | ( n8071 & n8224 ) ;
  assign n8226 = ~n8089 & n8093 ;
  assign n8227 = ( n8093 & ~n8101 ) | ( n8093 & n8226 ) | ( ~n8101 & n8226 ) ;
  assign n8228 = ~n8225 & n8227 ;
  assign n8229 = n8225 & ~n8227 ;
  assign n8230 = n8228 | n8229 ;
  assign n8231 = n8106 | n8230 ;
  assign n8232 = n8223 | n8231 ;
  assign n8233 = n8106 & n8230 ;
  assign n8234 = ( n8223 & n8230 ) | ( n8223 & n8233 ) | ( n8230 & n8233 ) ;
  assign n8235 = n8232 & ~n8234 ;
  assign n8236 = n8222 | n8235 ;
  assign n8237 = n8207 & n8236 ;
  assign n8238 = n8219 & n8232 ;
  assign n8239 = n8221 | n8234 ;
  assign n8240 = n8238 & ~n8239 ;
  assign n8241 = ( n8106 & n8225 ) | ( n8106 & n8227 ) | ( n8225 & n8227 ) ;
  assign n8242 = n8225 | n8227 ;
  assign n8243 = ( n8223 & n8241 ) | ( n8223 & n8242 ) | ( n8241 & n8242 ) ;
  assign n8244 = ( n8191 & n8212 ) | ( n8191 & n8214 ) | ( n8212 & n8214 ) ;
  assign n8245 = n8212 | n8214 ;
  assign n8246 = ( n8210 & n8244 ) | ( n8210 & n8245 ) | ( n8244 & n8245 ) ;
  assign n8247 = ~n8243 & n8246 ;
  assign n8248 = n8243 & ~n8246 ;
  assign n8249 = n8247 | n8248 ;
  assign n8250 = n8240 | n8249 ;
  assign n8251 = n8237 | n8250 ;
  assign n8252 = n8236 | n8240 ;
  assign n8253 = ( n8207 & n8240 ) | ( n8207 & n8252 ) | ( n8240 & n8252 ) ;
  assign n8254 = n8249 & n8253 ;
  assign n8255 = n8251 & ~n8254 ;
  assign n8256 = ( x574 & x575 ) | ( x574 & x576 ) | ( x575 & x576 ) ;
  assign n8257 = ( x571 & x572 ) | ( x571 & x573 ) | ( x572 & x573 ) ;
  assign n8258 = n8256 & ~n8257 ;
  assign n8259 = ~n8256 & n8257 ;
  assign n8260 = n8258 | n8259 ;
  assign n8261 = ~x571 & x572 ;
  assign n8262 = x571 & ~x572 ;
  assign n8263 = n8261 | n8262 ;
  assign n8264 = ~x573 & n8263 ;
  assign n8265 = x573 & ~n8263 ;
  assign n8266 = n8264 | n8265 ;
  assign n8267 = ~x574 & x575 ;
  assign n8268 = x574 & ~x575 ;
  assign n8269 = n8267 | n8268 ;
  assign n8270 = ~x576 & n8269 ;
  assign n8271 = x576 & ~n8269 ;
  assign n8272 = n8270 | n8271 ;
  assign n8273 = n8266 & n8272 ;
  assign n8274 = n8260 & ~n8273 ;
  assign n8275 = ~n8260 & n8273 ;
  assign n8276 = n8274 | n8275 ;
  assign n8277 = n8266 & ~n8272 ;
  assign n8278 = ~n8266 & n8272 ;
  assign n8279 = n8277 | n8278 ;
  assign n8280 = ( n8256 & n8257 ) | ( n8256 & n8273 ) | ( n8257 & n8273 ) ;
  assign n8281 = n8279 & n8280 ;
  assign n8282 = n8276 & ~n8281 ;
  assign n8283 = n8276 & n8280 ;
  assign n8284 = ~x577 & x578 ;
  assign n8285 = x577 & ~x578 ;
  assign n8286 = n8284 | n8285 ;
  assign n8287 = ~x579 & n8286 ;
  assign n8288 = x579 & ~n8286 ;
  assign n8289 = n8287 | n8288 ;
  assign n8290 = ~x580 & x581 ;
  assign n8291 = x580 & ~x581 ;
  assign n8292 = n8290 | n8291 ;
  assign n8293 = ~x582 & n8292 ;
  assign n8294 = x582 & ~n8292 ;
  assign n8295 = n8293 | n8294 ;
  assign n8296 = n8289 & ~n8295 ;
  assign n8297 = ~n8289 & n8295 ;
  assign n8298 = n8296 | n8297 ;
  assign n8299 = ( x580 & x581 ) | ( x580 & x582 ) | ( x581 & x582 ) ;
  assign n8300 = ( x577 & x578 ) | ( x577 & x579 ) | ( x578 & x579 ) ;
  assign n8301 = n8289 & n8295 ;
  assign n8302 = ( n8299 & n8300 ) | ( n8299 & n8301 ) | ( n8300 & n8301 ) ;
  assign n8303 = n8298 & n8302 ;
  assign n8304 = n8283 | n8303 ;
  assign n8305 = n8299 & ~n8300 ;
  assign n8306 = ~n8299 & n8300 ;
  assign n8307 = n8305 | n8306 ;
  assign n8308 = ~n8301 & n8307 ;
  assign n8309 = n8301 & ~n8307 ;
  assign n8310 = n8308 | n8309 ;
  assign n8311 = n8302 & n8310 ;
  assign n8312 = n8279 & n8298 ;
  assign n8313 = n8310 & n8312 ;
  assign n8314 = ~n8311 & n8313 ;
  assign n8315 = ~n8304 & n8314 ;
  assign n8316 = n8282 & n8315 ;
  assign n8317 = ~n8311 & n8312 ;
  assign n8318 = ~n8303 & n8310 ;
  assign n8319 = n8283 & ~n8318 ;
  assign n8320 = ( n8317 & n8318 ) | ( n8317 & ~n8319 ) | ( n8318 & ~n8319 ) ;
  assign n8321 = ( n8282 & n8316 ) | ( n8282 & ~n8320 ) | ( n8316 & ~n8320 ) ;
  assign n8322 = n8298 & ~n8302 ;
  assign n8323 = ( n8298 & ~n8310 ) | ( n8298 & n8322 ) | ( ~n8310 & n8322 ) ;
  assign n8324 = n8279 & ~n8280 ;
  assign n8325 = ( ~n8276 & n8279 ) | ( ~n8276 & n8324 ) | ( n8279 & n8324 ) ;
  assign n8326 = ~n8323 & n8325 ;
  assign n8327 = n8323 & ~n8325 ;
  assign n8328 = n8326 | n8327 ;
  assign n8329 = ( x568 & x569 ) | ( x568 & x570 ) | ( x569 & x570 ) ;
  assign n8330 = ( x565 & x566 ) | ( x565 & x567 ) | ( x566 & x567 ) ;
  assign n8331 = n8329 & ~n8330 ;
  assign n8332 = ~n8329 & n8330 ;
  assign n8333 = n8331 | n8332 ;
  assign n8334 = ~x565 & x566 ;
  assign n8335 = x565 & ~x566 ;
  assign n8336 = n8334 | n8335 ;
  assign n8337 = ~x567 & n8336 ;
  assign n8338 = x567 & ~n8336 ;
  assign n8339 = n8337 | n8338 ;
  assign n8340 = ~x568 & x569 ;
  assign n8341 = x568 & ~x569 ;
  assign n8342 = n8340 | n8341 ;
  assign n8343 = ~x570 & n8342 ;
  assign n8344 = x570 & ~n8342 ;
  assign n8345 = n8343 | n8344 ;
  assign n8346 = n8339 & n8345 ;
  assign n8347 = n8333 & ~n8346 ;
  assign n8348 = ~n8333 & n8346 ;
  assign n8349 = n8347 | n8348 ;
  assign n8350 = n8339 & ~n8345 ;
  assign n8351 = ~n8339 & n8345 ;
  assign n8352 = n8350 | n8351 ;
  assign n8353 = ( n8329 & n8330 ) | ( n8329 & n8346 ) | ( n8330 & n8346 ) ;
  assign n8354 = n8352 & ~n8353 ;
  assign n8355 = ( ~n8349 & n8352 ) | ( ~n8349 & n8354 ) | ( n8352 & n8354 ) ;
  assign n8356 = ~x559 & x560 ;
  assign n8357 = x559 & ~x560 ;
  assign n8358 = n8356 | n8357 ;
  assign n8359 = ~x561 & n8358 ;
  assign n8360 = x561 & ~n8358 ;
  assign n8361 = n8359 | n8360 ;
  assign n8362 = ~x562 & x563 ;
  assign n8363 = x562 & ~x563 ;
  assign n8364 = n8362 | n8363 ;
  assign n8365 = ~x564 & n8364 ;
  assign n8366 = x564 & ~n8364 ;
  assign n8367 = n8365 | n8366 ;
  assign n8368 = n8361 & ~n8367 ;
  assign n8369 = ~n8361 & n8367 ;
  assign n8370 = n8368 | n8369 ;
  assign n8371 = ( x562 & x563 ) | ( x562 & x564 ) | ( x563 & x564 ) ;
  assign n8372 = ( x559 & x560 ) | ( x559 & x561 ) | ( x560 & x561 ) ;
  assign n8373 = n8371 & ~n8372 ;
  assign n8374 = ~n8371 & n8372 ;
  assign n8375 = n8373 | n8374 ;
  assign n8376 = n8361 & n8367 ;
  assign n8377 = n8375 & ~n8376 ;
  assign n8378 = ~n8375 & n8376 ;
  assign n8379 = n8377 | n8378 ;
  assign n8380 = ( n8371 & n8372 ) | ( n8371 & n8376 ) | ( n8372 & n8376 ) ;
  assign n8381 = n8370 & ~n8380 ;
  assign n8382 = ( n8370 & ~n8379 ) | ( n8370 & n8381 ) | ( ~n8379 & n8381 ) ;
  assign n8383 = ~n8355 & n8382 ;
  assign n8384 = n8355 & ~n8382 ;
  assign n8385 = n8383 | n8384 ;
  assign n8386 = n8328 & n8385 ;
  assign n8387 = ( n8282 & ~n8283 ) | ( n8282 & n8318 ) | ( ~n8283 & n8318 ) ;
  assign n8388 = n8282 & n8318 ;
  assign n8389 = ( n8317 & n8387 ) | ( n8317 & n8388 ) | ( n8387 & n8388 ) ;
  assign n8390 = n8320 & ~n8389 ;
  assign n8391 = n8386 | n8390 ;
  assign n8392 = n8321 | n8391 ;
  assign n8393 = n8379 & n8380 ;
  assign n8394 = n8352 & n8353 ;
  assign n8395 = n8393 | n8394 ;
  assign n8396 = n8349 & n8353 ;
  assign n8397 = n8352 & n8370 ;
  assign n8398 = n8349 & n8397 ;
  assign n8399 = ~n8396 & n8398 ;
  assign n8400 = ~n8395 & n8399 ;
  assign n8401 = n8370 & n8380 ;
  assign n8402 = n8379 & ~n8401 ;
  assign n8403 = ~n8400 & n8402 ;
  assign n8404 = ~n8396 & n8397 ;
  assign n8405 = n8349 & ~n8394 ;
  assign n8406 = ( n8393 & n8402 ) | ( n8393 & n8405 ) | ( n8402 & n8405 ) ;
  assign n8407 = n8402 | n8405 ;
  assign n8408 = ( ~n8404 & n8406 ) | ( ~n8404 & n8407 ) | ( n8406 & n8407 ) ;
  assign n8409 = n8393 | n8405 ;
  assign n8410 = n8404 & ~n8409 ;
  assign n8411 = ( ~n8405 & n8408 ) | ( ~n8405 & n8410 ) | ( n8408 & n8410 ) ;
  assign n8412 = ( ~n8403 & n8408 ) | ( ~n8403 & n8411 ) | ( n8408 & n8411 ) ;
  assign n8413 = n8392 & n8412 ;
  assign n8414 = n8386 & n8390 ;
  assign n8415 = ( n8321 & n8386 ) | ( n8321 & n8414 ) | ( n8386 & n8414 ) ;
  assign n8416 = n8413 | n8415 ;
  assign n8417 = n8393 & ~n8405 ;
  assign n8418 = ( n8404 & n8405 ) | ( n8404 & ~n8417 ) | ( n8405 & ~n8417 ) ;
  assign n8419 = n8402 & n8418 ;
  assign n8420 = ~n8370 & n8380 ;
  assign n8421 = ( ~n8379 & n8380 ) | ( ~n8379 & n8420 ) | ( n8380 & n8420 ) ;
  assign n8422 = ~n8352 & n8353 ;
  assign n8423 = ( ~n8349 & n8353 ) | ( ~n8349 & n8422 ) | ( n8353 & n8422 ) ;
  assign n8424 = ~n8421 & n8423 ;
  assign n8425 = n8421 & ~n8423 ;
  assign n8426 = n8424 | n8425 ;
  assign n8427 = n8400 | n8426 ;
  assign n8428 = n8419 | n8427 ;
  assign n8429 = n8400 & n8426 ;
  assign n8430 = ( n8419 & n8426 ) | ( n8419 & n8429 ) | ( n8426 & n8429 ) ;
  assign n8431 = n8428 & ~n8430 ;
  assign n8432 = n8282 & n8320 ;
  assign n8433 = ~n8279 & n8280 ;
  assign n8434 = ( ~n8276 & n8280 ) | ( ~n8276 & n8433 ) | ( n8280 & n8433 ) ;
  assign n8435 = ~n8298 & n8302 ;
  assign n8436 = ( n8302 & ~n8310 ) | ( n8302 & n8435 ) | ( ~n8310 & n8435 ) ;
  assign n8437 = ~n8434 & n8436 ;
  assign n8438 = n8434 & ~n8436 ;
  assign n8439 = n8437 | n8438 ;
  assign n8440 = n8315 | n8439 ;
  assign n8441 = n8432 | n8440 ;
  assign n8442 = n8315 & n8439 ;
  assign n8443 = ( n8432 & n8439 ) | ( n8432 & n8442 ) | ( n8439 & n8442 ) ;
  assign n8444 = n8441 & ~n8443 ;
  assign n8445 = n8431 | n8444 ;
  assign n8446 = n8416 & n8445 ;
  assign n8447 = n8428 & n8441 ;
  assign n8448 = n8430 | n8443 ;
  assign n8449 = n8447 & ~n8448 ;
  assign n8450 = ( n8315 & n8434 ) | ( n8315 & n8436 ) | ( n8434 & n8436 ) ;
  assign n8451 = n8434 | n8436 ;
  assign n8452 = ( n8432 & n8450 ) | ( n8432 & n8451 ) | ( n8450 & n8451 ) ;
  assign n8453 = ( n8400 & n8421 ) | ( n8400 & n8423 ) | ( n8421 & n8423 ) ;
  assign n8454 = n8421 | n8423 ;
  assign n8455 = ( n8419 & n8453 ) | ( n8419 & n8454 ) | ( n8453 & n8454 ) ;
  assign n8456 = ~n8452 & n8455 ;
  assign n8457 = n8452 & ~n8455 ;
  assign n8458 = n8456 | n8457 ;
  assign n8459 = n8449 | n8458 ;
  assign n8460 = n8446 | n8459 ;
  assign n8461 = n8445 | n8449 ;
  assign n8462 = ( n8416 & n8449 ) | ( n8416 & n8461 ) | ( n8449 & n8461 ) ;
  assign n8463 = n8458 & n8462 ;
  assign n8464 = n8460 & ~n8463 ;
  assign n8465 = n8255 | n8464 ;
  assign n8466 = n8183 & ~n8206 ;
  assign n8467 = n8203 & ~n8466 ;
  assign n8468 = n8119 & ~n8176 ;
  assign n8469 = ~n8119 & n8176 ;
  assign n8470 = n8468 | n8469 ;
  assign n8471 = n8328 & ~n8385 ;
  assign n8472 = ~n8328 & n8385 ;
  assign n8473 = n8471 | n8472 ;
  assign n8474 = n8470 & n8473 ;
  assign n8475 = ~n8177 & n8183 ;
  assign n8476 = n8183 & ~n8203 ;
  assign n8477 = n8112 | n8181 ;
  assign n8478 = n8203 | n8477 ;
  assign n8479 = ( n8475 & n8476 ) | ( n8475 & ~n8478 ) | ( n8476 & ~n8478 ) ;
  assign n8480 = n8474 | n8479 ;
  assign n8481 = n8467 | n8480 ;
  assign n8482 = n8321 | n8390 ;
  assign n8483 = ( n8386 & n8412 ) | ( n8386 & ~n8482 ) | ( n8412 & ~n8482 ) ;
  assign n8484 = ( ~n8412 & n8482 ) | ( ~n8412 & n8483 ) | ( n8482 & n8483 ) ;
  assign n8485 = ( ~n8386 & n8483 ) | ( ~n8386 & n8484 ) | ( n8483 & n8484 ) ;
  assign n8486 = n8481 & n8485 ;
  assign n8487 = n8467 | n8479 ;
  assign n8488 = n8474 & n8487 ;
  assign n8489 = ( n8415 & ~n8431 ) | ( n8415 & n8444 ) | ( ~n8431 & n8444 ) ;
  assign n8490 = n8431 & ~n8444 ;
  assign n8491 = ( n8413 & n8489 ) | ( n8413 & ~n8490 ) | ( n8489 & ~n8490 ) ;
  assign n8492 = ( ~n8416 & n8431 ) | ( ~n8416 & n8491 ) | ( n8431 & n8491 ) ;
  assign n8493 = ( ~n8444 & n8491 ) | ( ~n8444 & n8492 ) | ( n8491 & n8492 ) ;
  assign n8494 = ( n8206 & ~n8222 ) | ( n8206 & n8235 ) | ( ~n8222 & n8235 ) ;
  assign n8495 = n8222 & ~n8235 ;
  assign n8496 = ( n8204 & n8494 ) | ( n8204 & ~n8495 ) | ( n8494 & ~n8495 ) ;
  assign n8497 = ( ~n8207 & n8222 ) | ( ~n8207 & n8496 ) | ( n8222 & n8496 ) ;
  assign n8498 = ( ~n8235 & n8496 ) | ( ~n8235 & n8497 ) | ( n8496 & n8497 ) ;
  assign n8499 = ( n8488 & n8493 ) | ( n8488 & n8498 ) | ( n8493 & n8498 ) ;
  assign n8500 = n8493 | n8498 ;
  assign n8501 = ( n8486 & n8499 ) | ( n8486 & n8500 ) | ( n8499 & n8500 ) ;
  assign n8502 = n8465 & n8501 ;
  assign n8503 = n8251 & n8460 ;
  assign n8504 = n8254 | n8463 ;
  assign n8505 = n8503 & ~n8504 ;
  assign n8506 = n8452 & n8455 ;
  assign n8507 = n8452 | n8455 ;
  assign n8508 = n8506 | n8507 ;
  assign n8509 = ( n8462 & n8506 ) | ( n8462 & n8508 ) | ( n8506 & n8508 ) ;
  assign n8510 = n8243 & n8246 ;
  assign n8511 = n8243 | n8246 ;
  assign n8512 = n8510 | n8511 ;
  assign n8513 = ( n8253 & n8510 ) | ( n8253 & n8512 ) | ( n8510 & n8512 ) ;
  assign n8514 = n8509 & n8513 ;
  assign n8515 = n8513 & ~n8514 ;
  assign n8516 = ( n8509 & ~n8514 ) | ( n8509 & n8515 ) | ( ~n8514 & n8515 ) ;
  assign n8517 = n8505 | n8516 ;
  assign n8518 = n8502 | n8517 ;
  assign n8519 = n8502 | n8505 ;
  assign n8520 = n8516 & n8519 ;
  assign n8521 = n8518 & ~n8520 ;
  assign n8522 = ( x646 & x647 ) | ( x646 & x648 ) | ( x647 & x648 ) ;
  assign n8523 = ( x643 & x644 ) | ( x643 & x645 ) | ( x644 & x645 ) ;
  assign n8524 = n8522 & ~n8523 ;
  assign n8525 = ~n8522 & n8523 ;
  assign n8526 = n8524 | n8525 ;
  assign n8527 = ~x643 & x644 ;
  assign n8528 = x643 & ~x644 ;
  assign n8529 = n8527 | n8528 ;
  assign n8530 = ~x645 & n8529 ;
  assign n8531 = x645 & ~n8529 ;
  assign n8532 = n8530 | n8531 ;
  assign n8533 = ~x646 & x647 ;
  assign n8534 = x646 & ~x647 ;
  assign n8535 = n8533 | n8534 ;
  assign n8536 = ~x648 & n8535 ;
  assign n8537 = x648 & ~n8535 ;
  assign n8538 = n8536 | n8537 ;
  assign n8539 = n8532 & n8538 ;
  assign n8540 = n8526 & ~n8539 ;
  assign n8541 = ~n8526 & n8539 ;
  assign n8542 = n8540 | n8541 ;
  assign n8543 = n8532 & ~n8538 ;
  assign n8544 = ~n8532 & n8538 ;
  assign n8545 = n8543 | n8544 ;
  assign n8546 = ( n8522 & n8523 ) | ( n8522 & n8539 ) | ( n8523 & n8539 ) ;
  assign n8547 = n8545 & n8546 ;
  assign n8548 = n8542 & ~n8547 ;
  assign n8549 = n8542 & n8546 ;
  assign n8550 = ~x649 & x650 ;
  assign n8551 = x649 & ~x650 ;
  assign n8552 = n8550 | n8551 ;
  assign n8553 = ~x651 & n8552 ;
  assign n8554 = x651 & ~n8552 ;
  assign n8555 = n8553 | n8554 ;
  assign n8556 = ~x652 & x653 ;
  assign n8557 = x652 & ~x653 ;
  assign n8558 = n8556 | n8557 ;
  assign n8559 = ~x654 & n8558 ;
  assign n8560 = x654 & ~n8558 ;
  assign n8561 = n8559 | n8560 ;
  assign n8562 = n8555 & ~n8561 ;
  assign n8563 = ~n8555 & n8561 ;
  assign n8564 = n8562 | n8563 ;
  assign n8565 = ( x652 & x653 ) | ( x652 & x654 ) | ( x653 & x654 ) ;
  assign n8566 = ( x649 & x650 ) | ( x649 & x651 ) | ( x650 & x651 ) ;
  assign n8567 = n8555 & n8561 ;
  assign n8568 = ( n8565 & n8566 ) | ( n8565 & n8567 ) | ( n8566 & n8567 ) ;
  assign n8569 = n8564 & n8568 ;
  assign n8570 = n8549 | n8569 ;
  assign n8571 = n8565 & ~n8566 ;
  assign n8572 = ~n8565 & n8566 ;
  assign n8573 = n8571 | n8572 ;
  assign n8574 = ~n8567 & n8573 ;
  assign n8575 = n8567 & ~n8573 ;
  assign n8576 = n8574 | n8575 ;
  assign n8577 = n8568 & n8576 ;
  assign n8578 = n8545 & n8564 ;
  assign n8579 = n8576 & n8578 ;
  assign n8580 = ~n8577 & n8579 ;
  assign n8581 = ~n8570 & n8580 ;
  assign n8582 = n8548 & n8581 ;
  assign n8583 = ~n8577 & n8578 ;
  assign n8584 = ~n8569 & n8576 ;
  assign n8585 = n8549 & ~n8584 ;
  assign n8586 = ( n8583 & n8584 ) | ( n8583 & ~n8585 ) | ( n8584 & ~n8585 ) ;
  assign n8587 = ( n8548 & n8582 ) | ( n8548 & ~n8586 ) | ( n8582 & ~n8586 ) ;
  assign n8588 = n8564 & ~n8568 ;
  assign n8589 = ( n8564 & ~n8576 ) | ( n8564 & n8588 ) | ( ~n8576 & n8588 ) ;
  assign n8590 = n8545 & ~n8546 ;
  assign n8591 = ( ~n8542 & n8545 ) | ( ~n8542 & n8590 ) | ( n8545 & n8590 ) ;
  assign n8592 = ~n8589 & n8591 ;
  assign n8593 = n8589 & ~n8591 ;
  assign n8594 = n8592 | n8593 ;
  assign n8595 = ( x640 & x641 ) | ( x640 & x642 ) | ( x641 & x642 ) ;
  assign n8596 = ( x637 & x638 ) | ( x637 & x639 ) | ( x638 & x639 ) ;
  assign n8597 = n8595 & ~n8596 ;
  assign n8598 = ~n8595 & n8596 ;
  assign n8599 = n8597 | n8598 ;
  assign n8600 = ~x637 & x638 ;
  assign n8601 = x637 & ~x638 ;
  assign n8602 = n8600 | n8601 ;
  assign n8603 = ~x639 & n8602 ;
  assign n8604 = x639 & ~n8602 ;
  assign n8605 = n8603 | n8604 ;
  assign n8606 = ~x640 & x641 ;
  assign n8607 = x640 & ~x641 ;
  assign n8608 = n8606 | n8607 ;
  assign n8609 = ~x642 & n8608 ;
  assign n8610 = x642 & ~n8608 ;
  assign n8611 = n8609 | n8610 ;
  assign n8612 = n8605 & n8611 ;
  assign n8613 = n8599 & ~n8612 ;
  assign n8614 = ~n8599 & n8612 ;
  assign n8615 = n8613 | n8614 ;
  assign n8616 = n8605 & ~n8611 ;
  assign n8617 = ~n8605 & n8611 ;
  assign n8618 = n8616 | n8617 ;
  assign n8619 = ( n8595 & n8596 ) | ( n8595 & n8612 ) | ( n8596 & n8612 ) ;
  assign n8620 = n8618 & ~n8619 ;
  assign n8621 = ( ~n8615 & n8618 ) | ( ~n8615 & n8620 ) | ( n8618 & n8620 ) ;
  assign n8622 = ~x631 & x632 ;
  assign n8623 = x631 & ~x632 ;
  assign n8624 = n8622 | n8623 ;
  assign n8625 = ~x633 & n8624 ;
  assign n8626 = x633 & ~n8624 ;
  assign n8627 = n8625 | n8626 ;
  assign n8628 = ~x634 & x635 ;
  assign n8629 = x634 & ~x635 ;
  assign n8630 = n8628 | n8629 ;
  assign n8631 = ~x636 & n8630 ;
  assign n8632 = x636 & ~n8630 ;
  assign n8633 = n8631 | n8632 ;
  assign n8634 = n8627 & ~n8633 ;
  assign n8635 = ~n8627 & n8633 ;
  assign n8636 = n8634 | n8635 ;
  assign n8637 = ( x634 & x635 ) | ( x634 & x636 ) | ( x635 & x636 ) ;
  assign n8638 = ( x631 & x632 ) | ( x631 & x633 ) | ( x632 & x633 ) ;
  assign n8639 = n8637 & ~n8638 ;
  assign n8640 = ~n8637 & n8638 ;
  assign n8641 = n8639 | n8640 ;
  assign n8642 = n8627 & n8633 ;
  assign n8643 = n8641 & ~n8642 ;
  assign n8644 = ~n8641 & n8642 ;
  assign n8645 = n8643 | n8644 ;
  assign n8646 = ( n8637 & n8638 ) | ( n8637 & n8642 ) | ( n8638 & n8642 ) ;
  assign n8647 = n8636 & ~n8646 ;
  assign n8648 = ( n8636 & ~n8645 ) | ( n8636 & n8647 ) | ( ~n8645 & n8647 ) ;
  assign n8649 = ~n8621 & n8648 ;
  assign n8650 = n8621 & ~n8648 ;
  assign n8651 = n8649 | n8650 ;
  assign n8652 = n8594 & n8651 ;
  assign n8653 = ( n8548 & ~n8549 ) | ( n8548 & n8584 ) | ( ~n8549 & n8584 ) ;
  assign n8654 = n8548 & n8584 ;
  assign n8655 = ( n8583 & n8653 ) | ( n8583 & n8654 ) | ( n8653 & n8654 ) ;
  assign n8656 = n8586 & ~n8655 ;
  assign n8657 = n8652 | n8656 ;
  assign n8658 = n8587 | n8657 ;
  assign n8659 = n8645 & n8646 ;
  assign n8660 = n8618 & n8619 ;
  assign n8661 = n8659 | n8660 ;
  assign n8662 = n8615 & n8619 ;
  assign n8663 = n8618 & n8636 ;
  assign n8664 = n8615 & n8663 ;
  assign n8665 = ~n8662 & n8664 ;
  assign n8666 = ~n8661 & n8665 ;
  assign n8667 = n8636 & n8646 ;
  assign n8668 = n8645 & ~n8667 ;
  assign n8669 = ~n8666 & n8668 ;
  assign n8670 = ~n8662 & n8663 ;
  assign n8671 = n8615 & ~n8660 ;
  assign n8672 = ( n8659 & n8668 ) | ( n8659 & n8671 ) | ( n8668 & n8671 ) ;
  assign n8673 = n8668 | n8671 ;
  assign n8674 = ( ~n8670 & n8672 ) | ( ~n8670 & n8673 ) | ( n8672 & n8673 ) ;
  assign n8675 = n8659 | n8671 ;
  assign n8676 = n8670 & ~n8675 ;
  assign n8677 = ( ~n8671 & n8674 ) | ( ~n8671 & n8676 ) | ( n8674 & n8676 ) ;
  assign n8678 = ( ~n8669 & n8674 ) | ( ~n8669 & n8677 ) | ( n8674 & n8677 ) ;
  assign n8679 = n8658 & n8678 ;
  assign n8680 = n8652 & n8656 ;
  assign n8681 = ( n8587 & n8652 ) | ( n8587 & n8680 ) | ( n8652 & n8680 ) ;
  assign n8682 = n8679 | n8681 ;
  assign n8683 = n8659 & ~n8671 ;
  assign n8684 = ( n8670 & n8671 ) | ( n8670 & ~n8683 ) | ( n8671 & ~n8683 ) ;
  assign n8685 = n8668 & n8684 ;
  assign n8686 = ~n8636 & n8646 ;
  assign n8687 = ( ~n8645 & n8646 ) | ( ~n8645 & n8686 ) | ( n8646 & n8686 ) ;
  assign n8688 = ~n8618 & n8619 ;
  assign n8689 = ( ~n8615 & n8619 ) | ( ~n8615 & n8688 ) | ( n8619 & n8688 ) ;
  assign n8690 = ~n8687 & n8689 ;
  assign n8691 = n8687 & ~n8689 ;
  assign n8692 = n8690 | n8691 ;
  assign n8693 = n8666 | n8692 ;
  assign n8694 = n8685 | n8693 ;
  assign n8695 = n8666 & n8692 ;
  assign n8696 = ( n8685 & n8692 ) | ( n8685 & n8695 ) | ( n8692 & n8695 ) ;
  assign n8697 = n8694 & ~n8696 ;
  assign n8698 = n8548 & n8586 ;
  assign n8699 = ~n8545 & n8546 ;
  assign n8700 = ( ~n8542 & n8546 ) | ( ~n8542 & n8699 ) | ( n8546 & n8699 ) ;
  assign n8701 = ~n8564 & n8568 ;
  assign n8702 = ( n8568 & ~n8576 ) | ( n8568 & n8701 ) | ( ~n8576 & n8701 ) ;
  assign n8703 = ~n8700 & n8702 ;
  assign n8704 = n8700 & ~n8702 ;
  assign n8705 = n8703 | n8704 ;
  assign n8706 = n8581 | n8705 ;
  assign n8707 = n8698 | n8706 ;
  assign n8708 = n8581 & n8705 ;
  assign n8709 = ( n8698 & n8705 ) | ( n8698 & n8708 ) | ( n8705 & n8708 ) ;
  assign n8710 = n8707 & ~n8709 ;
  assign n8711 = n8697 | n8710 ;
  assign n8712 = n8682 & n8711 ;
  assign n8713 = n8694 & n8707 ;
  assign n8714 = n8696 | n8709 ;
  assign n8715 = n8713 & ~n8714 ;
  assign n8716 = ( n8581 & n8700 ) | ( n8581 & n8702 ) | ( n8700 & n8702 ) ;
  assign n8717 = n8700 | n8702 ;
  assign n8718 = ( n8698 & n8716 ) | ( n8698 & n8717 ) | ( n8716 & n8717 ) ;
  assign n8719 = ( n8666 & n8687 ) | ( n8666 & n8689 ) | ( n8687 & n8689 ) ;
  assign n8720 = n8687 | n8689 ;
  assign n8721 = ( n8685 & n8719 ) | ( n8685 & n8720 ) | ( n8719 & n8720 ) ;
  assign n8722 = ~n8718 & n8721 ;
  assign n8723 = n8718 & ~n8721 ;
  assign n8724 = n8722 | n8723 ;
  assign n8725 = n8715 | n8724 ;
  assign n8726 = n8712 | n8725 ;
  assign n8727 = n8711 | n8715 ;
  assign n8728 = ( n8682 & n8715 ) | ( n8682 & n8727 ) | ( n8715 & n8727 ) ;
  assign n8729 = n8724 & n8728 ;
  assign n8730 = n8726 & ~n8729 ;
  assign n8731 = ( x622 & x623 ) | ( x622 & x624 ) | ( x623 & x624 ) ;
  assign n8732 = ( x619 & x620 ) | ( x619 & x621 ) | ( x620 & x621 ) ;
  assign n8733 = n8731 & ~n8732 ;
  assign n8734 = ~n8731 & n8732 ;
  assign n8735 = n8733 | n8734 ;
  assign n8736 = ~x619 & x620 ;
  assign n8737 = x619 & ~x620 ;
  assign n8738 = n8736 | n8737 ;
  assign n8739 = ~x621 & n8738 ;
  assign n8740 = x621 & ~n8738 ;
  assign n8741 = n8739 | n8740 ;
  assign n8742 = ~x622 & x623 ;
  assign n8743 = x622 & ~x623 ;
  assign n8744 = n8742 | n8743 ;
  assign n8745 = ~x624 & n8744 ;
  assign n8746 = x624 & ~n8744 ;
  assign n8747 = n8745 | n8746 ;
  assign n8748 = n8741 & n8747 ;
  assign n8749 = n8735 & ~n8748 ;
  assign n8750 = ~n8735 & n8748 ;
  assign n8751 = n8749 | n8750 ;
  assign n8752 = n8741 & ~n8747 ;
  assign n8753 = ~n8741 & n8747 ;
  assign n8754 = n8752 | n8753 ;
  assign n8755 = ( n8731 & n8732 ) | ( n8731 & n8748 ) | ( n8732 & n8748 ) ;
  assign n8756 = n8754 & n8755 ;
  assign n8757 = n8751 & ~n8756 ;
  assign n8758 = n8751 & n8755 ;
  assign n8759 = ~x625 & x626 ;
  assign n8760 = x625 & ~x626 ;
  assign n8761 = n8759 | n8760 ;
  assign n8762 = ~x627 & n8761 ;
  assign n8763 = x627 & ~n8761 ;
  assign n8764 = n8762 | n8763 ;
  assign n8765 = ~x628 & x629 ;
  assign n8766 = x628 & ~x629 ;
  assign n8767 = n8765 | n8766 ;
  assign n8768 = ~x630 & n8767 ;
  assign n8769 = x630 & ~n8767 ;
  assign n8770 = n8768 | n8769 ;
  assign n8771 = n8764 & ~n8770 ;
  assign n8772 = ~n8764 & n8770 ;
  assign n8773 = n8771 | n8772 ;
  assign n8774 = ( x628 & x629 ) | ( x628 & x630 ) | ( x629 & x630 ) ;
  assign n8775 = ( x625 & x626 ) | ( x625 & x627 ) | ( x626 & x627 ) ;
  assign n8776 = n8764 & n8770 ;
  assign n8777 = ( n8774 & n8775 ) | ( n8774 & n8776 ) | ( n8775 & n8776 ) ;
  assign n8778 = n8773 & n8777 ;
  assign n8779 = n8758 | n8778 ;
  assign n8780 = n8774 & ~n8775 ;
  assign n8781 = ~n8774 & n8775 ;
  assign n8782 = n8780 | n8781 ;
  assign n8783 = ~n8776 & n8782 ;
  assign n8784 = n8776 & ~n8782 ;
  assign n8785 = n8783 | n8784 ;
  assign n8786 = n8777 & n8785 ;
  assign n8787 = n8754 & n8773 ;
  assign n8788 = n8785 & n8787 ;
  assign n8789 = ~n8786 & n8788 ;
  assign n8790 = ~n8779 & n8789 ;
  assign n8791 = n8757 & n8790 ;
  assign n8792 = ~n8786 & n8787 ;
  assign n8793 = ~n8778 & n8785 ;
  assign n8794 = n8758 & ~n8793 ;
  assign n8795 = ( n8792 & n8793 ) | ( n8792 & ~n8794 ) | ( n8793 & ~n8794 ) ;
  assign n8796 = ( n8757 & n8791 ) | ( n8757 & ~n8795 ) | ( n8791 & ~n8795 ) ;
  assign n8797 = n8773 & ~n8777 ;
  assign n8798 = ( n8773 & ~n8785 ) | ( n8773 & n8797 ) | ( ~n8785 & n8797 ) ;
  assign n8799 = n8754 & ~n8755 ;
  assign n8800 = ( ~n8751 & n8754 ) | ( ~n8751 & n8799 ) | ( n8754 & n8799 ) ;
  assign n8801 = ~n8798 & n8800 ;
  assign n8802 = n8798 & ~n8800 ;
  assign n8803 = n8801 | n8802 ;
  assign n8804 = ( x616 & x617 ) | ( x616 & x618 ) | ( x617 & x618 ) ;
  assign n8805 = ( x613 & x614 ) | ( x613 & x615 ) | ( x614 & x615 ) ;
  assign n8806 = n8804 & ~n8805 ;
  assign n8807 = ~n8804 & n8805 ;
  assign n8808 = n8806 | n8807 ;
  assign n8809 = ~x613 & x614 ;
  assign n8810 = x613 & ~x614 ;
  assign n8811 = n8809 | n8810 ;
  assign n8812 = ~x615 & n8811 ;
  assign n8813 = x615 & ~n8811 ;
  assign n8814 = n8812 | n8813 ;
  assign n8815 = ~x616 & x617 ;
  assign n8816 = x616 & ~x617 ;
  assign n8817 = n8815 | n8816 ;
  assign n8818 = ~x618 & n8817 ;
  assign n8819 = x618 & ~n8817 ;
  assign n8820 = n8818 | n8819 ;
  assign n8821 = n8814 & n8820 ;
  assign n8822 = n8808 & ~n8821 ;
  assign n8823 = ~n8808 & n8821 ;
  assign n8824 = n8822 | n8823 ;
  assign n8825 = n8814 & ~n8820 ;
  assign n8826 = ~n8814 & n8820 ;
  assign n8827 = n8825 | n8826 ;
  assign n8828 = ( n8804 & n8805 ) | ( n8804 & n8821 ) | ( n8805 & n8821 ) ;
  assign n8829 = n8827 & ~n8828 ;
  assign n8830 = ( ~n8824 & n8827 ) | ( ~n8824 & n8829 ) | ( n8827 & n8829 ) ;
  assign n8831 = ~x607 & x608 ;
  assign n8832 = x607 & ~x608 ;
  assign n8833 = n8831 | n8832 ;
  assign n8834 = ~x609 & n8833 ;
  assign n8835 = x609 & ~n8833 ;
  assign n8836 = n8834 | n8835 ;
  assign n8837 = ~x610 & x611 ;
  assign n8838 = x610 & ~x611 ;
  assign n8839 = n8837 | n8838 ;
  assign n8840 = ~x612 & n8839 ;
  assign n8841 = x612 & ~n8839 ;
  assign n8842 = n8840 | n8841 ;
  assign n8843 = n8836 & ~n8842 ;
  assign n8844 = ~n8836 & n8842 ;
  assign n8845 = n8843 | n8844 ;
  assign n8846 = ( x610 & x611 ) | ( x610 & x612 ) | ( x611 & x612 ) ;
  assign n8847 = ( x607 & x608 ) | ( x607 & x609 ) | ( x608 & x609 ) ;
  assign n8848 = n8846 & ~n8847 ;
  assign n8849 = ~n8846 & n8847 ;
  assign n8850 = n8848 | n8849 ;
  assign n8851 = n8836 & n8842 ;
  assign n8852 = n8850 & ~n8851 ;
  assign n8853 = ~n8850 & n8851 ;
  assign n8854 = n8852 | n8853 ;
  assign n8855 = ( n8846 & n8847 ) | ( n8846 & n8851 ) | ( n8847 & n8851 ) ;
  assign n8856 = n8845 & ~n8855 ;
  assign n8857 = ( n8845 & ~n8854 ) | ( n8845 & n8856 ) | ( ~n8854 & n8856 ) ;
  assign n8858 = ~n8830 & n8857 ;
  assign n8859 = n8830 & ~n8857 ;
  assign n8860 = n8858 | n8859 ;
  assign n8861 = n8803 & n8860 ;
  assign n8862 = ( n8757 & ~n8758 ) | ( n8757 & n8793 ) | ( ~n8758 & n8793 ) ;
  assign n8863 = n8757 & n8793 ;
  assign n8864 = ( n8792 & n8862 ) | ( n8792 & n8863 ) | ( n8862 & n8863 ) ;
  assign n8865 = n8795 & ~n8864 ;
  assign n8866 = n8861 | n8865 ;
  assign n8867 = n8796 | n8866 ;
  assign n8868 = n8854 & n8855 ;
  assign n8869 = n8827 & n8828 ;
  assign n8870 = n8868 | n8869 ;
  assign n8871 = n8824 & n8828 ;
  assign n8872 = n8827 & n8845 ;
  assign n8873 = n8824 & n8872 ;
  assign n8874 = ~n8871 & n8873 ;
  assign n8875 = ~n8870 & n8874 ;
  assign n8876 = n8845 & n8855 ;
  assign n8877 = n8854 & ~n8876 ;
  assign n8878 = ~n8875 & n8877 ;
  assign n8879 = ~n8871 & n8872 ;
  assign n8880 = n8824 & ~n8869 ;
  assign n8881 = ( n8868 & n8877 ) | ( n8868 & n8880 ) | ( n8877 & n8880 ) ;
  assign n8882 = n8877 | n8880 ;
  assign n8883 = ( ~n8879 & n8881 ) | ( ~n8879 & n8882 ) | ( n8881 & n8882 ) ;
  assign n8884 = n8868 | n8880 ;
  assign n8885 = n8879 & ~n8884 ;
  assign n8886 = ( ~n8880 & n8883 ) | ( ~n8880 & n8885 ) | ( n8883 & n8885 ) ;
  assign n8887 = ( ~n8878 & n8883 ) | ( ~n8878 & n8886 ) | ( n8883 & n8886 ) ;
  assign n8888 = n8867 & n8887 ;
  assign n8889 = n8861 & n8865 ;
  assign n8890 = ( n8796 & n8861 ) | ( n8796 & n8889 ) | ( n8861 & n8889 ) ;
  assign n8891 = n8888 | n8890 ;
  assign n8892 = n8868 & ~n8880 ;
  assign n8893 = ( n8879 & n8880 ) | ( n8879 & ~n8892 ) | ( n8880 & ~n8892 ) ;
  assign n8894 = n8877 & n8893 ;
  assign n8895 = ~n8845 & n8855 ;
  assign n8896 = ( ~n8854 & n8855 ) | ( ~n8854 & n8895 ) | ( n8855 & n8895 ) ;
  assign n8897 = ~n8827 & n8828 ;
  assign n8898 = ( ~n8824 & n8828 ) | ( ~n8824 & n8897 ) | ( n8828 & n8897 ) ;
  assign n8899 = ~n8896 & n8898 ;
  assign n8900 = n8896 & ~n8898 ;
  assign n8901 = n8899 | n8900 ;
  assign n8902 = n8875 | n8901 ;
  assign n8903 = n8894 | n8902 ;
  assign n8904 = n8875 & n8901 ;
  assign n8905 = ( n8894 & n8901 ) | ( n8894 & n8904 ) | ( n8901 & n8904 ) ;
  assign n8906 = n8903 & ~n8905 ;
  assign n8907 = n8757 & n8795 ;
  assign n8908 = ~n8754 & n8755 ;
  assign n8909 = ( ~n8751 & n8755 ) | ( ~n8751 & n8908 ) | ( n8755 & n8908 ) ;
  assign n8910 = ~n8773 & n8777 ;
  assign n8911 = ( n8777 & ~n8785 ) | ( n8777 & n8910 ) | ( ~n8785 & n8910 ) ;
  assign n8912 = ~n8909 & n8911 ;
  assign n8913 = n8909 & ~n8911 ;
  assign n8914 = n8912 | n8913 ;
  assign n8915 = n8790 | n8914 ;
  assign n8916 = n8907 | n8915 ;
  assign n8917 = n8790 & n8914 ;
  assign n8918 = ( n8907 & n8914 ) | ( n8907 & n8917 ) | ( n8914 & n8917 ) ;
  assign n8919 = n8916 & ~n8918 ;
  assign n8920 = n8906 | n8919 ;
  assign n8921 = n8891 & n8920 ;
  assign n8922 = n8903 & n8916 ;
  assign n8923 = n8905 | n8918 ;
  assign n8924 = n8922 & ~n8923 ;
  assign n8925 = ( n8790 & n8909 ) | ( n8790 & n8911 ) | ( n8909 & n8911 ) ;
  assign n8926 = n8909 | n8911 ;
  assign n8927 = ( n8907 & n8925 ) | ( n8907 & n8926 ) | ( n8925 & n8926 ) ;
  assign n8928 = ( n8875 & n8896 ) | ( n8875 & n8898 ) | ( n8896 & n8898 ) ;
  assign n8929 = n8896 | n8898 ;
  assign n8930 = ( n8894 & n8928 ) | ( n8894 & n8929 ) | ( n8928 & n8929 ) ;
  assign n8931 = ~n8927 & n8930 ;
  assign n8932 = n8927 & ~n8930 ;
  assign n8933 = n8931 | n8932 ;
  assign n8934 = n8924 | n8933 ;
  assign n8935 = n8921 | n8934 ;
  assign n8936 = n8920 | n8924 ;
  assign n8937 = ( n8891 & n8924 ) | ( n8891 & n8936 ) | ( n8924 & n8936 ) ;
  assign n8938 = n8933 & n8937 ;
  assign n8939 = n8935 & ~n8938 ;
  assign n8940 = n8730 | n8939 ;
  assign n8941 = n8658 & ~n8681 ;
  assign n8942 = n8678 & ~n8941 ;
  assign n8943 = n8594 & ~n8651 ;
  assign n8944 = ~n8594 & n8651 ;
  assign n8945 = n8943 | n8944 ;
  assign n8946 = n8803 & ~n8860 ;
  assign n8947 = ~n8803 & n8860 ;
  assign n8948 = n8946 | n8947 ;
  assign n8949 = n8945 & n8948 ;
  assign n8950 = ~n8652 & n8658 ;
  assign n8951 = n8658 & ~n8678 ;
  assign n8952 = n8587 | n8656 ;
  assign n8953 = n8678 | n8952 ;
  assign n8954 = ( n8950 & n8951 ) | ( n8950 & ~n8953 ) | ( n8951 & ~n8953 ) ;
  assign n8955 = n8949 | n8954 ;
  assign n8956 = n8942 | n8955 ;
  assign n8957 = n8796 | n8865 ;
  assign n8958 = ( n8861 & n8887 ) | ( n8861 & ~n8957 ) | ( n8887 & ~n8957 ) ;
  assign n8959 = ( ~n8887 & n8957 ) | ( ~n8887 & n8958 ) | ( n8957 & n8958 ) ;
  assign n8960 = ( ~n8861 & n8958 ) | ( ~n8861 & n8959 ) | ( n8958 & n8959 ) ;
  assign n8961 = n8956 & n8960 ;
  assign n8962 = n8942 | n8954 ;
  assign n8963 = n8949 & n8962 ;
  assign n8964 = ( n8890 & ~n8906 ) | ( n8890 & n8919 ) | ( ~n8906 & n8919 ) ;
  assign n8965 = n8906 & ~n8919 ;
  assign n8966 = ( n8888 & n8964 ) | ( n8888 & ~n8965 ) | ( n8964 & ~n8965 ) ;
  assign n8967 = ( ~n8891 & n8906 ) | ( ~n8891 & n8966 ) | ( n8906 & n8966 ) ;
  assign n8968 = ( ~n8919 & n8966 ) | ( ~n8919 & n8967 ) | ( n8966 & n8967 ) ;
  assign n8969 = ( n8681 & ~n8697 ) | ( n8681 & n8710 ) | ( ~n8697 & n8710 ) ;
  assign n8970 = n8697 & ~n8710 ;
  assign n8971 = ( n8679 & n8969 ) | ( n8679 & ~n8970 ) | ( n8969 & ~n8970 ) ;
  assign n8972 = ( ~n8682 & n8697 ) | ( ~n8682 & n8971 ) | ( n8697 & n8971 ) ;
  assign n8973 = ( ~n8710 & n8971 ) | ( ~n8710 & n8972 ) | ( n8971 & n8972 ) ;
  assign n8974 = ( n8963 & n8968 ) | ( n8963 & n8973 ) | ( n8968 & n8973 ) ;
  assign n8975 = n8968 | n8973 ;
  assign n8976 = ( n8961 & n8974 ) | ( n8961 & n8975 ) | ( n8974 & n8975 ) ;
  assign n8977 = n8940 & n8976 ;
  assign n8978 = n8726 & n8935 ;
  assign n8979 = n8729 | n8938 ;
  assign n8980 = n8978 & ~n8979 ;
  assign n8981 = n8927 & n8930 ;
  assign n8982 = n8927 | n8930 ;
  assign n8983 = n8981 | n8982 ;
  assign n8984 = ( n8937 & n8981 ) | ( n8937 & n8983 ) | ( n8981 & n8983 ) ;
  assign n8985 = n8718 & n8721 ;
  assign n8986 = n8718 | n8721 ;
  assign n8987 = n8985 | n8986 ;
  assign n8988 = ( n8728 & n8985 ) | ( n8728 & n8987 ) | ( n8985 & n8987 ) ;
  assign n8989 = n8984 & n8988 ;
  assign n8990 = n8988 & ~n8989 ;
  assign n8991 = ( n8984 & ~n8989 ) | ( n8984 & n8990 ) | ( ~n8989 & n8990 ) ;
  assign n8992 = n8980 | n8991 ;
  assign n8993 = n8977 | n8992 ;
  assign n8994 = n8977 | n8980 ;
  assign n8995 = n8991 & n8994 ;
  assign n8996 = n8993 & ~n8995 ;
  assign n8997 = n8521 | n8996 ;
  assign n8998 = ( ~n8730 & n8939 ) | ( ~n8730 & n8976 ) | ( n8939 & n8976 ) ;
  assign n8999 = ( n8730 & ~n8976 ) | ( n8730 & n8998 ) | ( ~n8976 & n8998 ) ;
  assign n9000 = ( ~n8939 & n8998 ) | ( ~n8939 & n8999 ) | ( n8998 & n8999 ) ;
  assign n9001 = ( ~n8255 & n8464 ) | ( ~n8255 & n8501 ) | ( n8464 & n8501 ) ;
  assign n9002 = ( n8255 & ~n8501 ) | ( n8255 & n9001 ) | ( ~n8501 & n9001 ) ;
  assign n9003 = ( ~n8464 & n9001 ) | ( ~n8464 & n9002 ) | ( n9001 & n9002 ) ;
  assign n9004 = ~n8474 & n8487 ;
  assign n9005 = n8474 & ~n8479 ;
  assign n9006 = ~n8467 & n9005 ;
  assign n9007 = ~n8485 & n9006 ;
  assign n9008 = ( ~n8485 & n9004 ) | ( ~n8485 & n9007 ) | ( n9004 & n9007 ) ;
  assign n9009 = n8486 & ~n8488 ;
  assign n9010 = ( n8485 & n9008 ) | ( n8485 & ~n9009 ) | ( n9008 & ~n9009 ) ;
  assign n9011 = n8945 & ~n8948 ;
  assign n9012 = ~n8945 & n8948 ;
  assign n9013 = n9011 | n9012 ;
  assign n9014 = n8470 & ~n8473 ;
  assign n9015 = ~n8470 & n8473 ;
  assign n9016 = n9014 | n9015 ;
  assign n9017 = n9013 & n9016 ;
  assign n9018 = ~n8956 & n8960 ;
  assign n9019 = ( n8960 & n8963 ) | ( n8960 & n9018 ) | ( n8963 & n9018 ) ;
  assign n9020 = ~n8949 & n8962 ;
  assign n9021 = n8949 & ~n8954 ;
  assign n9022 = ~n8942 & n9021 ;
  assign n9023 = ~n8960 & n9022 ;
  assign n9024 = ( ~n8960 & n9020 ) | ( ~n8960 & n9023 ) | ( n9020 & n9023 ) ;
  assign n9025 = n9019 | n9024 ;
  assign n9026 = n9017 | n9025 ;
  assign n9027 = n9010 & n9026 ;
  assign n9028 = n9017 & n9025 ;
  assign n9030 = ( n8488 & ~n8493 ) | ( n8488 & n8498 ) | ( ~n8493 & n8498 ) ;
  assign n9031 = n8493 & ~n8498 ;
  assign n9032 = ( n8486 & n9030 ) | ( n8486 & ~n9031 ) | ( n9030 & ~n9031 ) ;
  assign n9029 = n8486 | n8488 ;
  assign n9033 = ( n8493 & ~n9029 ) | ( n8493 & n9032 ) | ( ~n9029 & n9032 ) ;
  assign n9034 = ( ~n8498 & n9032 ) | ( ~n8498 & n9033 ) | ( n9032 & n9033 ) ;
  assign n9036 = ( n8963 & ~n8968 ) | ( n8963 & n8973 ) | ( ~n8968 & n8973 ) ;
  assign n9037 = n8968 & ~n8973 ;
  assign n9038 = ( n8961 & n9036 ) | ( n8961 & ~n9037 ) | ( n9036 & ~n9037 ) ;
  assign n9035 = n8961 | n8963 ;
  assign n9039 = ( n8968 & ~n9035 ) | ( n8968 & n9038 ) | ( ~n9035 & n9038 ) ;
  assign n9040 = ( ~n8973 & n9038 ) | ( ~n8973 & n9039 ) | ( n9038 & n9039 ) ;
  assign n9041 = ( n9028 & n9034 ) | ( n9028 & n9040 ) | ( n9034 & n9040 ) ;
  assign n9042 = n9034 | n9040 ;
  assign n9043 = ( n9027 & n9041 ) | ( n9027 & n9042 ) | ( n9041 & n9042 ) ;
  assign n9044 = ( n9000 & n9003 ) | ( n9000 & n9043 ) | ( n9003 & n9043 ) ;
  assign n9045 = n8997 & n9044 ;
  assign n9046 = n8518 & n8993 ;
  assign n9047 = n8520 | n8995 ;
  assign n9048 = n9046 & ~n9047 ;
  assign n9057 = n8253 & n8511 ;
  assign n9058 = n8455 | n8510 ;
  assign n9059 = n8452 | n8510 ;
  assign n9060 = ( n8462 & n9058 ) | ( n8462 & n9059 ) | ( n9058 & n9059 ) ;
  assign n9061 = n9057 | n9060 ;
  assign n9062 = n8514 | n9061 ;
  assign n9063 = ( n8505 & n8514 ) | ( n8505 & n9062 ) | ( n8514 & n9062 ) ;
  assign n9064 = n8514 | n9062 ;
  assign n9065 = ( n8502 & n9063 ) | ( n8502 & n9064 ) | ( n9063 & n9064 ) ;
  assign n9049 = n8728 & n8986 ;
  assign n9050 = n8930 | n8985 ;
  assign n9051 = n8927 | n8985 ;
  assign n9052 = ( n8937 & n9050 ) | ( n8937 & n9051 ) | ( n9050 & n9051 ) ;
  assign n9053 = n9049 | n9052 ;
  assign n9054 = n8980 & n9053 ;
  assign n9055 = ( n8977 & n9053 ) | ( n8977 & n9054 ) | ( n9053 & n9054 ) ;
  assign n9056 = n8989 | n9055 ;
  assign n9066 = n9056 & n9065 ;
  assign n9067 = n9056 & ~n9066 ;
  assign n9068 = ( n9065 & ~n9066 ) | ( n9065 & n9067 ) | ( ~n9066 & n9067 ) ;
  assign n9069 = n9048 | n9068 ;
  assign n9070 = n9045 | n9069 ;
  assign n9071 = n9045 | n9048 ;
  assign n9072 = n9068 & n9071 ;
  assign n9073 = n9070 & ~n9072 ;
  assign n9074 = ( x502 & x503 ) | ( x502 & x504 ) | ( x503 & x504 ) ;
  assign n9075 = ( x499 & x500 ) | ( x499 & x501 ) | ( x500 & x501 ) ;
  assign n9076 = n9074 & ~n9075 ;
  assign n9077 = ~n9074 & n9075 ;
  assign n9078 = n9076 | n9077 ;
  assign n9079 = ~x499 & x500 ;
  assign n9080 = x499 & ~x500 ;
  assign n9081 = n9079 | n9080 ;
  assign n9082 = ~x501 & n9081 ;
  assign n9083 = x501 & ~n9081 ;
  assign n9084 = n9082 | n9083 ;
  assign n9085 = ~x502 & x503 ;
  assign n9086 = x502 & ~x503 ;
  assign n9087 = n9085 | n9086 ;
  assign n9088 = ~x504 & n9087 ;
  assign n9089 = x504 & ~n9087 ;
  assign n9090 = n9088 | n9089 ;
  assign n9091 = n9084 & n9090 ;
  assign n9092 = n9078 & ~n9091 ;
  assign n9093 = ~n9078 & n9091 ;
  assign n9094 = n9092 | n9093 ;
  assign n9095 = n9084 & ~n9090 ;
  assign n9096 = ~n9084 & n9090 ;
  assign n9097 = n9095 | n9096 ;
  assign n9098 = ( n9074 & n9075 ) | ( n9074 & n9091 ) | ( n9075 & n9091 ) ;
  assign n9099 = n9097 & n9098 ;
  assign n9100 = n9094 & ~n9099 ;
  assign n9101 = n9094 & n9098 ;
  assign n9102 = ~x505 & x506 ;
  assign n9103 = x505 & ~x506 ;
  assign n9104 = n9102 | n9103 ;
  assign n9105 = ~x507 & n9104 ;
  assign n9106 = x507 & ~n9104 ;
  assign n9107 = n9105 | n9106 ;
  assign n9108 = ~x508 & x509 ;
  assign n9109 = x508 & ~x509 ;
  assign n9110 = n9108 | n9109 ;
  assign n9111 = ~x510 & n9110 ;
  assign n9112 = x510 & ~n9110 ;
  assign n9113 = n9111 | n9112 ;
  assign n9114 = n9107 & ~n9113 ;
  assign n9115 = ~n9107 & n9113 ;
  assign n9116 = n9114 | n9115 ;
  assign n9117 = ( x508 & x509 ) | ( x508 & x510 ) | ( x509 & x510 ) ;
  assign n9118 = ( x505 & x506 ) | ( x505 & x507 ) | ( x506 & x507 ) ;
  assign n9119 = n9107 & n9113 ;
  assign n9120 = ( n9117 & n9118 ) | ( n9117 & n9119 ) | ( n9118 & n9119 ) ;
  assign n9121 = n9116 & n9120 ;
  assign n9122 = n9101 | n9121 ;
  assign n9123 = n9117 & ~n9118 ;
  assign n9124 = ~n9117 & n9118 ;
  assign n9125 = n9123 | n9124 ;
  assign n9126 = ~n9119 & n9125 ;
  assign n9127 = n9119 & ~n9125 ;
  assign n9128 = n9126 | n9127 ;
  assign n9129 = n9120 & n9128 ;
  assign n9130 = n9097 & n9116 ;
  assign n9131 = n9128 & n9130 ;
  assign n9132 = ~n9129 & n9131 ;
  assign n9133 = ~n9122 & n9132 ;
  assign n9134 = n9100 & n9133 ;
  assign n9135 = ~n9129 & n9130 ;
  assign n9136 = ~n9121 & n9128 ;
  assign n9137 = n9101 & ~n9136 ;
  assign n9138 = ( n9135 & n9136 ) | ( n9135 & ~n9137 ) | ( n9136 & ~n9137 ) ;
  assign n9139 = ( n9100 & n9134 ) | ( n9100 & ~n9138 ) | ( n9134 & ~n9138 ) ;
  assign n9140 = n9116 & ~n9120 ;
  assign n9141 = ( n9116 & ~n9128 ) | ( n9116 & n9140 ) | ( ~n9128 & n9140 ) ;
  assign n9142 = n9097 & ~n9098 ;
  assign n9143 = ( ~n9094 & n9097 ) | ( ~n9094 & n9142 ) | ( n9097 & n9142 ) ;
  assign n9144 = ~n9141 & n9143 ;
  assign n9145 = n9141 & ~n9143 ;
  assign n9146 = n9144 | n9145 ;
  assign n9147 = ( x496 & x497 ) | ( x496 & x498 ) | ( x497 & x498 ) ;
  assign n9148 = ( x493 & x494 ) | ( x493 & x495 ) | ( x494 & x495 ) ;
  assign n9149 = n9147 & ~n9148 ;
  assign n9150 = ~n9147 & n9148 ;
  assign n9151 = n9149 | n9150 ;
  assign n9152 = ~x493 & x494 ;
  assign n9153 = x493 & ~x494 ;
  assign n9154 = n9152 | n9153 ;
  assign n9155 = ~x495 & n9154 ;
  assign n9156 = x495 & ~n9154 ;
  assign n9157 = n9155 | n9156 ;
  assign n9158 = ~x496 & x497 ;
  assign n9159 = x496 & ~x497 ;
  assign n9160 = n9158 | n9159 ;
  assign n9161 = ~x498 & n9160 ;
  assign n9162 = x498 & ~n9160 ;
  assign n9163 = n9161 | n9162 ;
  assign n9164 = n9157 & n9163 ;
  assign n9165 = n9151 & ~n9164 ;
  assign n9166 = ~n9151 & n9164 ;
  assign n9167 = n9165 | n9166 ;
  assign n9168 = n9157 & ~n9163 ;
  assign n9169 = ~n9157 & n9163 ;
  assign n9170 = n9168 | n9169 ;
  assign n9171 = ( n9147 & n9148 ) | ( n9147 & n9164 ) | ( n9148 & n9164 ) ;
  assign n9172 = n9170 & ~n9171 ;
  assign n9173 = ( ~n9167 & n9170 ) | ( ~n9167 & n9172 ) | ( n9170 & n9172 ) ;
  assign n9174 = ~x487 & x488 ;
  assign n9175 = x487 & ~x488 ;
  assign n9176 = n9174 | n9175 ;
  assign n9177 = ~x489 & n9176 ;
  assign n9178 = x489 & ~n9176 ;
  assign n9179 = n9177 | n9178 ;
  assign n9180 = ~x490 & x491 ;
  assign n9181 = x490 & ~x491 ;
  assign n9182 = n9180 | n9181 ;
  assign n9183 = ~x492 & n9182 ;
  assign n9184 = x492 & ~n9182 ;
  assign n9185 = n9183 | n9184 ;
  assign n9186 = n9179 & ~n9185 ;
  assign n9187 = ~n9179 & n9185 ;
  assign n9188 = n9186 | n9187 ;
  assign n9189 = ( x490 & x491 ) | ( x490 & x492 ) | ( x491 & x492 ) ;
  assign n9190 = ( x487 & x488 ) | ( x487 & x489 ) | ( x488 & x489 ) ;
  assign n9191 = n9189 & ~n9190 ;
  assign n9192 = ~n9189 & n9190 ;
  assign n9193 = n9191 | n9192 ;
  assign n9194 = n9179 & n9185 ;
  assign n9195 = n9193 & ~n9194 ;
  assign n9196 = ~n9193 & n9194 ;
  assign n9197 = n9195 | n9196 ;
  assign n9198 = ( n9189 & n9190 ) | ( n9189 & n9194 ) | ( n9190 & n9194 ) ;
  assign n9199 = n9188 & ~n9198 ;
  assign n9200 = ( n9188 & ~n9197 ) | ( n9188 & n9199 ) | ( ~n9197 & n9199 ) ;
  assign n9201 = ~n9173 & n9200 ;
  assign n9202 = n9173 & ~n9200 ;
  assign n9203 = n9201 | n9202 ;
  assign n9204 = n9146 & n9203 ;
  assign n9205 = ( n9100 & ~n9101 ) | ( n9100 & n9136 ) | ( ~n9101 & n9136 ) ;
  assign n9206 = n9100 & n9136 ;
  assign n9207 = ( n9135 & n9205 ) | ( n9135 & n9206 ) | ( n9205 & n9206 ) ;
  assign n9208 = n9138 & ~n9207 ;
  assign n9209 = n9204 | n9208 ;
  assign n9210 = n9139 | n9209 ;
  assign n9211 = n9197 & n9198 ;
  assign n9212 = n9170 & n9171 ;
  assign n9213 = n9211 | n9212 ;
  assign n9214 = n9167 & n9171 ;
  assign n9215 = n9170 & n9188 ;
  assign n9216 = n9167 & n9215 ;
  assign n9217 = ~n9214 & n9216 ;
  assign n9218 = ~n9213 & n9217 ;
  assign n9219 = n9188 & n9198 ;
  assign n9220 = n9197 & ~n9219 ;
  assign n9221 = ~n9218 & n9220 ;
  assign n9222 = ~n9214 & n9215 ;
  assign n9223 = n9167 & ~n9212 ;
  assign n9224 = ( n9211 & n9220 ) | ( n9211 & n9223 ) | ( n9220 & n9223 ) ;
  assign n9225 = n9220 | n9223 ;
  assign n9226 = ( ~n9222 & n9224 ) | ( ~n9222 & n9225 ) | ( n9224 & n9225 ) ;
  assign n9227 = n9211 | n9223 ;
  assign n9228 = n9222 & ~n9227 ;
  assign n9229 = ( ~n9223 & n9226 ) | ( ~n9223 & n9228 ) | ( n9226 & n9228 ) ;
  assign n9230 = ( ~n9221 & n9226 ) | ( ~n9221 & n9229 ) | ( n9226 & n9229 ) ;
  assign n9231 = n9210 & n9230 ;
  assign n9232 = n9204 & n9208 ;
  assign n9233 = ( n9139 & n9204 ) | ( n9139 & n9232 ) | ( n9204 & n9232 ) ;
  assign n9234 = n9231 | n9233 ;
  assign n9235 = n9211 & ~n9223 ;
  assign n9236 = ( n9222 & n9223 ) | ( n9222 & ~n9235 ) | ( n9223 & ~n9235 ) ;
  assign n9237 = n9220 & n9236 ;
  assign n9238 = ~n9188 & n9198 ;
  assign n9239 = ( ~n9197 & n9198 ) | ( ~n9197 & n9238 ) | ( n9198 & n9238 ) ;
  assign n9240 = ~n9170 & n9171 ;
  assign n9241 = ( ~n9167 & n9171 ) | ( ~n9167 & n9240 ) | ( n9171 & n9240 ) ;
  assign n9242 = ~n9239 & n9241 ;
  assign n9243 = n9239 & ~n9241 ;
  assign n9244 = n9242 | n9243 ;
  assign n9245 = n9218 | n9244 ;
  assign n9246 = n9237 | n9245 ;
  assign n9247 = n9218 & n9244 ;
  assign n9248 = ( n9237 & n9244 ) | ( n9237 & n9247 ) | ( n9244 & n9247 ) ;
  assign n9249 = n9246 & ~n9248 ;
  assign n9250 = n9100 & n9138 ;
  assign n9251 = ~n9097 & n9098 ;
  assign n9252 = ( ~n9094 & n9098 ) | ( ~n9094 & n9251 ) | ( n9098 & n9251 ) ;
  assign n9253 = ~n9116 & n9120 ;
  assign n9254 = ( n9120 & ~n9128 ) | ( n9120 & n9253 ) | ( ~n9128 & n9253 ) ;
  assign n9255 = ~n9252 & n9254 ;
  assign n9256 = n9252 & ~n9254 ;
  assign n9257 = n9255 | n9256 ;
  assign n9258 = n9133 | n9257 ;
  assign n9259 = n9250 | n9258 ;
  assign n9260 = n9133 & n9257 ;
  assign n9261 = ( n9250 & n9257 ) | ( n9250 & n9260 ) | ( n9257 & n9260 ) ;
  assign n9262 = n9259 & ~n9261 ;
  assign n9263 = n9249 | n9262 ;
  assign n9264 = n9234 & n9263 ;
  assign n9265 = n9246 & n9259 ;
  assign n9266 = n9248 | n9261 ;
  assign n9267 = n9265 & ~n9266 ;
  assign n9268 = ( n9133 & n9252 ) | ( n9133 & n9254 ) | ( n9252 & n9254 ) ;
  assign n9269 = n9252 | n9254 ;
  assign n9270 = ( n9250 & n9268 ) | ( n9250 & n9269 ) | ( n9268 & n9269 ) ;
  assign n9271 = ( n9218 & n9239 ) | ( n9218 & n9241 ) | ( n9239 & n9241 ) ;
  assign n9272 = n9239 | n9241 ;
  assign n9273 = ( n9237 & n9271 ) | ( n9237 & n9272 ) | ( n9271 & n9272 ) ;
  assign n9274 = ~n9270 & n9273 ;
  assign n9275 = n9270 & ~n9273 ;
  assign n9276 = n9274 | n9275 ;
  assign n9277 = n9267 | n9276 ;
  assign n9278 = n9264 | n9277 ;
  assign n9279 = n9263 | n9267 ;
  assign n9280 = ( n9234 & n9267 ) | ( n9234 & n9279 ) | ( n9267 & n9279 ) ;
  assign n9281 = n9276 & n9280 ;
  assign n9282 = n9278 & ~n9281 ;
  assign n9283 = ( x478 & x479 ) | ( x478 & x480 ) | ( x479 & x480 ) ;
  assign n9284 = ( x475 & x476 ) | ( x475 & x477 ) | ( x476 & x477 ) ;
  assign n9285 = n9283 & ~n9284 ;
  assign n9286 = ~n9283 & n9284 ;
  assign n9287 = n9285 | n9286 ;
  assign n9288 = ~x475 & x476 ;
  assign n9289 = x475 & ~x476 ;
  assign n9290 = n9288 | n9289 ;
  assign n9291 = ~x477 & n9290 ;
  assign n9292 = x477 & ~n9290 ;
  assign n9293 = n9291 | n9292 ;
  assign n9294 = ~x478 & x479 ;
  assign n9295 = x478 & ~x479 ;
  assign n9296 = n9294 | n9295 ;
  assign n9297 = ~x480 & n9296 ;
  assign n9298 = x480 & ~n9296 ;
  assign n9299 = n9297 | n9298 ;
  assign n9300 = n9293 & n9299 ;
  assign n9301 = n9287 & ~n9300 ;
  assign n9302 = ~n9287 & n9300 ;
  assign n9303 = n9301 | n9302 ;
  assign n9304 = n9293 & ~n9299 ;
  assign n9305 = ~n9293 & n9299 ;
  assign n9306 = n9304 | n9305 ;
  assign n9307 = ( n9283 & n9284 ) | ( n9283 & n9300 ) | ( n9284 & n9300 ) ;
  assign n9308 = n9306 & n9307 ;
  assign n9309 = n9303 & ~n9308 ;
  assign n9310 = n9303 & n9307 ;
  assign n9311 = ~x481 & x482 ;
  assign n9312 = x481 & ~x482 ;
  assign n9313 = n9311 | n9312 ;
  assign n9314 = ~x483 & n9313 ;
  assign n9315 = x483 & ~n9313 ;
  assign n9316 = n9314 | n9315 ;
  assign n9317 = ~x484 & x485 ;
  assign n9318 = x484 & ~x485 ;
  assign n9319 = n9317 | n9318 ;
  assign n9320 = ~x486 & n9319 ;
  assign n9321 = x486 & ~n9319 ;
  assign n9322 = n9320 | n9321 ;
  assign n9323 = n9316 & ~n9322 ;
  assign n9324 = ~n9316 & n9322 ;
  assign n9325 = n9323 | n9324 ;
  assign n9326 = ( x484 & x485 ) | ( x484 & x486 ) | ( x485 & x486 ) ;
  assign n9327 = ( x481 & x482 ) | ( x481 & x483 ) | ( x482 & x483 ) ;
  assign n9328 = n9316 & n9322 ;
  assign n9329 = ( n9326 & n9327 ) | ( n9326 & n9328 ) | ( n9327 & n9328 ) ;
  assign n9330 = n9325 & n9329 ;
  assign n9331 = n9310 | n9330 ;
  assign n9332 = n9326 & ~n9327 ;
  assign n9333 = ~n9326 & n9327 ;
  assign n9334 = n9332 | n9333 ;
  assign n9335 = ~n9328 & n9334 ;
  assign n9336 = n9328 & ~n9334 ;
  assign n9337 = n9335 | n9336 ;
  assign n9338 = n9329 & n9337 ;
  assign n9339 = n9306 & n9325 ;
  assign n9340 = n9337 & n9339 ;
  assign n9341 = ~n9338 & n9340 ;
  assign n9342 = ~n9331 & n9341 ;
  assign n9343 = n9309 & n9342 ;
  assign n9344 = ~n9338 & n9339 ;
  assign n9345 = ~n9330 & n9337 ;
  assign n9346 = n9310 & ~n9345 ;
  assign n9347 = ( n9344 & n9345 ) | ( n9344 & ~n9346 ) | ( n9345 & ~n9346 ) ;
  assign n9348 = ( n9309 & n9343 ) | ( n9309 & ~n9347 ) | ( n9343 & ~n9347 ) ;
  assign n9349 = ( x472 & x473 ) | ( x472 & x474 ) | ( x473 & x474 ) ;
  assign n9350 = ( x469 & x470 ) | ( x469 & x471 ) | ( x470 & x471 ) ;
  assign n9351 = n9349 & ~n9350 ;
  assign n9352 = ~n9349 & n9350 ;
  assign n9353 = n9351 | n9352 ;
  assign n9354 = ~x469 & x470 ;
  assign n9355 = x469 & ~x470 ;
  assign n9356 = n9354 | n9355 ;
  assign n9357 = ~x471 & n9356 ;
  assign n9358 = x471 & ~n9356 ;
  assign n9359 = n9357 | n9358 ;
  assign n9360 = ~x472 & x473 ;
  assign n9361 = x472 & ~x473 ;
  assign n9362 = n9360 | n9361 ;
  assign n9363 = ~x474 & n9362 ;
  assign n9364 = x474 & ~n9362 ;
  assign n9365 = n9363 | n9364 ;
  assign n9366 = n9359 & n9365 ;
  assign n9367 = n9353 & ~n9366 ;
  assign n9368 = ~n9353 & n9366 ;
  assign n9369 = n9367 | n9368 ;
  assign n9370 = n9359 & ~n9365 ;
  assign n9371 = ~n9359 & n9365 ;
  assign n9372 = n9370 | n9371 ;
  assign n9373 = ( n9349 & n9350 ) | ( n9349 & n9366 ) | ( n9350 & n9366 ) ;
  assign n9374 = n9372 & ~n9373 ;
  assign n9375 = ( ~n9369 & n9372 ) | ( ~n9369 & n9374 ) | ( n9372 & n9374 ) ;
  assign n9376 = ~x466 & x467 ;
  assign n9377 = x466 & ~x467 ;
  assign n9378 = n9376 | n9377 ;
  assign n9379 = ~x468 & n9378 ;
  assign n9380 = x468 & ~n9378 ;
  assign n9381 = n9379 | n9380 ;
  assign n9382 = ~x463 & x464 ;
  assign n9383 = x463 & ~x464 ;
  assign n9384 = n9382 | n9383 ;
  assign n9385 = ~x465 & n9384 ;
  assign n9386 = x465 & ~n9384 ;
  assign n9387 = n9385 | n9386 ;
  assign n9388 = n9381 & ~n9387 ;
  assign n9389 = ~n9381 & n9387 ;
  assign n9390 = n9388 | n9389 ;
  assign n9391 = n9381 & n9387 ;
  assign n9392 = ( x466 & x467 ) | ( x466 & x468 ) | ( x467 & x468 ) ;
  assign n9393 = ( x463 & x464 ) | ( x463 & x465 ) | ( x464 & x465 ) ;
  assign n9394 = ~n9392 & n9393 ;
  assign n9395 = n9392 & ~n9393 ;
  assign n9396 = n9394 | n9395 ;
  assign n9397 = ~n9391 & n9396 ;
  assign n9398 = n9391 & ~n9396 ;
  assign n9399 = n9397 | n9398 ;
  assign n9400 = ( n9391 & n9392 ) | ( n9391 & n9393 ) | ( n9392 & n9393 ) ;
  assign n9401 = n9390 & ~n9400 ;
  assign n9402 = ( n9390 & ~n9399 ) | ( n9390 & n9401 ) | ( ~n9399 & n9401 ) ;
  assign n9403 = ~n9375 & n9402 ;
  assign n9404 = n9375 & ~n9402 ;
  assign n9405 = n9403 | n9404 ;
  assign n9406 = n9325 & ~n9329 ;
  assign n9407 = ( n9325 & ~n9337 ) | ( n9325 & n9406 ) | ( ~n9337 & n9406 ) ;
  assign n9408 = n9306 & ~n9307 ;
  assign n9409 = ( ~n9303 & n9306 ) | ( ~n9303 & n9408 ) | ( n9306 & n9408 ) ;
  assign n9410 = ~n9407 & n9409 ;
  assign n9411 = n9407 & ~n9409 ;
  assign n9412 = n9410 | n9411 ;
  assign n9413 = n9405 & n9412 ;
  assign n9414 = ( n9309 & ~n9310 ) | ( n9309 & n9345 ) | ( ~n9310 & n9345 ) ;
  assign n9415 = n9309 & n9345 ;
  assign n9416 = ( n9344 & n9414 ) | ( n9344 & n9415 ) | ( n9414 & n9415 ) ;
  assign n9417 = n9347 & ~n9416 ;
  assign n9418 = n9413 | n9417 ;
  assign n9419 = n9348 | n9418 ;
  assign n9420 = n9399 & n9400 ;
  assign n9421 = n9372 & n9373 ;
  assign n9422 = n9420 | n9421 ;
  assign n9423 = n9369 & n9373 ;
  assign n9424 = n9372 & n9390 ;
  assign n9425 = n9369 & n9424 ;
  assign n9426 = ~n9423 & n9425 ;
  assign n9427 = ~n9422 & n9426 ;
  assign n9428 = n9390 & n9400 ;
  assign n9429 = n9399 & ~n9428 ;
  assign n9430 = ~n9427 & n9429 ;
  assign n9431 = ~n9423 & n9424 ;
  assign n9432 = n9369 & ~n9421 ;
  assign n9433 = ( n9420 & n9429 ) | ( n9420 & n9432 ) | ( n9429 & n9432 ) ;
  assign n9434 = n9429 | n9432 ;
  assign n9435 = ( ~n9431 & n9433 ) | ( ~n9431 & n9434 ) | ( n9433 & n9434 ) ;
  assign n9436 = n9420 | n9432 ;
  assign n9437 = n9431 & ~n9436 ;
  assign n9438 = ( ~n9432 & n9435 ) | ( ~n9432 & n9437 ) | ( n9435 & n9437 ) ;
  assign n9439 = ( ~n9430 & n9435 ) | ( ~n9430 & n9438 ) | ( n9435 & n9438 ) ;
  assign n9440 = n9419 & n9439 ;
  assign n9441 = n9413 & n9417 ;
  assign n9442 = ( n9348 & n9413 ) | ( n9348 & n9441 ) | ( n9413 & n9441 ) ;
  assign n9443 = n9440 | n9442 ;
  assign n9444 = n9420 & ~n9432 ;
  assign n9445 = ( n9431 & n9432 ) | ( n9431 & ~n9444 ) | ( n9432 & ~n9444 ) ;
  assign n9446 = n9429 & n9445 ;
  assign n9447 = ~n9390 & n9400 ;
  assign n9448 = ( ~n9399 & n9400 ) | ( ~n9399 & n9447 ) | ( n9400 & n9447 ) ;
  assign n9449 = ~n9372 & n9373 ;
  assign n9450 = ( ~n9369 & n9373 ) | ( ~n9369 & n9449 ) | ( n9373 & n9449 ) ;
  assign n9451 = ~n9448 & n9450 ;
  assign n9452 = n9448 & ~n9450 ;
  assign n9453 = n9451 | n9452 ;
  assign n9454 = n9427 | n9453 ;
  assign n9455 = n9446 | n9454 ;
  assign n9456 = n9427 & n9453 ;
  assign n9457 = ( n9446 & n9453 ) | ( n9446 & n9456 ) | ( n9453 & n9456 ) ;
  assign n9458 = n9455 & ~n9457 ;
  assign n9459 = n9309 & n9347 ;
  assign n9460 = ~n9306 & n9307 ;
  assign n9461 = ( ~n9303 & n9307 ) | ( ~n9303 & n9460 ) | ( n9307 & n9460 ) ;
  assign n9462 = ~n9325 & n9329 ;
  assign n9463 = ( n9329 & ~n9337 ) | ( n9329 & n9462 ) | ( ~n9337 & n9462 ) ;
  assign n9464 = ~n9461 & n9463 ;
  assign n9465 = n9461 & ~n9463 ;
  assign n9466 = n9464 | n9465 ;
  assign n9467 = n9342 | n9466 ;
  assign n9468 = n9459 | n9467 ;
  assign n9469 = n9342 & n9466 ;
  assign n9470 = ( n9459 & n9466 ) | ( n9459 & n9469 ) | ( n9466 & n9469 ) ;
  assign n9471 = n9468 & ~n9470 ;
  assign n9472 = n9458 | n9471 ;
  assign n9473 = n9443 & n9472 ;
  assign n9474 = n9455 & n9468 ;
  assign n9475 = n9457 | n9470 ;
  assign n9476 = n9474 & ~n9475 ;
  assign n9477 = ( n9342 & n9461 ) | ( n9342 & n9463 ) | ( n9461 & n9463 ) ;
  assign n9478 = n9461 | n9463 ;
  assign n9479 = ( n9459 & n9477 ) | ( n9459 & n9478 ) | ( n9477 & n9478 ) ;
  assign n9480 = ( n9427 & n9448 ) | ( n9427 & n9450 ) | ( n9448 & n9450 ) ;
  assign n9481 = n9448 | n9450 ;
  assign n9482 = ( n9446 & n9480 ) | ( n9446 & n9481 ) | ( n9480 & n9481 ) ;
  assign n9483 = ~n9479 & n9482 ;
  assign n9484 = n9479 & ~n9482 ;
  assign n9485 = n9483 | n9484 ;
  assign n9486 = n9476 | n9485 ;
  assign n9487 = n9473 | n9486 ;
  assign n9488 = n9472 | n9476 ;
  assign n9489 = ( n9443 & n9476 ) | ( n9443 & n9488 ) | ( n9476 & n9488 ) ;
  assign n9490 = n9485 & n9489 ;
  assign n9491 = n9487 & ~n9490 ;
  assign n9492 = n9282 | n9491 ;
  assign n9493 = n9210 & ~n9233 ;
  assign n9494 = n9230 & ~n9493 ;
  assign n9495 = n9405 & ~n9412 ;
  assign n9496 = ~n9405 & n9412 ;
  assign n9497 = n9495 | n9496 ;
  assign n9498 = n9146 & ~n9203 ;
  assign n9499 = ~n9146 & n9203 ;
  assign n9500 = n9498 | n9499 ;
  assign n9501 = n9497 & n9500 ;
  assign n9502 = ~n9204 & n9210 ;
  assign n9503 = n9210 & ~n9230 ;
  assign n9504 = n9139 | n9208 ;
  assign n9505 = n9230 | n9504 ;
  assign n9506 = ( n9502 & n9503 ) | ( n9502 & ~n9505 ) | ( n9503 & ~n9505 ) ;
  assign n9507 = n9501 | n9506 ;
  assign n9508 = n9494 | n9507 ;
  assign n9509 = n9348 | n9417 ;
  assign n9510 = ( n9413 & n9439 ) | ( n9413 & ~n9509 ) | ( n9439 & ~n9509 ) ;
  assign n9511 = ( ~n9439 & n9509 ) | ( ~n9439 & n9510 ) | ( n9509 & n9510 ) ;
  assign n9512 = ( ~n9413 & n9510 ) | ( ~n9413 & n9511 ) | ( n9510 & n9511 ) ;
  assign n9513 = n9508 & n9512 ;
  assign n9514 = n9494 | n9506 ;
  assign n9515 = n9501 & n9514 ;
  assign n9516 = ( n9442 & ~n9458 ) | ( n9442 & n9471 ) | ( ~n9458 & n9471 ) ;
  assign n9517 = n9458 & ~n9471 ;
  assign n9518 = ( n9440 & n9516 ) | ( n9440 & ~n9517 ) | ( n9516 & ~n9517 ) ;
  assign n9519 = ( ~n9443 & n9458 ) | ( ~n9443 & n9518 ) | ( n9458 & n9518 ) ;
  assign n9520 = ( ~n9471 & n9518 ) | ( ~n9471 & n9519 ) | ( n9518 & n9519 ) ;
  assign n9521 = ( n9233 & ~n9249 ) | ( n9233 & n9262 ) | ( ~n9249 & n9262 ) ;
  assign n9522 = n9249 & ~n9262 ;
  assign n9523 = ( n9231 & n9521 ) | ( n9231 & ~n9522 ) | ( n9521 & ~n9522 ) ;
  assign n9524 = ( ~n9234 & n9249 ) | ( ~n9234 & n9523 ) | ( n9249 & n9523 ) ;
  assign n9525 = ( ~n9262 & n9523 ) | ( ~n9262 & n9524 ) | ( n9523 & n9524 ) ;
  assign n9526 = ( n9515 & n9520 ) | ( n9515 & n9525 ) | ( n9520 & n9525 ) ;
  assign n9527 = n9520 | n9525 ;
  assign n9528 = ( n9513 & n9526 ) | ( n9513 & n9527 ) | ( n9526 & n9527 ) ;
  assign n9529 = n9492 & n9528 ;
  assign n9530 = n9278 & n9487 ;
  assign n9531 = n9281 | n9490 ;
  assign n9532 = n9530 & ~n9531 ;
  assign n9533 = n9479 & n9482 ;
  assign n9534 = n9479 | n9482 ;
  assign n9535 = n9533 | n9534 ;
  assign n9536 = ( n9489 & n9533 ) | ( n9489 & n9535 ) | ( n9533 & n9535 ) ;
  assign n9537 = n9270 & n9273 ;
  assign n9538 = n9270 | n9273 ;
  assign n9539 = n9537 | n9538 ;
  assign n9540 = ( n9280 & n9537 ) | ( n9280 & n9539 ) | ( n9537 & n9539 ) ;
  assign n9541 = n9536 & n9540 ;
  assign n9542 = n9540 & ~n9541 ;
  assign n9543 = ( n9536 & ~n9541 ) | ( n9536 & n9542 ) | ( ~n9541 & n9542 ) ;
  assign n9544 = n9532 | n9543 ;
  assign n9545 = n9529 | n9544 ;
  assign n9546 = n9529 | n9532 ;
  assign n9547 = n9543 & n9546 ;
  assign n9548 = n9545 & ~n9547 ;
  assign n9549 = ( x550 & x551 ) | ( x550 & x552 ) | ( x551 & x552 ) ;
  assign n9550 = ( x547 & x548 ) | ( x547 & x549 ) | ( x548 & x549 ) ;
  assign n9551 = n9549 & ~n9550 ;
  assign n9552 = ~n9549 & n9550 ;
  assign n9553 = n9551 | n9552 ;
  assign n9554 = ~x547 & x548 ;
  assign n9555 = x547 & ~x548 ;
  assign n9556 = n9554 | n9555 ;
  assign n9557 = ~x549 & n9556 ;
  assign n9558 = x549 & ~n9556 ;
  assign n9559 = n9557 | n9558 ;
  assign n9560 = ~x550 & x551 ;
  assign n9561 = x550 & ~x551 ;
  assign n9562 = n9560 | n9561 ;
  assign n9563 = ~x552 & n9562 ;
  assign n9564 = x552 & ~n9562 ;
  assign n9565 = n9563 | n9564 ;
  assign n9566 = n9559 & n9565 ;
  assign n9567 = n9553 & ~n9566 ;
  assign n9568 = ~n9553 & n9566 ;
  assign n9569 = n9567 | n9568 ;
  assign n9570 = n9559 & ~n9565 ;
  assign n9571 = ~n9559 & n9565 ;
  assign n9572 = n9570 | n9571 ;
  assign n9573 = ( n9549 & n9550 ) | ( n9549 & n9566 ) | ( n9550 & n9566 ) ;
  assign n9574 = n9572 & n9573 ;
  assign n9575 = n9569 & ~n9574 ;
  assign n9576 = n9569 & n9573 ;
  assign n9577 = ~x553 & x554 ;
  assign n9578 = x553 & ~x554 ;
  assign n9579 = n9577 | n9578 ;
  assign n9580 = ~x555 & n9579 ;
  assign n9581 = x555 & ~n9579 ;
  assign n9582 = n9580 | n9581 ;
  assign n9583 = ~x556 & x557 ;
  assign n9584 = x556 & ~x557 ;
  assign n9585 = n9583 | n9584 ;
  assign n9586 = ~x558 & n9585 ;
  assign n9587 = x558 & ~n9585 ;
  assign n9588 = n9586 | n9587 ;
  assign n9589 = n9582 & ~n9588 ;
  assign n9590 = ~n9582 & n9588 ;
  assign n9591 = n9589 | n9590 ;
  assign n9592 = ( x556 & x557 ) | ( x556 & x558 ) | ( x557 & x558 ) ;
  assign n9593 = ( x553 & x554 ) | ( x553 & x555 ) | ( x554 & x555 ) ;
  assign n9594 = n9582 & n9588 ;
  assign n9595 = ( n9592 & n9593 ) | ( n9592 & n9594 ) | ( n9593 & n9594 ) ;
  assign n9596 = n9591 & n9595 ;
  assign n9597 = n9576 | n9596 ;
  assign n9598 = n9592 & ~n9593 ;
  assign n9599 = ~n9592 & n9593 ;
  assign n9600 = n9598 | n9599 ;
  assign n9601 = ~n9594 & n9600 ;
  assign n9602 = n9594 & ~n9600 ;
  assign n9603 = n9601 | n9602 ;
  assign n9604 = n9595 & n9603 ;
  assign n9605 = n9572 & n9591 ;
  assign n9606 = n9603 & n9605 ;
  assign n9607 = ~n9604 & n9606 ;
  assign n9608 = ~n9597 & n9607 ;
  assign n9609 = n9575 & n9608 ;
  assign n9610 = ~n9604 & n9605 ;
  assign n9611 = ~n9596 & n9603 ;
  assign n9612 = n9576 & ~n9611 ;
  assign n9613 = ( n9610 & n9611 ) | ( n9610 & ~n9612 ) | ( n9611 & ~n9612 ) ;
  assign n9614 = ( n9575 & n9609 ) | ( n9575 & ~n9613 ) | ( n9609 & ~n9613 ) ;
  assign n9615 = n9591 & ~n9595 ;
  assign n9616 = ( n9591 & ~n9603 ) | ( n9591 & n9615 ) | ( ~n9603 & n9615 ) ;
  assign n9617 = n9572 & ~n9573 ;
  assign n9618 = ( ~n9569 & n9572 ) | ( ~n9569 & n9617 ) | ( n9572 & n9617 ) ;
  assign n9619 = ~n9616 & n9618 ;
  assign n9620 = n9616 & ~n9618 ;
  assign n9621 = n9619 | n9620 ;
  assign n9622 = ( x544 & x545 ) | ( x544 & x546 ) | ( x545 & x546 ) ;
  assign n9623 = ( x541 & x542 ) | ( x541 & x543 ) | ( x542 & x543 ) ;
  assign n9624 = n9622 & ~n9623 ;
  assign n9625 = ~n9622 & n9623 ;
  assign n9626 = n9624 | n9625 ;
  assign n9627 = ~x541 & x542 ;
  assign n9628 = x541 & ~x542 ;
  assign n9629 = n9627 | n9628 ;
  assign n9630 = ~x543 & n9629 ;
  assign n9631 = x543 & ~n9629 ;
  assign n9632 = n9630 | n9631 ;
  assign n9633 = ~x544 & x545 ;
  assign n9634 = x544 & ~x545 ;
  assign n9635 = n9633 | n9634 ;
  assign n9636 = ~x546 & n9635 ;
  assign n9637 = x546 & ~n9635 ;
  assign n9638 = n9636 | n9637 ;
  assign n9639 = n9632 & n9638 ;
  assign n9640 = n9626 & ~n9639 ;
  assign n9641 = ~n9626 & n9639 ;
  assign n9642 = n9640 | n9641 ;
  assign n9643 = n9632 & ~n9638 ;
  assign n9644 = ~n9632 & n9638 ;
  assign n9645 = n9643 | n9644 ;
  assign n9646 = ( n9622 & n9623 ) | ( n9622 & n9639 ) | ( n9623 & n9639 ) ;
  assign n9647 = n9645 & ~n9646 ;
  assign n9648 = ( ~n9642 & n9645 ) | ( ~n9642 & n9647 ) | ( n9645 & n9647 ) ;
  assign n9649 = ~x535 & x536 ;
  assign n9650 = x535 & ~x536 ;
  assign n9651 = n9649 | n9650 ;
  assign n9652 = ~x537 & n9651 ;
  assign n9653 = x537 & ~n9651 ;
  assign n9654 = n9652 | n9653 ;
  assign n9655 = ~x538 & x539 ;
  assign n9656 = x538 & ~x539 ;
  assign n9657 = n9655 | n9656 ;
  assign n9658 = ~x540 & n9657 ;
  assign n9659 = x540 & ~n9657 ;
  assign n9660 = n9658 | n9659 ;
  assign n9661 = n9654 & ~n9660 ;
  assign n9662 = ~n9654 & n9660 ;
  assign n9663 = n9661 | n9662 ;
  assign n9664 = ( x538 & x539 ) | ( x538 & x540 ) | ( x539 & x540 ) ;
  assign n9665 = ( x535 & x536 ) | ( x535 & x537 ) | ( x536 & x537 ) ;
  assign n9666 = n9664 & ~n9665 ;
  assign n9667 = ~n9664 & n9665 ;
  assign n9668 = n9666 | n9667 ;
  assign n9669 = n9654 & n9660 ;
  assign n9670 = n9668 & ~n9669 ;
  assign n9671 = ~n9668 & n9669 ;
  assign n9672 = n9670 | n9671 ;
  assign n9673 = ( n9664 & n9665 ) | ( n9664 & n9669 ) | ( n9665 & n9669 ) ;
  assign n9674 = n9663 & ~n9673 ;
  assign n9675 = ( n9663 & ~n9672 ) | ( n9663 & n9674 ) | ( ~n9672 & n9674 ) ;
  assign n9676 = ~n9648 & n9675 ;
  assign n9677 = n9648 & ~n9675 ;
  assign n9678 = n9676 | n9677 ;
  assign n9679 = n9621 & n9678 ;
  assign n9680 = ( n9575 & ~n9576 ) | ( n9575 & n9611 ) | ( ~n9576 & n9611 ) ;
  assign n9681 = n9575 & n9611 ;
  assign n9682 = ( n9610 & n9680 ) | ( n9610 & n9681 ) | ( n9680 & n9681 ) ;
  assign n9683 = n9613 & ~n9682 ;
  assign n9684 = n9679 | n9683 ;
  assign n9685 = n9614 | n9684 ;
  assign n9686 = n9672 & n9673 ;
  assign n9687 = n9645 & n9646 ;
  assign n9688 = n9686 | n9687 ;
  assign n9689 = n9642 & n9646 ;
  assign n9690 = n9645 & n9663 ;
  assign n9691 = n9642 & n9690 ;
  assign n9692 = ~n9689 & n9691 ;
  assign n9693 = ~n9688 & n9692 ;
  assign n9694 = n9663 & n9673 ;
  assign n9695 = n9672 & ~n9694 ;
  assign n9696 = ~n9693 & n9695 ;
  assign n9697 = ~n9689 & n9690 ;
  assign n9698 = n9642 & ~n9687 ;
  assign n9699 = ( n9686 & n9695 ) | ( n9686 & n9698 ) | ( n9695 & n9698 ) ;
  assign n9700 = n9695 | n9698 ;
  assign n9701 = ( ~n9697 & n9699 ) | ( ~n9697 & n9700 ) | ( n9699 & n9700 ) ;
  assign n9702 = n9686 | n9698 ;
  assign n9703 = n9697 & ~n9702 ;
  assign n9704 = ( ~n9698 & n9701 ) | ( ~n9698 & n9703 ) | ( n9701 & n9703 ) ;
  assign n9705 = ( ~n9696 & n9701 ) | ( ~n9696 & n9704 ) | ( n9701 & n9704 ) ;
  assign n9706 = n9685 & n9705 ;
  assign n9707 = n9679 & n9683 ;
  assign n9708 = ( n9614 & n9679 ) | ( n9614 & n9707 ) | ( n9679 & n9707 ) ;
  assign n9709 = n9706 | n9708 ;
  assign n9710 = n9686 & ~n9698 ;
  assign n9711 = ( n9697 & n9698 ) | ( n9697 & ~n9710 ) | ( n9698 & ~n9710 ) ;
  assign n9712 = n9695 & n9711 ;
  assign n9713 = ~n9663 & n9673 ;
  assign n9714 = ( ~n9672 & n9673 ) | ( ~n9672 & n9713 ) | ( n9673 & n9713 ) ;
  assign n9715 = ~n9645 & n9646 ;
  assign n9716 = ( ~n9642 & n9646 ) | ( ~n9642 & n9715 ) | ( n9646 & n9715 ) ;
  assign n9717 = ~n9714 & n9716 ;
  assign n9718 = n9714 & ~n9716 ;
  assign n9719 = n9717 | n9718 ;
  assign n9720 = n9693 | n9719 ;
  assign n9721 = n9712 | n9720 ;
  assign n9722 = n9693 & n9719 ;
  assign n9723 = ( n9712 & n9719 ) | ( n9712 & n9722 ) | ( n9719 & n9722 ) ;
  assign n9724 = n9721 & ~n9723 ;
  assign n9725 = n9575 & n9613 ;
  assign n9726 = ~n9572 & n9573 ;
  assign n9727 = ( ~n9569 & n9573 ) | ( ~n9569 & n9726 ) | ( n9573 & n9726 ) ;
  assign n9728 = ~n9591 & n9595 ;
  assign n9729 = ( n9595 & ~n9603 ) | ( n9595 & n9728 ) | ( ~n9603 & n9728 ) ;
  assign n9730 = ~n9727 & n9729 ;
  assign n9731 = n9727 & ~n9729 ;
  assign n9732 = n9730 | n9731 ;
  assign n9733 = n9608 | n9732 ;
  assign n9734 = n9725 | n9733 ;
  assign n9735 = n9608 & n9732 ;
  assign n9736 = ( n9725 & n9732 ) | ( n9725 & n9735 ) | ( n9732 & n9735 ) ;
  assign n9737 = n9734 & ~n9736 ;
  assign n9738 = n9724 | n9737 ;
  assign n9739 = n9709 & n9738 ;
  assign n9740 = n9721 & n9734 ;
  assign n9741 = n9723 | n9736 ;
  assign n9742 = n9740 & ~n9741 ;
  assign n9743 = ( n9608 & n9727 ) | ( n9608 & n9729 ) | ( n9727 & n9729 ) ;
  assign n9744 = n9727 | n9729 ;
  assign n9745 = ( n9725 & n9743 ) | ( n9725 & n9744 ) | ( n9743 & n9744 ) ;
  assign n9746 = ( n9693 & n9714 ) | ( n9693 & n9716 ) | ( n9714 & n9716 ) ;
  assign n9747 = n9714 | n9716 ;
  assign n9748 = ( n9712 & n9746 ) | ( n9712 & n9747 ) | ( n9746 & n9747 ) ;
  assign n9749 = ~n9745 & n9748 ;
  assign n9750 = n9745 & ~n9748 ;
  assign n9751 = n9749 | n9750 ;
  assign n9752 = n9742 | n9751 ;
  assign n9753 = n9739 | n9752 ;
  assign n9754 = n9738 | n9742 ;
  assign n9755 = ( n9709 & n9742 ) | ( n9709 & n9754 ) | ( n9742 & n9754 ) ;
  assign n9756 = n9751 & n9755 ;
  assign n9757 = n9753 & ~n9756 ;
  assign n9758 = ( x526 & x527 ) | ( x526 & x528 ) | ( x527 & x528 ) ;
  assign n9759 = ( x523 & x524 ) | ( x523 & x525 ) | ( x524 & x525 ) ;
  assign n9760 = n9758 & ~n9759 ;
  assign n9761 = ~n9758 & n9759 ;
  assign n9762 = n9760 | n9761 ;
  assign n9763 = ~x523 & x524 ;
  assign n9764 = x523 & ~x524 ;
  assign n9765 = n9763 | n9764 ;
  assign n9766 = ~x525 & n9765 ;
  assign n9767 = x525 & ~n9765 ;
  assign n9768 = n9766 | n9767 ;
  assign n9769 = ~x526 & x527 ;
  assign n9770 = x526 & ~x527 ;
  assign n9771 = n9769 | n9770 ;
  assign n9772 = ~x528 & n9771 ;
  assign n9773 = x528 & ~n9771 ;
  assign n9774 = n9772 | n9773 ;
  assign n9775 = n9768 & n9774 ;
  assign n9776 = n9762 & ~n9775 ;
  assign n9777 = ~n9762 & n9775 ;
  assign n9778 = n9776 | n9777 ;
  assign n9779 = n9768 & ~n9774 ;
  assign n9780 = ~n9768 & n9774 ;
  assign n9781 = n9779 | n9780 ;
  assign n9782 = ( n9758 & n9759 ) | ( n9758 & n9775 ) | ( n9759 & n9775 ) ;
  assign n9783 = n9781 & n9782 ;
  assign n9784 = n9778 & ~n9783 ;
  assign n9785 = n9778 & n9782 ;
  assign n9786 = ~x529 & x530 ;
  assign n9787 = x529 & ~x530 ;
  assign n9788 = n9786 | n9787 ;
  assign n9789 = ~x531 & n9788 ;
  assign n9790 = x531 & ~n9788 ;
  assign n9791 = n9789 | n9790 ;
  assign n9792 = ~x532 & x533 ;
  assign n9793 = x532 & ~x533 ;
  assign n9794 = n9792 | n9793 ;
  assign n9795 = ~x534 & n9794 ;
  assign n9796 = x534 & ~n9794 ;
  assign n9797 = n9795 | n9796 ;
  assign n9798 = n9791 & ~n9797 ;
  assign n9799 = ~n9791 & n9797 ;
  assign n9800 = n9798 | n9799 ;
  assign n9801 = ( x532 & x533 ) | ( x532 & x534 ) | ( x533 & x534 ) ;
  assign n9802 = ( x529 & x530 ) | ( x529 & x531 ) | ( x530 & x531 ) ;
  assign n9803 = n9791 & n9797 ;
  assign n9804 = ( n9801 & n9802 ) | ( n9801 & n9803 ) | ( n9802 & n9803 ) ;
  assign n9805 = n9800 & n9804 ;
  assign n9806 = n9785 | n9805 ;
  assign n9807 = n9801 & ~n9802 ;
  assign n9808 = ~n9801 & n9802 ;
  assign n9809 = n9807 | n9808 ;
  assign n9810 = ~n9803 & n9809 ;
  assign n9811 = n9803 & ~n9809 ;
  assign n9812 = n9810 | n9811 ;
  assign n9813 = n9804 & n9812 ;
  assign n9814 = n9781 & n9800 ;
  assign n9815 = n9812 & n9814 ;
  assign n9816 = ~n9813 & n9815 ;
  assign n9817 = ~n9806 & n9816 ;
  assign n9818 = n9784 & n9817 ;
  assign n9819 = ~n9813 & n9814 ;
  assign n9820 = ~n9805 & n9812 ;
  assign n9821 = n9785 & ~n9820 ;
  assign n9822 = ( n9819 & n9820 ) | ( n9819 & ~n9821 ) | ( n9820 & ~n9821 ) ;
  assign n9823 = ( n9784 & n9818 ) | ( n9784 & ~n9822 ) | ( n9818 & ~n9822 ) ;
  assign n9824 = n9800 & ~n9804 ;
  assign n9825 = ( n9800 & ~n9812 ) | ( n9800 & n9824 ) | ( ~n9812 & n9824 ) ;
  assign n9826 = n9781 & ~n9782 ;
  assign n9827 = ( ~n9778 & n9781 ) | ( ~n9778 & n9826 ) | ( n9781 & n9826 ) ;
  assign n9828 = ~n9825 & n9827 ;
  assign n9829 = n9825 & ~n9827 ;
  assign n9830 = n9828 | n9829 ;
  assign n9831 = ( x520 & x521 ) | ( x520 & x522 ) | ( x521 & x522 ) ;
  assign n9832 = ( x517 & x518 ) | ( x517 & x519 ) | ( x518 & x519 ) ;
  assign n9833 = n9831 & ~n9832 ;
  assign n9834 = ~n9831 & n9832 ;
  assign n9835 = n9833 | n9834 ;
  assign n9836 = ~x517 & x518 ;
  assign n9837 = x517 & ~x518 ;
  assign n9838 = n9836 | n9837 ;
  assign n9839 = ~x519 & n9838 ;
  assign n9840 = x519 & ~n9838 ;
  assign n9841 = n9839 | n9840 ;
  assign n9842 = ~x520 & x521 ;
  assign n9843 = x520 & ~x521 ;
  assign n9844 = n9842 | n9843 ;
  assign n9845 = ~x522 & n9844 ;
  assign n9846 = x522 & ~n9844 ;
  assign n9847 = n9845 | n9846 ;
  assign n9848 = n9841 & n9847 ;
  assign n9849 = n9835 & ~n9848 ;
  assign n9850 = ~n9835 & n9848 ;
  assign n9851 = n9849 | n9850 ;
  assign n9852 = n9841 & ~n9847 ;
  assign n9853 = ~n9841 & n9847 ;
  assign n9854 = n9852 | n9853 ;
  assign n9855 = ( n9831 & n9832 ) | ( n9831 & n9848 ) | ( n9832 & n9848 ) ;
  assign n9856 = n9854 & ~n9855 ;
  assign n9857 = ( ~n9851 & n9854 ) | ( ~n9851 & n9856 ) | ( n9854 & n9856 ) ;
  assign n9858 = ~x511 & x512 ;
  assign n9859 = x511 & ~x512 ;
  assign n9860 = n9858 | n9859 ;
  assign n9861 = ~x513 & n9860 ;
  assign n9862 = x513 & ~n9860 ;
  assign n9863 = n9861 | n9862 ;
  assign n9864 = ~x514 & x515 ;
  assign n9865 = x514 & ~x515 ;
  assign n9866 = n9864 | n9865 ;
  assign n9867 = ~x516 & n9866 ;
  assign n9868 = x516 & ~n9866 ;
  assign n9869 = n9867 | n9868 ;
  assign n9870 = n9863 & ~n9869 ;
  assign n9871 = ~n9863 & n9869 ;
  assign n9872 = n9870 | n9871 ;
  assign n9873 = ( x514 & x515 ) | ( x514 & x516 ) | ( x515 & x516 ) ;
  assign n9874 = ( x511 & x512 ) | ( x511 & x513 ) | ( x512 & x513 ) ;
  assign n9875 = n9873 & ~n9874 ;
  assign n9876 = ~n9873 & n9874 ;
  assign n9877 = n9875 | n9876 ;
  assign n9878 = n9863 & n9869 ;
  assign n9879 = n9877 & ~n9878 ;
  assign n9880 = ~n9877 & n9878 ;
  assign n9881 = n9879 | n9880 ;
  assign n9882 = ( n9873 & n9874 ) | ( n9873 & n9878 ) | ( n9874 & n9878 ) ;
  assign n9883 = n9872 & ~n9882 ;
  assign n9884 = ( n9872 & ~n9881 ) | ( n9872 & n9883 ) | ( ~n9881 & n9883 ) ;
  assign n9885 = ~n9857 & n9884 ;
  assign n9886 = n9857 & ~n9884 ;
  assign n9887 = n9885 | n9886 ;
  assign n9888 = n9830 & n9887 ;
  assign n9889 = ( n9784 & ~n9785 ) | ( n9784 & n9820 ) | ( ~n9785 & n9820 ) ;
  assign n9890 = n9784 & n9820 ;
  assign n9891 = ( n9819 & n9889 ) | ( n9819 & n9890 ) | ( n9889 & n9890 ) ;
  assign n9892 = n9822 & ~n9891 ;
  assign n9893 = n9888 | n9892 ;
  assign n9894 = n9823 | n9893 ;
  assign n9895 = n9881 & n9882 ;
  assign n9896 = n9854 & n9855 ;
  assign n9897 = n9895 | n9896 ;
  assign n9898 = n9851 & n9855 ;
  assign n9899 = n9854 & n9872 ;
  assign n9900 = n9851 & n9899 ;
  assign n9901 = ~n9898 & n9900 ;
  assign n9902 = ~n9897 & n9901 ;
  assign n9903 = n9872 & n9882 ;
  assign n9904 = n9881 & ~n9903 ;
  assign n9905 = ~n9902 & n9904 ;
  assign n9906 = ~n9898 & n9899 ;
  assign n9907 = n9851 & ~n9896 ;
  assign n9908 = ( n9895 & n9904 ) | ( n9895 & n9907 ) | ( n9904 & n9907 ) ;
  assign n9909 = n9904 | n9907 ;
  assign n9910 = ( ~n9906 & n9908 ) | ( ~n9906 & n9909 ) | ( n9908 & n9909 ) ;
  assign n9911 = n9895 | n9907 ;
  assign n9912 = n9906 & ~n9911 ;
  assign n9913 = ( ~n9907 & n9910 ) | ( ~n9907 & n9912 ) | ( n9910 & n9912 ) ;
  assign n9914 = ( ~n9905 & n9910 ) | ( ~n9905 & n9913 ) | ( n9910 & n9913 ) ;
  assign n9915 = n9894 & n9914 ;
  assign n9916 = n9888 & n9892 ;
  assign n9917 = ( n9823 & n9888 ) | ( n9823 & n9916 ) | ( n9888 & n9916 ) ;
  assign n9918 = n9915 | n9917 ;
  assign n9919 = n9895 & ~n9907 ;
  assign n9920 = ( n9906 & n9907 ) | ( n9906 & ~n9919 ) | ( n9907 & ~n9919 ) ;
  assign n9921 = n9904 & n9920 ;
  assign n9922 = ~n9872 & n9882 ;
  assign n9923 = ( ~n9881 & n9882 ) | ( ~n9881 & n9922 ) | ( n9882 & n9922 ) ;
  assign n9924 = ~n9854 & n9855 ;
  assign n9925 = ( ~n9851 & n9855 ) | ( ~n9851 & n9924 ) | ( n9855 & n9924 ) ;
  assign n9926 = ~n9923 & n9925 ;
  assign n9927 = n9923 & ~n9925 ;
  assign n9928 = n9926 | n9927 ;
  assign n9929 = n9902 | n9928 ;
  assign n9930 = n9921 | n9929 ;
  assign n9931 = n9902 & n9928 ;
  assign n9932 = ( n9921 & n9928 ) | ( n9921 & n9931 ) | ( n9928 & n9931 ) ;
  assign n9933 = n9930 & ~n9932 ;
  assign n9934 = n9784 & n9822 ;
  assign n9935 = ~n9781 & n9782 ;
  assign n9936 = ( ~n9778 & n9782 ) | ( ~n9778 & n9935 ) | ( n9782 & n9935 ) ;
  assign n9937 = ~n9800 & n9804 ;
  assign n9938 = ( n9804 & ~n9812 ) | ( n9804 & n9937 ) | ( ~n9812 & n9937 ) ;
  assign n9939 = ~n9936 & n9938 ;
  assign n9940 = n9936 & ~n9938 ;
  assign n9941 = n9939 | n9940 ;
  assign n9942 = n9817 | n9941 ;
  assign n9943 = n9934 | n9942 ;
  assign n9944 = n9817 & n9941 ;
  assign n9945 = ( n9934 & n9941 ) | ( n9934 & n9944 ) | ( n9941 & n9944 ) ;
  assign n9946 = n9943 & ~n9945 ;
  assign n9947 = n9933 | n9946 ;
  assign n9948 = n9918 & n9947 ;
  assign n9949 = n9930 & n9943 ;
  assign n9950 = n9932 | n9945 ;
  assign n9951 = n9949 & ~n9950 ;
  assign n9952 = ( n9817 & n9936 ) | ( n9817 & n9938 ) | ( n9936 & n9938 ) ;
  assign n9953 = n9936 | n9938 ;
  assign n9954 = ( n9934 & n9952 ) | ( n9934 & n9953 ) | ( n9952 & n9953 ) ;
  assign n9955 = ( n9902 & n9923 ) | ( n9902 & n9925 ) | ( n9923 & n9925 ) ;
  assign n9956 = n9923 | n9925 ;
  assign n9957 = ( n9921 & n9955 ) | ( n9921 & n9956 ) | ( n9955 & n9956 ) ;
  assign n9958 = ~n9954 & n9957 ;
  assign n9959 = n9954 & ~n9957 ;
  assign n9960 = n9958 | n9959 ;
  assign n9961 = n9951 | n9960 ;
  assign n9962 = n9948 | n9961 ;
  assign n9963 = n9947 | n9951 ;
  assign n9964 = ( n9918 & n9951 ) | ( n9918 & n9963 ) | ( n9951 & n9963 ) ;
  assign n9965 = n9960 & n9964 ;
  assign n9966 = n9962 & ~n9965 ;
  assign n9967 = n9757 | n9966 ;
  assign n9968 = n9685 & ~n9708 ;
  assign n9969 = n9705 & ~n9968 ;
  assign n9970 = n9621 & ~n9678 ;
  assign n9971 = ~n9621 & n9678 ;
  assign n9972 = n9970 | n9971 ;
  assign n9973 = n9830 & ~n9887 ;
  assign n9974 = ~n9830 & n9887 ;
  assign n9975 = n9973 | n9974 ;
  assign n9976 = n9972 & n9975 ;
  assign n9977 = ~n9679 & n9685 ;
  assign n9978 = n9685 & ~n9705 ;
  assign n9979 = n9614 | n9683 ;
  assign n9980 = n9705 | n9979 ;
  assign n9981 = ( n9977 & n9978 ) | ( n9977 & ~n9980 ) | ( n9978 & ~n9980 ) ;
  assign n9982 = n9976 | n9981 ;
  assign n9983 = n9969 | n9982 ;
  assign n9984 = n9823 | n9892 ;
  assign n9985 = ( n9888 & n9914 ) | ( n9888 & ~n9984 ) | ( n9914 & ~n9984 ) ;
  assign n9986 = ( ~n9914 & n9984 ) | ( ~n9914 & n9985 ) | ( n9984 & n9985 ) ;
  assign n9987 = ( ~n9888 & n9985 ) | ( ~n9888 & n9986 ) | ( n9985 & n9986 ) ;
  assign n9988 = n9983 & n9987 ;
  assign n9989 = n9969 | n9981 ;
  assign n9990 = n9976 & n9989 ;
  assign n9991 = ( n9917 & ~n9933 ) | ( n9917 & n9946 ) | ( ~n9933 & n9946 ) ;
  assign n9992 = n9933 & ~n9946 ;
  assign n9993 = ( n9915 & n9991 ) | ( n9915 & ~n9992 ) | ( n9991 & ~n9992 ) ;
  assign n9994 = ( ~n9918 & n9933 ) | ( ~n9918 & n9993 ) | ( n9933 & n9993 ) ;
  assign n9995 = ( ~n9946 & n9993 ) | ( ~n9946 & n9994 ) | ( n9993 & n9994 ) ;
  assign n9996 = ( n9708 & ~n9724 ) | ( n9708 & n9737 ) | ( ~n9724 & n9737 ) ;
  assign n9997 = n9724 & ~n9737 ;
  assign n9998 = ( n9706 & n9996 ) | ( n9706 & ~n9997 ) | ( n9996 & ~n9997 ) ;
  assign n9999 = ( ~n9709 & n9724 ) | ( ~n9709 & n9998 ) | ( n9724 & n9998 ) ;
  assign n10000 = ( ~n9737 & n9998 ) | ( ~n9737 & n9999 ) | ( n9998 & n9999 ) ;
  assign n10001 = ( n9990 & n9995 ) | ( n9990 & n10000 ) | ( n9995 & n10000 ) ;
  assign n10002 = n9995 | n10000 ;
  assign n10003 = ( n9988 & n10001 ) | ( n9988 & n10002 ) | ( n10001 & n10002 ) ;
  assign n10004 = n9967 & n10003 ;
  assign n10005 = n9753 & n9962 ;
  assign n10006 = n9756 | n9965 ;
  assign n10007 = n10005 & ~n10006 ;
  assign n10008 = n9954 & n9957 ;
  assign n10009 = n9954 | n9957 ;
  assign n10010 = n10008 | n10009 ;
  assign n10011 = ( n9964 & n10008 ) | ( n9964 & n10010 ) | ( n10008 & n10010 ) ;
  assign n10012 = n9745 & n9748 ;
  assign n10013 = n9745 | n9748 ;
  assign n10014 = n10012 | n10013 ;
  assign n10015 = ( n9755 & n10012 ) | ( n9755 & n10014 ) | ( n10012 & n10014 ) ;
  assign n10016 = n10011 & n10015 ;
  assign n10017 = n10015 & ~n10016 ;
  assign n10018 = ( n10011 & ~n10016 ) | ( n10011 & n10017 ) | ( ~n10016 & n10017 ) ;
  assign n10019 = n10007 | n10018 ;
  assign n10020 = n10004 | n10019 ;
  assign n10021 = n10004 | n10007 ;
  assign n10022 = n10018 & n10021 ;
  assign n10023 = n10020 & ~n10022 ;
  assign n10024 = n9548 | n10023 ;
  assign n10025 = n9497 & ~n9500 ;
  assign n10026 = ~n9497 & n9500 ;
  assign n10027 = n10025 | n10026 ;
  assign n10028 = n9972 & ~n9975 ;
  assign n10029 = ~n9972 & n9975 ;
  assign n10030 = n10028 | n10029 ;
  assign n10031 = n10027 & n10030 ;
  assign n10032 = ~n9983 & n9987 ;
  assign n10033 = ( n9987 & n9990 ) | ( n9987 & n10032 ) | ( n9990 & n10032 ) ;
  assign n10034 = ~n9976 & n9989 ;
  assign n10035 = n9976 & ~n9981 ;
  assign n10036 = ~n9969 & n10035 ;
  assign n10037 = ~n9987 & n10036 ;
  assign n10038 = ( ~n9987 & n10034 ) | ( ~n9987 & n10037 ) | ( n10034 & n10037 ) ;
  assign n10039 = n10033 | n10038 ;
  assign n10040 = n10031 & n10039 ;
  assign n10041 = n10031 | n10034 ;
  assign n10042 = n9987 & ~n10031 ;
  assign n10043 = ( n10037 & n10041 ) | ( n10037 & ~n10042 ) | ( n10041 & ~n10042 ) ;
  assign n10044 = n10033 | n10043 ;
  assign n10045 = ~n9501 & n9514 ;
  assign n10046 = n9501 & ~n9506 ;
  assign n10047 = ~n9494 & n10046 ;
  assign n10048 = ~n9512 & n10047 ;
  assign n10049 = ( ~n9512 & n10045 ) | ( ~n9512 & n10048 ) | ( n10045 & n10048 ) ;
  assign n10050 = n9513 & ~n9515 ;
  assign n10051 = ( n9512 & n10049 ) | ( n9512 & ~n10050 ) | ( n10049 & ~n10050 ) ;
  assign n10052 = n10044 & n10051 ;
  assign n10053 = n10040 | n10052 ;
  assign n10055 = ( n9515 & ~n9520 ) | ( n9515 & n9525 ) | ( ~n9520 & n9525 ) ;
  assign n10056 = n9520 & ~n9525 ;
  assign n10057 = ( n9513 & n10055 ) | ( n9513 & ~n10056 ) | ( n10055 & ~n10056 ) ;
  assign n10054 = n9513 | n9515 ;
  assign n10058 = ( n9520 & ~n10054 ) | ( n9520 & n10057 ) | ( ~n10054 & n10057 ) ;
  assign n10059 = ( ~n9525 & n10057 ) | ( ~n9525 & n10058 ) | ( n10057 & n10058 ) ;
  assign n10061 = ( n9990 & ~n9995 ) | ( n9990 & n10000 ) | ( ~n9995 & n10000 ) ;
  assign n10062 = n9995 & ~n10000 ;
  assign n10063 = ( n9988 & n10061 ) | ( n9988 & ~n10062 ) | ( n10061 & ~n10062 ) ;
  assign n10060 = n9988 | n9990 ;
  assign n10064 = ( n9995 & ~n10060 ) | ( n9995 & n10063 ) | ( ~n10060 & n10063 ) ;
  assign n10065 = ( ~n10000 & n10063 ) | ( ~n10000 & n10064 ) | ( n10063 & n10064 ) ;
  assign n10066 = ( n10053 & n10059 ) | ( n10053 & n10065 ) | ( n10059 & n10065 ) ;
  assign n10067 = ( ~n9757 & n9966 ) | ( ~n9757 & n10003 ) | ( n9966 & n10003 ) ;
  assign n10068 = ( n9757 & ~n10003 ) | ( n9757 & n10067 ) | ( ~n10003 & n10067 ) ;
  assign n10069 = ( ~n9966 & n10067 ) | ( ~n9966 & n10068 ) | ( n10067 & n10068 ) ;
  assign n10070 = ( ~n9282 & n9491 ) | ( ~n9282 & n9528 ) | ( n9491 & n9528 ) ;
  assign n10071 = ( n9282 & ~n9528 ) | ( n9282 & n10070 ) | ( ~n9528 & n10070 ) ;
  assign n10072 = ( ~n9491 & n10070 ) | ( ~n9491 & n10071 ) | ( n10070 & n10071 ) ;
  assign n10073 = ( n10066 & n10069 ) | ( n10066 & n10072 ) | ( n10069 & n10072 ) ;
  assign n10074 = n10024 & n10073 ;
  assign n10075 = n9545 & n10020 ;
  assign n10076 = n9547 | n10022 ;
  assign n10077 = n10075 & ~n10076 ;
  assign n10086 = n9280 & n9538 ;
  assign n10087 = n9482 | n9537 ;
  assign n10088 = n9479 | n9537 ;
  assign n10089 = ( n9489 & n10087 ) | ( n9489 & n10088 ) | ( n10087 & n10088 ) ;
  assign n10090 = n10086 | n10089 ;
  assign n10091 = n9541 | n10090 ;
  assign n10092 = ( n9532 & n9541 ) | ( n9532 & n10091 ) | ( n9541 & n10091 ) ;
  assign n10093 = n9541 | n10091 ;
  assign n10094 = ( n9529 & n10092 ) | ( n9529 & n10093 ) | ( n10092 & n10093 ) ;
  assign n10078 = n9755 & n10013 ;
  assign n10079 = n9957 | n10012 ;
  assign n10080 = n9954 | n10012 ;
  assign n10081 = ( n9964 & n10079 ) | ( n9964 & n10080 ) | ( n10079 & n10080 ) ;
  assign n10082 = n10078 | n10081 ;
  assign n10083 = n10007 & n10082 ;
  assign n10084 = ( n10004 & n10082 ) | ( n10004 & n10083 ) | ( n10082 & n10083 ) ;
  assign n10085 = n10016 | n10084 ;
  assign n10095 = n10085 & n10094 ;
  assign n10096 = n10085 & ~n10095 ;
  assign n10097 = ( n10094 & ~n10095 ) | ( n10094 & n10096 ) | ( ~n10095 & n10096 ) ;
  assign n10098 = n10077 | n10097 ;
  assign n10099 = n10074 | n10098 ;
  assign n10100 = n10074 | n10077 ;
  assign n10101 = n10097 & n10100 ;
  assign n10102 = n10099 & ~n10101 ;
  assign n10103 = n9073 | n10102 ;
  assign n10104 = ( ~n9548 & n10023 ) | ( ~n9548 & n10073 ) | ( n10023 & n10073 ) ;
  assign n10105 = ( n9548 & ~n10073 ) | ( n9548 & n10104 ) | ( ~n10073 & n10104 ) ;
  assign n10106 = ( ~n10023 & n10104 ) | ( ~n10023 & n10105 ) | ( n10104 & n10105 ) ;
  assign n10107 = ( ~n8521 & n8996 ) | ( ~n8521 & n9044 ) | ( n8996 & n9044 ) ;
  assign n10108 = ( n8521 & ~n9044 ) | ( n8521 & n10107 ) | ( ~n9044 & n10107 ) ;
  assign n10109 = ( ~n8996 & n10107 ) | ( ~n8996 & n10108 ) | ( n10107 & n10108 ) ;
  assign n10110 = n10027 & ~n10030 ;
  assign n10111 = ~n10027 & n10030 ;
  assign n10112 = n10110 | n10111 ;
  assign n10113 = n9013 & ~n9016 ;
  assign n10114 = ~n9013 & n9016 ;
  assign n10115 = n10113 | n10114 ;
  assign n10116 = n10112 & n10115 ;
  assign n10117 = n9026 & ~n9028 ;
  assign n10118 = n9010 & ~n10117 ;
  assign n10119 = ~n9017 & n9025 ;
  assign n10120 = n9017 & ~n9025 ;
  assign n10121 = n10119 | n10120 ;
  assign n10122 = ~n9010 & n10121 ;
  assign n10123 = n10118 | n10122 ;
  assign n10124 = n10116 & n10123 ;
  assign n10125 = n9010 & ~n10116 ;
  assign n10126 = ( n10116 & n10121 ) | ( n10116 & ~n10125 ) | ( n10121 & ~n10125 ) ;
  assign n10127 = n10118 | n10126 ;
  assign n10128 = ( n10031 & ~n10039 ) | ( n10031 & n10051 ) | ( ~n10039 & n10051 ) ;
  assign n10129 = ( ~n10031 & n10039 ) | ( ~n10031 & n10128 ) | ( n10039 & n10128 ) ;
  assign n10130 = ( ~n10051 & n10128 ) | ( ~n10051 & n10129 ) | ( n10128 & n10129 ) ;
  assign n10131 = n10127 & n10130 ;
  assign n10132 = n10124 | n10131 ;
  assign n10133 = ( n10053 & ~n10059 ) | ( n10053 & n10065 ) | ( ~n10059 & n10065 ) ;
  assign n10134 = ( ~n10053 & n10059 ) | ( ~n10053 & n10133 ) | ( n10059 & n10133 ) ;
  assign n10135 = ( ~n10065 & n10133 ) | ( ~n10065 & n10134 ) | ( n10133 & n10134 ) ;
  assign n10137 = ( n9028 & ~n9034 ) | ( n9028 & n9040 ) | ( ~n9034 & n9040 ) ;
  assign n10138 = n9034 & ~n9040 ;
  assign n10139 = ( n9027 & n10137 ) | ( n9027 & ~n10138 ) | ( n10137 & ~n10138 ) ;
  assign n10136 = n9027 | n9028 ;
  assign n10140 = ( n9034 & ~n10136 ) | ( n9034 & n10139 ) | ( ~n10136 & n10139 ) ;
  assign n10141 = ( ~n9040 & n10139 ) | ( ~n9040 & n10140 ) | ( n10139 & n10140 ) ;
  assign n10142 = ( n10132 & n10135 ) | ( n10132 & n10141 ) | ( n10135 & n10141 ) ;
  assign n10143 = ( ~n9000 & n9003 ) | ( ~n9000 & n9043 ) | ( n9003 & n9043 ) ;
  assign n10144 = ( n9000 & ~n9043 ) | ( n9000 & n10143 ) | ( ~n9043 & n10143 ) ;
  assign n10145 = ( ~n9003 & n10143 ) | ( ~n9003 & n10144 ) | ( n10143 & n10144 ) ;
  assign n10146 = ( n10066 & ~n10069 ) | ( n10066 & n10072 ) | ( ~n10069 & n10072 ) ;
  assign n10147 = ( ~n10066 & n10069 ) | ( ~n10066 & n10146 ) | ( n10069 & n10146 ) ;
  assign n10148 = ( ~n10072 & n10146 ) | ( ~n10072 & n10147 ) | ( n10146 & n10147 ) ;
  assign n10149 = ( n10142 & n10145 ) | ( n10142 & n10148 ) | ( n10145 & n10148 ) ;
  assign n10150 = ( n10106 & n10109 ) | ( n10106 & n10149 ) | ( n10109 & n10149 ) ;
  assign n10151 = n10103 & n10150 ;
  assign n10152 = n9070 & n10099 ;
  assign n10153 = n9072 | n10101 ;
  assign n10154 = n10152 & ~n10153 ;
  assign n10162 = n9541 | n10016 ;
  assign n10163 = n10090 | n10162 ;
  assign n10164 = ( n9546 & n10162 ) | ( n9546 & n10163 ) | ( n10162 & n10163 ) ;
  assign n10165 = n10084 | n10164 ;
  assign n10166 = n10095 | n10165 ;
  assign n10167 = ( n10077 & n10095 ) | ( n10077 & n10166 ) | ( n10095 & n10166 ) ;
  assign n10168 = n10095 | n10166 ;
  assign n10169 = ( n10074 & n10167 ) | ( n10074 & n10168 ) | ( n10167 & n10168 ) ;
  assign n10155 = n8514 | n8989 ;
  assign n10156 = n9061 | n10155 ;
  assign n10157 = ( n8519 & n10155 ) | ( n8519 & n10156 ) | ( n10155 & n10156 ) ;
  assign n10158 = n9055 | n10157 ;
  assign n10159 = n9048 & n10158 ;
  assign n10160 = ( n9045 & n10158 ) | ( n9045 & n10159 ) | ( n10158 & n10159 ) ;
  assign n10161 = n9066 | n10160 ;
  assign n10170 = n10161 & n10169 ;
  assign n10171 = n10161 & ~n10170 ;
  assign n10172 = ( n10169 & ~n10170 ) | ( n10169 & n10171 ) | ( ~n10170 & n10171 ) ;
  assign n10173 = n10154 | n10172 ;
  assign n10174 = n10151 | n10173 ;
  assign n10175 = ~x787 & x788 ;
  assign n10176 = x787 & ~x788 ;
  assign n10177 = n10175 | n10176 ;
  assign n10178 = ~x789 & n10177 ;
  assign n10179 = x789 & ~n10177 ;
  assign n10180 = n10178 | n10179 ;
  assign n10181 = ~x790 & x791 ;
  assign n10182 = x790 & ~x791 ;
  assign n10183 = n10181 | n10182 ;
  assign n10184 = ~x792 & n10183 ;
  assign n10185 = x792 & ~n10183 ;
  assign n10186 = n10184 | n10185 ;
  assign n10187 = n10180 & n10186 ;
  assign n10188 = ( x790 & x791 ) | ( x790 & x792 ) | ( x791 & x792 ) ;
  assign n10189 = ( x787 & x788 ) | ( x787 & x789 ) | ( x788 & x789 ) ;
  assign n10190 = ~n10188 & n10189 ;
  assign n10191 = n10188 & ~n10189 ;
  assign n10192 = n10190 | n10191 ;
  assign n10193 = ~n10187 & n10192 ;
  assign n10194 = n10187 & ~n10192 ;
  assign n10195 = n10193 | n10194 ;
  assign n10196 = n10180 & ~n10186 ;
  assign n10197 = ~n10180 & n10186 ;
  assign n10198 = n10196 | n10197 ;
  assign n10199 = ( n10187 & n10188 ) | ( n10187 & n10189 ) | ( n10188 & n10189 ) ;
  assign n10200 = n10198 & n10199 ;
  assign n10201 = n10195 & ~n10200 ;
  assign n10202 = n10195 & n10199 ;
  assign n10203 = x793 & ~x794 ;
  assign n10204 = ~x793 & x794 ;
  assign n10205 = n10203 | n10204 ;
  assign n10206 = ~x795 & n10205 ;
  assign n10207 = x795 & ~n10205 ;
  assign n10208 = n10206 | n10207 ;
  assign n10209 = x796 & ~x797 ;
  assign n10210 = ~x796 & x797 ;
  assign n10211 = n10209 | n10210 ;
  assign n10212 = ~x798 & n10211 ;
  assign n10213 = x798 & ~n10211 ;
  assign n10214 = n10212 | n10213 ;
  assign n10215 = n10208 & ~n10214 ;
  assign n10216 = ~n10208 & n10214 ;
  assign n10217 = n10215 | n10216 ;
  assign n10218 = ( x796 & x797 ) | ( x796 & x798 ) | ( x797 & x798 ) ;
  assign n10219 = ( x793 & x794 ) | ( x793 & x795 ) | ( x794 & x795 ) ;
  assign n10220 = n10208 & n10214 ;
  assign n10221 = ( n10218 & n10219 ) | ( n10218 & n10220 ) | ( n10219 & n10220 ) ;
  assign n10222 = n10217 & n10221 ;
  assign n10223 = n10202 | n10222 ;
  assign n10224 = n10218 & ~n10219 ;
  assign n10225 = ~n10218 & n10219 ;
  assign n10226 = n10224 | n10225 ;
  assign n10227 = ~n10220 & n10226 ;
  assign n10228 = n10220 & ~n10226 ;
  assign n10229 = n10227 | n10228 ;
  assign n10230 = n10221 & n10229 ;
  assign n10231 = n10198 & n10217 ;
  assign n10232 = n10229 & n10231 ;
  assign n10233 = ~n10230 & n10232 ;
  assign n10234 = ~n10223 & n10233 ;
  assign n10235 = n10201 & n10234 ;
  assign n10236 = ~n10230 & n10231 ;
  assign n10237 = ~n10222 & n10229 ;
  assign n10238 = n10202 & ~n10237 ;
  assign n10239 = ( n10236 & n10237 ) | ( n10236 & ~n10238 ) | ( n10237 & ~n10238 ) ;
  assign n10240 = ( n10201 & n10235 ) | ( n10201 & ~n10239 ) | ( n10235 & ~n10239 ) ;
  assign n10241 = n10217 & ~n10221 ;
  assign n10242 = ( n10217 & ~n10229 ) | ( n10217 & n10241 ) | ( ~n10229 & n10241 ) ;
  assign n10243 = n10198 & ~n10199 ;
  assign n10244 = ( ~n10195 & n10198 ) | ( ~n10195 & n10243 ) | ( n10198 & n10243 ) ;
  assign n10245 = ~n10242 & n10244 ;
  assign n10246 = n10242 & ~n10244 ;
  assign n10247 = n10245 | n10246 ;
  assign n10248 = ( x784 & x785 ) | ( x784 & x786 ) | ( x785 & x786 ) ;
  assign n10249 = ( x781 & x782 ) | ( x781 & x783 ) | ( x782 & x783 ) ;
  assign n10250 = n10248 & ~n10249 ;
  assign n10251 = ~n10248 & n10249 ;
  assign n10252 = n10250 | n10251 ;
  assign n10253 = x781 & ~x782 ;
  assign n10254 = ~x781 & x782 ;
  assign n10255 = n10253 | n10254 ;
  assign n10256 = ~x783 & n10255 ;
  assign n10257 = x783 & ~n10255 ;
  assign n10258 = n10256 | n10257 ;
  assign n10259 = x784 & ~x785 ;
  assign n10260 = ~x784 & x785 ;
  assign n10261 = n10259 | n10260 ;
  assign n10262 = ~x786 & n10261 ;
  assign n10263 = x786 & ~n10261 ;
  assign n10264 = n10262 | n10263 ;
  assign n10265 = n10258 & n10264 ;
  assign n10266 = n10252 & ~n10265 ;
  assign n10267 = ~n10252 & n10265 ;
  assign n10268 = n10266 | n10267 ;
  assign n10269 = n10258 & ~n10264 ;
  assign n10270 = ~n10258 & n10264 ;
  assign n10271 = n10269 | n10270 ;
  assign n10272 = ( n10248 & n10249 ) | ( n10248 & n10265 ) | ( n10249 & n10265 ) ;
  assign n10273 = n10271 & ~n10272 ;
  assign n10274 = ( ~n10268 & n10271 ) | ( ~n10268 & n10273 ) | ( n10271 & n10273 ) ;
  assign n10275 = ~x775 & x776 ;
  assign n10276 = x775 & ~x776 ;
  assign n10277 = n10275 | n10276 ;
  assign n10278 = ~x777 & n10277 ;
  assign n10279 = x777 & ~n10277 ;
  assign n10280 = n10278 | n10279 ;
  assign n10281 = ~x778 & x779 ;
  assign n10282 = x778 & ~x779 ;
  assign n10283 = n10281 | n10282 ;
  assign n10284 = ~x780 & n10283 ;
  assign n10285 = x780 & ~n10283 ;
  assign n10286 = n10284 | n10285 ;
  assign n10287 = n10280 & n10286 ;
  assign n10288 = ( x778 & x779 ) | ( x778 & x780 ) | ( x779 & x780 ) ;
  assign n10289 = ( x775 & x776 ) | ( x775 & x777 ) | ( x776 & x777 ) ;
  assign n10290 = ~n10288 & n10289 ;
  assign n10291 = n10288 & ~n10289 ;
  assign n10292 = n10290 | n10291 ;
  assign n10293 = ~n10287 & n10292 ;
  assign n10294 = n10287 & ~n10292 ;
  assign n10295 = n10293 | n10294 ;
  assign n10296 = n10280 & ~n10286 ;
  assign n10297 = ~n10280 & n10286 ;
  assign n10298 = n10296 | n10297 ;
  assign n10299 = ( n10287 & n10288 ) | ( n10287 & n10289 ) | ( n10288 & n10289 ) ;
  assign n10300 = n10298 & ~n10299 ;
  assign n10301 = ( ~n10295 & n10298 ) | ( ~n10295 & n10300 ) | ( n10298 & n10300 ) ;
  assign n10302 = ~n10274 & n10301 ;
  assign n10303 = n10274 & ~n10301 ;
  assign n10304 = n10302 | n10303 ;
  assign n10305 = n10247 & n10304 ;
  assign n10306 = ( n10201 & ~n10202 ) | ( n10201 & n10237 ) | ( ~n10202 & n10237 ) ;
  assign n10307 = n10201 & n10237 ;
  assign n10308 = ( n10236 & n10306 ) | ( n10236 & n10307 ) | ( n10306 & n10307 ) ;
  assign n10309 = n10239 & ~n10308 ;
  assign n10310 = n10305 | n10309 ;
  assign n10311 = n10240 | n10310 ;
  assign n10312 = n10295 & n10299 ;
  assign n10313 = n10271 & n10272 ;
  assign n10314 = n10312 | n10313 ;
  assign n10315 = n10268 & n10272 ;
  assign n10316 = n10271 & n10298 ;
  assign n10317 = n10268 & n10316 ;
  assign n10318 = ~n10315 & n10317 ;
  assign n10319 = ~n10314 & n10318 ;
  assign n10320 = n10298 & n10299 ;
  assign n10321 = n10295 & ~n10320 ;
  assign n10322 = ~n10319 & n10321 ;
  assign n10323 = ~n10315 & n10316 ;
  assign n10324 = n10268 & ~n10313 ;
  assign n10325 = ( n10312 & n10321 ) | ( n10312 & n10324 ) | ( n10321 & n10324 ) ;
  assign n10326 = n10321 | n10324 ;
  assign n10327 = ( ~n10323 & n10325 ) | ( ~n10323 & n10326 ) | ( n10325 & n10326 ) ;
  assign n10328 = n10312 | n10324 ;
  assign n10329 = n10323 & ~n10328 ;
  assign n10330 = ( ~n10324 & n10327 ) | ( ~n10324 & n10329 ) | ( n10327 & n10329 ) ;
  assign n10331 = ( ~n10322 & n10327 ) | ( ~n10322 & n10330 ) | ( n10327 & n10330 ) ;
  assign n10332 = n10311 & n10331 ;
  assign n10333 = n10305 & n10309 ;
  assign n10334 = ( n10240 & n10305 ) | ( n10240 & n10333 ) | ( n10305 & n10333 ) ;
  assign n10335 = n10332 | n10334 ;
  assign n10336 = n10312 & ~n10324 ;
  assign n10337 = ( n10323 & n10324 ) | ( n10323 & ~n10336 ) | ( n10324 & ~n10336 ) ;
  assign n10338 = n10321 & n10337 ;
  assign n10339 = ~n10298 & n10299 ;
  assign n10340 = ( ~n10295 & n10299 ) | ( ~n10295 & n10339 ) | ( n10299 & n10339 ) ;
  assign n10341 = ~n10271 & n10272 ;
  assign n10342 = ( ~n10268 & n10272 ) | ( ~n10268 & n10341 ) | ( n10272 & n10341 ) ;
  assign n10343 = ~n10340 & n10342 ;
  assign n10344 = n10340 & ~n10342 ;
  assign n10345 = n10343 | n10344 ;
  assign n10346 = n10319 | n10345 ;
  assign n10347 = n10338 | n10346 ;
  assign n10348 = n10319 & n10345 ;
  assign n10349 = ( n10338 & n10345 ) | ( n10338 & n10348 ) | ( n10345 & n10348 ) ;
  assign n10350 = n10347 & ~n10349 ;
  assign n10351 = n10201 & n10239 ;
  assign n10352 = ~n10198 & n10199 ;
  assign n10353 = ( ~n10195 & n10199 ) | ( ~n10195 & n10352 ) | ( n10199 & n10352 ) ;
  assign n10354 = ~n10217 & n10221 ;
  assign n10355 = ( n10221 & ~n10229 ) | ( n10221 & n10354 ) | ( ~n10229 & n10354 ) ;
  assign n10356 = ~n10353 & n10355 ;
  assign n10357 = n10353 & ~n10355 ;
  assign n10358 = n10356 | n10357 ;
  assign n10359 = n10234 | n10358 ;
  assign n10360 = n10351 | n10359 ;
  assign n10361 = n10234 & n10358 ;
  assign n10362 = ( n10351 & n10358 ) | ( n10351 & n10361 ) | ( n10358 & n10361 ) ;
  assign n10363 = n10360 & ~n10362 ;
  assign n10364 = n10350 | n10363 ;
  assign n10365 = n10335 & n10364 ;
  assign n10366 = n10347 & n10360 ;
  assign n10367 = n10349 | n10362 ;
  assign n10368 = n10366 & ~n10367 ;
  assign n10369 = ( n10234 & n10353 ) | ( n10234 & n10355 ) | ( n10353 & n10355 ) ;
  assign n10370 = n10353 | n10355 ;
  assign n10371 = ( n10351 & n10369 ) | ( n10351 & n10370 ) | ( n10369 & n10370 ) ;
  assign n10372 = ( n10319 & n10340 ) | ( n10319 & n10342 ) | ( n10340 & n10342 ) ;
  assign n10373 = n10340 | n10342 ;
  assign n10374 = ( n10338 & n10372 ) | ( n10338 & n10373 ) | ( n10372 & n10373 ) ;
  assign n10375 = ~n10371 & n10374 ;
  assign n10376 = n10371 & ~n10374 ;
  assign n10377 = n10375 | n10376 ;
  assign n10378 = n10368 | n10377 ;
  assign n10379 = n10365 | n10378 ;
  assign n10380 = n10364 | n10368 ;
  assign n10381 = ( n10335 & n10368 ) | ( n10335 & n10380 ) | ( n10368 & n10380 ) ;
  assign n10382 = n10377 & n10381 ;
  assign n10383 = n10379 & ~n10382 ;
  assign n10384 = ( x766 & x767 ) | ( x766 & x768 ) | ( x767 & x768 ) ;
  assign n10385 = ( x763 & x764 ) | ( x763 & x765 ) | ( x764 & x765 ) ;
  assign n10386 = n10384 & ~n10385 ;
  assign n10387 = ~n10384 & n10385 ;
  assign n10388 = n10386 | n10387 ;
  assign n10389 = ~x763 & x764 ;
  assign n10390 = x763 & ~x764 ;
  assign n10391 = n10389 | n10390 ;
  assign n10392 = ~x765 & n10391 ;
  assign n10393 = x765 & ~n10391 ;
  assign n10394 = n10392 | n10393 ;
  assign n10395 = ~x766 & x767 ;
  assign n10396 = x766 & ~x767 ;
  assign n10397 = n10395 | n10396 ;
  assign n10398 = ~x768 & n10397 ;
  assign n10399 = x768 & ~n10397 ;
  assign n10400 = n10398 | n10399 ;
  assign n10401 = n10394 & n10400 ;
  assign n10402 = n10388 & ~n10401 ;
  assign n10403 = ~n10388 & n10401 ;
  assign n10404 = n10402 | n10403 ;
  assign n10405 = n10394 & ~n10400 ;
  assign n10406 = ~n10394 & n10400 ;
  assign n10407 = n10405 | n10406 ;
  assign n10408 = ( n10384 & n10385 ) | ( n10384 & n10401 ) | ( n10385 & n10401 ) ;
  assign n10409 = n10407 & n10408 ;
  assign n10410 = n10404 & ~n10409 ;
  assign n10411 = n10404 & n10408 ;
  assign n10412 = ~x769 & x770 ;
  assign n10413 = x769 & ~x770 ;
  assign n10414 = n10412 | n10413 ;
  assign n10415 = ~x771 & n10414 ;
  assign n10416 = x771 & ~n10414 ;
  assign n10417 = n10415 | n10416 ;
  assign n10418 = ~x772 & x773 ;
  assign n10419 = x772 & ~x773 ;
  assign n10420 = n10418 | n10419 ;
  assign n10421 = ~x774 & n10420 ;
  assign n10422 = x774 & ~n10420 ;
  assign n10423 = n10421 | n10422 ;
  assign n10424 = n10417 & ~n10423 ;
  assign n10425 = ~n10417 & n10423 ;
  assign n10426 = n10424 | n10425 ;
  assign n10427 = ( x772 & x773 ) | ( x772 & x774 ) | ( x773 & x774 ) ;
  assign n10428 = ( x769 & x770 ) | ( x769 & x771 ) | ( x770 & x771 ) ;
  assign n10429 = n10417 & n10423 ;
  assign n10430 = ( n10427 & n10428 ) | ( n10427 & n10429 ) | ( n10428 & n10429 ) ;
  assign n10431 = n10426 & n10430 ;
  assign n10432 = n10411 | n10431 ;
  assign n10433 = n10427 & ~n10428 ;
  assign n10434 = ~n10427 & n10428 ;
  assign n10435 = n10433 | n10434 ;
  assign n10436 = ~n10429 & n10435 ;
  assign n10437 = n10429 & ~n10435 ;
  assign n10438 = n10436 | n10437 ;
  assign n10439 = n10430 & n10438 ;
  assign n10440 = n10407 & n10426 ;
  assign n10441 = n10438 & n10440 ;
  assign n10442 = ~n10439 & n10441 ;
  assign n10443 = ~n10432 & n10442 ;
  assign n10444 = n10410 & n10443 ;
  assign n10445 = ~n10439 & n10440 ;
  assign n10446 = ~n10431 & n10438 ;
  assign n10447 = n10411 & ~n10446 ;
  assign n10448 = ( n10445 & n10446 ) | ( n10445 & ~n10447 ) | ( n10446 & ~n10447 ) ;
  assign n10449 = ( n10410 & n10444 ) | ( n10410 & ~n10448 ) | ( n10444 & ~n10448 ) ;
  assign n10450 = n10426 & ~n10430 ;
  assign n10451 = ( n10426 & ~n10438 ) | ( n10426 & n10450 ) | ( ~n10438 & n10450 ) ;
  assign n10452 = n10407 & ~n10408 ;
  assign n10453 = ( ~n10404 & n10407 ) | ( ~n10404 & n10452 ) | ( n10407 & n10452 ) ;
  assign n10454 = ~n10451 & n10453 ;
  assign n10455 = n10451 & ~n10453 ;
  assign n10456 = n10454 | n10455 ;
  assign n10457 = ( x760 & x761 ) | ( x760 & x762 ) | ( x761 & x762 ) ;
  assign n10458 = ( x757 & x758 ) | ( x757 & x759 ) | ( x758 & x759 ) ;
  assign n10459 = n10457 & ~n10458 ;
  assign n10460 = ~n10457 & n10458 ;
  assign n10461 = n10459 | n10460 ;
  assign n10462 = ~x757 & x758 ;
  assign n10463 = x757 & ~x758 ;
  assign n10464 = n10462 | n10463 ;
  assign n10465 = ~x759 & n10464 ;
  assign n10466 = x759 & ~n10464 ;
  assign n10467 = n10465 | n10466 ;
  assign n10468 = ~x760 & x761 ;
  assign n10469 = x760 & ~x761 ;
  assign n10470 = n10468 | n10469 ;
  assign n10471 = ~x762 & n10470 ;
  assign n10472 = x762 & ~n10470 ;
  assign n10473 = n10471 | n10472 ;
  assign n10474 = n10467 & n10473 ;
  assign n10475 = n10461 & ~n10474 ;
  assign n10476 = ~n10461 & n10474 ;
  assign n10477 = n10475 | n10476 ;
  assign n10478 = n10467 & ~n10473 ;
  assign n10479 = ~n10467 & n10473 ;
  assign n10480 = n10478 | n10479 ;
  assign n10481 = ( n10457 & n10458 ) | ( n10457 & n10474 ) | ( n10458 & n10474 ) ;
  assign n10482 = n10480 & ~n10481 ;
  assign n10483 = ( ~n10477 & n10480 ) | ( ~n10477 & n10482 ) | ( n10480 & n10482 ) ;
  assign n10484 = ~x751 & x752 ;
  assign n10485 = x751 & ~x752 ;
  assign n10486 = n10484 | n10485 ;
  assign n10487 = ~x753 & n10486 ;
  assign n10488 = x753 & ~n10486 ;
  assign n10489 = n10487 | n10488 ;
  assign n10490 = ~x754 & x755 ;
  assign n10491 = x754 & ~x755 ;
  assign n10492 = n10490 | n10491 ;
  assign n10493 = ~x756 & n10492 ;
  assign n10494 = x756 & ~n10492 ;
  assign n10495 = n10493 | n10494 ;
  assign n10496 = n10489 & ~n10495 ;
  assign n10497 = ~n10489 & n10495 ;
  assign n10498 = n10496 | n10497 ;
  assign n10499 = ( x754 & x755 ) | ( x754 & x756 ) | ( x755 & x756 ) ;
  assign n10500 = ( x751 & x752 ) | ( x751 & x753 ) | ( x752 & x753 ) ;
  assign n10501 = n10499 & ~n10500 ;
  assign n10502 = ~n10499 & n10500 ;
  assign n10503 = n10501 | n10502 ;
  assign n10504 = n10489 & n10495 ;
  assign n10505 = n10503 & ~n10504 ;
  assign n10506 = ~n10503 & n10504 ;
  assign n10507 = n10505 | n10506 ;
  assign n10508 = ( n10499 & n10500 ) | ( n10499 & n10504 ) | ( n10500 & n10504 ) ;
  assign n10509 = n10498 & ~n10508 ;
  assign n10510 = ( n10498 & ~n10507 ) | ( n10498 & n10509 ) | ( ~n10507 & n10509 ) ;
  assign n10511 = ~n10483 & n10510 ;
  assign n10512 = n10483 & ~n10510 ;
  assign n10513 = n10511 | n10512 ;
  assign n10514 = n10456 & n10513 ;
  assign n10515 = ( n10410 & ~n10411 ) | ( n10410 & n10446 ) | ( ~n10411 & n10446 ) ;
  assign n10516 = n10410 & n10446 ;
  assign n10517 = ( n10445 & n10515 ) | ( n10445 & n10516 ) | ( n10515 & n10516 ) ;
  assign n10518 = n10448 & ~n10517 ;
  assign n10519 = n10514 | n10518 ;
  assign n10520 = n10449 | n10519 ;
  assign n10521 = n10507 & n10508 ;
  assign n10522 = n10480 & n10481 ;
  assign n10523 = n10521 | n10522 ;
  assign n10524 = n10477 & n10481 ;
  assign n10525 = n10480 & n10498 ;
  assign n10526 = n10477 & n10525 ;
  assign n10527 = ~n10524 & n10526 ;
  assign n10528 = ~n10523 & n10527 ;
  assign n10529 = n10498 & n10508 ;
  assign n10530 = n10507 & ~n10529 ;
  assign n10531 = ~n10528 & n10530 ;
  assign n10532 = ~n10524 & n10525 ;
  assign n10533 = n10477 & ~n10522 ;
  assign n10534 = ( n10521 & n10530 ) | ( n10521 & n10533 ) | ( n10530 & n10533 ) ;
  assign n10535 = n10530 | n10533 ;
  assign n10536 = ( ~n10532 & n10534 ) | ( ~n10532 & n10535 ) | ( n10534 & n10535 ) ;
  assign n10537 = n10521 | n10533 ;
  assign n10538 = n10532 & ~n10537 ;
  assign n10539 = ( ~n10533 & n10536 ) | ( ~n10533 & n10538 ) | ( n10536 & n10538 ) ;
  assign n10540 = ( ~n10531 & n10536 ) | ( ~n10531 & n10539 ) | ( n10536 & n10539 ) ;
  assign n10541 = n10520 & n10540 ;
  assign n10542 = n10514 & n10518 ;
  assign n10543 = ( n10449 & n10514 ) | ( n10449 & n10542 ) | ( n10514 & n10542 ) ;
  assign n10544 = n10541 | n10543 ;
  assign n10545 = n10521 & ~n10533 ;
  assign n10546 = ( n10532 & n10533 ) | ( n10532 & ~n10545 ) | ( n10533 & ~n10545 ) ;
  assign n10547 = n10530 & n10546 ;
  assign n10548 = ~n10498 & n10508 ;
  assign n10549 = ( ~n10507 & n10508 ) | ( ~n10507 & n10548 ) | ( n10508 & n10548 ) ;
  assign n10550 = ~n10480 & n10481 ;
  assign n10551 = ( ~n10477 & n10481 ) | ( ~n10477 & n10550 ) | ( n10481 & n10550 ) ;
  assign n10552 = ~n10549 & n10551 ;
  assign n10553 = n10549 & ~n10551 ;
  assign n10554 = n10552 | n10553 ;
  assign n10555 = n10528 | n10554 ;
  assign n10556 = n10547 | n10555 ;
  assign n10557 = n10528 & n10554 ;
  assign n10558 = ( n10547 & n10554 ) | ( n10547 & n10557 ) | ( n10554 & n10557 ) ;
  assign n10559 = n10556 & ~n10558 ;
  assign n10560 = n10410 & n10448 ;
  assign n10561 = ~n10407 & n10408 ;
  assign n10562 = ( ~n10404 & n10408 ) | ( ~n10404 & n10561 ) | ( n10408 & n10561 ) ;
  assign n10563 = ~n10426 & n10430 ;
  assign n10564 = ( n10430 & ~n10438 ) | ( n10430 & n10563 ) | ( ~n10438 & n10563 ) ;
  assign n10565 = ~n10562 & n10564 ;
  assign n10566 = n10562 & ~n10564 ;
  assign n10567 = n10565 | n10566 ;
  assign n10568 = n10443 | n10567 ;
  assign n10569 = n10560 | n10568 ;
  assign n10570 = n10443 & n10567 ;
  assign n10571 = ( n10560 & n10567 ) | ( n10560 & n10570 ) | ( n10567 & n10570 ) ;
  assign n10572 = n10569 & ~n10571 ;
  assign n10573 = n10559 | n10572 ;
  assign n10574 = n10544 & n10573 ;
  assign n10575 = n10556 & n10569 ;
  assign n10576 = n10558 | n10571 ;
  assign n10577 = n10575 & ~n10576 ;
  assign n10578 = ( n10443 & n10562 ) | ( n10443 & n10564 ) | ( n10562 & n10564 ) ;
  assign n10579 = n10562 | n10564 ;
  assign n10580 = ( n10560 & n10578 ) | ( n10560 & n10579 ) | ( n10578 & n10579 ) ;
  assign n10581 = ( n10528 & n10549 ) | ( n10528 & n10551 ) | ( n10549 & n10551 ) ;
  assign n10582 = n10549 | n10551 ;
  assign n10583 = ( n10547 & n10581 ) | ( n10547 & n10582 ) | ( n10581 & n10582 ) ;
  assign n10584 = ~n10580 & n10583 ;
  assign n10585 = n10580 & ~n10583 ;
  assign n10586 = n10584 | n10585 ;
  assign n10587 = n10577 | n10586 ;
  assign n10588 = n10574 | n10587 ;
  assign n10589 = n10573 | n10577 ;
  assign n10590 = ( n10544 & n10577 ) | ( n10544 & n10589 ) | ( n10577 & n10589 ) ;
  assign n10591 = n10586 & n10590 ;
  assign n10592 = n10588 & ~n10591 ;
  assign n10593 = n10383 | n10592 ;
  assign n10594 = n10311 & ~n10334 ;
  assign n10595 = n10331 & ~n10594 ;
  assign n10596 = n10247 & ~n10304 ;
  assign n10597 = ~n10247 & n10304 ;
  assign n10598 = n10596 | n10597 ;
  assign n10599 = n10456 & ~n10513 ;
  assign n10600 = ~n10456 & n10513 ;
  assign n10601 = n10599 | n10600 ;
  assign n10602 = n10598 & n10601 ;
  assign n10603 = ~n10305 & n10311 ;
  assign n10604 = n10311 & ~n10331 ;
  assign n10605 = n10240 | n10309 ;
  assign n10606 = n10331 | n10605 ;
  assign n10607 = ( n10603 & n10604 ) | ( n10603 & ~n10606 ) | ( n10604 & ~n10606 ) ;
  assign n10608 = n10602 | n10607 ;
  assign n10609 = n10595 | n10608 ;
  assign n10610 = n10449 | n10518 ;
  assign n10611 = ( n10514 & n10540 ) | ( n10514 & ~n10610 ) | ( n10540 & ~n10610 ) ;
  assign n10612 = ( ~n10540 & n10610 ) | ( ~n10540 & n10611 ) | ( n10610 & n10611 ) ;
  assign n10613 = ( ~n10514 & n10611 ) | ( ~n10514 & n10612 ) | ( n10611 & n10612 ) ;
  assign n10614 = n10609 & n10613 ;
  assign n10615 = n10595 | n10607 ;
  assign n10616 = n10602 & n10615 ;
  assign n10617 = ( n10543 & ~n10559 ) | ( n10543 & n10572 ) | ( ~n10559 & n10572 ) ;
  assign n10618 = n10559 & ~n10572 ;
  assign n10619 = ( n10541 & n10617 ) | ( n10541 & ~n10618 ) | ( n10617 & ~n10618 ) ;
  assign n10620 = ( ~n10544 & n10559 ) | ( ~n10544 & n10619 ) | ( n10559 & n10619 ) ;
  assign n10621 = ( ~n10572 & n10619 ) | ( ~n10572 & n10620 ) | ( n10619 & n10620 ) ;
  assign n10622 = ( n10334 & ~n10350 ) | ( n10334 & n10363 ) | ( ~n10350 & n10363 ) ;
  assign n10623 = n10350 & ~n10363 ;
  assign n10624 = ( n10332 & n10622 ) | ( n10332 & ~n10623 ) | ( n10622 & ~n10623 ) ;
  assign n10625 = ( ~n10335 & n10350 ) | ( ~n10335 & n10624 ) | ( n10350 & n10624 ) ;
  assign n10626 = ( ~n10363 & n10624 ) | ( ~n10363 & n10625 ) | ( n10624 & n10625 ) ;
  assign n10627 = ( n10616 & n10621 ) | ( n10616 & n10626 ) | ( n10621 & n10626 ) ;
  assign n10628 = n10621 | n10626 ;
  assign n10629 = ( n10614 & n10627 ) | ( n10614 & n10628 ) | ( n10627 & n10628 ) ;
  assign n10630 = n10593 & n10629 ;
  assign n10631 = n10379 & n10588 ;
  assign n10632 = n10382 | n10591 ;
  assign n10633 = n10631 & ~n10632 ;
  assign n10634 = n10580 & n10583 ;
  assign n10635 = n10580 | n10583 ;
  assign n10636 = n10634 | n10635 ;
  assign n10637 = ( n10590 & n10634 ) | ( n10590 & n10636 ) | ( n10634 & n10636 ) ;
  assign n10638 = n10371 & n10374 ;
  assign n10639 = n10371 | n10374 ;
  assign n10640 = n10638 | n10639 ;
  assign n10641 = ( n10381 & n10638 ) | ( n10381 & n10640 ) | ( n10638 & n10640 ) ;
  assign n10642 = n10637 & n10641 ;
  assign n10643 = n10641 & ~n10642 ;
  assign n10644 = ( n10637 & ~n10642 ) | ( n10637 & n10643 ) | ( ~n10642 & n10643 ) ;
  assign n10645 = n10633 | n10644 ;
  assign n10646 = n10630 | n10645 ;
  assign n10647 = n10630 | n10633 ;
  assign n10648 = n10644 & n10647 ;
  assign n10649 = n10646 & ~n10648 ;
  assign n10650 = ~x835 & x836 ;
  assign n10651 = x835 & ~x836 ;
  assign n10652 = n10650 | n10651 ;
  assign n10653 = ~x837 & n10652 ;
  assign n10654 = x837 & ~n10652 ;
  assign n10655 = n10653 | n10654 ;
  assign n10656 = ~x838 & x839 ;
  assign n10657 = x838 & ~x839 ;
  assign n10658 = n10656 | n10657 ;
  assign n10659 = ~x840 & n10658 ;
  assign n10660 = x840 & ~n10658 ;
  assign n10661 = n10659 | n10660 ;
  assign n10662 = n10655 & n10661 ;
  assign n10663 = ( x838 & x839 ) | ( x838 & x840 ) | ( x839 & x840 ) ;
  assign n10664 = ( x835 & x836 ) | ( x835 & x837 ) | ( x836 & x837 ) ;
  assign n10665 = ~n10663 & n10664 ;
  assign n10666 = n10663 & ~n10664 ;
  assign n10667 = n10665 | n10666 ;
  assign n10668 = ~n10662 & n10667 ;
  assign n10669 = n10662 & ~n10667 ;
  assign n10670 = n10668 | n10669 ;
  assign n10671 = n10655 & ~n10661 ;
  assign n10672 = ~n10655 & n10661 ;
  assign n10673 = n10671 | n10672 ;
  assign n10674 = ( n10662 & n10663 ) | ( n10662 & n10664 ) | ( n10663 & n10664 ) ;
  assign n10675 = n10673 & n10674 ;
  assign n10676 = n10670 & ~n10675 ;
  assign n10677 = n10670 & n10674 ;
  assign n10678 = x841 & ~x842 ;
  assign n10679 = ~x841 & x842 ;
  assign n10680 = n10678 | n10679 ;
  assign n10681 = ~x843 & n10680 ;
  assign n10682 = x843 & ~n10680 ;
  assign n10683 = n10681 | n10682 ;
  assign n10684 = x844 & ~x845 ;
  assign n10685 = ~x844 & x845 ;
  assign n10686 = n10684 | n10685 ;
  assign n10687 = ~x846 & n10686 ;
  assign n10688 = x846 & ~n10686 ;
  assign n10689 = n10687 | n10688 ;
  assign n10690 = n10683 & ~n10689 ;
  assign n10691 = ~n10683 & n10689 ;
  assign n10692 = n10690 | n10691 ;
  assign n10693 = ( x844 & x845 ) | ( x844 & x846 ) | ( x845 & x846 ) ;
  assign n10694 = ( x841 & x842 ) | ( x841 & x843 ) | ( x842 & x843 ) ;
  assign n10695 = n10683 & n10689 ;
  assign n10696 = ( n10693 & n10694 ) | ( n10693 & n10695 ) | ( n10694 & n10695 ) ;
  assign n10697 = n10692 & n10696 ;
  assign n10698 = n10677 | n10697 ;
  assign n10699 = n10693 & ~n10694 ;
  assign n10700 = ~n10693 & n10694 ;
  assign n10701 = n10699 | n10700 ;
  assign n10702 = ~n10695 & n10701 ;
  assign n10703 = n10695 & ~n10701 ;
  assign n10704 = n10702 | n10703 ;
  assign n10705 = n10696 & n10704 ;
  assign n10706 = n10673 & n10692 ;
  assign n10707 = n10704 & n10706 ;
  assign n10708 = ~n10705 & n10707 ;
  assign n10709 = ~n10698 & n10708 ;
  assign n10710 = n10676 & n10709 ;
  assign n10711 = ~n10705 & n10706 ;
  assign n10712 = ~n10697 & n10704 ;
  assign n10713 = n10677 & ~n10712 ;
  assign n10714 = ( n10711 & n10712 ) | ( n10711 & ~n10713 ) | ( n10712 & ~n10713 ) ;
  assign n10715 = ( n10676 & n10710 ) | ( n10676 & ~n10714 ) | ( n10710 & ~n10714 ) ;
  assign n10716 = n10692 & ~n10696 ;
  assign n10717 = ( n10692 & ~n10704 ) | ( n10692 & n10716 ) | ( ~n10704 & n10716 ) ;
  assign n10718 = n10673 & ~n10674 ;
  assign n10719 = ( ~n10670 & n10673 ) | ( ~n10670 & n10718 ) | ( n10673 & n10718 ) ;
  assign n10720 = ~n10717 & n10719 ;
  assign n10721 = n10717 & ~n10719 ;
  assign n10722 = n10720 | n10721 ;
  assign n10723 = ( x832 & x833 ) | ( x832 & x834 ) | ( x833 & x834 ) ;
  assign n10724 = ( x829 & x830 ) | ( x829 & x831 ) | ( x830 & x831 ) ;
  assign n10725 = n10723 & ~n10724 ;
  assign n10726 = ~n10723 & n10724 ;
  assign n10727 = n10725 | n10726 ;
  assign n10728 = x829 & ~x830 ;
  assign n10729 = ~x829 & x830 ;
  assign n10730 = n10728 | n10729 ;
  assign n10731 = ~x831 & n10730 ;
  assign n10732 = x831 & ~n10730 ;
  assign n10733 = n10731 | n10732 ;
  assign n10734 = x832 & ~x833 ;
  assign n10735 = ~x832 & x833 ;
  assign n10736 = n10734 | n10735 ;
  assign n10737 = ~x834 & n10736 ;
  assign n10738 = x834 & ~n10736 ;
  assign n10739 = n10737 | n10738 ;
  assign n10740 = n10733 & n10739 ;
  assign n10741 = n10727 & ~n10740 ;
  assign n10742 = ~n10727 & n10740 ;
  assign n10743 = n10741 | n10742 ;
  assign n10744 = n10733 & ~n10739 ;
  assign n10745 = ~n10733 & n10739 ;
  assign n10746 = n10744 | n10745 ;
  assign n10747 = ( n10723 & n10724 ) | ( n10723 & n10740 ) | ( n10724 & n10740 ) ;
  assign n10748 = n10746 & ~n10747 ;
  assign n10749 = ( ~n10743 & n10746 ) | ( ~n10743 & n10748 ) | ( n10746 & n10748 ) ;
  assign n10750 = ~x823 & x824 ;
  assign n10751 = x823 & ~x824 ;
  assign n10752 = n10750 | n10751 ;
  assign n10753 = ~x825 & n10752 ;
  assign n10754 = x825 & ~n10752 ;
  assign n10755 = n10753 | n10754 ;
  assign n10756 = ~x826 & x827 ;
  assign n10757 = x826 & ~x827 ;
  assign n10758 = n10756 | n10757 ;
  assign n10759 = ~x828 & n10758 ;
  assign n10760 = x828 & ~n10758 ;
  assign n10761 = n10759 | n10760 ;
  assign n10762 = n10755 & n10761 ;
  assign n10763 = ( x826 & x827 ) | ( x826 & x828 ) | ( x827 & x828 ) ;
  assign n10764 = ( x823 & x824 ) | ( x823 & x825 ) | ( x824 & x825 ) ;
  assign n10765 = ~n10763 & n10764 ;
  assign n10766 = n10763 & ~n10764 ;
  assign n10767 = n10765 | n10766 ;
  assign n10768 = ~n10762 & n10767 ;
  assign n10769 = n10762 & ~n10767 ;
  assign n10770 = n10768 | n10769 ;
  assign n10771 = n10755 & ~n10761 ;
  assign n10772 = ~n10755 & n10761 ;
  assign n10773 = n10771 | n10772 ;
  assign n10774 = ( n10762 & n10763 ) | ( n10762 & n10764 ) | ( n10763 & n10764 ) ;
  assign n10775 = n10773 & ~n10774 ;
  assign n10776 = ( ~n10770 & n10773 ) | ( ~n10770 & n10775 ) | ( n10773 & n10775 ) ;
  assign n10777 = ~n10749 & n10776 ;
  assign n10778 = n10749 & ~n10776 ;
  assign n10779 = n10777 | n10778 ;
  assign n10780 = n10722 & n10779 ;
  assign n10781 = ( n10676 & ~n10677 ) | ( n10676 & n10712 ) | ( ~n10677 & n10712 ) ;
  assign n10782 = n10676 & n10712 ;
  assign n10783 = ( n10711 & n10781 ) | ( n10711 & n10782 ) | ( n10781 & n10782 ) ;
  assign n10784 = n10714 & ~n10783 ;
  assign n10785 = n10780 | n10784 ;
  assign n10786 = n10715 | n10785 ;
  assign n10787 = n10770 & n10774 ;
  assign n10788 = n10746 & n10747 ;
  assign n10789 = n10787 | n10788 ;
  assign n10790 = n10743 & n10747 ;
  assign n10791 = n10746 & n10773 ;
  assign n10792 = n10743 & n10791 ;
  assign n10793 = ~n10790 & n10792 ;
  assign n10794 = ~n10789 & n10793 ;
  assign n10795 = n10773 & n10774 ;
  assign n10796 = n10770 & ~n10795 ;
  assign n10797 = ~n10794 & n10796 ;
  assign n10798 = ~n10790 & n10791 ;
  assign n10799 = n10743 & ~n10788 ;
  assign n10800 = ( n10787 & n10796 ) | ( n10787 & n10799 ) | ( n10796 & n10799 ) ;
  assign n10801 = n10796 | n10799 ;
  assign n10802 = ( ~n10798 & n10800 ) | ( ~n10798 & n10801 ) | ( n10800 & n10801 ) ;
  assign n10803 = n10787 | n10799 ;
  assign n10804 = n10798 & ~n10803 ;
  assign n10805 = ( ~n10799 & n10802 ) | ( ~n10799 & n10804 ) | ( n10802 & n10804 ) ;
  assign n10806 = ( ~n10797 & n10802 ) | ( ~n10797 & n10805 ) | ( n10802 & n10805 ) ;
  assign n10807 = n10786 & n10806 ;
  assign n10808 = n10780 & n10784 ;
  assign n10809 = ( n10715 & n10780 ) | ( n10715 & n10808 ) | ( n10780 & n10808 ) ;
  assign n10810 = n10807 | n10809 ;
  assign n10811 = n10787 & ~n10799 ;
  assign n10812 = ( n10798 & n10799 ) | ( n10798 & ~n10811 ) | ( n10799 & ~n10811 ) ;
  assign n10813 = n10796 & n10812 ;
  assign n10814 = ~n10773 & n10774 ;
  assign n10815 = ( ~n10770 & n10774 ) | ( ~n10770 & n10814 ) | ( n10774 & n10814 ) ;
  assign n10816 = ~n10746 & n10747 ;
  assign n10817 = ( ~n10743 & n10747 ) | ( ~n10743 & n10816 ) | ( n10747 & n10816 ) ;
  assign n10818 = ~n10815 & n10817 ;
  assign n10819 = n10815 & ~n10817 ;
  assign n10820 = n10818 | n10819 ;
  assign n10821 = n10794 | n10820 ;
  assign n10822 = n10813 | n10821 ;
  assign n10823 = n10794 & n10820 ;
  assign n10824 = ( n10813 & n10820 ) | ( n10813 & n10823 ) | ( n10820 & n10823 ) ;
  assign n10825 = n10822 & ~n10824 ;
  assign n10826 = n10676 & n10714 ;
  assign n10827 = ~n10673 & n10674 ;
  assign n10828 = ( ~n10670 & n10674 ) | ( ~n10670 & n10827 ) | ( n10674 & n10827 ) ;
  assign n10829 = ~n10692 & n10696 ;
  assign n10830 = ( n10696 & ~n10704 ) | ( n10696 & n10829 ) | ( ~n10704 & n10829 ) ;
  assign n10831 = ~n10828 & n10830 ;
  assign n10832 = n10828 & ~n10830 ;
  assign n10833 = n10831 | n10832 ;
  assign n10834 = n10709 | n10833 ;
  assign n10835 = n10826 | n10834 ;
  assign n10836 = n10709 & n10833 ;
  assign n10837 = ( n10826 & n10833 ) | ( n10826 & n10836 ) | ( n10833 & n10836 ) ;
  assign n10838 = n10835 & ~n10837 ;
  assign n10839 = n10825 | n10838 ;
  assign n10840 = n10810 & n10839 ;
  assign n10841 = n10822 & n10835 ;
  assign n10842 = n10824 | n10837 ;
  assign n10843 = n10841 & ~n10842 ;
  assign n10844 = ( n10709 & n10828 ) | ( n10709 & n10830 ) | ( n10828 & n10830 ) ;
  assign n10845 = n10828 | n10830 ;
  assign n10846 = ( n10826 & n10844 ) | ( n10826 & n10845 ) | ( n10844 & n10845 ) ;
  assign n10847 = ( n10794 & n10815 ) | ( n10794 & n10817 ) | ( n10815 & n10817 ) ;
  assign n10848 = n10815 | n10817 ;
  assign n10849 = ( n10813 & n10847 ) | ( n10813 & n10848 ) | ( n10847 & n10848 ) ;
  assign n10850 = ~n10846 & n10849 ;
  assign n10851 = n10846 & ~n10849 ;
  assign n10852 = n10850 | n10851 ;
  assign n10853 = n10843 | n10852 ;
  assign n10854 = n10840 | n10853 ;
  assign n10855 = n10839 | n10843 ;
  assign n10856 = ( n10810 & n10843 ) | ( n10810 & n10855 ) | ( n10843 & n10855 ) ;
  assign n10857 = n10852 & n10856 ;
  assign n10858 = n10854 & ~n10857 ;
  assign n10859 = ~x811 & x812 ;
  assign n10860 = x811 & ~x812 ;
  assign n10861 = n10859 | n10860 ;
  assign n10862 = ~x813 & n10861 ;
  assign n10863 = x813 & ~n10861 ;
  assign n10864 = n10862 | n10863 ;
  assign n10865 = ~x814 & x815 ;
  assign n10866 = x814 & ~x815 ;
  assign n10867 = n10865 | n10866 ;
  assign n10868 = ~x816 & n10867 ;
  assign n10869 = x816 & ~n10867 ;
  assign n10870 = n10868 | n10869 ;
  assign n10871 = n10864 & n10870 ;
  assign n10872 = ( x814 & x815 ) | ( x814 & x816 ) | ( x815 & x816 ) ;
  assign n10873 = ( x811 & x812 ) | ( x811 & x813 ) | ( x812 & x813 ) ;
  assign n10874 = ~n10872 & n10873 ;
  assign n10875 = n10872 & ~n10873 ;
  assign n10876 = n10874 | n10875 ;
  assign n10877 = ~n10871 & n10876 ;
  assign n10878 = n10871 & ~n10876 ;
  assign n10879 = n10877 | n10878 ;
  assign n10880 = n10864 & ~n10870 ;
  assign n10881 = ~n10864 & n10870 ;
  assign n10882 = n10880 | n10881 ;
  assign n10883 = ( n10871 & n10872 ) | ( n10871 & n10873 ) | ( n10872 & n10873 ) ;
  assign n10884 = n10882 & n10883 ;
  assign n10885 = n10879 & ~n10884 ;
  assign n10886 = n10879 & n10883 ;
  assign n10887 = x817 & ~x818 ;
  assign n10888 = ~x817 & x818 ;
  assign n10889 = n10887 | n10888 ;
  assign n10890 = ~x819 & n10889 ;
  assign n10891 = x819 & ~n10889 ;
  assign n10892 = n10890 | n10891 ;
  assign n10893 = x820 & ~x821 ;
  assign n10894 = ~x820 & x821 ;
  assign n10895 = n10893 | n10894 ;
  assign n10896 = ~x822 & n10895 ;
  assign n10897 = x822 & ~n10895 ;
  assign n10898 = n10896 | n10897 ;
  assign n10899 = n10892 & ~n10898 ;
  assign n10900 = ~n10892 & n10898 ;
  assign n10901 = n10899 | n10900 ;
  assign n10902 = ( x820 & x821 ) | ( x820 & x822 ) | ( x821 & x822 ) ;
  assign n10903 = ( x817 & x818 ) | ( x817 & x819 ) | ( x818 & x819 ) ;
  assign n10904 = n10892 & n10898 ;
  assign n10905 = ( n10902 & n10903 ) | ( n10902 & n10904 ) | ( n10903 & n10904 ) ;
  assign n10906 = n10901 & n10905 ;
  assign n10907 = n10886 | n10906 ;
  assign n10908 = n10902 & ~n10903 ;
  assign n10909 = ~n10902 & n10903 ;
  assign n10910 = n10908 | n10909 ;
  assign n10911 = ~n10904 & n10910 ;
  assign n10912 = n10904 & ~n10910 ;
  assign n10913 = n10911 | n10912 ;
  assign n10914 = n10905 & n10913 ;
  assign n10915 = n10882 & n10901 ;
  assign n10916 = n10913 & n10915 ;
  assign n10917 = ~n10914 & n10916 ;
  assign n10918 = ~n10907 & n10917 ;
  assign n10919 = n10885 & n10918 ;
  assign n10920 = ~n10914 & n10915 ;
  assign n10921 = ~n10906 & n10913 ;
  assign n10922 = n10886 & ~n10921 ;
  assign n10923 = ( n10920 & n10921 ) | ( n10920 & ~n10922 ) | ( n10921 & ~n10922 ) ;
  assign n10924 = ( n10885 & n10919 ) | ( n10885 & ~n10923 ) | ( n10919 & ~n10923 ) ;
  assign n10925 = n10901 & ~n10905 ;
  assign n10926 = ( n10901 & ~n10913 ) | ( n10901 & n10925 ) | ( ~n10913 & n10925 ) ;
  assign n10927 = n10882 & ~n10883 ;
  assign n10928 = ( ~n10879 & n10882 ) | ( ~n10879 & n10927 ) | ( n10882 & n10927 ) ;
  assign n10929 = ~n10926 & n10928 ;
  assign n10930 = n10926 & ~n10928 ;
  assign n10931 = n10929 | n10930 ;
  assign n10932 = ( x808 & x809 ) | ( x808 & x810 ) | ( x809 & x810 ) ;
  assign n10933 = ( x805 & x806 ) | ( x805 & x807 ) | ( x806 & x807 ) ;
  assign n10934 = n10932 & ~n10933 ;
  assign n10935 = ~n10932 & n10933 ;
  assign n10936 = n10934 | n10935 ;
  assign n10937 = ~x805 & x806 ;
  assign n10938 = x805 & ~x806 ;
  assign n10939 = n10937 | n10938 ;
  assign n10940 = ~x807 & n10939 ;
  assign n10941 = x807 & ~n10939 ;
  assign n10942 = n10940 | n10941 ;
  assign n10943 = ~x808 & x809 ;
  assign n10944 = x808 & ~x809 ;
  assign n10945 = n10943 | n10944 ;
  assign n10946 = ~x810 & n10945 ;
  assign n10947 = x810 & ~n10945 ;
  assign n10948 = n10946 | n10947 ;
  assign n10949 = n10942 & n10948 ;
  assign n10950 = n10936 & ~n10949 ;
  assign n10951 = ~n10936 & n10949 ;
  assign n10952 = n10950 | n10951 ;
  assign n10953 = n10942 & ~n10948 ;
  assign n10954 = ~n10942 & n10948 ;
  assign n10955 = n10953 | n10954 ;
  assign n10956 = ( n10932 & n10933 ) | ( n10932 & n10949 ) | ( n10933 & n10949 ) ;
  assign n10957 = n10955 & ~n10956 ;
  assign n10958 = ( ~n10952 & n10955 ) | ( ~n10952 & n10957 ) | ( n10955 & n10957 ) ;
  assign n10959 = ~x799 & x800 ;
  assign n10960 = x799 & ~x800 ;
  assign n10961 = n10959 | n10960 ;
  assign n10962 = ~x801 & n10961 ;
  assign n10963 = x801 & ~n10961 ;
  assign n10964 = n10962 | n10963 ;
  assign n10965 = ~x802 & x803 ;
  assign n10966 = x802 & ~x803 ;
  assign n10967 = n10965 | n10966 ;
  assign n10968 = ~x804 & n10967 ;
  assign n10969 = x804 & ~n10967 ;
  assign n10970 = n10968 | n10969 ;
  assign n10971 = n10964 & ~n10970 ;
  assign n10972 = ~n10964 & n10970 ;
  assign n10973 = n10971 | n10972 ;
  assign n10974 = ( x802 & x803 ) | ( x802 & x804 ) | ( x803 & x804 ) ;
  assign n10975 = ( x799 & x800 ) | ( x799 & x801 ) | ( x800 & x801 ) ;
  assign n10976 = n10974 & ~n10975 ;
  assign n10977 = ~n10974 & n10975 ;
  assign n10978 = n10976 | n10977 ;
  assign n10979 = n10964 & n10970 ;
  assign n10980 = n10978 & ~n10979 ;
  assign n10981 = ~n10978 & n10979 ;
  assign n10982 = n10980 | n10981 ;
  assign n10983 = ( n10974 & n10975 ) | ( n10974 & n10979 ) | ( n10975 & n10979 ) ;
  assign n10984 = n10973 & ~n10983 ;
  assign n10985 = ( n10973 & ~n10982 ) | ( n10973 & n10984 ) | ( ~n10982 & n10984 ) ;
  assign n10986 = ~n10958 & n10985 ;
  assign n10987 = n10958 & ~n10985 ;
  assign n10988 = n10986 | n10987 ;
  assign n10989 = n10931 & n10988 ;
  assign n10990 = ( n10885 & ~n10886 ) | ( n10885 & n10921 ) | ( ~n10886 & n10921 ) ;
  assign n10991 = n10885 & n10921 ;
  assign n10992 = ( n10920 & n10990 ) | ( n10920 & n10991 ) | ( n10990 & n10991 ) ;
  assign n10993 = n10923 & ~n10992 ;
  assign n10994 = n10989 | n10993 ;
  assign n10995 = n10924 | n10994 ;
  assign n10996 = n10982 & n10983 ;
  assign n10997 = n10955 & n10956 ;
  assign n10998 = n10996 | n10997 ;
  assign n10999 = n10952 & n10956 ;
  assign n11000 = n10955 & n10973 ;
  assign n11001 = n10952 & n11000 ;
  assign n11002 = ~n10999 & n11001 ;
  assign n11003 = ~n10998 & n11002 ;
  assign n11004 = n10973 & n10983 ;
  assign n11005 = n10982 & ~n11004 ;
  assign n11006 = ~n11003 & n11005 ;
  assign n11007 = ~n10999 & n11000 ;
  assign n11008 = n10952 & ~n10997 ;
  assign n11009 = ( n10996 & n11005 ) | ( n10996 & n11008 ) | ( n11005 & n11008 ) ;
  assign n11010 = n11005 | n11008 ;
  assign n11011 = ( ~n11007 & n11009 ) | ( ~n11007 & n11010 ) | ( n11009 & n11010 ) ;
  assign n11012 = n10996 | n11008 ;
  assign n11013 = n11007 & ~n11012 ;
  assign n11014 = ( ~n11008 & n11011 ) | ( ~n11008 & n11013 ) | ( n11011 & n11013 ) ;
  assign n11015 = ( ~n11006 & n11011 ) | ( ~n11006 & n11014 ) | ( n11011 & n11014 ) ;
  assign n11016 = n10995 & n11015 ;
  assign n11017 = n10989 & n10993 ;
  assign n11018 = ( n10924 & n10989 ) | ( n10924 & n11017 ) | ( n10989 & n11017 ) ;
  assign n11019 = n11016 | n11018 ;
  assign n11020 = n10996 & ~n11008 ;
  assign n11021 = ( n11007 & n11008 ) | ( n11007 & ~n11020 ) | ( n11008 & ~n11020 ) ;
  assign n11022 = n11005 & n11021 ;
  assign n11023 = ~n10973 & n10983 ;
  assign n11024 = ( ~n10982 & n10983 ) | ( ~n10982 & n11023 ) | ( n10983 & n11023 ) ;
  assign n11025 = ~n10955 & n10956 ;
  assign n11026 = ( ~n10952 & n10956 ) | ( ~n10952 & n11025 ) | ( n10956 & n11025 ) ;
  assign n11027 = ~n11024 & n11026 ;
  assign n11028 = n11024 & ~n11026 ;
  assign n11029 = n11027 | n11028 ;
  assign n11030 = n11003 | n11029 ;
  assign n11031 = n11022 | n11030 ;
  assign n11032 = n11003 & n11029 ;
  assign n11033 = ( n11022 & n11029 ) | ( n11022 & n11032 ) | ( n11029 & n11032 ) ;
  assign n11034 = n11031 & ~n11033 ;
  assign n11035 = n10885 & n10923 ;
  assign n11036 = ~n10882 & n10883 ;
  assign n11037 = ( ~n10879 & n10883 ) | ( ~n10879 & n11036 ) | ( n10883 & n11036 ) ;
  assign n11038 = ~n10901 & n10905 ;
  assign n11039 = ( n10905 & ~n10913 ) | ( n10905 & n11038 ) | ( ~n10913 & n11038 ) ;
  assign n11040 = ~n11037 & n11039 ;
  assign n11041 = n11037 & ~n11039 ;
  assign n11042 = n11040 | n11041 ;
  assign n11043 = n10918 | n11042 ;
  assign n11044 = n11035 | n11043 ;
  assign n11045 = n10918 & n11042 ;
  assign n11046 = ( n11035 & n11042 ) | ( n11035 & n11045 ) | ( n11042 & n11045 ) ;
  assign n11047 = n11044 & ~n11046 ;
  assign n11048 = n11034 | n11047 ;
  assign n11049 = n11019 & n11048 ;
  assign n11050 = n11031 & n11044 ;
  assign n11051 = n11033 | n11046 ;
  assign n11052 = n11050 & ~n11051 ;
  assign n11053 = ( n10918 & n11037 ) | ( n10918 & n11039 ) | ( n11037 & n11039 ) ;
  assign n11054 = n11037 | n11039 ;
  assign n11055 = ( n11035 & n11053 ) | ( n11035 & n11054 ) | ( n11053 & n11054 ) ;
  assign n11056 = ( n11003 & n11024 ) | ( n11003 & n11026 ) | ( n11024 & n11026 ) ;
  assign n11057 = n11024 | n11026 ;
  assign n11058 = ( n11022 & n11056 ) | ( n11022 & n11057 ) | ( n11056 & n11057 ) ;
  assign n11059 = ~n11055 & n11058 ;
  assign n11060 = n11055 & ~n11058 ;
  assign n11061 = n11059 | n11060 ;
  assign n11062 = n11052 | n11061 ;
  assign n11063 = n11049 | n11062 ;
  assign n11064 = n11048 | n11052 ;
  assign n11065 = ( n11019 & n11052 ) | ( n11019 & n11064 ) | ( n11052 & n11064 ) ;
  assign n11066 = n11061 & n11065 ;
  assign n11067 = n11063 & ~n11066 ;
  assign n11068 = n10858 | n11067 ;
  assign n11069 = n10786 & ~n10809 ;
  assign n11070 = n10806 & ~n11069 ;
  assign n11071 = n10722 & ~n10779 ;
  assign n11072 = ~n10722 & n10779 ;
  assign n11073 = n11071 | n11072 ;
  assign n11074 = n10931 & ~n10988 ;
  assign n11075 = ~n10931 & n10988 ;
  assign n11076 = n11074 | n11075 ;
  assign n11077 = n11073 & n11076 ;
  assign n11078 = ~n10780 & n10786 ;
  assign n11079 = n10786 & ~n10806 ;
  assign n11080 = n10715 | n10784 ;
  assign n11081 = n10806 | n11080 ;
  assign n11082 = ( n11078 & n11079 ) | ( n11078 & ~n11081 ) | ( n11079 & ~n11081 ) ;
  assign n11083 = n11077 | n11082 ;
  assign n11084 = n11070 | n11083 ;
  assign n11085 = n10924 | n10993 ;
  assign n11086 = ( n10989 & n11015 ) | ( n10989 & ~n11085 ) | ( n11015 & ~n11085 ) ;
  assign n11087 = ( ~n11015 & n11085 ) | ( ~n11015 & n11086 ) | ( n11085 & n11086 ) ;
  assign n11088 = ( ~n10989 & n11086 ) | ( ~n10989 & n11087 ) | ( n11086 & n11087 ) ;
  assign n11089 = n11084 & n11088 ;
  assign n11090 = n11070 | n11082 ;
  assign n11091 = n11077 & n11090 ;
  assign n11092 = ( n11018 & ~n11034 ) | ( n11018 & n11047 ) | ( ~n11034 & n11047 ) ;
  assign n11093 = n11034 & ~n11047 ;
  assign n11094 = ( n11016 & n11092 ) | ( n11016 & ~n11093 ) | ( n11092 & ~n11093 ) ;
  assign n11095 = ( ~n11019 & n11034 ) | ( ~n11019 & n11094 ) | ( n11034 & n11094 ) ;
  assign n11096 = ( ~n11047 & n11094 ) | ( ~n11047 & n11095 ) | ( n11094 & n11095 ) ;
  assign n11097 = ( n10809 & ~n10825 ) | ( n10809 & n10838 ) | ( ~n10825 & n10838 ) ;
  assign n11098 = n10825 & ~n10838 ;
  assign n11099 = ( n10807 & n11097 ) | ( n10807 & ~n11098 ) | ( n11097 & ~n11098 ) ;
  assign n11100 = ( ~n10810 & n10825 ) | ( ~n10810 & n11099 ) | ( n10825 & n11099 ) ;
  assign n11101 = ( ~n10838 & n11099 ) | ( ~n10838 & n11100 ) | ( n11099 & n11100 ) ;
  assign n11102 = ( n11091 & n11096 ) | ( n11091 & n11101 ) | ( n11096 & n11101 ) ;
  assign n11103 = n11096 | n11101 ;
  assign n11104 = ( n11089 & n11102 ) | ( n11089 & n11103 ) | ( n11102 & n11103 ) ;
  assign n11105 = n11068 & n11104 ;
  assign n11106 = n10854 & n11063 ;
  assign n11107 = n10857 | n11066 ;
  assign n11108 = n11106 & ~n11107 ;
  assign n11109 = n11055 & n11058 ;
  assign n11110 = n11055 | n11058 ;
  assign n11111 = n11109 | n11110 ;
  assign n11112 = ( n11065 & n11109 ) | ( n11065 & n11111 ) | ( n11109 & n11111 ) ;
  assign n11113 = n10846 & n10849 ;
  assign n11114 = n10846 | n10849 ;
  assign n11115 = n11113 | n11114 ;
  assign n11116 = ( n10856 & n11113 ) | ( n10856 & n11115 ) | ( n11113 & n11115 ) ;
  assign n11117 = n11112 & n11116 ;
  assign n11118 = n11116 & ~n11117 ;
  assign n11119 = ( n11112 & ~n11117 ) | ( n11112 & n11118 ) | ( ~n11117 & n11118 ) ;
  assign n11120 = n11108 | n11119 ;
  assign n11121 = n11105 | n11120 ;
  assign n11122 = n11105 | n11108 ;
  assign n11123 = n11119 & n11122 ;
  assign n11124 = n11121 & ~n11123 ;
  assign n11125 = n10649 | n11124 ;
  assign n11126 = ( ~n10858 & n11067 ) | ( ~n10858 & n11104 ) | ( n11067 & n11104 ) ;
  assign n11127 = ( n10858 & ~n11104 ) | ( n10858 & n11126 ) | ( ~n11104 & n11126 ) ;
  assign n11128 = ( ~n11067 & n11126 ) | ( ~n11067 & n11127 ) | ( n11126 & n11127 ) ;
  assign n11129 = ( ~n10383 & n10592 ) | ( ~n10383 & n10629 ) | ( n10592 & n10629 ) ;
  assign n11130 = ( n10383 & ~n10629 ) | ( n10383 & n11129 ) | ( ~n10629 & n11129 ) ;
  assign n11131 = ( ~n10592 & n11129 ) | ( ~n10592 & n11130 ) | ( n11129 & n11130 ) ;
  assign n11132 = ~n10602 & n10615 ;
  assign n11133 = n10602 & ~n10607 ;
  assign n11134 = ~n10595 & n11133 ;
  assign n11135 = ~n10613 & n11134 ;
  assign n11136 = ( ~n10613 & n11132 ) | ( ~n10613 & n11135 ) | ( n11132 & n11135 ) ;
  assign n11137 = n10614 & ~n10616 ;
  assign n11138 = ( n10613 & n11136 ) | ( n10613 & ~n11137 ) | ( n11136 & ~n11137 ) ;
  assign n11139 = n11073 & ~n11076 ;
  assign n11140 = ~n11073 & n11076 ;
  assign n11141 = n11139 | n11140 ;
  assign n11142 = n10598 & ~n10601 ;
  assign n11143 = ~n10598 & n10601 ;
  assign n11144 = n11142 | n11143 ;
  assign n11145 = n11141 & n11144 ;
  assign n11146 = ~n11084 & n11088 ;
  assign n11147 = ( n11088 & n11091 ) | ( n11088 & n11146 ) | ( n11091 & n11146 ) ;
  assign n11148 = ~n11077 & n11090 ;
  assign n11149 = n11077 & ~n11082 ;
  assign n11150 = ~n11070 & n11149 ;
  assign n11151 = ~n11088 & n11150 ;
  assign n11152 = ( ~n11088 & n11148 ) | ( ~n11088 & n11151 ) | ( n11148 & n11151 ) ;
  assign n11153 = n11147 | n11152 ;
  assign n11154 = n11145 | n11153 ;
  assign n11155 = n11138 & n11154 ;
  assign n11156 = n11145 & n11153 ;
  assign n11158 = ( n10616 & ~n10621 ) | ( n10616 & n10626 ) | ( ~n10621 & n10626 ) ;
  assign n11159 = n10621 & ~n10626 ;
  assign n11160 = ( n10614 & n11158 ) | ( n10614 & ~n11159 ) | ( n11158 & ~n11159 ) ;
  assign n11157 = n10614 | n10616 ;
  assign n11161 = ( n10621 & ~n11157 ) | ( n10621 & n11160 ) | ( ~n11157 & n11160 ) ;
  assign n11162 = ( ~n10626 & n11160 ) | ( ~n10626 & n11161 ) | ( n11160 & n11161 ) ;
  assign n11164 = ( n11091 & ~n11096 ) | ( n11091 & n11101 ) | ( ~n11096 & n11101 ) ;
  assign n11165 = n11096 & ~n11101 ;
  assign n11166 = ( n11089 & n11164 ) | ( n11089 & ~n11165 ) | ( n11164 & ~n11165 ) ;
  assign n11163 = n11089 | n11091 ;
  assign n11167 = ( n11096 & ~n11163 ) | ( n11096 & n11166 ) | ( ~n11163 & n11166 ) ;
  assign n11168 = ( ~n11101 & n11166 ) | ( ~n11101 & n11167 ) | ( n11166 & n11167 ) ;
  assign n11169 = ( n11156 & n11162 ) | ( n11156 & n11168 ) | ( n11162 & n11168 ) ;
  assign n11170 = n11162 | n11168 ;
  assign n11171 = ( n11155 & n11169 ) | ( n11155 & n11170 ) | ( n11169 & n11170 ) ;
  assign n11172 = ( n11128 & n11131 ) | ( n11128 & n11171 ) | ( n11131 & n11171 ) ;
  assign n11173 = n11125 & n11172 ;
  assign n11174 = n10646 & n11121 ;
  assign n11175 = n10648 | n11123 ;
  assign n11176 = n11174 & ~n11175 ;
  assign n11185 = n10381 & n10639 ;
  assign n11186 = n10583 | n10638 ;
  assign n11187 = n10580 | n10638 ;
  assign n11188 = ( n10590 & n11186 ) | ( n10590 & n11187 ) | ( n11186 & n11187 ) ;
  assign n11189 = n11185 | n11188 ;
  assign n11190 = n10642 | n11189 ;
  assign n11191 = ( n10633 & n10642 ) | ( n10633 & n11190 ) | ( n10642 & n11190 ) ;
  assign n11192 = n10642 | n11190 ;
  assign n11193 = ( n10630 & n11191 ) | ( n10630 & n11192 ) | ( n11191 & n11192 ) ;
  assign n11177 = n10856 & n11114 ;
  assign n11178 = n11058 | n11113 ;
  assign n11179 = n11055 | n11113 ;
  assign n11180 = ( n11065 & n11178 ) | ( n11065 & n11179 ) | ( n11178 & n11179 ) ;
  assign n11181 = n11177 | n11180 ;
  assign n11182 = n11108 & n11181 ;
  assign n11183 = ( n11105 & n11181 ) | ( n11105 & n11182 ) | ( n11181 & n11182 ) ;
  assign n11184 = n11117 | n11183 ;
  assign n11194 = n11184 & n11193 ;
  assign n11195 = n11184 & ~n11194 ;
  assign n11196 = ( n11193 & ~n11194 ) | ( n11193 & n11195 ) | ( ~n11194 & n11195 ) ;
  assign n11197 = n11176 | n11196 ;
  assign n11198 = n11173 | n11197 ;
  assign n11199 = n11173 | n11176 ;
  assign n11200 = n11196 & n11199 ;
  assign n11201 = n11198 & ~n11200 ;
  assign n11202 = ( x694 & x695 ) | ( x694 & x696 ) | ( x695 & x696 ) ;
  assign n11203 = ( x691 & x692 ) | ( x691 & x693 ) | ( x692 & x693 ) ;
  assign n11204 = n11202 & ~n11203 ;
  assign n11205 = ~n11202 & n11203 ;
  assign n11206 = n11204 | n11205 ;
  assign n11207 = ~x691 & x692 ;
  assign n11208 = x691 & ~x692 ;
  assign n11209 = n11207 | n11208 ;
  assign n11210 = ~x693 & n11209 ;
  assign n11211 = x693 & ~n11209 ;
  assign n11212 = n11210 | n11211 ;
  assign n11213 = ~x694 & x695 ;
  assign n11214 = x694 & ~x695 ;
  assign n11215 = n11213 | n11214 ;
  assign n11216 = ~x696 & n11215 ;
  assign n11217 = x696 & ~n11215 ;
  assign n11218 = n11216 | n11217 ;
  assign n11219 = n11212 & n11218 ;
  assign n11220 = n11206 & ~n11219 ;
  assign n11221 = ~n11206 & n11219 ;
  assign n11222 = n11220 | n11221 ;
  assign n11223 = n11212 & ~n11218 ;
  assign n11224 = ~n11212 & n11218 ;
  assign n11225 = n11223 | n11224 ;
  assign n11226 = ( n11202 & n11203 ) | ( n11202 & n11219 ) | ( n11203 & n11219 ) ;
  assign n11227 = n11225 & n11226 ;
  assign n11228 = n11222 & ~n11227 ;
  assign n11229 = n11222 & n11226 ;
  assign n11230 = ~x697 & x698 ;
  assign n11231 = x697 & ~x698 ;
  assign n11232 = n11230 | n11231 ;
  assign n11233 = ~x699 & n11232 ;
  assign n11234 = x699 & ~n11232 ;
  assign n11235 = n11233 | n11234 ;
  assign n11236 = ~x700 & x701 ;
  assign n11237 = x700 & ~x701 ;
  assign n11238 = n11236 | n11237 ;
  assign n11239 = ~x702 & n11238 ;
  assign n11240 = x702 & ~n11238 ;
  assign n11241 = n11239 | n11240 ;
  assign n11242 = n11235 & ~n11241 ;
  assign n11243 = ~n11235 & n11241 ;
  assign n11244 = n11242 | n11243 ;
  assign n11245 = ( x700 & x701 ) | ( x700 & x702 ) | ( x701 & x702 ) ;
  assign n11246 = ( x697 & x698 ) | ( x697 & x699 ) | ( x698 & x699 ) ;
  assign n11247 = n11235 & n11241 ;
  assign n11248 = ( n11245 & n11246 ) | ( n11245 & n11247 ) | ( n11246 & n11247 ) ;
  assign n11249 = n11244 & n11248 ;
  assign n11250 = n11229 | n11249 ;
  assign n11251 = n11245 & ~n11246 ;
  assign n11252 = ~n11245 & n11246 ;
  assign n11253 = n11251 | n11252 ;
  assign n11254 = ~n11247 & n11253 ;
  assign n11255 = n11247 & ~n11253 ;
  assign n11256 = n11254 | n11255 ;
  assign n11257 = n11248 & n11256 ;
  assign n11258 = n11225 & n11244 ;
  assign n11259 = n11256 & n11258 ;
  assign n11260 = ~n11257 & n11259 ;
  assign n11261 = ~n11250 & n11260 ;
  assign n11262 = n11228 & n11261 ;
  assign n11263 = ~n11257 & n11258 ;
  assign n11264 = ~n11249 & n11256 ;
  assign n11265 = n11229 & ~n11264 ;
  assign n11266 = ( n11263 & n11264 ) | ( n11263 & ~n11265 ) | ( n11264 & ~n11265 ) ;
  assign n11267 = ( n11228 & n11262 ) | ( n11228 & ~n11266 ) | ( n11262 & ~n11266 ) ;
  assign n11268 = n11244 & ~n11248 ;
  assign n11269 = ( n11244 & ~n11256 ) | ( n11244 & n11268 ) | ( ~n11256 & n11268 ) ;
  assign n11270 = n11225 & ~n11226 ;
  assign n11271 = ( ~n11222 & n11225 ) | ( ~n11222 & n11270 ) | ( n11225 & n11270 ) ;
  assign n11272 = ~n11269 & n11271 ;
  assign n11273 = n11269 & ~n11271 ;
  assign n11274 = n11272 | n11273 ;
  assign n11275 = ( x688 & x689 ) | ( x688 & x690 ) | ( x689 & x690 ) ;
  assign n11276 = ( x685 & x686 ) | ( x685 & x687 ) | ( x686 & x687 ) ;
  assign n11277 = n11275 & ~n11276 ;
  assign n11278 = ~n11275 & n11276 ;
  assign n11279 = n11277 | n11278 ;
  assign n11280 = ~x685 & x686 ;
  assign n11281 = x685 & ~x686 ;
  assign n11282 = n11280 | n11281 ;
  assign n11283 = ~x687 & n11282 ;
  assign n11284 = x687 & ~n11282 ;
  assign n11285 = n11283 | n11284 ;
  assign n11286 = ~x688 & x689 ;
  assign n11287 = x688 & ~x689 ;
  assign n11288 = n11286 | n11287 ;
  assign n11289 = ~x690 & n11288 ;
  assign n11290 = x690 & ~n11288 ;
  assign n11291 = n11289 | n11290 ;
  assign n11292 = n11285 & n11291 ;
  assign n11293 = n11279 & ~n11292 ;
  assign n11294 = ~n11279 & n11292 ;
  assign n11295 = n11293 | n11294 ;
  assign n11296 = n11285 & ~n11291 ;
  assign n11297 = ~n11285 & n11291 ;
  assign n11298 = n11296 | n11297 ;
  assign n11299 = ( n11275 & n11276 ) | ( n11275 & n11292 ) | ( n11276 & n11292 ) ;
  assign n11300 = n11298 & ~n11299 ;
  assign n11301 = ( ~n11295 & n11298 ) | ( ~n11295 & n11300 ) | ( n11298 & n11300 ) ;
  assign n11302 = ~x679 & x680 ;
  assign n11303 = x679 & ~x680 ;
  assign n11304 = n11302 | n11303 ;
  assign n11305 = ~x681 & n11304 ;
  assign n11306 = x681 & ~n11304 ;
  assign n11307 = n11305 | n11306 ;
  assign n11308 = ~x682 & x683 ;
  assign n11309 = x682 & ~x683 ;
  assign n11310 = n11308 | n11309 ;
  assign n11311 = ~x684 & n11310 ;
  assign n11312 = x684 & ~n11310 ;
  assign n11313 = n11311 | n11312 ;
  assign n11314 = n11307 & ~n11313 ;
  assign n11315 = ~n11307 & n11313 ;
  assign n11316 = n11314 | n11315 ;
  assign n11317 = ( x682 & x683 ) | ( x682 & x684 ) | ( x683 & x684 ) ;
  assign n11318 = ( x679 & x680 ) | ( x679 & x681 ) | ( x680 & x681 ) ;
  assign n11319 = n11317 & ~n11318 ;
  assign n11320 = ~n11317 & n11318 ;
  assign n11321 = n11319 | n11320 ;
  assign n11322 = n11307 & n11313 ;
  assign n11323 = n11321 & ~n11322 ;
  assign n11324 = ~n11321 & n11322 ;
  assign n11325 = n11323 | n11324 ;
  assign n11326 = ( n11317 & n11318 ) | ( n11317 & n11322 ) | ( n11318 & n11322 ) ;
  assign n11327 = n11316 & ~n11326 ;
  assign n11328 = ( n11316 & ~n11325 ) | ( n11316 & n11327 ) | ( ~n11325 & n11327 ) ;
  assign n11329 = ~n11301 & n11328 ;
  assign n11330 = n11301 & ~n11328 ;
  assign n11331 = n11329 | n11330 ;
  assign n11332 = n11274 & n11331 ;
  assign n11333 = ( n11228 & ~n11229 ) | ( n11228 & n11264 ) | ( ~n11229 & n11264 ) ;
  assign n11334 = n11228 & n11264 ;
  assign n11335 = ( n11263 & n11333 ) | ( n11263 & n11334 ) | ( n11333 & n11334 ) ;
  assign n11336 = n11266 & ~n11335 ;
  assign n11337 = n11332 | n11336 ;
  assign n11338 = n11267 | n11337 ;
  assign n11339 = n11325 & n11326 ;
  assign n11340 = n11298 & n11299 ;
  assign n11341 = n11339 | n11340 ;
  assign n11342 = n11295 & n11299 ;
  assign n11343 = n11298 & n11316 ;
  assign n11344 = n11295 & n11343 ;
  assign n11345 = ~n11342 & n11344 ;
  assign n11346 = ~n11341 & n11345 ;
  assign n11347 = n11316 & n11326 ;
  assign n11348 = n11325 & ~n11347 ;
  assign n11349 = ~n11346 & n11348 ;
  assign n11350 = ~n11342 & n11343 ;
  assign n11351 = n11295 & ~n11340 ;
  assign n11352 = ( n11339 & n11348 ) | ( n11339 & n11351 ) | ( n11348 & n11351 ) ;
  assign n11353 = n11348 | n11351 ;
  assign n11354 = ( ~n11350 & n11352 ) | ( ~n11350 & n11353 ) | ( n11352 & n11353 ) ;
  assign n11355 = n11339 | n11351 ;
  assign n11356 = n11350 & ~n11355 ;
  assign n11357 = ( ~n11351 & n11354 ) | ( ~n11351 & n11356 ) | ( n11354 & n11356 ) ;
  assign n11358 = ( ~n11349 & n11354 ) | ( ~n11349 & n11357 ) | ( n11354 & n11357 ) ;
  assign n11359 = n11338 & n11358 ;
  assign n11360 = n11332 & n11336 ;
  assign n11361 = ( n11267 & n11332 ) | ( n11267 & n11360 ) | ( n11332 & n11360 ) ;
  assign n11362 = n11359 | n11361 ;
  assign n11363 = n11339 & ~n11351 ;
  assign n11364 = ( n11350 & n11351 ) | ( n11350 & ~n11363 ) | ( n11351 & ~n11363 ) ;
  assign n11365 = n11348 & n11364 ;
  assign n11366 = ~n11316 & n11326 ;
  assign n11367 = ( ~n11325 & n11326 ) | ( ~n11325 & n11366 ) | ( n11326 & n11366 ) ;
  assign n11368 = ~n11298 & n11299 ;
  assign n11369 = ( ~n11295 & n11299 ) | ( ~n11295 & n11368 ) | ( n11299 & n11368 ) ;
  assign n11370 = ~n11367 & n11369 ;
  assign n11371 = n11367 & ~n11369 ;
  assign n11372 = n11370 | n11371 ;
  assign n11373 = n11346 | n11372 ;
  assign n11374 = n11365 | n11373 ;
  assign n11375 = n11346 & n11372 ;
  assign n11376 = ( n11365 & n11372 ) | ( n11365 & n11375 ) | ( n11372 & n11375 ) ;
  assign n11377 = n11374 & ~n11376 ;
  assign n11378 = n11228 & n11266 ;
  assign n11379 = ~n11225 & n11226 ;
  assign n11380 = ( ~n11222 & n11226 ) | ( ~n11222 & n11379 ) | ( n11226 & n11379 ) ;
  assign n11381 = ~n11244 & n11248 ;
  assign n11382 = ( n11248 & ~n11256 ) | ( n11248 & n11381 ) | ( ~n11256 & n11381 ) ;
  assign n11383 = ~n11380 & n11382 ;
  assign n11384 = n11380 & ~n11382 ;
  assign n11385 = n11383 | n11384 ;
  assign n11386 = n11261 | n11385 ;
  assign n11387 = n11378 | n11386 ;
  assign n11388 = n11261 & n11385 ;
  assign n11389 = ( n11378 & n11385 ) | ( n11378 & n11388 ) | ( n11385 & n11388 ) ;
  assign n11390 = n11387 & ~n11389 ;
  assign n11391 = n11377 | n11390 ;
  assign n11392 = n11362 & n11391 ;
  assign n11393 = n11374 & n11387 ;
  assign n11394 = n11376 | n11389 ;
  assign n11395 = n11393 & ~n11394 ;
  assign n11396 = ( n11261 & n11380 ) | ( n11261 & n11382 ) | ( n11380 & n11382 ) ;
  assign n11397 = n11380 | n11382 ;
  assign n11398 = ( n11378 & n11396 ) | ( n11378 & n11397 ) | ( n11396 & n11397 ) ;
  assign n11399 = ( n11346 & n11367 ) | ( n11346 & n11369 ) | ( n11367 & n11369 ) ;
  assign n11400 = n11367 | n11369 ;
  assign n11401 = ( n11365 & n11399 ) | ( n11365 & n11400 ) | ( n11399 & n11400 ) ;
  assign n11402 = ~n11398 & n11401 ;
  assign n11403 = n11398 & ~n11401 ;
  assign n11404 = n11402 | n11403 ;
  assign n11405 = n11395 | n11404 ;
  assign n11406 = n11392 | n11405 ;
  assign n11407 = n11391 | n11395 ;
  assign n11408 = ( n11362 & n11395 ) | ( n11362 & n11407 ) | ( n11395 & n11407 ) ;
  assign n11409 = n11404 & n11408 ;
  assign n11410 = n11406 & ~n11409 ;
  assign n11411 = ( x670 & x671 ) | ( x670 & x672 ) | ( x671 & x672 ) ;
  assign n11412 = ( x667 & x668 ) | ( x667 & x669 ) | ( x668 & x669 ) ;
  assign n11413 = n11411 & ~n11412 ;
  assign n11414 = ~n11411 & n11412 ;
  assign n11415 = n11413 | n11414 ;
  assign n11416 = ~x667 & x668 ;
  assign n11417 = x667 & ~x668 ;
  assign n11418 = n11416 | n11417 ;
  assign n11419 = ~x669 & n11418 ;
  assign n11420 = x669 & ~n11418 ;
  assign n11421 = n11419 | n11420 ;
  assign n11422 = ~x670 & x671 ;
  assign n11423 = x670 & ~x671 ;
  assign n11424 = n11422 | n11423 ;
  assign n11425 = ~x672 & n11424 ;
  assign n11426 = x672 & ~n11424 ;
  assign n11427 = n11425 | n11426 ;
  assign n11428 = n11421 & n11427 ;
  assign n11429 = n11415 & ~n11428 ;
  assign n11430 = ~n11415 & n11428 ;
  assign n11431 = n11429 | n11430 ;
  assign n11432 = n11421 & ~n11427 ;
  assign n11433 = ~n11421 & n11427 ;
  assign n11434 = n11432 | n11433 ;
  assign n11435 = ( n11411 & n11412 ) | ( n11411 & n11428 ) | ( n11412 & n11428 ) ;
  assign n11436 = n11434 & n11435 ;
  assign n11437 = n11431 & ~n11436 ;
  assign n11438 = n11431 & n11435 ;
  assign n11439 = ~x673 & x674 ;
  assign n11440 = x673 & ~x674 ;
  assign n11441 = n11439 | n11440 ;
  assign n11442 = ~x675 & n11441 ;
  assign n11443 = x675 & ~n11441 ;
  assign n11444 = n11442 | n11443 ;
  assign n11445 = ~x676 & x677 ;
  assign n11446 = x676 & ~x677 ;
  assign n11447 = n11445 | n11446 ;
  assign n11448 = ~x678 & n11447 ;
  assign n11449 = x678 & ~n11447 ;
  assign n11450 = n11448 | n11449 ;
  assign n11451 = n11444 & ~n11450 ;
  assign n11452 = ~n11444 & n11450 ;
  assign n11453 = n11451 | n11452 ;
  assign n11454 = ( x676 & x677 ) | ( x676 & x678 ) | ( x677 & x678 ) ;
  assign n11455 = ( x673 & x674 ) | ( x673 & x675 ) | ( x674 & x675 ) ;
  assign n11456 = n11444 & n11450 ;
  assign n11457 = ( n11454 & n11455 ) | ( n11454 & n11456 ) | ( n11455 & n11456 ) ;
  assign n11458 = n11453 & n11457 ;
  assign n11459 = n11438 | n11458 ;
  assign n11460 = n11454 & ~n11455 ;
  assign n11461 = ~n11454 & n11455 ;
  assign n11462 = n11460 | n11461 ;
  assign n11463 = ~n11456 & n11462 ;
  assign n11464 = n11456 & ~n11462 ;
  assign n11465 = n11463 | n11464 ;
  assign n11466 = n11457 & n11465 ;
  assign n11467 = n11434 & n11453 ;
  assign n11468 = n11465 & n11467 ;
  assign n11469 = ~n11466 & n11468 ;
  assign n11470 = ~n11459 & n11469 ;
  assign n11471 = n11437 & n11470 ;
  assign n11472 = ~n11466 & n11467 ;
  assign n11473 = ~n11458 & n11465 ;
  assign n11474 = n11438 & ~n11473 ;
  assign n11475 = ( n11472 & n11473 ) | ( n11472 & ~n11474 ) | ( n11473 & ~n11474 ) ;
  assign n11476 = ( n11437 & n11471 ) | ( n11437 & ~n11475 ) | ( n11471 & ~n11475 ) ;
  assign n11477 = n11453 & ~n11457 ;
  assign n11478 = ( n11453 & ~n11465 ) | ( n11453 & n11477 ) | ( ~n11465 & n11477 ) ;
  assign n11479 = n11434 & ~n11435 ;
  assign n11480 = ( ~n11431 & n11434 ) | ( ~n11431 & n11479 ) | ( n11434 & n11479 ) ;
  assign n11481 = ~n11478 & n11480 ;
  assign n11482 = n11478 & ~n11480 ;
  assign n11483 = n11481 | n11482 ;
  assign n11484 = ( x664 & x665 ) | ( x664 & x666 ) | ( x665 & x666 ) ;
  assign n11485 = ( x661 & x662 ) | ( x661 & x663 ) | ( x662 & x663 ) ;
  assign n11486 = n11484 & ~n11485 ;
  assign n11487 = ~n11484 & n11485 ;
  assign n11488 = n11486 | n11487 ;
  assign n11489 = ~x661 & x662 ;
  assign n11490 = x661 & ~x662 ;
  assign n11491 = n11489 | n11490 ;
  assign n11492 = ~x663 & n11491 ;
  assign n11493 = x663 & ~n11491 ;
  assign n11494 = n11492 | n11493 ;
  assign n11495 = ~x664 & x665 ;
  assign n11496 = x664 & ~x665 ;
  assign n11497 = n11495 | n11496 ;
  assign n11498 = ~x666 & n11497 ;
  assign n11499 = x666 & ~n11497 ;
  assign n11500 = n11498 | n11499 ;
  assign n11501 = n11494 & n11500 ;
  assign n11502 = n11488 & ~n11501 ;
  assign n11503 = ~n11488 & n11501 ;
  assign n11504 = n11502 | n11503 ;
  assign n11505 = n11494 & ~n11500 ;
  assign n11506 = ~n11494 & n11500 ;
  assign n11507 = n11505 | n11506 ;
  assign n11508 = ( n11484 & n11485 ) | ( n11484 & n11501 ) | ( n11485 & n11501 ) ;
  assign n11509 = n11507 & ~n11508 ;
  assign n11510 = ( ~n11504 & n11507 ) | ( ~n11504 & n11509 ) | ( n11507 & n11509 ) ;
  assign n11511 = ~x655 & x656 ;
  assign n11512 = x655 & ~x656 ;
  assign n11513 = n11511 | n11512 ;
  assign n11514 = ~x657 & n11513 ;
  assign n11515 = x657 & ~n11513 ;
  assign n11516 = n11514 | n11515 ;
  assign n11517 = ~x658 & x659 ;
  assign n11518 = x658 & ~x659 ;
  assign n11519 = n11517 | n11518 ;
  assign n11520 = ~x660 & n11519 ;
  assign n11521 = x660 & ~n11519 ;
  assign n11522 = n11520 | n11521 ;
  assign n11523 = n11516 & ~n11522 ;
  assign n11524 = ~n11516 & n11522 ;
  assign n11525 = n11523 | n11524 ;
  assign n11526 = ( x658 & x659 ) | ( x658 & x660 ) | ( x659 & x660 ) ;
  assign n11527 = ( x655 & x656 ) | ( x655 & x657 ) | ( x656 & x657 ) ;
  assign n11528 = n11526 & ~n11527 ;
  assign n11529 = ~n11526 & n11527 ;
  assign n11530 = n11528 | n11529 ;
  assign n11531 = n11516 & n11522 ;
  assign n11532 = n11530 & ~n11531 ;
  assign n11533 = ~n11530 & n11531 ;
  assign n11534 = n11532 | n11533 ;
  assign n11535 = ( n11526 & n11527 ) | ( n11526 & n11531 ) | ( n11527 & n11531 ) ;
  assign n11536 = n11525 & ~n11535 ;
  assign n11537 = ( n11525 & ~n11534 ) | ( n11525 & n11536 ) | ( ~n11534 & n11536 ) ;
  assign n11538 = ~n11510 & n11537 ;
  assign n11539 = n11510 & ~n11537 ;
  assign n11540 = n11538 | n11539 ;
  assign n11541 = n11483 & n11540 ;
  assign n11542 = ( n11437 & ~n11438 ) | ( n11437 & n11473 ) | ( ~n11438 & n11473 ) ;
  assign n11543 = n11437 & n11473 ;
  assign n11544 = ( n11472 & n11542 ) | ( n11472 & n11543 ) | ( n11542 & n11543 ) ;
  assign n11545 = n11475 & ~n11544 ;
  assign n11546 = n11541 | n11545 ;
  assign n11547 = n11476 | n11546 ;
  assign n11548 = n11534 & n11535 ;
  assign n11549 = n11507 & n11508 ;
  assign n11550 = n11548 | n11549 ;
  assign n11551 = n11504 & n11508 ;
  assign n11552 = n11507 & n11525 ;
  assign n11553 = n11504 & n11552 ;
  assign n11554 = ~n11551 & n11553 ;
  assign n11555 = ~n11550 & n11554 ;
  assign n11556 = n11525 & n11535 ;
  assign n11557 = n11534 & ~n11556 ;
  assign n11558 = ~n11555 & n11557 ;
  assign n11559 = ~n11551 & n11552 ;
  assign n11560 = n11504 & ~n11549 ;
  assign n11561 = ( n11548 & n11557 ) | ( n11548 & n11560 ) | ( n11557 & n11560 ) ;
  assign n11562 = n11557 | n11560 ;
  assign n11563 = ( ~n11559 & n11561 ) | ( ~n11559 & n11562 ) | ( n11561 & n11562 ) ;
  assign n11564 = n11548 | n11560 ;
  assign n11565 = n11559 & ~n11564 ;
  assign n11566 = ( ~n11560 & n11563 ) | ( ~n11560 & n11565 ) | ( n11563 & n11565 ) ;
  assign n11567 = ( ~n11558 & n11563 ) | ( ~n11558 & n11566 ) | ( n11563 & n11566 ) ;
  assign n11568 = n11547 & n11567 ;
  assign n11569 = n11541 & n11545 ;
  assign n11570 = ( n11476 & n11541 ) | ( n11476 & n11569 ) | ( n11541 & n11569 ) ;
  assign n11571 = n11568 | n11570 ;
  assign n11572 = n11548 & ~n11560 ;
  assign n11573 = ( n11559 & n11560 ) | ( n11559 & ~n11572 ) | ( n11560 & ~n11572 ) ;
  assign n11574 = n11557 & n11573 ;
  assign n11575 = ~n11525 & n11535 ;
  assign n11576 = ( ~n11534 & n11535 ) | ( ~n11534 & n11575 ) | ( n11535 & n11575 ) ;
  assign n11577 = ~n11507 & n11508 ;
  assign n11578 = ( ~n11504 & n11508 ) | ( ~n11504 & n11577 ) | ( n11508 & n11577 ) ;
  assign n11579 = ~n11576 & n11578 ;
  assign n11580 = n11576 & ~n11578 ;
  assign n11581 = n11579 | n11580 ;
  assign n11582 = n11555 | n11581 ;
  assign n11583 = n11574 | n11582 ;
  assign n11584 = n11555 & n11581 ;
  assign n11585 = ( n11574 & n11581 ) | ( n11574 & n11584 ) | ( n11581 & n11584 ) ;
  assign n11586 = n11583 & ~n11585 ;
  assign n11587 = n11437 & n11475 ;
  assign n11588 = ~n11434 & n11435 ;
  assign n11589 = ( ~n11431 & n11435 ) | ( ~n11431 & n11588 ) | ( n11435 & n11588 ) ;
  assign n11590 = ~n11453 & n11457 ;
  assign n11591 = ( n11457 & ~n11465 ) | ( n11457 & n11590 ) | ( ~n11465 & n11590 ) ;
  assign n11592 = ~n11589 & n11591 ;
  assign n11593 = n11589 & ~n11591 ;
  assign n11594 = n11592 | n11593 ;
  assign n11595 = n11470 | n11594 ;
  assign n11596 = n11587 | n11595 ;
  assign n11597 = n11470 & n11594 ;
  assign n11598 = ( n11587 & n11594 ) | ( n11587 & n11597 ) | ( n11594 & n11597 ) ;
  assign n11599 = n11596 & ~n11598 ;
  assign n11600 = n11586 | n11599 ;
  assign n11601 = n11571 & n11600 ;
  assign n11602 = n11583 & n11596 ;
  assign n11603 = n11585 | n11598 ;
  assign n11604 = n11602 & ~n11603 ;
  assign n11605 = ( n11470 & n11589 ) | ( n11470 & n11591 ) | ( n11589 & n11591 ) ;
  assign n11606 = n11589 | n11591 ;
  assign n11607 = ( n11587 & n11605 ) | ( n11587 & n11606 ) | ( n11605 & n11606 ) ;
  assign n11608 = ( n11555 & n11576 ) | ( n11555 & n11578 ) | ( n11576 & n11578 ) ;
  assign n11609 = n11576 | n11578 ;
  assign n11610 = ( n11574 & n11608 ) | ( n11574 & n11609 ) | ( n11608 & n11609 ) ;
  assign n11611 = ~n11607 & n11610 ;
  assign n11612 = n11607 & ~n11610 ;
  assign n11613 = n11611 | n11612 ;
  assign n11614 = n11604 | n11613 ;
  assign n11615 = n11601 | n11614 ;
  assign n11616 = n11600 | n11604 ;
  assign n11617 = ( n11571 & n11604 ) | ( n11571 & n11616 ) | ( n11604 & n11616 ) ;
  assign n11618 = n11613 & n11617 ;
  assign n11619 = n11615 & ~n11618 ;
  assign n11620 = n11410 | n11619 ;
  assign n11621 = n11338 & ~n11361 ;
  assign n11622 = n11358 & ~n11621 ;
  assign n11623 = n11274 & ~n11331 ;
  assign n11624 = ~n11274 & n11331 ;
  assign n11625 = n11623 | n11624 ;
  assign n11626 = n11483 & ~n11540 ;
  assign n11627 = ~n11483 & n11540 ;
  assign n11628 = n11626 | n11627 ;
  assign n11629 = n11625 & n11628 ;
  assign n11630 = ~n11332 & n11338 ;
  assign n11631 = n11338 & ~n11358 ;
  assign n11632 = n11267 | n11336 ;
  assign n11633 = n11358 | n11632 ;
  assign n11634 = ( n11630 & n11631 ) | ( n11630 & ~n11633 ) | ( n11631 & ~n11633 ) ;
  assign n11635 = n11629 | n11634 ;
  assign n11636 = n11622 | n11635 ;
  assign n11637 = n11476 | n11545 ;
  assign n11638 = ( n11541 & n11567 ) | ( n11541 & ~n11637 ) | ( n11567 & ~n11637 ) ;
  assign n11639 = ( ~n11567 & n11637 ) | ( ~n11567 & n11638 ) | ( n11637 & n11638 ) ;
  assign n11640 = ( ~n11541 & n11638 ) | ( ~n11541 & n11639 ) | ( n11638 & n11639 ) ;
  assign n11641 = n11636 & n11640 ;
  assign n11642 = n11622 | n11634 ;
  assign n11643 = n11629 & n11642 ;
  assign n11644 = ( n11570 & ~n11586 ) | ( n11570 & n11599 ) | ( ~n11586 & n11599 ) ;
  assign n11645 = n11586 & ~n11599 ;
  assign n11646 = ( n11568 & n11644 ) | ( n11568 & ~n11645 ) | ( n11644 & ~n11645 ) ;
  assign n11647 = ( ~n11571 & n11586 ) | ( ~n11571 & n11646 ) | ( n11586 & n11646 ) ;
  assign n11648 = ( ~n11599 & n11646 ) | ( ~n11599 & n11647 ) | ( n11646 & n11647 ) ;
  assign n11649 = ( n11361 & ~n11377 ) | ( n11361 & n11390 ) | ( ~n11377 & n11390 ) ;
  assign n11650 = n11377 & ~n11390 ;
  assign n11651 = ( n11359 & n11649 ) | ( n11359 & ~n11650 ) | ( n11649 & ~n11650 ) ;
  assign n11652 = ( ~n11362 & n11377 ) | ( ~n11362 & n11651 ) | ( n11377 & n11651 ) ;
  assign n11653 = ( ~n11390 & n11651 ) | ( ~n11390 & n11652 ) | ( n11651 & n11652 ) ;
  assign n11654 = ( n11643 & n11648 ) | ( n11643 & n11653 ) | ( n11648 & n11653 ) ;
  assign n11655 = n11648 | n11653 ;
  assign n11656 = ( n11641 & n11654 ) | ( n11641 & n11655 ) | ( n11654 & n11655 ) ;
  assign n11657 = n11620 & n11656 ;
  assign n11658 = n11406 & n11615 ;
  assign n11659 = n11409 | n11618 ;
  assign n11660 = n11658 & ~n11659 ;
  assign n11661 = n11607 & n11610 ;
  assign n11662 = n11607 | n11610 ;
  assign n11663 = n11661 | n11662 ;
  assign n11664 = ( n11617 & n11661 ) | ( n11617 & n11663 ) | ( n11661 & n11663 ) ;
  assign n11665 = n11398 & n11401 ;
  assign n11666 = n11398 | n11401 ;
  assign n11667 = n11665 | n11666 ;
  assign n11668 = ( n11408 & n11665 ) | ( n11408 & n11667 ) | ( n11665 & n11667 ) ;
  assign n11669 = n11664 & n11668 ;
  assign n11670 = n11668 & ~n11669 ;
  assign n11671 = ( n11664 & ~n11669 ) | ( n11664 & n11670 ) | ( ~n11669 & n11670 ) ;
  assign n11672 = n11660 | n11671 ;
  assign n11673 = n11657 | n11672 ;
  assign n11674 = n11657 | n11660 ;
  assign n11675 = n11671 & n11674 ;
  assign n11676 = n11673 & ~n11675 ;
  assign n11677 = ~x739 & x740 ;
  assign n11678 = x739 & ~x740 ;
  assign n11679 = n11677 | n11678 ;
  assign n11680 = ~x741 & n11679 ;
  assign n11681 = x741 & ~n11679 ;
  assign n11682 = n11680 | n11681 ;
  assign n11683 = ~x742 & x743 ;
  assign n11684 = x742 & ~x743 ;
  assign n11685 = n11683 | n11684 ;
  assign n11686 = ~x744 & n11685 ;
  assign n11687 = x744 & ~n11685 ;
  assign n11688 = n11686 | n11687 ;
  assign n11689 = n11682 & n11688 ;
  assign n11690 = ( x742 & x743 ) | ( x742 & x744 ) | ( x743 & x744 ) ;
  assign n11691 = ( x739 & x740 ) | ( x739 & x741 ) | ( x740 & x741 ) ;
  assign n11692 = ~n11690 & n11691 ;
  assign n11693 = n11690 & ~n11691 ;
  assign n11694 = n11692 | n11693 ;
  assign n11695 = ~n11689 & n11694 ;
  assign n11696 = n11689 & ~n11694 ;
  assign n11697 = n11695 | n11696 ;
  assign n11698 = n11682 & ~n11688 ;
  assign n11699 = ~n11682 & n11688 ;
  assign n11700 = n11698 | n11699 ;
  assign n11701 = ( n11689 & n11690 ) | ( n11689 & n11691 ) | ( n11690 & n11691 ) ;
  assign n11702 = n11700 & n11701 ;
  assign n11703 = n11697 & ~n11702 ;
  assign n11704 = n11697 & n11701 ;
  assign n11705 = x745 & ~x746 ;
  assign n11706 = ~x745 & x746 ;
  assign n11707 = n11705 | n11706 ;
  assign n11708 = ~x747 & n11707 ;
  assign n11709 = x747 & ~n11707 ;
  assign n11710 = n11708 | n11709 ;
  assign n11711 = x748 & ~x749 ;
  assign n11712 = ~x748 & x749 ;
  assign n11713 = n11711 | n11712 ;
  assign n11714 = ~x750 & n11713 ;
  assign n11715 = x750 & ~n11713 ;
  assign n11716 = n11714 | n11715 ;
  assign n11717 = n11710 & ~n11716 ;
  assign n11718 = ~n11710 & n11716 ;
  assign n11719 = n11717 | n11718 ;
  assign n11720 = ( x748 & x749 ) | ( x748 & x750 ) | ( x749 & x750 ) ;
  assign n11721 = ( x745 & x746 ) | ( x745 & x747 ) | ( x746 & x747 ) ;
  assign n11722 = n11710 & n11716 ;
  assign n11723 = ( n11720 & n11721 ) | ( n11720 & n11722 ) | ( n11721 & n11722 ) ;
  assign n11724 = n11719 & n11723 ;
  assign n11725 = n11704 | n11724 ;
  assign n11726 = n11720 & ~n11721 ;
  assign n11727 = ~n11720 & n11721 ;
  assign n11728 = n11726 | n11727 ;
  assign n11729 = ~n11722 & n11728 ;
  assign n11730 = n11722 & ~n11728 ;
  assign n11731 = n11729 | n11730 ;
  assign n11732 = n11723 & n11731 ;
  assign n11733 = n11700 & n11719 ;
  assign n11734 = n11731 & n11733 ;
  assign n11735 = ~n11732 & n11734 ;
  assign n11736 = ~n11725 & n11735 ;
  assign n11737 = n11703 & n11736 ;
  assign n11738 = ~n11732 & n11733 ;
  assign n11739 = ~n11724 & n11731 ;
  assign n11740 = n11704 & ~n11739 ;
  assign n11741 = ( n11738 & n11739 ) | ( n11738 & ~n11740 ) | ( n11739 & ~n11740 ) ;
  assign n11742 = ( n11703 & n11737 ) | ( n11703 & ~n11741 ) | ( n11737 & ~n11741 ) ;
  assign n11743 = n11719 & ~n11723 ;
  assign n11744 = ( n11719 & ~n11731 ) | ( n11719 & n11743 ) | ( ~n11731 & n11743 ) ;
  assign n11745 = n11700 & ~n11701 ;
  assign n11746 = ( ~n11697 & n11700 ) | ( ~n11697 & n11745 ) | ( n11700 & n11745 ) ;
  assign n11747 = ~n11744 & n11746 ;
  assign n11748 = n11744 & ~n11746 ;
  assign n11749 = n11747 | n11748 ;
  assign n11750 = ( x736 & x737 ) | ( x736 & x738 ) | ( x737 & x738 ) ;
  assign n11751 = ( x733 & x734 ) | ( x733 & x735 ) | ( x734 & x735 ) ;
  assign n11752 = n11750 & ~n11751 ;
  assign n11753 = ~n11750 & n11751 ;
  assign n11754 = n11752 | n11753 ;
  assign n11755 = x733 & ~x734 ;
  assign n11756 = ~x733 & x734 ;
  assign n11757 = n11755 | n11756 ;
  assign n11758 = ~x735 & n11757 ;
  assign n11759 = x735 & ~n11757 ;
  assign n11760 = n11758 | n11759 ;
  assign n11761 = x736 & ~x737 ;
  assign n11762 = ~x736 & x737 ;
  assign n11763 = n11761 | n11762 ;
  assign n11764 = ~x738 & n11763 ;
  assign n11765 = x738 & ~n11763 ;
  assign n11766 = n11764 | n11765 ;
  assign n11767 = n11760 & n11766 ;
  assign n11768 = n11754 & ~n11767 ;
  assign n11769 = ~n11754 & n11767 ;
  assign n11770 = n11768 | n11769 ;
  assign n11771 = n11760 & ~n11766 ;
  assign n11772 = ~n11760 & n11766 ;
  assign n11773 = n11771 | n11772 ;
  assign n11774 = ( n11750 & n11751 ) | ( n11750 & n11767 ) | ( n11751 & n11767 ) ;
  assign n11775 = n11773 & ~n11774 ;
  assign n11776 = ( ~n11770 & n11773 ) | ( ~n11770 & n11775 ) | ( n11773 & n11775 ) ;
  assign n11777 = ~x727 & x728 ;
  assign n11778 = x727 & ~x728 ;
  assign n11779 = n11777 | n11778 ;
  assign n11780 = ~x729 & n11779 ;
  assign n11781 = x729 & ~n11779 ;
  assign n11782 = n11780 | n11781 ;
  assign n11783 = ~x730 & x731 ;
  assign n11784 = x730 & ~x731 ;
  assign n11785 = n11783 | n11784 ;
  assign n11786 = ~x732 & n11785 ;
  assign n11787 = x732 & ~n11785 ;
  assign n11788 = n11786 | n11787 ;
  assign n11789 = n11782 & n11788 ;
  assign n11790 = ( x730 & x731 ) | ( x730 & x732 ) | ( x731 & x732 ) ;
  assign n11791 = ( x727 & x728 ) | ( x727 & x729 ) | ( x728 & x729 ) ;
  assign n11792 = ~n11790 & n11791 ;
  assign n11793 = n11790 & ~n11791 ;
  assign n11794 = n11792 | n11793 ;
  assign n11795 = ~n11789 & n11794 ;
  assign n11796 = n11789 & ~n11794 ;
  assign n11797 = n11795 | n11796 ;
  assign n11798 = n11782 & ~n11788 ;
  assign n11799 = ~n11782 & n11788 ;
  assign n11800 = n11798 | n11799 ;
  assign n11801 = ( n11789 & n11790 ) | ( n11789 & n11791 ) | ( n11790 & n11791 ) ;
  assign n11802 = n11800 & ~n11801 ;
  assign n11803 = ( ~n11797 & n11800 ) | ( ~n11797 & n11802 ) | ( n11800 & n11802 ) ;
  assign n11804 = ~n11776 & n11803 ;
  assign n11805 = n11776 & ~n11803 ;
  assign n11806 = n11804 | n11805 ;
  assign n11807 = n11749 & n11806 ;
  assign n11808 = ( n11703 & ~n11704 ) | ( n11703 & n11739 ) | ( ~n11704 & n11739 ) ;
  assign n11809 = n11703 & n11739 ;
  assign n11810 = ( n11738 & n11808 ) | ( n11738 & n11809 ) | ( n11808 & n11809 ) ;
  assign n11811 = n11741 & ~n11810 ;
  assign n11812 = n11807 | n11811 ;
  assign n11813 = n11742 | n11812 ;
  assign n11814 = n11797 & n11801 ;
  assign n11815 = n11773 & n11774 ;
  assign n11816 = n11814 | n11815 ;
  assign n11817 = n11770 & n11774 ;
  assign n11818 = n11773 & n11800 ;
  assign n11819 = n11770 & n11818 ;
  assign n11820 = ~n11817 & n11819 ;
  assign n11821 = ~n11816 & n11820 ;
  assign n11822 = n11800 & n11801 ;
  assign n11823 = n11797 & ~n11822 ;
  assign n11824 = ~n11821 & n11823 ;
  assign n11825 = ~n11817 & n11818 ;
  assign n11826 = n11770 & ~n11815 ;
  assign n11827 = ( n11814 & n11823 ) | ( n11814 & n11826 ) | ( n11823 & n11826 ) ;
  assign n11828 = n11823 | n11826 ;
  assign n11829 = ( ~n11825 & n11827 ) | ( ~n11825 & n11828 ) | ( n11827 & n11828 ) ;
  assign n11830 = n11814 | n11826 ;
  assign n11831 = n11825 & ~n11830 ;
  assign n11832 = ( ~n11826 & n11829 ) | ( ~n11826 & n11831 ) | ( n11829 & n11831 ) ;
  assign n11833 = ( ~n11824 & n11829 ) | ( ~n11824 & n11832 ) | ( n11829 & n11832 ) ;
  assign n11834 = n11813 & n11833 ;
  assign n11835 = n11807 & n11811 ;
  assign n11836 = ( n11742 & n11807 ) | ( n11742 & n11835 ) | ( n11807 & n11835 ) ;
  assign n11837 = n11834 | n11836 ;
  assign n11838 = n11814 & ~n11826 ;
  assign n11839 = ( n11825 & n11826 ) | ( n11825 & ~n11838 ) | ( n11826 & ~n11838 ) ;
  assign n11840 = n11823 & n11839 ;
  assign n11841 = ~n11800 & n11801 ;
  assign n11842 = ( ~n11797 & n11801 ) | ( ~n11797 & n11841 ) | ( n11801 & n11841 ) ;
  assign n11843 = ~n11773 & n11774 ;
  assign n11844 = ( ~n11770 & n11774 ) | ( ~n11770 & n11843 ) | ( n11774 & n11843 ) ;
  assign n11845 = ~n11842 & n11844 ;
  assign n11846 = n11842 & ~n11844 ;
  assign n11847 = n11845 | n11846 ;
  assign n11848 = n11821 | n11847 ;
  assign n11849 = n11840 | n11848 ;
  assign n11850 = n11821 & n11847 ;
  assign n11851 = ( n11840 & n11847 ) | ( n11840 & n11850 ) | ( n11847 & n11850 ) ;
  assign n11852 = n11849 & ~n11851 ;
  assign n11853 = n11703 & n11741 ;
  assign n11854 = ~n11700 & n11701 ;
  assign n11855 = ( ~n11697 & n11701 ) | ( ~n11697 & n11854 ) | ( n11701 & n11854 ) ;
  assign n11856 = ~n11719 & n11723 ;
  assign n11857 = ( n11723 & ~n11731 ) | ( n11723 & n11856 ) | ( ~n11731 & n11856 ) ;
  assign n11858 = ~n11855 & n11857 ;
  assign n11859 = n11855 & ~n11857 ;
  assign n11860 = n11858 | n11859 ;
  assign n11861 = n11736 | n11860 ;
  assign n11862 = n11853 | n11861 ;
  assign n11863 = n11736 & n11860 ;
  assign n11864 = ( n11853 & n11860 ) | ( n11853 & n11863 ) | ( n11860 & n11863 ) ;
  assign n11865 = n11862 & ~n11864 ;
  assign n11866 = n11852 | n11865 ;
  assign n11867 = n11837 & n11866 ;
  assign n11868 = n11849 & n11862 ;
  assign n11869 = n11851 | n11864 ;
  assign n11870 = n11868 & ~n11869 ;
  assign n11871 = ( n11736 & n11855 ) | ( n11736 & n11857 ) | ( n11855 & n11857 ) ;
  assign n11872 = n11855 | n11857 ;
  assign n11873 = ( n11853 & n11871 ) | ( n11853 & n11872 ) | ( n11871 & n11872 ) ;
  assign n11874 = ( n11821 & n11842 ) | ( n11821 & n11844 ) | ( n11842 & n11844 ) ;
  assign n11875 = n11842 | n11844 ;
  assign n11876 = ( n11840 & n11874 ) | ( n11840 & n11875 ) | ( n11874 & n11875 ) ;
  assign n11877 = ~n11873 & n11876 ;
  assign n11878 = n11873 & ~n11876 ;
  assign n11879 = n11877 | n11878 ;
  assign n11880 = n11870 | n11879 ;
  assign n11881 = n11867 | n11880 ;
  assign n11882 = n11866 | n11870 ;
  assign n11883 = ( n11837 & n11870 ) | ( n11837 & n11882 ) | ( n11870 & n11882 ) ;
  assign n11884 = n11879 & n11883 ;
  assign n11885 = n11881 & ~n11884 ;
  assign n11886 = ~x715 & x716 ;
  assign n11887 = x715 & ~x716 ;
  assign n11888 = n11886 | n11887 ;
  assign n11889 = ~x717 & n11888 ;
  assign n11890 = x717 & ~n11888 ;
  assign n11891 = n11889 | n11890 ;
  assign n11892 = ~x718 & x719 ;
  assign n11893 = x718 & ~x719 ;
  assign n11894 = n11892 | n11893 ;
  assign n11895 = ~x720 & n11894 ;
  assign n11896 = x720 & ~n11894 ;
  assign n11897 = n11895 | n11896 ;
  assign n11898 = n11891 & n11897 ;
  assign n11899 = ( x718 & x719 ) | ( x718 & x720 ) | ( x719 & x720 ) ;
  assign n11900 = ( x715 & x716 ) | ( x715 & x717 ) | ( x716 & x717 ) ;
  assign n11901 = ~n11899 & n11900 ;
  assign n11902 = n11899 & ~n11900 ;
  assign n11903 = n11901 | n11902 ;
  assign n11904 = ~n11898 & n11903 ;
  assign n11905 = n11898 & ~n11903 ;
  assign n11906 = n11904 | n11905 ;
  assign n11907 = n11891 & ~n11897 ;
  assign n11908 = ~n11891 & n11897 ;
  assign n11909 = n11907 | n11908 ;
  assign n11910 = ( n11898 & n11899 ) | ( n11898 & n11900 ) | ( n11899 & n11900 ) ;
  assign n11911 = n11909 & n11910 ;
  assign n11912 = n11906 & ~n11911 ;
  assign n11913 = n11906 & n11910 ;
  assign n11914 = x721 & ~x722 ;
  assign n11915 = ~x721 & x722 ;
  assign n11916 = n11914 | n11915 ;
  assign n11917 = ~x723 & n11916 ;
  assign n11918 = x723 & ~n11916 ;
  assign n11919 = n11917 | n11918 ;
  assign n11920 = x724 & ~x725 ;
  assign n11921 = ~x724 & x725 ;
  assign n11922 = n11920 | n11921 ;
  assign n11923 = ~x726 & n11922 ;
  assign n11924 = x726 & ~n11922 ;
  assign n11925 = n11923 | n11924 ;
  assign n11926 = n11919 & ~n11925 ;
  assign n11927 = ~n11919 & n11925 ;
  assign n11928 = n11926 | n11927 ;
  assign n11929 = ( x724 & x725 ) | ( x724 & x726 ) | ( x725 & x726 ) ;
  assign n11930 = ( x721 & x722 ) | ( x721 & x723 ) | ( x722 & x723 ) ;
  assign n11931 = n11919 & n11925 ;
  assign n11932 = ( n11929 & n11930 ) | ( n11929 & n11931 ) | ( n11930 & n11931 ) ;
  assign n11933 = n11928 & n11932 ;
  assign n11934 = n11913 | n11933 ;
  assign n11935 = n11929 & ~n11930 ;
  assign n11936 = ~n11929 & n11930 ;
  assign n11937 = n11935 | n11936 ;
  assign n11938 = ~n11931 & n11937 ;
  assign n11939 = n11931 & ~n11937 ;
  assign n11940 = n11938 | n11939 ;
  assign n11941 = n11932 & n11940 ;
  assign n11942 = n11909 & n11928 ;
  assign n11943 = n11940 & n11942 ;
  assign n11944 = ~n11941 & n11943 ;
  assign n11945 = ~n11934 & n11944 ;
  assign n11946 = n11912 & n11945 ;
  assign n11947 = ~n11941 & n11942 ;
  assign n11948 = ~n11933 & n11940 ;
  assign n11949 = n11913 & ~n11948 ;
  assign n11950 = ( n11947 & n11948 ) | ( n11947 & ~n11949 ) | ( n11948 & ~n11949 ) ;
  assign n11951 = ( n11912 & n11946 ) | ( n11912 & ~n11950 ) | ( n11946 & ~n11950 ) ;
  assign n11952 = n11928 & ~n11932 ;
  assign n11953 = ( n11928 & ~n11940 ) | ( n11928 & n11952 ) | ( ~n11940 & n11952 ) ;
  assign n11954 = n11909 & ~n11910 ;
  assign n11955 = ( ~n11906 & n11909 ) | ( ~n11906 & n11954 ) | ( n11909 & n11954 ) ;
  assign n11956 = ~n11953 & n11955 ;
  assign n11957 = n11953 & ~n11955 ;
  assign n11958 = n11956 | n11957 ;
  assign n11959 = ( x712 & x713 ) | ( x712 & x714 ) | ( x713 & x714 ) ;
  assign n11960 = ( x709 & x710 ) | ( x709 & x711 ) | ( x710 & x711 ) ;
  assign n11961 = n11959 & ~n11960 ;
  assign n11962 = ~n11959 & n11960 ;
  assign n11963 = n11961 | n11962 ;
  assign n11964 = ~x709 & x710 ;
  assign n11965 = x709 & ~x710 ;
  assign n11966 = n11964 | n11965 ;
  assign n11967 = ~x711 & n11966 ;
  assign n11968 = x711 & ~n11966 ;
  assign n11969 = n11967 | n11968 ;
  assign n11970 = ~x712 & x713 ;
  assign n11971 = x712 & ~x713 ;
  assign n11972 = n11970 | n11971 ;
  assign n11973 = ~x714 & n11972 ;
  assign n11974 = x714 & ~n11972 ;
  assign n11975 = n11973 | n11974 ;
  assign n11976 = n11969 & n11975 ;
  assign n11977 = n11963 & ~n11976 ;
  assign n11978 = ~n11963 & n11976 ;
  assign n11979 = n11977 | n11978 ;
  assign n11980 = n11969 & ~n11975 ;
  assign n11981 = ~n11969 & n11975 ;
  assign n11982 = n11980 | n11981 ;
  assign n11983 = ( n11959 & n11960 ) | ( n11959 & n11976 ) | ( n11960 & n11976 ) ;
  assign n11984 = n11982 & ~n11983 ;
  assign n11985 = ( ~n11979 & n11982 ) | ( ~n11979 & n11984 ) | ( n11982 & n11984 ) ;
  assign n11986 = ~x703 & x704 ;
  assign n11987 = x703 & ~x704 ;
  assign n11988 = n11986 | n11987 ;
  assign n11989 = ~x705 & n11988 ;
  assign n11990 = x705 & ~n11988 ;
  assign n11991 = n11989 | n11990 ;
  assign n11992 = ~x706 & x707 ;
  assign n11993 = x706 & ~x707 ;
  assign n11994 = n11992 | n11993 ;
  assign n11995 = ~x708 & n11994 ;
  assign n11996 = x708 & ~n11994 ;
  assign n11997 = n11995 | n11996 ;
  assign n11998 = n11991 & ~n11997 ;
  assign n11999 = ~n11991 & n11997 ;
  assign n12000 = n11998 | n11999 ;
  assign n12001 = ( x706 & x707 ) | ( x706 & x708 ) | ( x707 & x708 ) ;
  assign n12002 = ( x703 & x704 ) | ( x703 & x705 ) | ( x704 & x705 ) ;
  assign n12003 = n12001 & ~n12002 ;
  assign n12004 = ~n12001 & n12002 ;
  assign n12005 = n12003 | n12004 ;
  assign n12006 = n11991 & n11997 ;
  assign n12007 = n12005 & ~n12006 ;
  assign n12008 = ~n12005 & n12006 ;
  assign n12009 = n12007 | n12008 ;
  assign n12010 = ( n12001 & n12002 ) | ( n12001 & n12006 ) | ( n12002 & n12006 ) ;
  assign n12011 = n12000 & ~n12010 ;
  assign n12012 = ( n12000 & ~n12009 ) | ( n12000 & n12011 ) | ( ~n12009 & n12011 ) ;
  assign n12013 = ~n11985 & n12012 ;
  assign n12014 = n11985 & ~n12012 ;
  assign n12015 = n12013 | n12014 ;
  assign n12016 = n11958 & n12015 ;
  assign n12017 = ( n11912 & ~n11913 ) | ( n11912 & n11948 ) | ( ~n11913 & n11948 ) ;
  assign n12018 = n11912 & n11948 ;
  assign n12019 = ( n11947 & n12017 ) | ( n11947 & n12018 ) | ( n12017 & n12018 ) ;
  assign n12020 = n11950 & ~n12019 ;
  assign n12021 = n12016 | n12020 ;
  assign n12022 = n11951 | n12021 ;
  assign n12023 = n12009 & n12010 ;
  assign n12024 = n11982 & n11983 ;
  assign n12025 = n12023 | n12024 ;
  assign n12026 = n11979 & n11983 ;
  assign n12027 = n11982 & n12000 ;
  assign n12028 = n11979 & n12027 ;
  assign n12029 = ~n12026 & n12028 ;
  assign n12030 = ~n12025 & n12029 ;
  assign n12031 = n12000 & n12010 ;
  assign n12032 = n12009 & ~n12031 ;
  assign n12033 = ~n12030 & n12032 ;
  assign n12034 = ~n12026 & n12027 ;
  assign n12035 = n11979 & ~n12024 ;
  assign n12036 = ( n12023 & n12032 ) | ( n12023 & n12035 ) | ( n12032 & n12035 ) ;
  assign n12037 = n12032 | n12035 ;
  assign n12038 = ( ~n12034 & n12036 ) | ( ~n12034 & n12037 ) | ( n12036 & n12037 ) ;
  assign n12039 = n12023 | n12035 ;
  assign n12040 = n12034 & ~n12039 ;
  assign n12041 = ( ~n12035 & n12038 ) | ( ~n12035 & n12040 ) | ( n12038 & n12040 ) ;
  assign n12042 = ( ~n12033 & n12038 ) | ( ~n12033 & n12041 ) | ( n12038 & n12041 ) ;
  assign n12043 = n12022 & n12042 ;
  assign n12044 = n12016 & n12020 ;
  assign n12045 = ( n11951 & n12016 ) | ( n11951 & n12044 ) | ( n12016 & n12044 ) ;
  assign n12046 = n12043 | n12045 ;
  assign n12047 = n12023 & ~n12035 ;
  assign n12048 = ( n12034 & n12035 ) | ( n12034 & ~n12047 ) | ( n12035 & ~n12047 ) ;
  assign n12049 = n12032 & n12048 ;
  assign n12050 = ~n12000 & n12010 ;
  assign n12051 = ( ~n12009 & n12010 ) | ( ~n12009 & n12050 ) | ( n12010 & n12050 ) ;
  assign n12052 = ~n11982 & n11983 ;
  assign n12053 = ( ~n11979 & n11983 ) | ( ~n11979 & n12052 ) | ( n11983 & n12052 ) ;
  assign n12054 = ~n12051 & n12053 ;
  assign n12055 = n12051 & ~n12053 ;
  assign n12056 = n12054 | n12055 ;
  assign n12057 = n12030 | n12056 ;
  assign n12058 = n12049 | n12057 ;
  assign n12059 = n12030 & n12056 ;
  assign n12060 = ( n12049 & n12056 ) | ( n12049 & n12059 ) | ( n12056 & n12059 ) ;
  assign n12061 = n12058 & ~n12060 ;
  assign n12062 = n11912 & n11950 ;
  assign n12063 = ~n11909 & n11910 ;
  assign n12064 = ( ~n11906 & n11910 ) | ( ~n11906 & n12063 ) | ( n11910 & n12063 ) ;
  assign n12065 = ~n11928 & n11932 ;
  assign n12066 = ( n11932 & ~n11940 ) | ( n11932 & n12065 ) | ( ~n11940 & n12065 ) ;
  assign n12067 = ~n12064 & n12066 ;
  assign n12068 = n12064 & ~n12066 ;
  assign n12069 = n12067 | n12068 ;
  assign n12070 = n11945 | n12069 ;
  assign n12071 = n12062 | n12070 ;
  assign n12072 = n11945 & n12069 ;
  assign n12073 = ( n12062 & n12069 ) | ( n12062 & n12072 ) | ( n12069 & n12072 ) ;
  assign n12074 = n12071 & ~n12073 ;
  assign n12075 = n12061 | n12074 ;
  assign n12076 = n12046 & n12075 ;
  assign n12077 = n12058 & n12071 ;
  assign n12078 = n12060 | n12073 ;
  assign n12079 = n12077 & ~n12078 ;
  assign n12080 = ( n11945 & n12064 ) | ( n11945 & n12066 ) | ( n12064 & n12066 ) ;
  assign n12081 = n12064 | n12066 ;
  assign n12082 = ( n12062 & n12080 ) | ( n12062 & n12081 ) | ( n12080 & n12081 ) ;
  assign n12083 = ( n12030 & n12051 ) | ( n12030 & n12053 ) | ( n12051 & n12053 ) ;
  assign n12084 = n12051 | n12053 ;
  assign n12085 = ( n12049 & n12083 ) | ( n12049 & n12084 ) | ( n12083 & n12084 ) ;
  assign n12086 = ~n12082 & n12085 ;
  assign n12087 = n12082 & ~n12085 ;
  assign n12088 = n12086 | n12087 ;
  assign n12089 = n12079 | n12088 ;
  assign n12090 = n12076 | n12089 ;
  assign n12091 = n12075 | n12079 ;
  assign n12092 = ( n12046 & n12079 ) | ( n12046 & n12091 ) | ( n12079 & n12091 ) ;
  assign n12093 = n12088 & n12092 ;
  assign n12094 = n12090 & ~n12093 ;
  assign n12095 = n11885 | n12094 ;
  assign n12096 = n11813 & ~n11836 ;
  assign n12097 = n11833 & ~n12096 ;
  assign n12098 = n11749 & ~n11806 ;
  assign n12099 = ~n11749 & n11806 ;
  assign n12100 = n12098 | n12099 ;
  assign n12101 = n11958 & ~n12015 ;
  assign n12102 = ~n11958 & n12015 ;
  assign n12103 = n12101 | n12102 ;
  assign n12104 = n12100 & n12103 ;
  assign n12105 = ~n11807 & n11813 ;
  assign n12106 = n11813 & ~n11833 ;
  assign n12107 = n11742 | n11811 ;
  assign n12108 = n11833 | n12107 ;
  assign n12109 = ( n12105 & n12106 ) | ( n12105 & ~n12108 ) | ( n12106 & ~n12108 ) ;
  assign n12110 = n12104 | n12109 ;
  assign n12111 = n12097 | n12110 ;
  assign n12112 = n11951 | n12020 ;
  assign n12113 = ( n12016 & n12042 ) | ( n12016 & ~n12112 ) | ( n12042 & ~n12112 ) ;
  assign n12114 = ( ~n12042 & n12112 ) | ( ~n12042 & n12113 ) | ( n12112 & n12113 ) ;
  assign n12115 = ( ~n12016 & n12113 ) | ( ~n12016 & n12114 ) | ( n12113 & n12114 ) ;
  assign n12116 = n12111 & n12115 ;
  assign n12117 = n12097 | n12109 ;
  assign n12118 = n12104 & n12117 ;
  assign n12119 = ( n12045 & ~n12061 ) | ( n12045 & n12074 ) | ( ~n12061 & n12074 ) ;
  assign n12120 = n12061 & ~n12074 ;
  assign n12121 = ( n12043 & n12119 ) | ( n12043 & ~n12120 ) | ( n12119 & ~n12120 ) ;
  assign n12122 = ( ~n12046 & n12061 ) | ( ~n12046 & n12121 ) | ( n12061 & n12121 ) ;
  assign n12123 = ( ~n12074 & n12121 ) | ( ~n12074 & n12122 ) | ( n12121 & n12122 ) ;
  assign n12124 = ( n11836 & ~n11852 ) | ( n11836 & n11865 ) | ( ~n11852 & n11865 ) ;
  assign n12125 = n11852 & ~n11865 ;
  assign n12126 = ( n11834 & n12124 ) | ( n11834 & ~n12125 ) | ( n12124 & ~n12125 ) ;
  assign n12127 = ( ~n11837 & n11852 ) | ( ~n11837 & n12126 ) | ( n11852 & n12126 ) ;
  assign n12128 = ( ~n11865 & n12126 ) | ( ~n11865 & n12127 ) | ( n12126 & n12127 ) ;
  assign n12129 = ( n12118 & n12123 ) | ( n12118 & n12128 ) | ( n12123 & n12128 ) ;
  assign n12130 = n12123 | n12128 ;
  assign n12131 = ( n12116 & n12129 ) | ( n12116 & n12130 ) | ( n12129 & n12130 ) ;
  assign n12132 = n12095 & n12131 ;
  assign n12133 = n11881 & n12090 ;
  assign n12134 = n11884 | n12093 ;
  assign n12135 = n12133 & ~n12134 ;
  assign n12136 = n12082 & n12085 ;
  assign n12137 = n12082 | n12085 ;
  assign n12138 = n12136 | n12137 ;
  assign n12139 = ( n12092 & n12136 ) | ( n12092 & n12138 ) | ( n12136 & n12138 ) ;
  assign n12140 = n11873 & n11876 ;
  assign n12141 = n11873 | n11876 ;
  assign n12142 = n12140 | n12141 ;
  assign n12143 = ( n11883 & n12140 ) | ( n11883 & n12142 ) | ( n12140 & n12142 ) ;
  assign n12144 = n12139 & n12143 ;
  assign n12145 = n12143 & ~n12144 ;
  assign n12146 = ( n12139 & ~n12144 ) | ( n12139 & n12145 ) | ( ~n12144 & n12145 ) ;
  assign n12147 = n12135 | n12146 ;
  assign n12148 = n12132 | n12147 ;
  assign n12149 = n12132 | n12135 ;
  assign n12150 = n12146 & n12149 ;
  assign n12151 = n12148 & ~n12150 ;
  assign n12152 = n11676 | n12151 ;
  assign n12153 = n12100 & ~n12103 ;
  assign n12154 = ~n12100 & n12103 ;
  assign n12155 = n12153 | n12154 ;
  assign n12156 = n11625 & ~n11628 ;
  assign n12157 = ~n11625 & n11628 ;
  assign n12158 = n12156 | n12157 ;
  assign n12159 = n12155 & n12158 ;
  assign n12160 = ~n12111 & n12115 ;
  assign n12161 = ( n12115 & n12118 ) | ( n12115 & n12160 ) | ( n12118 & n12160 ) ;
  assign n12162 = ~n12104 & n12117 ;
  assign n12163 = n12104 & ~n12109 ;
  assign n12164 = ~n12097 & n12163 ;
  assign n12165 = ~n12115 & n12164 ;
  assign n12166 = ( ~n12115 & n12162 ) | ( ~n12115 & n12165 ) | ( n12162 & n12165 ) ;
  assign n12167 = n12161 | n12166 ;
  assign n12168 = n12159 & n12167 ;
  assign n12169 = n12159 | n12162 ;
  assign n12170 = n12115 & ~n12159 ;
  assign n12171 = ( n12165 & n12169 ) | ( n12165 & ~n12170 ) | ( n12169 & ~n12170 ) ;
  assign n12172 = n12161 | n12171 ;
  assign n12173 = ~n11629 & n11642 ;
  assign n12174 = n11629 & ~n11634 ;
  assign n12175 = ~n11622 & n12174 ;
  assign n12176 = ~n11640 & n12175 ;
  assign n12177 = ( ~n11640 & n12173 ) | ( ~n11640 & n12176 ) | ( n12173 & n12176 ) ;
  assign n12178 = n11641 & ~n11643 ;
  assign n12179 = ( n11640 & n12177 ) | ( n11640 & ~n12178 ) | ( n12177 & ~n12178 ) ;
  assign n12180 = n12172 & n12179 ;
  assign n12181 = n12168 | n12180 ;
  assign n12183 = ( n11643 & ~n11648 ) | ( n11643 & n11653 ) | ( ~n11648 & n11653 ) ;
  assign n12184 = n11648 & ~n11653 ;
  assign n12185 = ( n11641 & n12183 ) | ( n11641 & ~n12184 ) | ( n12183 & ~n12184 ) ;
  assign n12182 = n11641 | n11643 ;
  assign n12186 = ( n11648 & ~n12182 ) | ( n11648 & n12185 ) | ( ~n12182 & n12185 ) ;
  assign n12187 = ( ~n11653 & n12185 ) | ( ~n11653 & n12186 ) | ( n12185 & n12186 ) ;
  assign n12189 = ( n12118 & ~n12123 ) | ( n12118 & n12128 ) | ( ~n12123 & n12128 ) ;
  assign n12190 = n12123 & ~n12128 ;
  assign n12191 = ( n12116 & n12189 ) | ( n12116 & ~n12190 ) | ( n12189 & ~n12190 ) ;
  assign n12188 = n12116 | n12118 ;
  assign n12192 = ( n12123 & ~n12188 ) | ( n12123 & n12191 ) | ( ~n12188 & n12191 ) ;
  assign n12193 = ( ~n12128 & n12191 ) | ( ~n12128 & n12192 ) | ( n12191 & n12192 ) ;
  assign n12194 = ( n12181 & n12187 ) | ( n12181 & n12193 ) | ( n12187 & n12193 ) ;
  assign n12195 = ( ~n11885 & n12094 ) | ( ~n11885 & n12131 ) | ( n12094 & n12131 ) ;
  assign n12196 = ( n11885 & ~n12131 ) | ( n11885 & n12195 ) | ( ~n12131 & n12195 ) ;
  assign n12197 = ( ~n12094 & n12195 ) | ( ~n12094 & n12196 ) | ( n12195 & n12196 ) ;
  assign n12198 = ( ~n11410 & n11619 ) | ( ~n11410 & n11656 ) | ( n11619 & n11656 ) ;
  assign n12199 = ( n11410 & ~n11656 ) | ( n11410 & n12198 ) | ( ~n11656 & n12198 ) ;
  assign n12200 = ( ~n11619 & n12198 ) | ( ~n11619 & n12199 ) | ( n12198 & n12199 ) ;
  assign n12201 = ( n12194 & n12197 ) | ( n12194 & n12200 ) | ( n12197 & n12200 ) ;
  assign n12202 = n12152 & n12201 ;
  assign n12203 = n11673 & n12148 ;
  assign n12204 = n11675 | n12150 ;
  assign n12205 = n12203 & ~n12204 ;
  assign n12214 = n11408 & n11666 ;
  assign n12215 = n11610 | n11665 ;
  assign n12216 = n11607 | n11665 ;
  assign n12217 = ( n11617 & n12215 ) | ( n11617 & n12216 ) | ( n12215 & n12216 ) ;
  assign n12218 = n12214 | n12217 ;
  assign n12219 = n11669 | n12218 ;
  assign n12220 = ( n11660 & n11669 ) | ( n11660 & n12219 ) | ( n11669 & n12219 ) ;
  assign n12221 = n11669 | n12219 ;
  assign n12222 = ( n11657 & n12220 ) | ( n11657 & n12221 ) | ( n12220 & n12221 ) ;
  assign n12206 = n11883 & n12141 ;
  assign n12207 = n12085 | n12140 ;
  assign n12208 = n12082 | n12140 ;
  assign n12209 = ( n12092 & n12207 ) | ( n12092 & n12208 ) | ( n12207 & n12208 ) ;
  assign n12210 = n12206 | n12209 ;
  assign n12211 = n12135 & n12210 ;
  assign n12212 = ( n12132 & n12210 ) | ( n12132 & n12211 ) | ( n12210 & n12211 ) ;
  assign n12213 = n12144 | n12212 ;
  assign n12223 = n12213 & n12222 ;
  assign n12224 = n12213 & ~n12223 ;
  assign n12225 = ( n12222 & ~n12223 ) | ( n12222 & n12224 ) | ( ~n12223 & n12224 ) ;
  assign n12226 = n12205 | n12225 ;
  assign n12227 = n12202 | n12226 ;
  assign n12228 = n12202 | n12205 ;
  assign n12229 = n12225 & n12228 ;
  assign n12230 = n12227 & ~n12229 ;
  assign n12231 = n11201 | n12230 ;
  assign n12232 = ( ~n11676 & n12151 ) | ( ~n11676 & n12201 ) | ( n12151 & n12201 ) ;
  assign n12233 = ( n11676 & ~n12201 ) | ( n11676 & n12232 ) | ( ~n12201 & n12232 ) ;
  assign n12234 = ( ~n12151 & n12232 ) | ( ~n12151 & n12233 ) | ( n12232 & n12233 ) ;
  assign n12235 = ( ~n10649 & n11124 ) | ( ~n10649 & n11172 ) | ( n11124 & n11172 ) ;
  assign n12236 = ( n10649 & ~n11172 ) | ( n10649 & n12235 ) | ( ~n11172 & n12235 ) ;
  assign n12237 = ( ~n11124 & n12235 ) | ( ~n11124 & n12236 ) | ( n12235 & n12236 ) ;
  assign n12238 = n11141 & ~n11144 ;
  assign n12239 = ~n11141 & n11144 ;
  assign n12240 = n12238 | n12239 ;
  assign n12241 = n12155 & ~n12158 ;
  assign n12242 = ~n12155 & n12158 ;
  assign n12243 = n12241 | n12242 ;
  assign n12244 = n12240 & n12243 ;
  assign n12245 = n11154 & ~n11156 ;
  assign n12246 = n11138 & ~n12245 ;
  assign n12247 = ~n11145 & n11153 ;
  assign n12248 = n11145 & ~n11153 ;
  assign n12249 = n12247 | n12248 ;
  assign n12250 = ~n11138 & n12249 ;
  assign n12251 = n12246 | n12250 ;
  assign n12252 = n12244 & n12251 ;
  assign n12253 = n11138 & ~n12244 ;
  assign n12254 = ( n12244 & n12249 ) | ( n12244 & ~n12253 ) | ( n12249 & ~n12253 ) ;
  assign n12255 = n12246 | n12254 ;
  assign n12256 = ( n12159 & ~n12167 ) | ( n12159 & n12179 ) | ( ~n12167 & n12179 ) ;
  assign n12257 = ( ~n12159 & n12167 ) | ( ~n12159 & n12256 ) | ( n12167 & n12256 ) ;
  assign n12258 = ( ~n12179 & n12256 ) | ( ~n12179 & n12257 ) | ( n12256 & n12257 ) ;
  assign n12259 = n12255 & n12258 ;
  assign n12260 = n12252 | n12259 ;
  assign n12261 = ( n12181 & ~n12187 ) | ( n12181 & n12193 ) | ( ~n12187 & n12193 ) ;
  assign n12262 = ( ~n12181 & n12187 ) | ( ~n12181 & n12261 ) | ( n12187 & n12261 ) ;
  assign n12263 = ( ~n12193 & n12261 ) | ( ~n12193 & n12262 ) | ( n12261 & n12262 ) ;
  assign n12265 = ( n11156 & ~n11162 ) | ( n11156 & n11168 ) | ( ~n11162 & n11168 ) ;
  assign n12266 = n11162 & ~n11168 ;
  assign n12267 = ( n11155 & n12265 ) | ( n11155 & ~n12266 ) | ( n12265 & ~n12266 ) ;
  assign n12264 = n11155 | n11156 ;
  assign n12268 = ( n11162 & ~n12264 ) | ( n11162 & n12267 ) | ( ~n12264 & n12267 ) ;
  assign n12269 = ( ~n11168 & n12267 ) | ( ~n11168 & n12268 ) | ( n12267 & n12268 ) ;
  assign n12270 = ( n12260 & n12263 ) | ( n12260 & n12269 ) | ( n12263 & n12269 ) ;
  assign n12271 = ( ~n11128 & n11131 ) | ( ~n11128 & n11171 ) | ( n11131 & n11171 ) ;
  assign n12272 = ( n11128 & ~n11171 ) | ( n11128 & n12271 ) | ( ~n11171 & n12271 ) ;
  assign n12273 = ( ~n11131 & n12271 ) | ( ~n11131 & n12272 ) | ( n12271 & n12272 ) ;
  assign n12274 = ( n12194 & ~n12197 ) | ( n12194 & n12200 ) | ( ~n12197 & n12200 ) ;
  assign n12275 = ( ~n12194 & n12197 ) | ( ~n12194 & n12274 ) | ( n12197 & n12274 ) ;
  assign n12276 = ( ~n12200 & n12274 ) | ( ~n12200 & n12275 ) | ( n12274 & n12275 ) ;
  assign n12277 = ( n12270 & n12273 ) | ( n12270 & n12276 ) | ( n12273 & n12276 ) ;
  assign n12278 = ( n12234 & n12237 ) | ( n12234 & n12277 ) | ( n12237 & n12277 ) ;
  assign n12279 = n12231 & n12278 ;
  assign n12280 = n11198 & n12227 ;
  assign n12281 = n11200 | n12229 ;
  assign n12282 = n12280 & ~n12281 ;
  assign n12290 = n11669 | n12144 ;
  assign n12291 = n12218 | n12290 ;
  assign n12292 = ( n11674 & n12290 ) | ( n11674 & n12291 ) | ( n12290 & n12291 ) ;
  assign n12293 = n12212 | n12292 ;
  assign n12294 = n12223 | n12293 ;
  assign n12295 = ( n12205 & n12223 ) | ( n12205 & n12294 ) | ( n12223 & n12294 ) ;
  assign n12296 = n12223 | n12294 ;
  assign n12297 = ( n12202 & n12295 ) | ( n12202 & n12296 ) | ( n12295 & n12296 ) ;
  assign n12283 = n10642 | n11117 ;
  assign n12284 = n11189 | n12283 ;
  assign n12285 = ( n10647 & n12283 ) | ( n10647 & n12284 ) | ( n12283 & n12284 ) ;
  assign n12286 = n11183 | n12285 ;
  assign n12287 = n11176 & n12286 ;
  assign n12288 = ( n11173 & n12286 ) | ( n11173 & n12287 ) | ( n12286 & n12287 ) ;
  assign n12289 = n11194 | n12288 ;
  assign n12298 = n12289 & n12297 ;
  assign n12299 = n12289 & ~n12298 ;
  assign n12300 = ( n12297 & ~n12298 ) | ( n12297 & n12299 ) | ( ~n12298 & n12299 ) ;
  assign n12301 = n12282 | n12300 ;
  assign n12302 = n12279 | n12301 ;
  assign n12303 = n10174 & n12302 ;
  assign n12304 = n10151 | n10154 ;
  assign n12305 = n10172 & n12304 ;
  assign n12306 = n12279 | n12282 ;
  assign n12307 = n12300 & n12306 ;
  assign n12308 = n12305 | n12307 ;
  assign n12309 = n12303 & ~n12308 ;
  assign n12310 = n10174 & ~n12305 ;
  assign n12311 = n12302 & ~n12307 ;
  assign n12312 = n12310 | n12311 ;
  assign n12313 = ( ~n11201 & n12230 ) | ( ~n11201 & n12278 ) | ( n12230 & n12278 ) ;
  assign n12314 = ( n11201 & ~n12278 ) | ( n11201 & n12313 ) | ( ~n12278 & n12313 ) ;
  assign n12315 = ( ~n12230 & n12313 ) | ( ~n12230 & n12314 ) | ( n12313 & n12314 ) ;
  assign n12316 = ( ~n9073 & n10102 ) | ( ~n9073 & n10150 ) | ( n10102 & n10150 ) ;
  assign n12317 = ( n9073 & ~n10150 ) | ( n9073 & n12316 ) | ( ~n10150 & n12316 ) ;
  assign n12318 = ( ~n10102 & n12316 ) | ( ~n10102 & n12317 ) | ( n12316 & n12317 ) ;
  assign n12319 = n10112 & ~n10115 ;
  assign n12320 = ~n10112 & n10115 ;
  assign n12321 = n12319 | n12320 ;
  assign n12322 = n12240 & ~n12243 ;
  assign n12323 = ~n12240 & n12243 ;
  assign n12324 = n12322 | n12323 ;
  assign n12325 = n12321 & n12324 ;
  assign n12326 = ~n12255 & n12258 ;
  assign n12327 = ( n12252 & n12258 ) | ( n12252 & n12326 ) | ( n12258 & n12326 ) ;
  assign n12328 = ~n12244 & n12251 ;
  assign n12329 = n11138 & n12244 ;
  assign n12330 = ( n12244 & ~n12249 ) | ( n12244 & n12329 ) | ( ~n12249 & n12329 ) ;
  assign n12331 = ~n12246 & n12330 ;
  assign n12332 = ~n12258 & n12331 ;
  assign n12333 = ( ~n12258 & n12328 ) | ( ~n12258 & n12332 ) | ( n12328 & n12332 ) ;
  assign n12334 = n12327 | n12333 ;
  assign n12335 = n12325 & n12334 ;
  assign n12336 = n12325 | n12333 ;
  assign n12337 = n12327 | n12336 ;
  assign n12338 = ~n10116 & n10123 ;
  assign n12339 = n9010 & n10116 ;
  assign n12340 = ( n10116 & ~n10121 ) | ( n10116 & n12339 ) | ( ~n10121 & n12339 ) ;
  assign n12341 = ~n10118 & n12340 ;
  assign n12342 = ~n10130 & n12341 ;
  assign n12343 = ( ~n10130 & n12338 ) | ( ~n10130 & n12342 ) | ( n12338 & n12342 ) ;
  assign n12344 = ~n10124 & n10131 ;
  assign n12345 = ( n10130 & n12343 ) | ( n10130 & ~n12344 ) | ( n12343 & ~n12344 ) ;
  assign n12346 = n12337 & n12345 ;
  assign n12347 = n12335 | n12346 ;
  assign n12348 = ( n10132 & ~n10135 ) | ( n10132 & n10141 ) | ( ~n10135 & n10141 ) ;
  assign n12349 = ( ~n10132 & n10135 ) | ( ~n10132 & n12348 ) | ( n10135 & n12348 ) ;
  assign n12350 = ( ~n10141 & n12348 ) | ( ~n10141 & n12349 ) | ( n12348 & n12349 ) ;
  assign n12351 = ( n12260 & ~n12263 ) | ( n12260 & n12269 ) | ( ~n12263 & n12269 ) ;
  assign n12352 = ( ~n12260 & n12263 ) | ( ~n12260 & n12351 ) | ( n12263 & n12351 ) ;
  assign n12353 = ( ~n12269 & n12351 ) | ( ~n12269 & n12352 ) | ( n12351 & n12352 ) ;
  assign n12354 = ( n12347 & n12350 ) | ( n12347 & n12353 ) | ( n12350 & n12353 ) ;
  assign n12355 = ( n10106 & ~n10109 ) | ( n10106 & n10149 ) | ( ~n10109 & n10149 ) ;
  assign n12356 = ( ~n10106 & n10109 ) | ( ~n10106 & n10149 ) | ( n10109 & n10149 ) ;
  assign n12357 = ( ~n10149 & n12355 ) | ( ~n10149 & n12356 ) | ( n12355 & n12356 ) ;
  assign n12358 = ( n12234 & ~n12237 ) | ( n12234 & n12277 ) | ( ~n12237 & n12277 ) ;
  assign n12359 = ( ~n12234 & n12237 ) | ( ~n12234 & n12277 ) | ( n12237 & n12277 ) ;
  assign n12360 = ( ~n12277 & n12358 ) | ( ~n12277 & n12359 ) | ( n12358 & n12359 ) ;
  assign n12361 = ( n10142 & ~n10145 ) | ( n10142 & n10148 ) | ( ~n10145 & n10148 ) ;
  assign n12362 = ( ~n10142 & n10145 ) | ( ~n10142 & n12361 ) | ( n10145 & n12361 ) ;
  assign n12363 = ( ~n10148 & n12361 ) | ( ~n10148 & n12362 ) | ( n12361 & n12362 ) ;
  assign n12364 = ( n12357 & n12360 ) | ( n12357 & n12363 ) | ( n12360 & n12363 ) ;
  assign n12365 = ( n12270 & ~n12273 ) | ( n12270 & n12276 ) | ( ~n12273 & n12276 ) ;
  assign n12366 = ( ~n12270 & n12273 ) | ( ~n12270 & n12365 ) | ( n12273 & n12365 ) ;
  assign n12367 = ( ~n12276 & n12365 ) | ( ~n12276 & n12366 ) | ( n12365 & n12366 ) ;
  assign n12368 = ( n12357 & n12360 ) | ( n12357 & n12367 ) | ( n12360 & n12367 ) ;
  assign n12369 = ( n12354 & n12364 ) | ( n12354 & n12368 ) | ( n12364 & n12368 ) ;
  assign n12370 = ( n12315 & n12318 ) | ( n12315 & n12369 ) | ( n12318 & n12369 ) ;
  assign n12371 = n12312 & n12370 ;
  assign n12372 = n12309 | n12371 ;
  assign n12380 = n9066 | n10095 ;
  assign n12381 = n10165 | n12380 ;
  assign n12382 = ( n10100 & n12380 ) | ( n10100 & n12381 ) | ( n12380 & n12381 ) ;
  assign n12383 = n10160 | n12382 ;
  assign n12384 = n10170 | n12383 ;
  assign n12385 = ( n10154 & n10170 ) | ( n10154 & n12384 ) | ( n10170 & n12384 ) ;
  assign n12386 = n10170 | n12384 ;
  assign n12387 = ( n10151 & n12385 ) | ( n10151 & n12386 ) | ( n12385 & n12386 ) ;
  assign n12373 = n11194 | n12223 ;
  assign n12374 = n12293 | n12373 ;
  assign n12375 = ( n12228 & n12373 ) | ( n12228 & n12374 ) | ( n12373 & n12374 ) ;
  assign n12376 = n12288 | n12375 ;
  assign n12377 = n12282 & n12376 ;
  assign n12378 = ( n12279 & n12376 ) | ( n12279 & n12377 ) | ( n12376 & n12377 ) ;
  assign n12379 = n12298 | n12378 ;
  assign n12388 = n12379 & n12387 ;
  assign n12389 = n12379 & ~n12388 ;
  assign n12390 = ( n12387 & ~n12388 ) | ( n12387 & n12389 ) | ( ~n12388 & n12389 ) ;
  assign n12391 = n12372 & n12390 ;
  assign n12392 = n12309 | n12390 ;
  assign n12393 = n12371 | n12392 ;
  assign n12394 = ~n12391 & n12393 ;
  assign n12395 = ~n8007 & n12394 ;
  assign n12396 = ( ~n8045 & n12394 ) | ( ~n8045 & n12395 ) | ( n12394 & n12395 ) ;
  assign n12397 = n8046 & n12396 ;
  assign n12398 = n8007 & n8045 ;
  assign n12399 = n8046 & ~n12398 ;
  assign n12400 = n12394 | n12399 ;
  assign n12401 = ~n3612 & n7934 ;
  assign n12402 = n3612 & ~n7934 ;
  assign n12403 = n12401 | n12402 ;
  assign n12404 = n8006 | n12403 ;
  assign n12405 = ( ~n12310 & n12311 ) | ( ~n12310 & n12370 ) | ( n12311 & n12370 ) ;
  assign n12406 = ( n12310 & ~n12370 ) | ( n12310 & n12405 ) | ( ~n12370 & n12405 ) ;
  assign n12407 = ( ~n12311 & n12405 ) | ( ~n12311 & n12406 ) | ( n12405 & n12406 ) ;
  assign n12408 = ~n8006 & n12407 ;
  assign n12409 = ( ~n12403 & n12407 ) | ( ~n12403 & n12408 ) | ( n12407 & n12408 ) ;
  assign n12410 = n12404 & n12409 ;
  assign n12411 = n8006 & n12403 ;
  assign n12412 = n12404 & ~n12411 ;
  assign n12413 = n12407 | n12412 ;
  assign n12414 = n7942 & n7945 ;
  assign n12415 = ~n7942 & n7945 ;
  assign n12416 = ( n7942 & ~n12414 ) | ( n7942 & n12415 ) | ( ~n12414 & n12415 ) ;
  assign n12417 = n8005 | n12416 ;
  assign n12418 = ( n12315 & ~n12318 ) | ( n12315 & n12369 ) | ( ~n12318 & n12369 ) ;
  assign n12419 = ( ~n12315 & n12318 ) | ( ~n12315 & n12418 ) | ( n12318 & n12418 ) ;
  assign n12420 = ( ~n12369 & n12418 ) | ( ~n12369 & n12419 ) | ( n12418 & n12419 ) ;
  assign n12421 = ~n8005 & n12420 ;
  assign n12422 = ( ~n12416 & n12420 ) | ( ~n12416 & n12421 ) | ( n12420 & n12421 ) ;
  assign n12423 = n12417 & n12422 ;
  assign n12424 = n8005 & n12416 ;
  assign n12425 = n12417 & ~n12424 ;
  assign n12426 = n12420 | n12425 ;
  assign n12427 = ~n7952 & n8004 ;
  assign n12428 = n7952 & ~n8004 ;
  assign n12429 = n12427 | n12428 ;
  assign n12430 = n7998 | n12429 ;
  assign n12431 = ( n12354 & n12363 ) | ( n12354 & n12367 ) | ( n12363 & n12367 ) ;
  assign n12432 = ( n12357 & ~n12360 ) | ( n12357 & n12363 ) | ( ~n12360 & n12363 ) ;
  assign n12433 = ( n12357 & ~n12360 ) | ( n12357 & n12367 ) | ( ~n12360 & n12367 ) ;
  assign n12434 = ( n12354 & n12432 ) | ( n12354 & n12433 ) | ( n12432 & n12433 ) ;
  assign n12435 = ( ~n12357 & n12360 ) | ( ~n12357 & n12434 ) | ( n12360 & n12434 ) ;
  assign n12436 = ( ~n12431 & n12434 ) | ( ~n12431 & n12435 ) | ( n12434 & n12435 ) ;
  assign n12437 = ~n7998 & n12436 ;
  assign n12438 = ( ~n12429 & n12436 ) | ( ~n12429 & n12437 ) | ( n12436 & n12437 ) ;
  assign n12439 = n12430 & n12438 ;
  assign n12440 = n7998 & n12429 ;
  assign n12441 = n12430 & ~n12440 ;
  assign n12442 = n12436 | n12441 ;
  assign n12443 = n7961 & n7997 ;
  assign n12444 = n7997 & ~n12443 ;
  assign n12445 = ~n7994 & n12443 ;
  assign n12446 = n7961 | n7994 ;
  assign n12447 = ( n12444 & ~n12445 ) | ( n12444 & n12446 ) | ( ~n12445 & n12446 ) ;
  assign n12448 = n7994 & ~n12443 ;
  assign n12449 = n7961 & n7994 ;
  assign n12450 = ( n12444 & n12448 ) | ( n12444 & n12449 ) | ( n12448 & n12449 ) ;
  assign n12451 = n12447 & ~n12450 ;
  assign n12452 = ( n12354 & n12363 ) | ( n12354 & ~n12367 ) | ( n12363 & ~n12367 ) ;
  assign n12453 = ( ~n12354 & n12367 ) | ( ~n12354 & n12452 ) | ( n12367 & n12452 ) ;
  assign n12454 = ( ~n12363 & n12452 ) | ( ~n12363 & n12453 ) | ( n12452 & n12453 ) ;
  assign n12455 = n12451 | n12454 ;
  assign n12456 = ~n7967 & n7993 ;
  assign n12457 = n7967 & ~n7993 ;
  assign n12458 = n12456 | n12457 ;
  assign n12459 = n7990 | n12458 ;
  assign n12460 = n7990 & n12458 ;
  assign n12461 = n12459 & ~n12460 ;
  assign n12462 = ( n12347 & ~n12350 ) | ( n12347 & n12353 ) | ( ~n12350 & n12353 ) ;
  assign n12463 = ( ~n12347 & n12350 ) | ( ~n12347 & n12462 ) | ( n12350 & n12462 ) ;
  assign n12464 = ( ~n12353 & n12462 ) | ( ~n12353 & n12463 ) | ( n12462 & n12463 ) ;
  assign n12465 = ( n7990 & n12458 ) | ( n7990 & ~n12464 ) | ( n12458 & ~n12464 ) ;
  assign n12466 = ~n7985 & n7988 ;
  assign n12467 = ( n7982 & n7988 ) | ( n7982 & n12466 ) | ( n7988 & n12466 ) ;
  assign n12468 = ~n7974 & n7981 ;
  assign n12469 = n7905 & n7974 ;
  assign n12470 = ( n7974 & ~n7979 ) | ( n7974 & n12469 ) | ( ~n7979 & n12469 ) ;
  assign n12471 = ~n7976 & n12470 ;
  assign n12472 = ~n7988 & n12471 ;
  assign n12473 = ( ~n7988 & n12468 ) | ( ~n7988 & n12472 ) | ( n12468 & n12472 ) ;
  assign n12474 = n12467 | n12473 ;
  assign n12475 = ( n12325 & ~n12334 ) | ( n12325 & n12345 ) | ( ~n12334 & n12345 ) ;
  assign n12476 = ( ~n12325 & n12334 ) | ( ~n12325 & n12475 ) | ( n12334 & n12475 ) ;
  assign n12477 = ( ~n12345 & n12475 ) | ( ~n12345 & n12476 ) | ( n12475 & n12476 ) ;
  assign n12478 = n12464 & n12477 ;
  assign n12479 = n12321 & ~n12324 ;
  assign n12480 = ~n12321 & n12324 ;
  assign n12481 = n12479 | n12480 ;
  assign n12482 = n7970 & ~n7973 ;
  assign n12483 = ~n7970 & n7973 ;
  assign n12484 = n12482 | n12483 ;
  assign n12485 = n12481 & n12484 ;
  assign n12486 = n12464 & n12485 ;
  assign n12487 = ( n12474 & n12478 ) | ( n12474 & n12486 ) | ( n12478 & n12486 ) ;
  assign n12488 = ( n12459 & ~n12465 ) | ( n12459 & n12487 ) | ( ~n12465 & n12487 ) ;
  assign n12489 = ( n12474 & n12477 ) | ( n12474 & n12485 ) | ( n12477 & n12485 ) ;
  assign n12490 = ( n12459 & ~n12465 ) | ( n12459 & n12489 ) | ( ~n12465 & n12489 ) ;
  assign n12491 = ( n12461 & n12488 ) | ( n12461 & n12490 ) | ( n12488 & n12490 ) ;
  assign n12492 = ( ~n7994 & n12443 ) | ( ~n7994 & n12454 ) | ( n12443 & n12454 ) ;
  assign n12493 = ( n7961 & n7994 ) | ( n7961 & ~n12454 ) | ( n7994 & ~n12454 ) ;
  assign n12494 = ( n12444 & ~n12492 ) | ( n12444 & n12493 ) | ( ~n12492 & n12493 ) ;
  assign n12495 = ( n12447 & n12491 ) | ( n12447 & ~n12494 ) | ( n12491 & ~n12494 ) ;
  assign n12496 = n12447 & ~n12494 ;
  assign n12497 = ( n12455 & n12495 ) | ( n12455 & n12496 ) | ( n12495 & n12496 ) ;
  assign n12498 = ( n12439 & n12442 ) | ( n12439 & n12497 ) | ( n12442 & n12497 ) ;
  assign n12499 = ( n12423 & n12426 ) | ( n12423 & n12498 ) | ( n12426 & n12498 ) ;
  assign n12500 = ( n12410 & n12413 ) | ( n12410 & n12499 ) | ( n12413 & n12499 ) ;
  assign n12501 = n12400 & n12500 ;
  assign n12502 = n12397 | n12501 ;
  assign n12503 = n8007 & n8044 ;
  assign n12504 = n5736 | n7867 ;
  assign n12505 = n8024 | n12504 ;
  assign n12506 = ( n7872 & n12504 ) | ( n7872 & n12505 ) | ( n12504 & n12505 ) ;
  assign n12507 = n8019 | n12506 ;
  assign n12508 = n8010 & n12507 ;
  assign n12509 = ( n8012 & n12507 ) | ( n8012 & n12508 ) | ( n12507 & n12508 ) ;
  assign n12510 = n3523 | n8029 ;
  assign n12511 = n8029 | n8033 ;
  assign n12512 = ( n3610 & n12510 ) | ( n3610 & n12511 ) | ( n12510 & n12511 ) ;
  assign n12513 = n12509 | n12512 ;
  assign n12514 = n8029 | n12509 ;
  assign n12515 = n8034 & n12514 ;
  assign n12516 = n12513 & ~n12515 ;
  assign n12517 = n8042 | n12516 ;
  assign n12518 = n12503 | n12517 ;
  assign n12522 = n10170 | n12298 ;
  assign n12523 = n12383 | n12522 ;
  assign n12524 = ( n12304 & n12522 ) | ( n12304 & n12523 ) | ( n12522 & n12523 ) ;
  assign n12525 = n12378 | n12524 ;
  assign n12526 = n12388 | n12525 ;
  assign n12527 = ( n12309 & n12388 ) | ( n12309 & n12526 ) | ( n12388 & n12526 ) ;
  assign n12528 = n12388 | n12526 ;
  assign n12529 = ( n12371 & n12527 ) | ( n12371 & n12528 ) | ( n12527 & n12528 ) ;
  assign n12531 = n12518 & n12529 ;
  assign n12532 = n12513 | n12515 ;
  assign n12533 = ( n8042 & n12515 ) | ( n8042 & n12532 ) | ( n12515 & n12532 ) ;
  assign n12534 = n12515 | n12532 ;
  assign n12535 = ( n12503 & n12533 ) | ( n12503 & n12534 ) | ( n12533 & n12534 ) ;
  assign n12519 = n8042 & n12516 ;
  assign n12520 = ( n12503 & n12516 ) | ( n12503 & n12519 ) | ( n12516 & n12519 ) ;
  assign n12536 = n12520 & n12535 ;
  assign n12537 = ( ~n12531 & n12535 ) | ( ~n12531 & n12536 ) | ( n12535 & n12536 ) ;
  assign n12521 = n12518 & ~n12520 ;
  assign n12530 = n12521 | n12529 ;
  assign n12538 = ~n12530 & n12537 ;
  assign n12539 = ( ~n12502 & n12537 ) | ( ~n12502 & n12538 ) | ( n12537 & n12538 ) ;
  assign n12540 = ~n12520 & n12531 ;
  assign n12541 = n12530 | n12540 ;
  assign n12542 = ~n12535 & n12541 ;
  assign n12543 = ~n12535 & n12540 ;
  assign n12544 = ( n12502 & n12542 ) | ( n12502 & n12543 ) | ( n12542 & n12543 ) ;
  assign n12545 = n12539 | n12544 ;
  assign n12546 = ~n12521 & n12529 ;
  assign n12547 = n12518 & ~n12529 ;
  assign n12548 = ~n12520 & n12547 ;
  assign n12549 = n12546 | n12548 ;
  assign n12550 = n12502 & n12549 ;
  assign n12551 = n12397 | n12549 ;
  assign n12552 = n12501 | n12551 ;
  assign n12553 = ~n12550 & n12552 ;
  assign n12554 = ~n12451 & n12454 ;
  assign n12555 = n12450 | n12454 ;
  assign n12556 = n12447 & ~n12555 ;
  assign n12557 = n12554 | n12556 ;
  assign n12558 = n12491 | n12557 ;
  assign n12559 = n12491 & n12557 ;
  assign n12560 = n12481 & ~n12482 ;
  assign n12561 = ~n12483 & n12560 ;
  assign n12562 = ~n12481 & n12484 ;
  assign n12563 = n12561 | n12562 ;
  assign n12564 = x1000 & n12563 ;
  assign n12565 = ~n12461 & n12464 ;
  assign n12566 = n7990 | n12464 ;
  assign n12567 = ( n12458 & n12464 ) | ( n12458 & n12566 ) | ( n12464 & n12566 ) ;
  assign n12568 = n12459 & ~n12567 ;
  assign n12569 = n12489 & n12568 ;
  assign n12570 = ( n12489 & n12565 ) | ( n12489 & n12569 ) | ( n12565 & n12569 ) ;
  assign n12571 = n12564 & ~n12570 ;
  assign n12572 = n12474 & ~n12485 ;
  assign n12573 = ~n12474 & n12485 ;
  assign n12574 = n12572 | n12573 ;
  assign n12575 = ~n12477 & n12574 ;
  assign n12576 = n12474 & n12485 ;
  assign n12577 = n12473 | n12485 ;
  assign n12578 = n12467 | n12577 ;
  assign n12579 = ~n12576 & n12578 ;
  assign n12580 = n12477 & ~n12579 ;
  assign n12581 = n12575 | n12580 ;
  assign n12582 = n12489 | n12568 ;
  assign n12583 = n12565 | n12582 ;
  assign n12584 = n12581 & n12583 ;
  assign n12585 = n12571 & n12584 ;
  assign n12586 = ~n12559 & n12585 ;
  assign n12587 = n12558 & n12586 ;
  assign n12588 = ( n12436 & n12441 ) | ( n12436 & ~n12497 ) | ( n12441 & ~n12497 ) ;
  assign n12589 = ( ~n12441 & n12497 ) | ( ~n12441 & n12588 ) | ( n12497 & n12588 ) ;
  assign n12590 = ( ~n12436 & n12588 ) | ( ~n12436 & n12589 ) | ( n12588 & n12589 ) ;
  assign n12591 = n12587 & n12590 ;
  assign n12592 = ( n12420 & n12425 ) | ( n12420 & n12498 ) | ( n12425 & n12498 ) ;
  assign n12593 = ( n12425 & n12498 ) | ( n12425 & ~n12592 ) | ( n12498 & ~n12592 ) ;
  assign n12594 = ( n12420 & ~n12592 ) | ( n12420 & n12593 ) | ( ~n12592 & n12593 ) ;
  assign n12595 = n12591 & n12594 ;
  assign n12596 = ( n12407 & n12412 ) | ( n12407 & n12499 ) | ( n12412 & n12499 ) ;
  assign n12597 = ( n12412 & n12499 ) | ( n12412 & ~n12596 ) | ( n12499 & ~n12596 ) ;
  assign n12598 = ( n12407 & ~n12596 ) | ( n12407 & n12597 ) | ( ~n12596 & n12597 ) ;
  assign n12599 = n12595 & n12598 ;
  assign n12600 = ( n12394 & n12399 ) | ( n12394 & n12500 ) | ( n12399 & n12500 ) ;
  assign n12601 = ( n12399 & n12500 ) | ( n12399 & ~n12600 ) | ( n12500 & ~n12600 ) ;
  assign n12602 = ( n12394 & ~n12600 ) | ( n12394 & n12601 ) | ( ~n12600 & n12601 ) ;
  assign n12603 = n12599 & n12602 ;
  assign n12604 = n12553 & n12603 ;
  assign n12605 = ~n12545 & n12604 ;
  assign n12606 = n12545 & ~n12604 ;
  assign n12607 = n12605 | n12606 ;
  assign n12608 = n12553 | n12603 ;
  assign n12609 = ~n12604 & n12608 ;
  assign n12610 = n12599 | n12602 ;
  assign n12611 = ~n12603 & n12610 ;
  assign n12612 = n12558 & ~n12559 ;
  assign n12613 = n12585 | n12612 ;
  assign n12614 = ~n12570 & n12583 ;
  assign n12615 = n12564 & n12581 ;
  assign n12616 = n12614 | n12615 ;
  assign n12617 = ~n12585 & n12616 ;
  assign n12618 = ( n12564 & n12575 ) | ( n12564 & n12580 ) | ( n12575 & n12580 ) ;
  assign n12619 = ( n12564 & n12575 ) | ( n12564 & ~n12618 ) | ( n12575 & ~n12618 ) ;
  assign n12620 = ( n12580 & ~n12618 ) | ( n12580 & n12619 ) | ( ~n12618 & n12619 ) ;
  assign n12621 = n12617 | n12620 ;
  assign n12622 = ~n12587 & n12621 ;
  assign n12623 = n12613 & n12622 ;
  assign n12624 = n12587 | n12590 ;
  assign n12625 = ~n12591 & n12624 ;
  assign n12626 = n12623 | n12625 ;
  assign n12627 = n12591 | n12594 ;
  assign n12628 = ~n12595 & n12627 ;
  assign n12629 = n12626 & n12628 ;
  assign n12630 = n12595 | n12598 ;
  assign n12631 = ~n12599 & n12630 ;
  assign n12632 = n12629 & n12631 ;
  assign n12633 = n12611 & n12632 ;
  assign n12634 = n12609 & n12633 ;
  assign n12635 = n12607 & n12634 ;
  assign n12636 = n12535 & n12541 ;
  assign n12637 = n12535 & n12540 ;
  assign n12638 = ( n12502 & n12636 ) | ( n12502 & n12637 ) | ( n12636 & n12637 ) ;
  assign n12639 = n12545 & ~n12638 ;
  assign n12640 = n12604 & n12639 ;
  assign n12641 = n12535 & n12599 ;
  assign n12642 = ~n12550 & n12602 ;
  assign n12643 = n12641 & n12642 ;
  assign n12644 = ( n12502 & n12540 ) | ( n12502 & n12541 ) | ( n12540 & n12541 ) ;
  assign n12645 = n12552 & n12644 ;
  assign n12646 = n12545 & n12645 ;
  assign n12647 = n12643 & n12646 ;
  assign n12648 = n12640 | n12647 ;
  assign n12649 = ~n12545 & n12638 ;
  assign n12650 = ( ~n12604 & n12638 ) | ( ~n12604 & n12649 ) | ( n12638 & n12649 ) ;
  assign n12651 = n12648 | n12650 ;
  assign n12652 = n12635 | n12651 ;
  assign n12653 = n12633 & ~n12634 ;
  assign n12654 = n12611 | n12632 ;
  assign n12655 = ~n12633 & n12654 ;
  assign n12656 = ~n12629 & n12631 ;
  assign n12657 = n12655 & n12656 ;
  assign n12658 = ~n12587 & n12613 ;
  assign n12659 = ( x1000 & n12481 ) | ( x1000 & ~n12484 ) | ( n12481 & ~n12484 ) ;
  assign n12660 = ( ~n12481 & n12484 ) | ( ~n12481 & n12659 ) | ( n12484 & n12659 ) ;
  assign n12661 = ( ~x1000 & n12659 ) | ( ~x1000 & n12660 ) | ( n12659 & n12660 ) ;
  assign n12662 = n12618 & n12661 ;
  assign n12663 = ~n12580 & n12661 ;
  assign n12664 = ( ~n12619 & n12662 ) | ( ~n12619 & n12663 ) | ( n12662 & n12663 ) ;
  assign n12665 = n12620 | n12664 ;
  assign n12666 = ( n12617 & n12664 ) | ( n12617 & n12665 ) | ( n12664 & n12665 ) ;
  assign n12667 = n12621 & n12666 ;
  assign n12668 = ~n12658 & n12667 ;
  assign n12669 = ( ~n12623 & n12658 ) | ( ~n12623 & n12668 ) | ( n12658 & n12668 ) ;
  assign n12670 = ( n12623 & n12625 ) | ( n12623 & n12669 ) | ( n12625 & n12669 ) ;
  assign n12671 = n12628 & n12670 ;
  assign n12672 = n12611 & ~n12632 ;
  assign n12673 = ( n12611 & n12671 ) | ( n12611 & n12672 ) | ( n12671 & n12672 ) ;
  assign n12674 = n12655 | n12673 ;
  assign n12675 = n12671 | n12673 ;
  assign n12676 = ( n12657 & n12674 ) | ( n12657 & n12675 ) | ( n12674 & n12675 ) ;
  assign n12677 = n12653 & n12676 ;
  assign n12678 = n12609 & ~n12634 ;
  assign n12679 = ( n12609 & n12676 ) | ( n12609 & n12678 ) | ( n12676 & n12678 ) ;
  assign n12680 = n12677 | n12679 ;
  assign n12681 = n12634 & ~n12635 ;
  assign n12682 = n12680 & n12681 ;
  assign n12683 = n12635 & ~n12653 ;
  assign n12684 = ( n12635 & ~n12676 ) | ( n12635 & n12683 ) | ( ~n12676 & n12683 ) ;
  assign n12685 = ~n12679 & n12684 ;
  assign n12686 = n12607 | n12635 ;
  assign n12687 = ( n12635 & ~n12685 ) | ( n12635 & n12686 ) | ( ~n12685 & n12686 ) ;
  assign n12688 = n12682 | n12687 ;
  assign n12689 = n12640 | n12650 ;
  assign n12690 = n12647 & n12689 ;
  assign n12691 = ( n12635 & n12647 ) | ( n12635 & n12690 ) | ( n12647 & n12690 ) ;
  assign n12692 = n12652 & ~n12691 ;
  assign n12693 = ( n12635 & n12640 ) | ( n12635 & n12650 ) | ( n12640 & n12650 ) ;
  assign n12694 = n12635 & ~n12693 ;
  assign n12695 = n12692 | n12694 ;
  assign n12696 = ~n12652 & n12695 ;
  assign n12697 = ( n12652 & n12688 ) | ( n12652 & ~n12696 ) | ( n12688 & ~n12696 ) ;
  assign y0 = n12697 ;
endmodule
