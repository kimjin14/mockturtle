module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 ;
  assign n513 = ~x304 & x432 ;
  assign n514 = ~x311 & x439 ;
  assign n515 = ~x310 & x438 ;
  assign n516 = n514 | n515 ;
  assign n517 = ~x309 & x437 ;
  assign n518 = ~x308 & x436 ;
  assign n519 = n517 | n518 ;
  assign n520 = n516 | n519 ;
  assign n521 = ~x305 & x433 ;
  assign n522 = ~x307 & x435 ;
  assign n523 = ~x306 & x434 ;
  assign n524 = n522 | n523 ;
  assign n525 = n521 | n524 ;
  assign n526 = n520 | n525 ;
  assign n527 = n513 | n526 ;
  assign n528 = ~x303 & x431 ;
  assign n529 = ~x302 & x430 ;
  assign n530 = n528 | n529 ;
  assign n531 = ~x300 & x428 ;
  assign n532 = ~x301 & x429 ;
  assign n533 = n531 | n532 ;
  assign n534 = n530 | n533 ;
  assign n535 = ~x299 & x427 ;
  assign n536 = ~x298 & x426 ;
  assign n537 = n535 | n536 ;
  assign n538 = ~x297 & x425 ;
  assign n539 = ~x296 & x424 ;
  assign n540 = n538 | n539 ;
  assign n541 = n537 | n540 ;
  assign n542 = n534 | n541 ;
  assign n543 = ~x288 & x416 ;
  assign n544 = ~x295 & x423 ;
  assign n545 = ~x294 & x422 ;
  assign n546 = n544 | n545 ;
  assign n547 = ~x292 & x420 ;
  assign n548 = ~x293 & x421 ;
  assign n549 = n547 | n548 ;
  assign n550 = n546 | n549 ;
  assign n551 = ~x289 & x417 ;
  assign n552 = ~x291 & x419 ;
  assign n553 = ~x290 & x418 ;
  assign n554 = n552 | n553 ;
  assign n555 = n551 | n554 ;
  assign n556 = n550 | n555 ;
  assign n557 = n543 | n556 ;
  assign n558 = ~x285 & x413 ;
  assign n559 = x284 & ~x412 ;
  assign n560 = ~n558 & n559 ;
  assign n561 = ~x282 & x410 ;
  assign n562 = ( ~x283 & x411 ) | ( ~x283 & n561 ) | ( x411 & n561 ) ;
  assign n563 = ~x284 & x412 ;
  assign n564 = n558 | n563 ;
  assign n565 = ( ~n560 & n562 ) | ( ~n560 & n564 ) | ( n562 & n564 ) ;
  assign n566 = ~x287 & x415 ;
  assign n567 = ~x286 & x414 ;
  assign n568 = n566 | n567 ;
  assign n569 = x285 & ~x413 ;
  assign n570 = ~n567 & n569 ;
  assign n571 = x286 & ~x414 ;
  assign n572 = ~n566 & n571 ;
  assign n573 = ( ~n566 & n570 ) | ( ~n566 & n572 ) | ( n570 & n572 ) ;
  assign n574 = ( n565 & n568 ) | ( n565 & ~n573 ) | ( n568 & ~n573 ) ;
  assign n575 = x287 & ~x415 ;
  assign n576 = ( n557 & n574 ) | ( n557 & ~n575 ) | ( n574 & ~n575 ) ;
  assign n577 = n557 | n576 ;
  assign n578 = x294 & ~x422 ;
  assign n579 = ~n544 & n578 ;
  assign n580 = n550 & ~n579 ;
  assign n581 = x288 & ~x416 ;
  assign n582 = ( x289 & ~x417 ) | ( x289 & n581 ) | ( ~x417 & n581 ) ;
  assign n583 = ( x290 & ~x418 ) | ( x290 & n582 ) | ( ~x418 & n582 ) ;
  assign n584 = ( x291 & ~x419 ) | ( x291 & n583 ) | ( ~x419 & n583 ) ;
  assign n585 = ( n579 & ~n580 ) | ( n579 & n584 ) | ( ~n580 & n584 ) ;
  assign n586 = x292 & ~x420 ;
  assign n587 = ( x293 & ~x421 ) | ( x293 & n586 ) | ( ~x421 & n586 ) ;
  assign n588 = ~n545 & n587 ;
  assign n589 = ( x295 & ~x423 ) | ( x295 & n588 ) | ( ~x423 & n588 ) ;
  assign n590 = n585 | n589 ;
  assign n591 = ~n542 & n590 ;
  assign n592 = ( n542 & n577 ) | ( n542 & ~n591 ) | ( n577 & ~n591 ) ;
  assign n593 = x296 & ~x424 ;
  assign n594 = ( x297 & ~x425 ) | ( x297 & n593 ) | ( ~x425 & n593 ) ;
  assign n595 = ( x298 & ~x426 ) | ( x298 & n594 ) | ( ~x426 & n594 ) ;
  assign n596 = ( x299 & ~x427 ) | ( x299 & n595 ) | ( ~x427 & n595 ) ;
  assign n597 = ~n534 & n596 ;
  assign n598 = x303 & ~x431 ;
  assign n599 = x302 & ~x430 ;
  assign n600 = ~n528 & n599 ;
  assign n601 = x300 & ~x428 ;
  assign n602 = ( x301 & ~x429 ) | ( x301 & n601 ) | ( ~x429 & n601 ) ;
  assign n603 = ~n530 & n602 ;
  assign n604 = n600 | n603 ;
  assign n605 = n598 | n604 ;
  assign n606 = n597 | n605 ;
  assign n607 = ~n527 & n606 ;
  assign n608 = ( n527 & n592 ) | ( n527 & ~n607 ) | ( n592 & ~n607 ) ;
  assign n609 = ~x327 & x455 ;
  assign n610 = x326 & ~x454 ;
  assign n611 = ~n609 & n610 ;
  assign n612 = ~x326 & x454 ;
  assign n613 = n609 | n612 ;
  assign n614 = ~x325 & x453 ;
  assign n615 = ~x324 & x452 ;
  assign n616 = n614 | n615 ;
  assign n617 = n613 | n616 ;
  assign n618 = ~x323 & x451 ;
  assign n619 = ~x322 & x450 ;
  assign n620 = n618 | n619 ;
  assign n621 = ~x321 & x449 ;
  assign n622 = ~x320 & x448 ;
  assign n623 = n621 | n622 ;
  assign n624 = n620 | n623 ;
  assign n625 = n617 | n624 ;
  assign n626 = x320 & ~x448 ;
  assign n627 = ( x321 & ~x449 ) | ( x321 & n626 ) | ( ~x449 & n626 ) ;
  assign n628 = ( x322 & ~x450 ) | ( x322 & n627 ) | ( ~x450 & n627 ) ;
  assign n629 = ( x323 & ~x451 ) | ( x323 & n628 ) | ( ~x451 & n628 ) ;
  assign n630 = ( n617 & n625 ) | ( n617 & ~n629 ) | ( n625 & ~n629 ) ;
  assign n631 = ~n611 & n630 ;
  assign n632 = ~x335 & x463 ;
  assign n633 = ~x334 & x462 ;
  assign n634 = n632 | n633 ;
  assign n635 = ~x333 & x461 ;
  assign n636 = ~x332 & x460 ;
  assign n637 = n635 | n636 ;
  assign n638 = n634 | n637 ;
  assign n639 = ~x331 & x459 ;
  assign n640 = ~x330 & x458 ;
  assign n641 = n639 | n640 ;
  assign n642 = ~x329 & x457 ;
  assign n643 = ~x328 & x456 ;
  assign n644 = n642 | n643 ;
  assign n645 = n641 | n644 ;
  assign n646 = x324 & ~x452 ;
  assign n647 = ( x325 & ~x453 ) | ( x325 & n646 ) | ( ~x453 & n646 ) ;
  assign n648 = ~n612 & n647 ;
  assign n649 = ( x327 & ~x455 ) | ( x327 & n648 ) | ( ~x455 & n648 ) ;
  assign n650 = ~n645 & n649 ;
  assign n651 = x328 & ~x456 ;
  assign n652 = ( x329 & ~x457 ) | ( x329 & n651 ) | ( ~x457 & n651 ) ;
  assign n653 = ( x330 & ~x458 ) | ( x330 & n652 ) | ( ~x458 & n652 ) ;
  assign n654 = ( x331 & ~x459 ) | ( x331 & n653 ) | ( ~x459 & n653 ) ;
  assign n655 = ~n638 & n654 ;
  assign n656 = ( ~n638 & n650 ) | ( ~n638 & n655 ) | ( n650 & n655 ) ;
  assign n657 = n638 | n645 ;
  assign n658 = ( n638 & ~n654 ) | ( n638 & n657 ) | ( ~n654 & n657 ) ;
  assign n659 = ( n631 & ~n656 ) | ( n631 & n658 ) | ( ~n656 & n658 ) ;
  assign n660 = ~n611 & n617 ;
  assign n661 = ( n611 & n629 ) | ( n611 & ~n660 ) | ( n629 & ~n660 ) ;
  assign n662 = ( n656 & ~n658 ) | ( n656 & n661 ) | ( ~n658 & n661 ) ;
  assign n663 = ~x319 & x447 ;
  assign n664 = ~x318 & x446 ;
  assign n665 = n663 | n664 ;
  assign n666 = x316 & ~x444 ;
  assign n667 = ( x317 & ~x445 ) | ( x317 & n666 ) | ( ~x445 & n666 ) ;
  assign n668 = ~n665 & n667 ;
  assign n669 = x318 & ~x446 ;
  assign n670 = ~n663 & n669 ;
  assign n671 = n668 | n670 ;
  assign n672 = ~x317 & x445 ;
  assign n673 = ~x316 & x444 ;
  assign n674 = n672 | n673 ;
  assign n675 = n665 | n674 ;
  assign n676 = ~x315 & x443 ;
  assign n677 = ~x314 & x442 ;
  assign n678 = n676 | n677 ;
  assign n679 = ~x313 & x441 ;
  assign n680 = ~x312 & x440 ;
  assign n681 = n679 | n680 ;
  assign n682 = n678 | n681 ;
  assign n683 = n675 | n682 ;
  assign n684 = x319 & ~x447 ;
  assign n685 = x312 & ~x440 ;
  assign n686 = ( x313 & ~x441 ) | ( x313 & n685 ) | ( ~x441 & n685 ) ;
  assign n687 = ( x314 & ~x442 ) | ( x314 & n686 ) | ( ~x442 & n686 ) ;
  assign n688 = ( x315 & ~x443 ) | ( x315 & n687 ) | ( ~x443 & n687 ) ;
  assign n689 = ~n675 & n688 ;
  assign n690 = n684 | n689 ;
  assign n691 = ( n671 & n683 ) | ( n671 & ~n690 ) | ( n683 & ~n690 ) ;
  assign n692 = ~n671 & n691 ;
  assign n693 = ( n659 & ~n662 ) | ( n659 & n692 ) | ( ~n662 & n692 ) ;
  assign n694 = ~x343 & x471 ;
  assign n695 = ~x342 & x470 ;
  assign n696 = n694 | n695 ;
  assign n697 = ~x341 & x469 ;
  assign n698 = ~x340 & x468 ;
  assign n699 = n697 | n698 ;
  assign n700 = n696 | n699 ;
  assign n701 = ~x336 & x464 ;
  assign n702 = ~x339 & x467 ;
  assign n703 = ~x338 & x466 ;
  assign n704 = n702 | n703 ;
  assign n705 = ~x337 & x465 ;
  assign n706 = x335 & ~x463 ;
  assign n707 = ~n705 & n706 ;
  assign n708 = ~n704 & n707 ;
  assign n709 = ~n701 & n708 ;
  assign n710 = n701 | n705 ;
  assign n711 = n704 | n710 ;
  assign n712 = x332 & ~x460 ;
  assign n713 = ( x333 & ~x461 ) | ( x333 & n712 ) | ( ~x461 & n712 ) ;
  assign n714 = ( x334 & ~x462 ) | ( x334 & n713 ) | ( ~x462 & n713 ) ;
  assign n715 = ~n632 & n714 ;
  assign n716 = ( n709 & ~n711 ) | ( n709 & n715 ) | ( ~n711 & n715 ) ;
  assign n717 = x336 & ~x464 ;
  assign n718 = ( x337 & ~x465 ) | ( x337 & n717 ) | ( ~x465 & n717 ) ;
  assign n719 = ( x338 & ~x466 ) | ( x338 & n718 ) | ( ~x466 & n718 ) ;
  assign n720 = ( x339 & ~x467 ) | ( x339 & n719 ) | ( ~x467 & n719 ) ;
  assign n721 = ~n700 & n720 ;
  assign n722 = ( ~n700 & n716 ) | ( ~n700 & n721 ) | ( n716 & n721 ) ;
  assign n723 = x343 & ~x471 ;
  assign n724 = x340 & ~x468 ;
  assign n725 = ( x341 & ~x469 ) | ( x341 & n724 ) | ( ~x469 & n724 ) ;
  assign n726 = ( x342 & ~x470 ) | ( x342 & n725 ) | ( ~x470 & n725 ) ;
  assign n727 = ~n694 & n726 ;
  assign n728 = n723 | n727 ;
  assign n729 = n722 | n728 ;
  assign n730 = ~x351 & x479 ;
  assign n731 = x350 & ~x478 ;
  assign n732 = ~n730 & n731 ;
  assign n733 = ~x350 & x478 ;
  assign n734 = n730 | n733 ;
  assign n735 = ~x349 & x477 ;
  assign n736 = ~x348 & x476 ;
  assign n737 = n735 | n736 ;
  assign n738 = n734 | n737 ;
  assign n739 = ~x347 & x475 ;
  assign n740 = ~x346 & x474 ;
  assign n741 = n739 | n740 ;
  assign n742 = ~x345 & x473 ;
  assign n743 = ~x344 & x472 ;
  assign n744 = n742 | n743 ;
  assign n745 = n741 | n744 ;
  assign n746 = n738 | n745 ;
  assign n747 = x344 & ~x472 ;
  assign n748 = ( x345 & ~x473 ) | ( x345 & n747 ) | ( ~x473 & n747 ) ;
  assign n749 = ( x346 & ~x474 ) | ( x346 & n748 ) | ( ~x474 & n748 ) ;
  assign n750 = ( x347 & ~x475 ) | ( x347 & n749 ) | ( ~x475 & n749 ) ;
  assign n751 = ( n738 & n746 ) | ( n738 & ~n750 ) | ( n746 & ~n750 ) ;
  assign n752 = ~n732 & n751 ;
  assign n753 = ~x355 & x483 ;
  assign n754 = ~x354 & x482 ;
  assign n755 = n753 | n754 ;
  assign n756 = ~x352 & x480 ;
  assign n757 = ~x353 & x481 ;
  assign n758 = n756 | n757 ;
  assign n759 = n755 | n758 ;
  assign n760 = x348 & ~x476 ;
  assign n761 = ( x349 & ~x477 ) | ( x349 & n760 ) | ( ~x477 & n760 ) ;
  assign n762 = ~n733 & n761 ;
  assign n763 = ( x351 & ~x479 ) | ( x351 & n762 ) | ( ~x479 & n762 ) ;
  assign n764 = ~n759 & n763 ;
  assign n765 = ( n752 & n759 ) | ( n752 & ~n764 ) | ( n759 & ~n764 ) ;
  assign n766 = ~n732 & n738 ;
  assign n767 = ( n732 & n750 ) | ( n732 & ~n766 ) | ( n750 & ~n766 ) ;
  assign n768 = ( ~n759 & n764 ) | ( ~n759 & n767 ) | ( n764 & n767 ) ;
  assign n769 = ( n729 & ~n765 ) | ( n729 & n768 ) | ( ~n765 & n768 ) ;
  assign n770 = n700 | n711 ;
  assign n771 = ( n700 & ~n720 ) | ( n700 & n770 ) | ( ~n720 & n770 ) ;
  assign n772 = ~n727 & n771 ;
  assign n773 = n723 & ~n745 ;
  assign n774 = n750 | n773 ;
  assign n775 = ~n738 & n774 ;
  assign n776 = ( n751 & n772 ) | ( n751 & ~n775 ) | ( n772 & ~n775 ) ;
  assign n777 = ( n732 & ~n734 ) | ( n732 & n761 ) | ( ~n734 & n761 ) ;
  assign n778 = ( ~n759 & n764 ) | ( ~n759 & n777 ) | ( n764 & n777 ) ;
  assign n779 = ( n759 & n776 ) | ( n759 & ~n778 ) | ( n776 & ~n778 ) ;
  assign n780 = ( n693 & ~n769 ) | ( n693 & n779 ) | ( ~n769 & n779 ) ;
  assign n781 = x304 & ~x432 ;
  assign n782 = ( x305 & ~x433 ) | ( x305 & n781 ) | ( ~x433 & n781 ) ;
  assign n783 = ( x306 & ~x434 ) | ( x306 & n782 ) | ( ~x434 & n782 ) ;
  assign n784 = ( x307 & ~x435 ) | ( x307 & n783 ) | ( ~x435 & n783 ) ;
  assign n785 = ~n520 & n784 ;
  assign n786 = x308 & ~x436 ;
  assign n787 = ( x309 & ~x437 ) | ( x309 & n786 ) | ( ~x437 & n786 ) ;
  assign n788 = ( x310 & ~x438 ) | ( x310 & n787 ) | ( ~x438 & n787 ) ;
  assign n789 = ( x311 & ~x439 ) | ( x311 & n788 ) | ( ~x439 & n788 ) ;
  assign n790 = ~n683 & n789 ;
  assign n791 = ( ~n683 & n785 ) | ( ~n683 & n790 ) | ( n785 & n790 ) ;
  assign n792 = n671 | n689 ;
  assign n793 = n791 | n792 ;
  assign n794 = ~n624 & n684 ;
  assign n795 = n629 | n794 ;
  assign n796 = ( n611 & ~n660 ) | ( n611 & n795 ) | ( ~n660 & n795 ) ;
  assign n797 = ( n656 & ~n658 ) | ( n656 & n796 ) | ( ~n658 & n796 ) ;
  assign n798 = ( ~n659 & n793 ) | ( ~n659 & n797 ) | ( n793 & n797 ) ;
  assign n799 = ( n769 & ~n779 ) | ( n769 & n798 ) | ( ~n779 & n798 ) ;
  assign n800 = ( n608 & n780 ) | ( n608 & ~n799 ) | ( n780 & ~n799 ) ;
  assign n801 = x383 & ~x511 ;
  assign n802 = x380 & ~x508 ;
  assign n803 = ( x381 & ~x509 ) | ( x381 & n802 ) | ( ~x509 & n802 ) ;
  assign n804 = ( x382 & ~x510 ) | ( x382 & n803 ) | ( ~x510 & n803 ) ;
  assign n805 = ~n801 & n804 ;
  assign n806 = ~x382 & x510 ;
  assign n807 = ~x381 & x509 ;
  assign n808 = n806 | n807 ;
  assign n809 = ~x380 & x508 ;
  assign n810 = n808 | n809 ;
  assign n811 = ( x383 & ~x511 ) | ( x383 & n810 ) | ( ~x511 & n810 ) ;
  assign n812 = ~n805 & n811 ;
  assign n813 = x384 & n812 ;
  assign n814 = ~x383 & x511 ;
  assign n815 = n805 | n814 ;
  assign n816 = x384 & ~n815 ;
  assign n817 = ~x379 & x507 ;
  assign n818 = ~x378 & x506 ;
  assign n819 = n817 | n818 ;
  assign n820 = ~x377 & x505 ;
  assign n821 = ~x376 & x504 ;
  assign n822 = n820 | n821 ;
  assign n823 = n819 | n822 ;
  assign n824 = x376 & ~x504 ;
  assign n825 = ( x377 & ~x505 ) | ( x377 & n824 ) | ( ~x505 & n824 ) ;
  assign n826 = ( x378 & ~x506 ) | ( x378 & n825 ) | ( ~x506 & n825 ) ;
  assign n827 = ( x379 & ~x507 ) | ( x379 & n826 ) | ( ~x507 & n826 ) ;
  assign n828 = n823 & ~n827 ;
  assign n829 = ~x375 & x503 ;
  assign n830 = x374 & ~x502 ;
  assign n831 = ~n829 & n830 ;
  assign n832 = ~x374 & x502 ;
  assign n833 = n829 | n832 ;
  assign n834 = ~x373 & x501 ;
  assign n835 = ~x372 & x500 ;
  assign n836 = n834 | n835 ;
  assign n837 = n833 | n836 ;
  assign n838 = ~x369 & x497 ;
  assign n839 = ~x371 & x499 ;
  assign n840 = ~x370 & x498 ;
  assign n841 = n839 | n840 ;
  assign n842 = ~x368 & x496 ;
  assign n843 = n841 | n842 ;
  assign n844 = n838 | n843 ;
  assign n845 = n837 | n844 ;
  assign n846 = x368 & ~x496 ;
  assign n847 = ( x369 & ~x497 ) | ( x369 & n846 ) | ( ~x497 & n846 ) ;
  assign n848 = ( x370 & ~x498 ) | ( x370 & n847 ) | ( ~x498 & n847 ) ;
  assign n849 = ( x371 & ~x499 ) | ( x371 & n848 ) | ( ~x499 & n848 ) ;
  assign n850 = ( n837 & n845 ) | ( n837 & ~n849 ) | ( n845 & ~n849 ) ;
  assign n851 = ~n831 & n850 ;
  assign n852 = x375 & ~x503 ;
  assign n853 = x372 & ~x500 ;
  assign n854 = ( x373 & ~x501 ) | ( x373 & n853 ) | ( ~x501 & n853 ) ;
  assign n855 = ~n833 & n854 ;
  assign n856 = n852 | n855 ;
  assign n857 = ~n823 & n856 ;
  assign n858 = n827 | n857 ;
  assign n859 = ( n828 & n851 ) | ( n828 & ~n858 ) | ( n851 & ~n858 ) ;
  assign n860 = ~n831 & n837 ;
  assign n861 = ( n831 & n849 ) | ( n831 & ~n860 ) | ( n849 & ~n860 ) ;
  assign n862 = ( ~n828 & n858 ) | ( ~n828 & n861 ) | ( n858 & n861 ) ;
  assign n863 = x367 & ~x495 ;
  assign n864 = ~x367 & x495 ;
  assign n865 = ~x366 & x494 ;
  assign n866 = n864 | n865 ;
  assign n867 = x364 & ~x492 ;
  assign n868 = ( x365 & ~x493 ) | ( x365 & n867 ) | ( ~x493 & n867 ) ;
  assign n869 = ~n866 & n868 ;
  assign n870 = x366 & ~x494 ;
  assign n871 = ~n864 & n870 ;
  assign n872 = n869 | n871 ;
  assign n873 = ~x359 & x487 ;
  assign n874 = ~x358 & x486 ;
  assign n875 = n873 | n874 ;
  assign n876 = x356 & ~x484 ;
  assign n877 = ( x357 & ~x485 ) | ( x357 & n876 ) | ( ~x485 & n876 ) ;
  assign n878 = ~n875 & n877 ;
  assign n879 = ~x357 & x485 ;
  assign n880 = ~x356 & x484 ;
  assign n881 = n879 | n880 ;
  assign n882 = n875 | n881 ;
  assign n883 = x358 & ~x486 ;
  assign n884 = ~n873 & n883 ;
  assign n885 = n882 & ~n884 ;
  assign n886 = ~n878 & n885 ;
  assign n887 = ~x363 & x491 ;
  assign n888 = ~x362 & x490 ;
  assign n889 = n887 | n888 ;
  assign n890 = ~x361 & x489 ;
  assign n891 = ~x360 & x488 ;
  assign n892 = n890 | n891 ;
  assign n893 = n889 | n892 ;
  assign n894 = x360 & ~x488 ;
  assign n895 = ( x361 & ~x489 ) | ( x361 & n894 ) | ( ~x489 & n894 ) ;
  assign n896 = ( x362 & ~x490 ) | ( x362 & n895 ) | ( ~x490 & n895 ) ;
  assign n897 = ( x363 & ~x491 ) | ( x363 & n896 ) | ( ~x491 & n896 ) ;
  assign n898 = n893 & ~n897 ;
  assign n899 = x359 & ~x487 ;
  assign n900 = ( n897 & ~n898 ) | ( n897 & n899 ) | ( ~n898 & n899 ) ;
  assign n901 = ( n886 & n898 ) | ( n886 & ~n900 ) | ( n898 & ~n900 ) ;
  assign n902 = ~x365 & x493 ;
  assign n903 = ~x364 & x492 ;
  assign n904 = n902 | n903 ;
  assign n905 = n866 | n904 ;
  assign n906 = ( ~n872 & n901 ) | ( ~n872 & n905 ) | ( n901 & n905 ) ;
  assign n907 = ~n872 & n906 ;
  assign n908 = ~n863 & n907 ;
  assign n909 = ( n859 & ~n862 ) | ( n859 & n908 ) | ( ~n862 & n908 ) ;
  assign n910 = ( n813 & n816 ) | ( n813 & n909 ) | ( n816 & n909 ) ;
  assign n911 = x352 & ~x480 ;
  assign n912 = ( x353 & ~x481 ) | ( x353 & n911 ) | ( ~x481 & n911 ) ;
  assign n913 = ( x354 & ~x482 ) | ( x354 & n912 ) | ( ~x482 & n912 ) ;
  assign n914 = ( x355 & ~x483 ) | ( x355 & n913 ) | ( ~x483 & n913 ) ;
  assign n915 = ( n884 & ~n885 ) | ( n884 & n914 ) | ( ~n885 & n914 ) ;
  assign n916 = n878 | n899 ;
  assign n917 = n915 | n916 ;
  assign n918 = n898 | n905 ;
  assign n919 = n863 | n872 ;
  assign n920 = ~n838 & n919 ;
  assign n921 = ( n838 & n918 ) | ( n838 & ~n920 ) | ( n918 & ~n920 ) ;
  assign n922 = n897 & ~n905 ;
  assign n923 = ( ~n838 & n920 ) | ( ~n838 & n922 ) | ( n920 & n922 ) ;
  assign n924 = ( n917 & ~n921 ) | ( n917 & n923 ) | ( ~n921 & n923 ) ;
  assign n925 = n837 | n843 ;
  assign n926 = n855 | n861 ;
  assign n927 = n925 & ~n926 ;
  assign n928 = ( n828 & ~n858 ) | ( n828 & n927 ) | ( ~n858 & n927 ) ;
  assign n929 = ( n862 & n924 ) | ( n862 & ~n928 ) | ( n924 & ~n928 ) ;
  assign n930 = ( n813 & n816 ) | ( n813 & ~n929 ) | ( n816 & ~n929 ) ;
  assign n931 = ( n800 & n910 ) | ( n800 & n930 ) | ( n910 & n930 ) ;
  assign n932 = x283 & ~x411 ;
  assign n933 = ~n563 & n932 ;
  assign n934 = x282 & ~x410 ;
  assign n935 = ~n562 & n934 ;
  assign n936 = ( ~n563 & n933 ) | ( ~n563 & n935 ) | ( n933 & n935 ) ;
  assign n937 = ( ~n558 & n560 ) | ( ~n558 & n936 ) | ( n560 & n936 ) ;
  assign n938 = n569 | n937 ;
  assign n939 = ( ~n568 & n572 ) | ( ~n568 & n938 ) | ( n572 & n938 ) ;
  assign n940 = n575 | n939 ;
  assign n941 = ~n557 & n940 ;
  assign n942 = n590 | n941 ;
  assign n943 = n542 & ~n604 ;
  assign n944 = ( n604 & n942 ) | ( n604 & ~n943 ) | ( n942 & ~n943 ) ;
  assign n945 = n597 | n944 ;
  assign n946 = ( ~n527 & n598 ) | ( ~n527 & n945 ) | ( n598 & n945 ) ;
  assign n947 = ~n527 & n946 ;
  assign n948 = ( ~n780 & n799 ) | ( ~n780 & n947 ) | ( n799 & n947 ) ;
  assign n949 = ( n910 & n930 ) | ( n910 & ~n948 ) | ( n930 & ~n948 ) ;
  assign n950 = ~x277 & x405 ;
  assign n951 = x276 & ~x404 ;
  assign n952 = ~n950 & n951 ;
  assign n953 = ~x274 & x402 ;
  assign n954 = ( ~x275 & x403 ) | ( ~x275 & n953 ) | ( x403 & n953 ) ;
  assign n955 = ~x276 & x404 ;
  assign n956 = n950 | n955 ;
  assign n957 = ( ~n952 & n954 ) | ( ~n952 & n956 ) | ( n954 & n956 ) ;
  assign n958 = ~x279 & x407 ;
  assign n959 = ~x278 & x406 ;
  assign n960 = x277 & ~x405 ;
  assign n961 = ~n959 & n960 ;
  assign n962 = x278 & ~x406 ;
  assign n963 = ~n958 & n962 ;
  assign n964 = ( ~n958 & n961 ) | ( ~n958 & n963 ) | ( n961 & n963 ) ;
  assign n965 = x279 & ~x407 ;
  assign n966 = x280 & ~x408 ;
  assign n967 = ( ~x408 & n965 ) | ( ~x408 & n966 ) | ( n965 & n966 ) ;
  assign n968 = ( ~x408 & n964 ) | ( ~x408 & n967 ) | ( n964 & n967 ) ;
  assign n969 = n958 | n959 ;
  assign n970 = ~n965 & n969 ;
  assign n971 = ( x408 & ~n966 ) | ( x408 & n970 ) | ( ~n966 & n970 ) ;
  assign n972 = ( n957 & ~n968 ) | ( n957 & n971 ) | ( ~n968 & n971 ) ;
  assign n973 = x275 & ~x403 ;
  assign n974 = ~n955 & n973 ;
  assign n975 = x274 & ~x402 ;
  assign n976 = ~n954 & n975 ;
  assign n977 = ( ~n955 & n974 ) | ( ~n955 & n976 ) | ( n974 & n976 ) ;
  assign n978 = ( ~n950 & n952 ) | ( ~n950 & n977 ) | ( n952 & n977 ) ;
  assign n979 = n960 | n978 ;
  assign n980 = ( ~x408 & n963 ) | ( ~x408 & n967 ) | ( n963 & n967 ) ;
  assign n981 = ( ~n971 & n979 ) | ( ~n971 & n980 ) | ( n979 & n980 ) ;
  assign n982 = ~x269 & x397 ;
  assign n983 = x268 & ~x396 ;
  assign n984 = ~n982 & n983 ;
  assign n985 = ~x266 & x394 ;
  assign n986 = ( ~x267 & x395 ) | ( ~x267 & n985 ) | ( x395 & n985 ) ;
  assign n987 = ~x268 & x396 ;
  assign n988 = n982 | n987 ;
  assign n989 = ( ~n984 & n986 ) | ( ~n984 & n988 ) | ( n986 & n988 ) ;
  assign n990 = x271 & ~x399 ;
  assign n991 = ~x271 & x399 ;
  assign n992 = ~x270 & x398 ;
  assign n993 = x269 & ~x397 ;
  assign n994 = ~n992 & n993 ;
  assign n995 = x270 & ~x398 ;
  assign n996 = ~n991 & n995 ;
  assign n997 = ( ~n991 & n994 ) | ( ~n991 & n996 ) | ( n994 & n996 ) ;
  assign n998 = n990 | n997 ;
  assign n999 = ( ~x271 & x399 ) | ( ~x271 & n992 ) | ( x399 & n992 ) ;
  assign n1000 = ( n989 & ~n998 ) | ( n989 & n999 ) | ( ~n998 & n999 ) ;
  assign n1001 = x272 & ~n1000 ;
  assign n1002 = x272 & ~n999 ;
  assign n1003 = x272 & n990 ;
  assign n1004 = ( x272 & n996 ) | ( x272 & n1003 ) | ( n996 & n1003 ) ;
  assign n1005 = x267 & ~x395 ;
  assign n1006 = ~n987 & n1005 ;
  assign n1007 = x266 & ~x394 ;
  assign n1008 = ~n986 & n1007 ;
  assign n1009 = ( ~n987 & n1006 ) | ( ~n987 & n1008 ) | ( n1006 & n1008 ) ;
  assign n1010 = ( ~n982 & n984 ) | ( ~n982 & n1009 ) | ( n984 & n1009 ) ;
  assign n1011 = n993 | n1010 ;
  assign n1012 = ( n1002 & n1004 ) | ( n1002 & n1011 ) | ( n1004 & n1011 ) ;
  assign n1013 = x263 & ~x391 ;
  assign n1014 = x264 | n1013 ;
  assign n1015 = x262 & ~x390 ;
  assign n1016 = ~x262 & x390 ;
  assign n1017 = ( ~x263 & x391 ) | ( ~x263 & n1016 ) | ( x391 & n1016 ) ;
  assign n1018 = n1015 & ~n1017 ;
  assign n1019 = n1014 | n1018 ;
  assign n1020 = ~x392 & n1019 ;
  assign n1021 = x260 & ~x388 ;
  assign n1022 = x259 & ~x387 ;
  assign n1023 = ( ~x259 & x387 ) | ( ~x259 & n1022 ) | ( x387 & n1022 ) ;
  assign n1024 = ( x388 & ~n1021 ) | ( x388 & n1023 ) | ( ~n1021 & n1023 ) ;
  assign n1025 = ( ~x388 & n1021 ) | ( ~x388 & n1022 ) | ( n1021 & n1022 ) ;
  assign n1026 = x256 & ~x384 ;
  assign n1027 = ( x257 & ~x385 ) | ( x257 & n1026 ) | ( ~x385 & n1026 ) ;
  assign n1028 = ( x258 & ~x386 ) | ( x258 & n1027 ) | ( ~x386 & n1027 ) ;
  assign n1029 = ( ~n1024 & n1025 ) | ( ~n1024 & n1028 ) | ( n1025 & n1028 ) ;
  assign n1030 = ( x259 & ~x387 ) | ( x259 & n1028 ) | ( ~x387 & n1028 ) ;
  assign n1031 = x260 & n1030 ;
  assign n1032 = n1029 | n1031 ;
  assign n1033 = ( x261 & ~x389 ) | ( x261 & n1032 ) | ( ~x389 & n1032 ) ;
  assign n1034 = ( x392 & n1017 ) | ( x392 & ~n1020 ) | ( n1017 & ~n1020 ) ;
  assign n1035 = ( n1020 & n1033 ) | ( n1020 & ~n1034 ) | ( n1033 & ~n1034 ) ;
  assign n1036 = x264 & ~n1017 ;
  assign n1037 = x264 & n1013 ;
  assign n1038 = ( x264 & n1018 ) | ( x264 & n1037 ) | ( n1018 & n1037 ) ;
  assign n1039 = ( n1033 & n1036 ) | ( n1033 & n1038 ) | ( n1036 & n1038 ) ;
  assign n1040 = n1035 | n1039 ;
  assign n1041 = ( x265 & ~x393 ) | ( x265 & n1040 ) | ( ~x393 & n1040 ) ;
  assign n1042 = ( n1001 & n1012 ) | ( n1001 & n1041 ) | ( n1012 & n1041 ) ;
  assign n1043 = x272 & ~x400 ;
  assign n1044 = ( x400 & n1000 ) | ( x400 & ~n1043 ) | ( n1000 & ~n1043 ) ;
  assign n1045 = ( x400 & n999 ) | ( x400 & ~n1043 ) | ( n999 & ~n1043 ) ;
  assign n1046 = ( ~x400 & n990 ) | ( ~x400 & n1043 ) | ( n990 & n1043 ) ;
  assign n1047 = ( ~x400 & n996 ) | ( ~x400 & n1046 ) | ( n996 & n1046 ) ;
  assign n1048 = ( n1011 & ~n1045 ) | ( n1011 & n1047 ) | ( ~n1045 & n1047 ) ;
  assign n1049 = ( n1041 & ~n1044 ) | ( n1041 & n1048 ) | ( ~n1044 & n1048 ) ;
  assign n1050 = n1042 | n1049 ;
  assign n1051 = ( x273 & ~x401 ) | ( x273 & n1050 ) | ( ~x401 & n1050 ) ;
  assign n1052 = ( ~n972 & n981 ) | ( ~n972 & n1051 ) | ( n981 & n1051 ) ;
  assign n1053 = x280 & n965 ;
  assign n1054 = ( x280 & n963 ) | ( x280 & n1053 ) | ( n963 & n1053 ) ;
  assign n1055 = ( x280 & ~n969 ) | ( x280 & n1053 ) | ( ~n969 & n1053 ) ;
  assign n1056 = ( n979 & n1054 ) | ( n979 & n1055 ) | ( n1054 & n1055 ) ;
  assign n1057 = ( x280 & n964 ) | ( x280 & n1053 ) | ( n964 & n1053 ) ;
  assign n1058 = ( ~n957 & n1055 ) | ( ~n957 & n1057 ) | ( n1055 & n1057 ) ;
  assign n1059 = ( n1051 & n1056 ) | ( n1051 & n1058 ) | ( n1056 & n1058 ) ;
  assign n1060 = n1052 | n1059 ;
  assign n1061 = ( x281 & ~x409 ) | ( x281 & n1060 ) | ( ~x409 & n1060 ) ;
  assign n1062 = ( n931 & n949 ) | ( n931 & ~n1061 ) | ( n949 & ~n1061 ) ;
  assign n1063 = x256 & ~n812 ;
  assign n1064 = x256 & n815 ;
  assign n1065 = ( ~n909 & n1063 ) | ( ~n909 & n1064 ) | ( n1063 & n1064 ) ;
  assign n1066 = ( n929 & n1063 ) | ( n929 & n1064 ) | ( n1063 & n1064 ) ;
  assign n1067 = ( ~n800 & n1065 ) | ( ~n800 & n1066 ) | ( n1065 & n1066 ) ;
  assign n1068 = ( n948 & n1065 ) | ( n948 & n1066 ) | ( n1065 & n1066 ) ;
  assign n1069 = ( n1061 & n1067 ) | ( n1061 & n1068 ) | ( n1067 & n1068 ) ;
  assign n1070 = n1062 | n1069 ;
  assign n1071 = ~x48 & x176 ;
  assign n1072 = ~x55 & x183 ;
  assign n1073 = ~x54 & x182 ;
  assign n1074 = n1072 | n1073 ;
  assign n1075 = ~x53 & x181 ;
  assign n1076 = ~x52 & x180 ;
  assign n1077 = n1075 | n1076 ;
  assign n1078 = n1074 | n1077 ;
  assign n1079 = ~x49 & x177 ;
  assign n1080 = ~x51 & x179 ;
  assign n1081 = ~x50 & x178 ;
  assign n1082 = n1080 | n1081 ;
  assign n1083 = n1079 | n1082 ;
  assign n1084 = n1078 | n1083 ;
  assign n1085 = n1071 | n1084 ;
  assign n1086 = ~x47 & x175 ;
  assign n1087 = ~x46 & x174 ;
  assign n1088 = n1086 | n1087 ;
  assign n1089 = ~x44 & x172 ;
  assign n1090 = ~x45 & x173 ;
  assign n1091 = n1089 | n1090 ;
  assign n1092 = n1088 | n1091 ;
  assign n1093 = ~x43 & x171 ;
  assign n1094 = ~x42 & x170 ;
  assign n1095 = n1093 | n1094 ;
  assign n1096 = ~x41 & x169 ;
  assign n1097 = ~x40 & x168 ;
  assign n1098 = n1096 | n1097 ;
  assign n1099 = n1095 | n1098 ;
  assign n1100 = n1092 | n1099 ;
  assign n1101 = ~x32 & x160 ;
  assign n1102 = ~x39 & x167 ;
  assign n1103 = ~x38 & x166 ;
  assign n1104 = n1102 | n1103 ;
  assign n1105 = ~x36 & x164 ;
  assign n1106 = ~x37 & x165 ;
  assign n1107 = n1105 | n1106 ;
  assign n1108 = n1104 | n1107 ;
  assign n1109 = ~x33 & x161 ;
  assign n1110 = ~x35 & x163 ;
  assign n1111 = ~x34 & x162 ;
  assign n1112 = n1110 | n1111 ;
  assign n1113 = n1109 | n1112 ;
  assign n1114 = n1108 | n1113 ;
  assign n1115 = n1101 | n1114 ;
  assign n1116 = ~x29 & x157 ;
  assign n1117 = x28 & ~x156 ;
  assign n1118 = ~n1116 & n1117 ;
  assign n1119 = ~x26 & x154 ;
  assign n1120 = ( ~x27 & x155 ) | ( ~x27 & n1119 ) | ( x155 & n1119 ) ;
  assign n1121 = ~x28 & x156 ;
  assign n1122 = n1116 | n1121 ;
  assign n1123 = ( ~n1118 & n1120 ) | ( ~n1118 & n1122 ) | ( n1120 & n1122 ) ;
  assign n1124 = ~x31 & x159 ;
  assign n1125 = ~x30 & x158 ;
  assign n1126 = n1124 | n1125 ;
  assign n1127 = x29 & ~x157 ;
  assign n1128 = ~n1125 & n1127 ;
  assign n1129 = x30 & ~x158 ;
  assign n1130 = ~n1124 & n1129 ;
  assign n1131 = ( ~n1124 & n1128 ) | ( ~n1124 & n1130 ) | ( n1128 & n1130 ) ;
  assign n1132 = ( n1123 & n1126 ) | ( n1123 & ~n1131 ) | ( n1126 & ~n1131 ) ;
  assign n1133 = x31 & ~x159 ;
  assign n1134 = ( n1115 & n1132 ) | ( n1115 & ~n1133 ) | ( n1132 & ~n1133 ) ;
  assign n1135 = n1115 | n1134 ;
  assign n1136 = x38 & ~x166 ;
  assign n1137 = ~n1102 & n1136 ;
  assign n1138 = n1108 & ~n1137 ;
  assign n1139 = x32 & ~x160 ;
  assign n1140 = ( x33 & ~x161 ) | ( x33 & n1139 ) | ( ~x161 & n1139 ) ;
  assign n1141 = ( x34 & ~x162 ) | ( x34 & n1140 ) | ( ~x162 & n1140 ) ;
  assign n1142 = ( x35 & ~x163 ) | ( x35 & n1141 ) | ( ~x163 & n1141 ) ;
  assign n1143 = ( n1137 & ~n1138 ) | ( n1137 & n1142 ) | ( ~n1138 & n1142 ) ;
  assign n1144 = x36 & ~x164 ;
  assign n1145 = ( x37 & ~x165 ) | ( x37 & n1144 ) | ( ~x165 & n1144 ) ;
  assign n1146 = ~n1103 & n1145 ;
  assign n1147 = ( x39 & ~x167 ) | ( x39 & n1146 ) | ( ~x167 & n1146 ) ;
  assign n1148 = n1143 | n1147 ;
  assign n1149 = ~n1100 & n1148 ;
  assign n1150 = ( n1100 & n1135 ) | ( n1100 & ~n1149 ) | ( n1135 & ~n1149 ) ;
  assign n1151 = x40 & ~x168 ;
  assign n1152 = ( x41 & ~x169 ) | ( x41 & n1151 ) | ( ~x169 & n1151 ) ;
  assign n1153 = ( x42 & ~x170 ) | ( x42 & n1152 ) | ( ~x170 & n1152 ) ;
  assign n1154 = ( x43 & ~x171 ) | ( x43 & n1153 ) | ( ~x171 & n1153 ) ;
  assign n1155 = ~n1092 & n1154 ;
  assign n1156 = x47 & ~x175 ;
  assign n1157 = x46 & ~x174 ;
  assign n1158 = ~n1086 & n1157 ;
  assign n1159 = x44 & ~x172 ;
  assign n1160 = ( x45 & ~x173 ) | ( x45 & n1159 ) | ( ~x173 & n1159 ) ;
  assign n1161 = ~n1088 & n1160 ;
  assign n1162 = n1158 | n1161 ;
  assign n1163 = n1156 | n1162 ;
  assign n1164 = n1155 | n1163 ;
  assign n1165 = ~n1085 & n1164 ;
  assign n1166 = ( n1085 & n1150 ) | ( n1085 & ~n1165 ) | ( n1150 & ~n1165 ) ;
  assign n1167 = ~x71 & x199 ;
  assign n1168 = x70 & ~x198 ;
  assign n1169 = ~n1167 & n1168 ;
  assign n1170 = ~x70 & x198 ;
  assign n1171 = n1167 | n1170 ;
  assign n1172 = ~x69 & x197 ;
  assign n1173 = ~x68 & x196 ;
  assign n1174 = n1172 | n1173 ;
  assign n1175 = n1171 | n1174 ;
  assign n1176 = ~x67 & x195 ;
  assign n1177 = ~x66 & x194 ;
  assign n1178 = n1176 | n1177 ;
  assign n1179 = ~x65 & x193 ;
  assign n1180 = ~x64 & x192 ;
  assign n1181 = n1179 | n1180 ;
  assign n1182 = n1178 | n1181 ;
  assign n1183 = n1175 | n1182 ;
  assign n1184 = x64 & ~x192 ;
  assign n1185 = ( x65 & ~x193 ) | ( x65 & n1184 ) | ( ~x193 & n1184 ) ;
  assign n1186 = ( x66 & ~x194 ) | ( x66 & n1185 ) | ( ~x194 & n1185 ) ;
  assign n1187 = ( x67 & ~x195 ) | ( x67 & n1186 ) | ( ~x195 & n1186 ) ;
  assign n1188 = ( n1175 & n1183 ) | ( n1175 & ~n1187 ) | ( n1183 & ~n1187 ) ;
  assign n1189 = ~n1169 & n1188 ;
  assign n1190 = ~x79 & x207 ;
  assign n1191 = ~x78 & x206 ;
  assign n1192 = n1190 | n1191 ;
  assign n1193 = ~x77 & x205 ;
  assign n1194 = ~x76 & x204 ;
  assign n1195 = n1193 | n1194 ;
  assign n1196 = n1192 | n1195 ;
  assign n1197 = ~x75 & x203 ;
  assign n1198 = ~x74 & x202 ;
  assign n1199 = n1197 | n1198 ;
  assign n1200 = ~x73 & x201 ;
  assign n1201 = ~x72 & x200 ;
  assign n1202 = n1200 | n1201 ;
  assign n1203 = n1199 | n1202 ;
  assign n1204 = x68 & ~x196 ;
  assign n1205 = ( x69 & ~x197 ) | ( x69 & n1204 ) | ( ~x197 & n1204 ) ;
  assign n1206 = ~n1170 & n1205 ;
  assign n1207 = ( x71 & ~x199 ) | ( x71 & n1206 ) | ( ~x199 & n1206 ) ;
  assign n1208 = ~n1203 & n1207 ;
  assign n1209 = x72 & ~x200 ;
  assign n1210 = ( x73 & ~x201 ) | ( x73 & n1209 ) | ( ~x201 & n1209 ) ;
  assign n1211 = ( x74 & ~x202 ) | ( x74 & n1210 ) | ( ~x202 & n1210 ) ;
  assign n1212 = ( x75 & ~x203 ) | ( x75 & n1211 ) | ( ~x203 & n1211 ) ;
  assign n1213 = ~n1196 & n1212 ;
  assign n1214 = ( ~n1196 & n1208 ) | ( ~n1196 & n1213 ) | ( n1208 & n1213 ) ;
  assign n1215 = n1196 | n1203 ;
  assign n1216 = ( n1196 & ~n1212 ) | ( n1196 & n1215 ) | ( ~n1212 & n1215 ) ;
  assign n1217 = ( n1189 & ~n1214 ) | ( n1189 & n1216 ) | ( ~n1214 & n1216 ) ;
  assign n1218 = ~n1169 & n1175 ;
  assign n1219 = ( n1169 & n1187 ) | ( n1169 & ~n1218 ) | ( n1187 & ~n1218 ) ;
  assign n1220 = ( n1214 & ~n1216 ) | ( n1214 & n1219 ) | ( ~n1216 & n1219 ) ;
  assign n1221 = ~x63 & x191 ;
  assign n1222 = ~x62 & x190 ;
  assign n1223 = n1221 | n1222 ;
  assign n1224 = x60 & ~x188 ;
  assign n1225 = ( x61 & ~x189 ) | ( x61 & n1224 ) | ( ~x189 & n1224 ) ;
  assign n1226 = ~n1223 & n1225 ;
  assign n1227 = x62 & ~x190 ;
  assign n1228 = ~n1221 & n1227 ;
  assign n1229 = n1226 | n1228 ;
  assign n1230 = ~x61 & x189 ;
  assign n1231 = ~x60 & x188 ;
  assign n1232 = n1230 | n1231 ;
  assign n1233 = n1223 | n1232 ;
  assign n1234 = ~x59 & x187 ;
  assign n1235 = ~x58 & x186 ;
  assign n1236 = n1234 | n1235 ;
  assign n1237 = ~x57 & x185 ;
  assign n1238 = ~x56 & x184 ;
  assign n1239 = n1237 | n1238 ;
  assign n1240 = n1236 | n1239 ;
  assign n1241 = n1233 | n1240 ;
  assign n1242 = x63 & ~x191 ;
  assign n1243 = x56 & ~x184 ;
  assign n1244 = ( x57 & ~x185 ) | ( x57 & n1243 ) | ( ~x185 & n1243 ) ;
  assign n1245 = ( x58 & ~x186 ) | ( x58 & n1244 ) | ( ~x186 & n1244 ) ;
  assign n1246 = ( x59 & ~x187 ) | ( x59 & n1245 ) | ( ~x187 & n1245 ) ;
  assign n1247 = ~n1233 & n1246 ;
  assign n1248 = n1242 | n1247 ;
  assign n1249 = ( n1229 & n1241 ) | ( n1229 & ~n1248 ) | ( n1241 & ~n1248 ) ;
  assign n1250 = ~n1229 & n1249 ;
  assign n1251 = ( n1217 & ~n1220 ) | ( n1217 & n1250 ) | ( ~n1220 & n1250 ) ;
  assign n1252 = ~x87 & x215 ;
  assign n1253 = ~x86 & x214 ;
  assign n1254 = n1252 | n1253 ;
  assign n1255 = ~x85 & x213 ;
  assign n1256 = ~x84 & x212 ;
  assign n1257 = n1255 | n1256 ;
  assign n1258 = n1254 | n1257 ;
  assign n1259 = ~x80 & x208 ;
  assign n1260 = ~x83 & x211 ;
  assign n1261 = ~x82 & x210 ;
  assign n1262 = n1260 | n1261 ;
  assign n1263 = ~x81 & x209 ;
  assign n1264 = x79 & ~x207 ;
  assign n1265 = ~n1263 & n1264 ;
  assign n1266 = ~n1262 & n1265 ;
  assign n1267 = ~n1259 & n1266 ;
  assign n1268 = n1259 | n1263 ;
  assign n1269 = n1262 | n1268 ;
  assign n1270 = x76 & ~x204 ;
  assign n1271 = ( x77 & ~x205 ) | ( x77 & n1270 ) | ( ~x205 & n1270 ) ;
  assign n1272 = ( x78 & ~x206 ) | ( x78 & n1271 ) | ( ~x206 & n1271 ) ;
  assign n1273 = ~n1190 & n1272 ;
  assign n1274 = ( n1267 & ~n1269 ) | ( n1267 & n1273 ) | ( ~n1269 & n1273 ) ;
  assign n1275 = x80 & ~x208 ;
  assign n1276 = ( x81 & ~x209 ) | ( x81 & n1275 ) | ( ~x209 & n1275 ) ;
  assign n1277 = ( x82 & ~x210 ) | ( x82 & n1276 ) | ( ~x210 & n1276 ) ;
  assign n1278 = ( x83 & ~x211 ) | ( x83 & n1277 ) | ( ~x211 & n1277 ) ;
  assign n1279 = ~n1258 & n1278 ;
  assign n1280 = ( ~n1258 & n1274 ) | ( ~n1258 & n1279 ) | ( n1274 & n1279 ) ;
  assign n1281 = x87 & ~x215 ;
  assign n1282 = x84 & ~x212 ;
  assign n1283 = ( x85 & ~x213 ) | ( x85 & n1282 ) | ( ~x213 & n1282 ) ;
  assign n1284 = ( x86 & ~x214 ) | ( x86 & n1283 ) | ( ~x214 & n1283 ) ;
  assign n1285 = ~n1252 & n1284 ;
  assign n1286 = n1281 | n1285 ;
  assign n1287 = n1280 | n1286 ;
  assign n1288 = ~x95 & x223 ;
  assign n1289 = x94 & ~x222 ;
  assign n1290 = ~n1288 & n1289 ;
  assign n1291 = ~x94 & x222 ;
  assign n1292 = n1288 | n1291 ;
  assign n1293 = ~x93 & x221 ;
  assign n1294 = ~x92 & x220 ;
  assign n1295 = n1293 | n1294 ;
  assign n1296 = n1292 | n1295 ;
  assign n1297 = ~x91 & x219 ;
  assign n1298 = ~x90 & x218 ;
  assign n1299 = n1297 | n1298 ;
  assign n1300 = ~x89 & x217 ;
  assign n1301 = ~x88 & x216 ;
  assign n1302 = n1300 | n1301 ;
  assign n1303 = n1299 | n1302 ;
  assign n1304 = n1296 | n1303 ;
  assign n1305 = x88 & ~x216 ;
  assign n1306 = ( x89 & ~x217 ) | ( x89 & n1305 ) | ( ~x217 & n1305 ) ;
  assign n1307 = ( x90 & ~x218 ) | ( x90 & n1306 ) | ( ~x218 & n1306 ) ;
  assign n1308 = ( x91 & ~x219 ) | ( x91 & n1307 ) | ( ~x219 & n1307 ) ;
  assign n1309 = ( n1296 & n1304 ) | ( n1296 & ~n1308 ) | ( n1304 & ~n1308 ) ;
  assign n1310 = ~n1290 & n1309 ;
  assign n1311 = ~x99 & x227 ;
  assign n1312 = ~x98 & x226 ;
  assign n1313 = n1311 | n1312 ;
  assign n1314 = ~x96 & x224 ;
  assign n1315 = ~x97 & x225 ;
  assign n1316 = n1314 | n1315 ;
  assign n1317 = n1313 | n1316 ;
  assign n1318 = x92 & ~x220 ;
  assign n1319 = ( x93 & ~x221 ) | ( x93 & n1318 ) | ( ~x221 & n1318 ) ;
  assign n1320 = ~n1291 & n1319 ;
  assign n1321 = ( x95 & ~x223 ) | ( x95 & n1320 ) | ( ~x223 & n1320 ) ;
  assign n1322 = ~n1317 & n1321 ;
  assign n1323 = ( n1310 & n1317 ) | ( n1310 & ~n1322 ) | ( n1317 & ~n1322 ) ;
  assign n1324 = ~n1290 & n1296 ;
  assign n1325 = ( n1290 & n1308 ) | ( n1290 & ~n1324 ) | ( n1308 & ~n1324 ) ;
  assign n1326 = ( ~n1317 & n1322 ) | ( ~n1317 & n1325 ) | ( n1322 & n1325 ) ;
  assign n1327 = ( n1287 & ~n1323 ) | ( n1287 & n1326 ) | ( ~n1323 & n1326 ) ;
  assign n1328 = n1258 | n1269 ;
  assign n1329 = ( n1258 & ~n1278 ) | ( n1258 & n1328 ) | ( ~n1278 & n1328 ) ;
  assign n1330 = ~n1285 & n1329 ;
  assign n1331 = n1281 & ~n1303 ;
  assign n1332 = n1308 | n1331 ;
  assign n1333 = ~n1296 & n1332 ;
  assign n1334 = ( n1309 & n1330 ) | ( n1309 & ~n1333 ) | ( n1330 & ~n1333 ) ;
  assign n1335 = ( n1290 & ~n1292 ) | ( n1290 & n1319 ) | ( ~n1292 & n1319 ) ;
  assign n1336 = ( ~n1317 & n1322 ) | ( ~n1317 & n1335 ) | ( n1322 & n1335 ) ;
  assign n1337 = ( n1317 & n1334 ) | ( n1317 & ~n1336 ) | ( n1334 & ~n1336 ) ;
  assign n1338 = ( n1251 & ~n1327 ) | ( n1251 & n1337 ) | ( ~n1327 & n1337 ) ;
  assign n1339 = x48 & ~x176 ;
  assign n1340 = ( x49 & ~x177 ) | ( x49 & n1339 ) | ( ~x177 & n1339 ) ;
  assign n1341 = ( x50 & ~x178 ) | ( x50 & n1340 ) | ( ~x178 & n1340 ) ;
  assign n1342 = ( x51 & ~x179 ) | ( x51 & n1341 ) | ( ~x179 & n1341 ) ;
  assign n1343 = ~n1078 & n1342 ;
  assign n1344 = x52 & ~x180 ;
  assign n1345 = ( x53 & ~x181 ) | ( x53 & n1344 ) | ( ~x181 & n1344 ) ;
  assign n1346 = ( x54 & ~x182 ) | ( x54 & n1345 ) | ( ~x182 & n1345 ) ;
  assign n1347 = ( x55 & ~x183 ) | ( x55 & n1346 ) | ( ~x183 & n1346 ) ;
  assign n1348 = ~n1241 & n1347 ;
  assign n1349 = ( ~n1241 & n1343 ) | ( ~n1241 & n1348 ) | ( n1343 & n1348 ) ;
  assign n1350 = n1229 | n1247 ;
  assign n1351 = n1349 | n1350 ;
  assign n1352 = ~n1182 & n1242 ;
  assign n1353 = n1187 | n1352 ;
  assign n1354 = ( n1169 & ~n1218 ) | ( n1169 & n1353 ) | ( ~n1218 & n1353 ) ;
  assign n1355 = ( n1214 & ~n1216 ) | ( n1214 & n1354 ) | ( ~n1216 & n1354 ) ;
  assign n1356 = ( ~n1217 & n1351 ) | ( ~n1217 & n1355 ) | ( n1351 & n1355 ) ;
  assign n1357 = ( n1327 & ~n1337 ) | ( n1327 & n1356 ) | ( ~n1337 & n1356 ) ;
  assign n1358 = ( n1166 & n1338 ) | ( n1166 & ~n1357 ) | ( n1338 & ~n1357 ) ;
  assign n1359 = x127 & ~x255 ;
  assign n1360 = x124 & ~x252 ;
  assign n1361 = ( x125 & ~x253 ) | ( x125 & n1360 ) | ( ~x253 & n1360 ) ;
  assign n1362 = ( x126 & ~x254 ) | ( x126 & n1361 ) | ( ~x254 & n1361 ) ;
  assign n1363 = ~n1359 & n1362 ;
  assign n1364 = ~x126 & x254 ;
  assign n1365 = ~x125 & x253 ;
  assign n1366 = n1364 | n1365 ;
  assign n1367 = ~x124 & x252 ;
  assign n1368 = n1366 | n1367 ;
  assign n1369 = ( x127 & ~x255 ) | ( x127 & n1368 ) | ( ~x255 & n1368 ) ;
  assign n1370 = ~n1363 & n1369 ;
  assign n1371 = x239 & n1370 ;
  assign n1372 = ~x127 & x255 ;
  assign n1373 = n1363 | n1372 ;
  assign n1374 = x239 & ~n1373 ;
  assign n1375 = ~x123 & x251 ;
  assign n1376 = ~x122 & x250 ;
  assign n1377 = n1375 | n1376 ;
  assign n1378 = ~x121 & x249 ;
  assign n1379 = ~x120 & x248 ;
  assign n1380 = n1378 | n1379 ;
  assign n1381 = n1377 | n1380 ;
  assign n1382 = x120 & ~x248 ;
  assign n1383 = ( x121 & ~x249 ) | ( x121 & n1382 ) | ( ~x249 & n1382 ) ;
  assign n1384 = ( x122 & ~x250 ) | ( x122 & n1383 ) | ( ~x250 & n1383 ) ;
  assign n1385 = ( x123 & ~x251 ) | ( x123 & n1384 ) | ( ~x251 & n1384 ) ;
  assign n1386 = n1381 & ~n1385 ;
  assign n1387 = ~x119 & x247 ;
  assign n1388 = x118 & ~x246 ;
  assign n1389 = ~n1387 & n1388 ;
  assign n1390 = ~x118 & x246 ;
  assign n1391 = n1387 | n1390 ;
  assign n1392 = ~x117 & x245 ;
  assign n1393 = ~x116 & x244 ;
  assign n1394 = n1392 | n1393 ;
  assign n1395 = n1391 | n1394 ;
  assign n1396 = ~x113 & x241 ;
  assign n1397 = ~x115 & x243 ;
  assign n1398 = ~x114 & x242 ;
  assign n1399 = n1397 | n1398 ;
  assign n1400 = ~x112 & x240 ;
  assign n1401 = n1399 | n1400 ;
  assign n1402 = n1396 | n1401 ;
  assign n1403 = n1395 | n1402 ;
  assign n1404 = x112 & ~x240 ;
  assign n1405 = ( x113 & ~x241 ) | ( x113 & n1404 ) | ( ~x241 & n1404 ) ;
  assign n1406 = ( x114 & ~x242 ) | ( x114 & n1405 ) | ( ~x242 & n1405 ) ;
  assign n1407 = ( x115 & ~x243 ) | ( x115 & n1406 ) | ( ~x243 & n1406 ) ;
  assign n1408 = ( n1395 & n1403 ) | ( n1395 & ~n1407 ) | ( n1403 & ~n1407 ) ;
  assign n1409 = ~n1389 & n1408 ;
  assign n1410 = x119 & ~x247 ;
  assign n1411 = x116 & ~x244 ;
  assign n1412 = ( x117 & ~x245 ) | ( x117 & n1411 ) | ( ~x245 & n1411 ) ;
  assign n1413 = ~n1391 & n1412 ;
  assign n1414 = n1410 | n1413 ;
  assign n1415 = ~n1381 & n1414 ;
  assign n1416 = n1385 | n1415 ;
  assign n1417 = ( n1386 & n1409 ) | ( n1386 & ~n1416 ) | ( n1409 & ~n1416 ) ;
  assign n1418 = ~n1389 & n1395 ;
  assign n1419 = ( n1389 & n1407 ) | ( n1389 & ~n1418 ) | ( n1407 & ~n1418 ) ;
  assign n1420 = ( ~n1386 & n1416 ) | ( ~n1386 & n1419 ) | ( n1416 & n1419 ) ;
  assign n1421 = x111 & ~x239 ;
  assign n1422 = ~x111 & x239 ;
  assign n1423 = ~x110 & x238 ;
  assign n1424 = n1422 | n1423 ;
  assign n1425 = x108 & ~x236 ;
  assign n1426 = ( x109 & ~x237 ) | ( x109 & n1425 ) | ( ~x237 & n1425 ) ;
  assign n1427 = ~n1424 & n1426 ;
  assign n1428 = x110 & ~x238 ;
  assign n1429 = ~n1422 & n1428 ;
  assign n1430 = n1427 | n1429 ;
  assign n1431 = ~x103 & x231 ;
  assign n1432 = ~x102 & x230 ;
  assign n1433 = n1431 | n1432 ;
  assign n1434 = x100 & ~x228 ;
  assign n1435 = ( x101 & ~x229 ) | ( x101 & n1434 ) | ( ~x229 & n1434 ) ;
  assign n1436 = ~n1433 & n1435 ;
  assign n1437 = ~x101 & x229 ;
  assign n1438 = ~x100 & x228 ;
  assign n1439 = n1437 | n1438 ;
  assign n1440 = n1433 | n1439 ;
  assign n1441 = x102 & ~x230 ;
  assign n1442 = ~n1431 & n1441 ;
  assign n1443 = n1440 & ~n1442 ;
  assign n1444 = ~n1436 & n1443 ;
  assign n1445 = ~x107 & x235 ;
  assign n1446 = ~x106 & x234 ;
  assign n1447 = n1445 | n1446 ;
  assign n1448 = ~x105 & x233 ;
  assign n1449 = ~x104 & x232 ;
  assign n1450 = n1448 | n1449 ;
  assign n1451 = n1447 | n1450 ;
  assign n1452 = x104 & ~x232 ;
  assign n1453 = ( x105 & ~x233 ) | ( x105 & n1452 ) | ( ~x233 & n1452 ) ;
  assign n1454 = ( x106 & ~x234 ) | ( x106 & n1453 ) | ( ~x234 & n1453 ) ;
  assign n1455 = ( x107 & ~x235 ) | ( x107 & n1454 ) | ( ~x235 & n1454 ) ;
  assign n1456 = n1451 & ~n1455 ;
  assign n1457 = x103 & ~x231 ;
  assign n1458 = ( n1455 & ~n1456 ) | ( n1455 & n1457 ) | ( ~n1456 & n1457 ) ;
  assign n1459 = ( n1444 & n1456 ) | ( n1444 & ~n1458 ) | ( n1456 & ~n1458 ) ;
  assign n1460 = ~x109 & x237 ;
  assign n1461 = ~x108 & x236 ;
  assign n1462 = n1460 | n1461 ;
  assign n1463 = n1424 | n1462 ;
  assign n1464 = ( ~n1430 & n1459 ) | ( ~n1430 & n1463 ) | ( n1459 & n1463 ) ;
  assign n1465 = ~n1430 & n1464 ;
  assign n1466 = ~n1421 & n1465 ;
  assign n1467 = ( n1417 & ~n1420 ) | ( n1417 & n1466 ) | ( ~n1420 & n1466 ) ;
  assign n1468 = ( n1371 & n1374 ) | ( n1371 & n1467 ) | ( n1374 & n1467 ) ;
  assign n1469 = x96 & ~x224 ;
  assign n1470 = ( x97 & ~x225 ) | ( x97 & n1469 ) | ( ~x225 & n1469 ) ;
  assign n1471 = ( x98 & ~x226 ) | ( x98 & n1470 ) | ( ~x226 & n1470 ) ;
  assign n1472 = ( x99 & ~x227 ) | ( x99 & n1471 ) | ( ~x227 & n1471 ) ;
  assign n1473 = ( n1442 & ~n1443 ) | ( n1442 & n1472 ) | ( ~n1443 & n1472 ) ;
  assign n1474 = n1436 | n1457 ;
  assign n1475 = n1473 | n1474 ;
  assign n1476 = n1456 | n1463 ;
  assign n1477 = n1421 | n1430 ;
  assign n1478 = ~n1396 & n1477 ;
  assign n1479 = ( n1396 & n1476 ) | ( n1396 & ~n1478 ) | ( n1476 & ~n1478 ) ;
  assign n1480 = n1455 & ~n1463 ;
  assign n1481 = ( ~n1396 & n1478 ) | ( ~n1396 & n1480 ) | ( n1478 & n1480 ) ;
  assign n1482 = ( n1475 & ~n1479 ) | ( n1475 & n1481 ) | ( ~n1479 & n1481 ) ;
  assign n1483 = n1395 | n1401 ;
  assign n1484 = n1413 | n1419 ;
  assign n1485 = n1483 & ~n1484 ;
  assign n1486 = ( n1386 & ~n1416 ) | ( n1386 & n1485 ) | ( ~n1416 & n1485 ) ;
  assign n1487 = ( n1420 & n1482 ) | ( n1420 & ~n1486 ) | ( n1482 & ~n1486 ) ;
  assign n1488 = ( n1371 & n1374 ) | ( n1371 & ~n1487 ) | ( n1374 & ~n1487 ) ;
  assign n1489 = ( n1358 & n1468 ) | ( n1358 & n1488 ) | ( n1468 & n1488 ) ;
  assign n1490 = x27 & ~x155 ;
  assign n1491 = ~n1121 & n1490 ;
  assign n1492 = x26 & ~x154 ;
  assign n1493 = ~n1120 & n1492 ;
  assign n1494 = ( ~n1121 & n1491 ) | ( ~n1121 & n1493 ) | ( n1491 & n1493 ) ;
  assign n1495 = ( ~n1116 & n1118 ) | ( ~n1116 & n1494 ) | ( n1118 & n1494 ) ;
  assign n1496 = n1127 | n1495 ;
  assign n1497 = ( ~n1126 & n1130 ) | ( ~n1126 & n1496 ) | ( n1130 & n1496 ) ;
  assign n1498 = n1133 | n1497 ;
  assign n1499 = ~n1115 & n1498 ;
  assign n1500 = n1148 | n1499 ;
  assign n1501 = n1100 & ~n1162 ;
  assign n1502 = ( n1162 & n1500 ) | ( n1162 & ~n1501 ) | ( n1500 & ~n1501 ) ;
  assign n1503 = n1155 | n1502 ;
  assign n1504 = ( ~n1085 & n1156 ) | ( ~n1085 & n1503 ) | ( n1156 & n1503 ) ;
  assign n1505 = ~n1085 & n1504 ;
  assign n1506 = ( ~n1338 & n1357 ) | ( ~n1338 & n1505 ) | ( n1357 & n1505 ) ;
  assign n1507 = ( n1468 & n1488 ) | ( n1468 & ~n1506 ) | ( n1488 & ~n1506 ) ;
  assign n1508 = ~x21 & x149 ;
  assign n1509 = x20 & ~x148 ;
  assign n1510 = ~n1508 & n1509 ;
  assign n1511 = ~x18 & x146 ;
  assign n1512 = ( ~x19 & x147 ) | ( ~x19 & n1511 ) | ( x147 & n1511 ) ;
  assign n1513 = ~x20 & x148 ;
  assign n1514 = n1508 | n1513 ;
  assign n1515 = ( ~n1510 & n1512 ) | ( ~n1510 & n1514 ) | ( n1512 & n1514 ) ;
  assign n1516 = ~x23 & x151 ;
  assign n1517 = ~x22 & x150 ;
  assign n1518 = x21 & ~x149 ;
  assign n1519 = ~n1517 & n1518 ;
  assign n1520 = x22 & ~x150 ;
  assign n1521 = ~n1516 & n1520 ;
  assign n1522 = ( ~n1516 & n1519 ) | ( ~n1516 & n1521 ) | ( n1519 & n1521 ) ;
  assign n1523 = x23 & ~x151 ;
  assign n1524 = x24 & ~x152 ;
  assign n1525 = ( ~x152 & n1523 ) | ( ~x152 & n1524 ) | ( n1523 & n1524 ) ;
  assign n1526 = ( ~x152 & n1522 ) | ( ~x152 & n1525 ) | ( n1522 & n1525 ) ;
  assign n1527 = n1516 | n1517 ;
  assign n1528 = ~n1523 & n1527 ;
  assign n1529 = ( x152 & ~n1524 ) | ( x152 & n1528 ) | ( ~n1524 & n1528 ) ;
  assign n1530 = ( n1515 & ~n1526 ) | ( n1515 & n1529 ) | ( ~n1526 & n1529 ) ;
  assign n1531 = x19 & ~x147 ;
  assign n1532 = ~n1513 & n1531 ;
  assign n1533 = x18 & ~x146 ;
  assign n1534 = ~n1512 & n1533 ;
  assign n1535 = ( ~n1513 & n1532 ) | ( ~n1513 & n1534 ) | ( n1532 & n1534 ) ;
  assign n1536 = ( ~n1508 & n1510 ) | ( ~n1508 & n1535 ) | ( n1510 & n1535 ) ;
  assign n1537 = n1518 | n1536 ;
  assign n1538 = ( ~x152 & n1521 ) | ( ~x152 & n1525 ) | ( n1521 & n1525 ) ;
  assign n1539 = ( ~n1529 & n1537 ) | ( ~n1529 & n1538 ) | ( n1537 & n1538 ) ;
  assign n1540 = ~x13 & x141 ;
  assign n1541 = x12 & ~x140 ;
  assign n1542 = ~n1540 & n1541 ;
  assign n1543 = ~x10 & x138 ;
  assign n1544 = ( ~x11 & x139 ) | ( ~x11 & n1543 ) | ( x139 & n1543 ) ;
  assign n1545 = ~x12 & x140 ;
  assign n1546 = n1540 | n1545 ;
  assign n1547 = ( ~n1542 & n1544 ) | ( ~n1542 & n1546 ) | ( n1544 & n1546 ) ;
  assign n1548 = x15 & ~x143 ;
  assign n1549 = ~x15 & x143 ;
  assign n1550 = ~x14 & x142 ;
  assign n1551 = x13 & ~x141 ;
  assign n1552 = ~n1550 & n1551 ;
  assign n1553 = x14 & ~x142 ;
  assign n1554 = ~n1549 & n1553 ;
  assign n1555 = ( ~n1549 & n1552 ) | ( ~n1549 & n1554 ) | ( n1552 & n1554 ) ;
  assign n1556 = n1548 | n1555 ;
  assign n1557 = ( ~x15 & x143 ) | ( ~x15 & n1550 ) | ( x143 & n1550 ) ;
  assign n1558 = ( n1547 & ~n1556 ) | ( n1547 & n1557 ) | ( ~n1556 & n1557 ) ;
  assign n1559 = x16 & ~n1558 ;
  assign n1560 = x16 & ~n1557 ;
  assign n1561 = x16 & n1548 ;
  assign n1562 = ( x16 & n1554 ) | ( x16 & n1561 ) | ( n1554 & n1561 ) ;
  assign n1563 = x11 & ~x139 ;
  assign n1564 = ~n1545 & n1563 ;
  assign n1565 = x10 & ~x138 ;
  assign n1566 = ~n1544 & n1565 ;
  assign n1567 = ( ~n1545 & n1564 ) | ( ~n1545 & n1566 ) | ( n1564 & n1566 ) ;
  assign n1568 = ( ~n1540 & n1542 ) | ( ~n1540 & n1567 ) | ( n1542 & n1567 ) ;
  assign n1569 = n1551 | n1568 ;
  assign n1570 = ( n1560 & n1562 ) | ( n1560 & n1569 ) | ( n1562 & n1569 ) ;
  assign n1571 = x7 & ~x135 ;
  assign n1572 = x8 | n1571 ;
  assign n1573 = x6 & ~x134 ;
  assign n1574 = ~x6 & x134 ;
  assign n1575 = ( ~x7 & x135 ) | ( ~x7 & n1574 ) | ( x135 & n1574 ) ;
  assign n1576 = n1573 & ~n1575 ;
  assign n1577 = n1572 | n1576 ;
  assign n1578 = ~x136 & n1577 ;
  assign n1579 = x0 & ~x128 ;
  assign n1580 = ( x1 & ~x129 ) | ( x1 & n1579 ) | ( ~x129 & n1579 ) ;
  assign n1581 = ( x2 & ~x130 ) | ( x2 & n1580 ) | ( ~x130 & n1580 ) ;
  assign n1582 = ( x3 & ~x131 ) | ( x3 & n1581 ) | ( ~x131 & n1581 ) ;
  assign n1583 = ( x4 & ~x132 ) | ( x4 & n1582 ) | ( ~x132 & n1582 ) ;
  assign n1584 = ( x5 & ~x133 ) | ( x5 & n1583 ) | ( ~x133 & n1583 ) ;
  assign n1585 = ( x136 & n1575 ) | ( x136 & ~n1578 ) | ( n1575 & ~n1578 ) ;
  assign n1586 = ( n1578 & n1584 ) | ( n1578 & ~n1585 ) | ( n1584 & ~n1585 ) ;
  assign n1587 = x8 & ~n1575 ;
  assign n1588 = x8 & n1571 ;
  assign n1589 = ( x8 & n1576 ) | ( x8 & n1588 ) | ( n1576 & n1588 ) ;
  assign n1590 = ( n1584 & n1587 ) | ( n1584 & n1589 ) | ( n1587 & n1589 ) ;
  assign n1591 = n1586 | n1590 ;
  assign n1592 = ( x9 & ~x137 ) | ( x9 & n1591 ) | ( ~x137 & n1591 ) ;
  assign n1593 = ( n1559 & n1570 ) | ( n1559 & n1592 ) | ( n1570 & n1592 ) ;
  assign n1594 = x16 & ~x144 ;
  assign n1595 = ( x144 & n1558 ) | ( x144 & ~n1594 ) | ( n1558 & ~n1594 ) ;
  assign n1596 = ( x144 & n1557 ) | ( x144 & ~n1594 ) | ( n1557 & ~n1594 ) ;
  assign n1597 = ( ~x144 & n1548 ) | ( ~x144 & n1594 ) | ( n1548 & n1594 ) ;
  assign n1598 = ( ~x144 & n1554 ) | ( ~x144 & n1597 ) | ( n1554 & n1597 ) ;
  assign n1599 = ( n1569 & ~n1596 ) | ( n1569 & n1598 ) | ( ~n1596 & n1598 ) ;
  assign n1600 = ( n1592 & ~n1595 ) | ( n1592 & n1599 ) | ( ~n1595 & n1599 ) ;
  assign n1601 = n1593 | n1600 ;
  assign n1602 = ( x17 & ~x145 ) | ( x17 & n1601 ) | ( ~x145 & n1601 ) ;
  assign n1603 = ( ~n1530 & n1539 ) | ( ~n1530 & n1602 ) | ( n1539 & n1602 ) ;
  assign n1604 = x24 & n1523 ;
  assign n1605 = ( x24 & n1521 ) | ( x24 & n1604 ) | ( n1521 & n1604 ) ;
  assign n1606 = ( x24 & ~n1527 ) | ( x24 & n1604 ) | ( ~n1527 & n1604 ) ;
  assign n1607 = ( n1537 & n1605 ) | ( n1537 & n1606 ) | ( n1605 & n1606 ) ;
  assign n1608 = ( x24 & n1522 ) | ( x24 & n1604 ) | ( n1522 & n1604 ) ;
  assign n1609 = ( ~n1515 & n1606 ) | ( ~n1515 & n1608 ) | ( n1606 & n1608 ) ;
  assign n1610 = ( n1602 & n1607 ) | ( n1602 & n1609 ) | ( n1607 & n1609 ) ;
  assign n1611 = n1603 | n1610 ;
  assign n1612 = ( x25 & ~x153 ) | ( x25 & n1611 ) | ( ~x153 & n1611 ) ;
  assign n1613 = ( n1489 & n1507 ) | ( n1489 & ~n1612 ) | ( n1507 & ~n1612 ) ;
  assign n1614 = x111 & ~n1370 ;
  assign n1615 = x111 & n1373 ;
  assign n1616 = ( ~n1467 & n1614 ) | ( ~n1467 & n1615 ) | ( n1614 & n1615 ) ;
  assign n1617 = ( n1487 & n1614 ) | ( n1487 & n1615 ) | ( n1614 & n1615 ) ;
  assign n1618 = ( ~n1358 & n1616 ) | ( ~n1358 & n1617 ) | ( n1616 & n1617 ) ;
  assign n1619 = ( n1506 & n1616 ) | ( n1506 & n1617 ) | ( n1616 & n1617 ) ;
  assign n1620 = ( n1612 & n1618 ) | ( n1612 & n1619 ) | ( n1618 & n1619 ) ;
  assign n1621 = n1613 | n1620 ;
  assign n1622 = x495 & n812 ;
  assign n1623 = x495 & ~n815 ;
  assign n1624 = ( n909 & n1622 ) | ( n909 & n1623 ) | ( n1622 & n1623 ) ;
  assign n1625 = ( ~n929 & n1622 ) | ( ~n929 & n1623 ) | ( n1622 & n1623 ) ;
  assign n1626 = ( n800 & n1624 ) | ( n800 & n1625 ) | ( n1624 & n1625 ) ;
  assign n1627 = ( ~n948 & n1624 ) | ( ~n948 & n1625 ) | ( n1624 & n1625 ) ;
  assign n1628 = ( ~n1061 & n1626 ) | ( ~n1061 & n1627 ) | ( n1626 & n1627 ) ;
  assign n1629 = x367 & ~n812 ;
  assign n1630 = x367 & n815 ;
  assign n1631 = ( ~n909 & n1629 ) | ( ~n909 & n1630 ) | ( n1629 & n1630 ) ;
  assign n1632 = ( n929 & n1629 ) | ( n929 & n1630 ) | ( n1629 & n1630 ) ;
  assign n1633 = ( ~n800 & n1631 ) | ( ~n800 & n1632 ) | ( n1631 & n1632 ) ;
  assign n1634 = ( n948 & n1631 ) | ( n948 & n1632 ) | ( n1631 & n1632 ) ;
  assign n1635 = ( n1061 & n1633 ) | ( n1061 & n1634 ) | ( n1633 & n1634 ) ;
  assign n1636 = n1628 | n1635 ;
  assign n1637 = ~n1621 & n1636 ;
  assign n1638 = x494 & n812 ;
  assign n1639 = x494 & ~n815 ;
  assign n1640 = ( n909 & n1638 ) | ( n909 & n1639 ) | ( n1638 & n1639 ) ;
  assign n1641 = ( ~n929 & n1638 ) | ( ~n929 & n1639 ) | ( n1638 & n1639 ) ;
  assign n1642 = ( n800 & n1640 ) | ( n800 & n1641 ) | ( n1640 & n1641 ) ;
  assign n1643 = ( ~n948 & n1640 ) | ( ~n948 & n1641 ) | ( n1640 & n1641 ) ;
  assign n1644 = ( ~n1061 & n1642 ) | ( ~n1061 & n1643 ) | ( n1642 & n1643 ) ;
  assign n1645 = x366 & ~n812 ;
  assign n1646 = x366 & n815 ;
  assign n1647 = ( ~n909 & n1645 ) | ( ~n909 & n1646 ) | ( n1645 & n1646 ) ;
  assign n1648 = ( n929 & n1645 ) | ( n929 & n1646 ) | ( n1645 & n1646 ) ;
  assign n1649 = ( ~n800 & n1647 ) | ( ~n800 & n1648 ) | ( n1647 & n1648 ) ;
  assign n1650 = ( n948 & n1647 ) | ( n948 & n1648 ) | ( n1647 & n1648 ) ;
  assign n1651 = ( n1061 & n1649 ) | ( n1061 & n1650 ) | ( n1649 & n1650 ) ;
  assign n1652 = n1644 | n1651 ;
  assign n1653 = x238 & n1370 ;
  assign n1654 = x238 & ~n1373 ;
  assign n1655 = ( n1467 & n1653 ) | ( n1467 & n1654 ) | ( n1653 & n1654 ) ;
  assign n1656 = ( ~n1487 & n1653 ) | ( ~n1487 & n1654 ) | ( n1653 & n1654 ) ;
  assign n1657 = ( n1358 & n1655 ) | ( n1358 & n1656 ) | ( n1655 & n1656 ) ;
  assign n1658 = ( ~n1506 & n1655 ) | ( ~n1506 & n1656 ) | ( n1655 & n1656 ) ;
  assign n1659 = ( ~n1612 & n1657 ) | ( ~n1612 & n1658 ) | ( n1657 & n1658 ) ;
  assign n1660 = x110 & ~n1370 ;
  assign n1661 = x110 & n1373 ;
  assign n1662 = ( ~n1467 & n1660 ) | ( ~n1467 & n1661 ) | ( n1660 & n1661 ) ;
  assign n1663 = ( n1487 & n1660 ) | ( n1487 & n1661 ) | ( n1660 & n1661 ) ;
  assign n1664 = ( ~n1358 & n1662 ) | ( ~n1358 & n1663 ) | ( n1662 & n1663 ) ;
  assign n1665 = ( n1506 & n1662 ) | ( n1506 & n1663 ) | ( n1662 & n1663 ) ;
  assign n1666 = ( n1612 & n1664 ) | ( n1612 & n1665 ) | ( n1664 & n1665 ) ;
  assign n1667 = n1659 | n1666 ;
  assign n1668 = ~n1652 & n1667 ;
  assign n1669 = ~n1637 & n1668 ;
  assign n1670 = n1652 & ~n1667 ;
  assign n1671 = n1637 | n1670 ;
  assign n1672 = x237 & n1370 ;
  assign n1673 = x237 & ~n1373 ;
  assign n1674 = ( n1467 & n1672 ) | ( n1467 & n1673 ) | ( n1672 & n1673 ) ;
  assign n1675 = ( ~n1487 & n1672 ) | ( ~n1487 & n1673 ) | ( n1672 & n1673 ) ;
  assign n1676 = ( n1358 & n1674 ) | ( n1358 & n1675 ) | ( n1674 & n1675 ) ;
  assign n1677 = ( ~n1506 & n1674 ) | ( ~n1506 & n1675 ) | ( n1674 & n1675 ) ;
  assign n1678 = ( ~n1612 & n1676 ) | ( ~n1612 & n1677 ) | ( n1676 & n1677 ) ;
  assign n1679 = x109 & ~n1370 ;
  assign n1680 = x109 & n1373 ;
  assign n1681 = ( ~n1467 & n1679 ) | ( ~n1467 & n1680 ) | ( n1679 & n1680 ) ;
  assign n1682 = ( n1487 & n1679 ) | ( n1487 & n1680 ) | ( n1679 & n1680 ) ;
  assign n1683 = ( ~n1358 & n1681 ) | ( ~n1358 & n1682 ) | ( n1681 & n1682 ) ;
  assign n1684 = ( n1506 & n1681 ) | ( n1506 & n1682 ) | ( n1681 & n1682 ) ;
  assign n1685 = ( n1612 & n1683 ) | ( n1612 & n1684 ) | ( n1683 & n1684 ) ;
  assign n1686 = n1678 | n1685 ;
  assign n1687 = x493 & n812 ;
  assign n1688 = x493 & ~n815 ;
  assign n1689 = ( n909 & n1687 ) | ( n909 & n1688 ) | ( n1687 & n1688 ) ;
  assign n1690 = ( ~n929 & n1687 ) | ( ~n929 & n1688 ) | ( n1687 & n1688 ) ;
  assign n1691 = ( n800 & n1689 ) | ( n800 & n1690 ) | ( n1689 & n1690 ) ;
  assign n1692 = ( ~n948 & n1689 ) | ( ~n948 & n1690 ) | ( n1689 & n1690 ) ;
  assign n1693 = ( ~n1061 & n1691 ) | ( ~n1061 & n1692 ) | ( n1691 & n1692 ) ;
  assign n1694 = x365 & ~n812 ;
  assign n1695 = x365 & n815 ;
  assign n1696 = ( ~n909 & n1694 ) | ( ~n909 & n1695 ) | ( n1694 & n1695 ) ;
  assign n1697 = ( n929 & n1694 ) | ( n929 & n1695 ) | ( n1694 & n1695 ) ;
  assign n1698 = ( ~n800 & n1696 ) | ( ~n800 & n1697 ) | ( n1696 & n1697 ) ;
  assign n1699 = ( n948 & n1696 ) | ( n948 & n1697 ) | ( n1696 & n1697 ) ;
  assign n1700 = ( n1061 & n1698 ) | ( n1061 & n1699 ) | ( n1698 & n1699 ) ;
  assign n1701 = n1693 | n1700 ;
  assign n1702 = ~n1686 & n1701 ;
  assign n1703 = x236 & n1370 ;
  assign n1704 = x236 & ~n1373 ;
  assign n1705 = ( n1467 & n1703 ) | ( n1467 & n1704 ) | ( n1703 & n1704 ) ;
  assign n1706 = ( ~n1487 & n1703 ) | ( ~n1487 & n1704 ) | ( n1703 & n1704 ) ;
  assign n1707 = ( n1358 & n1705 ) | ( n1358 & n1706 ) | ( n1705 & n1706 ) ;
  assign n1708 = ( ~n1506 & n1705 ) | ( ~n1506 & n1706 ) | ( n1705 & n1706 ) ;
  assign n1709 = ( ~n1612 & n1707 ) | ( ~n1612 & n1708 ) | ( n1707 & n1708 ) ;
  assign n1710 = x108 & ~n1370 ;
  assign n1711 = x108 & n1373 ;
  assign n1712 = ( ~n1467 & n1710 ) | ( ~n1467 & n1711 ) | ( n1710 & n1711 ) ;
  assign n1713 = ( n1487 & n1710 ) | ( n1487 & n1711 ) | ( n1710 & n1711 ) ;
  assign n1714 = ( ~n1358 & n1712 ) | ( ~n1358 & n1713 ) | ( n1712 & n1713 ) ;
  assign n1715 = ( n1506 & n1712 ) | ( n1506 & n1713 ) | ( n1712 & n1713 ) ;
  assign n1716 = ( n1612 & n1714 ) | ( n1612 & n1715 ) | ( n1714 & n1715 ) ;
  assign n1717 = n1709 | n1716 ;
  assign n1718 = x492 & n812 ;
  assign n1719 = x492 & ~n815 ;
  assign n1720 = ( n909 & n1718 ) | ( n909 & n1719 ) | ( n1718 & n1719 ) ;
  assign n1721 = ( ~n929 & n1718 ) | ( ~n929 & n1719 ) | ( n1718 & n1719 ) ;
  assign n1722 = ( n800 & n1720 ) | ( n800 & n1721 ) | ( n1720 & n1721 ) ;
  assign n1723 = ( ~n948 & n1720 ) | ( ~n948 & n1721 ) | ( n1720 & n1721 ) ;
  assign n1724 = ( ~n1061 & n1722 ) | ( ~n1061 & n1723 ) | ( n1722 & n1723 ) ;
  assign n1725 = x364 & ~n812 ;
  assign n1726 = x364 & n815 ;
  assign n1727 = ( ~n909 & n1725 ) | ( ~n909 & n1726 ) | ( n1725 & n1726 ) ;
  assign n1728 = ( n929 & n1725 ) | ( n929 & n1726 ) | ( n1725 & n1726 ) ;
  assign n1729 = ( ~n800 & n1727 ) | ( ~n800 & n1728 ) | ( n1727 & n1728 ) ;
  assign n1730 = ( n948 & n1727 ) | ( n948 & n1728 ) | ( n1727 & n1728 ) ;
  assign n1731 = ( n1061 & n1729 ) | ( n1061 & n1730 ) | ( n1729 & n1730 ) ;
  assign n1732 = n1724 | n1731 ;
  assign n1733 = ~n1717 & n1732 ;
  assign n1734 = n1702 | n1733 ;
  assign n1735 = n1671 | n1734 ;
  assign n1736 = ~n1669 & n1735 ;
  assign n1737 = x235 & n1370 ;
  assign n1738 = x235 & ~n1373 ;
  assign n1739 = ( n1467 & n1737 ) | ( n1467 & n1738 ) | ( n1737 & n1738 ) ;
  assign n1740 = ( ~n1487 & n1737 ) | ( ~n1487 & n1738 ) | ( n1737 & n1738 ) ;
  assign n1741 = ( n1358 & n1739 ) | ( n1358 & n1740 ) | ( n1739 & n1740 ) ;
  assign n1742 = ( ~n1506 & n1739 ) | ( ~n1506 & n1740 ) | ( n1739 & n1740 ) ;
  assign n1743 = ( ~n1612 & n1741 ) | ( ~n1612 & n1742 ) | ( n1741 & n1742 ) ;
  assign n1744 = x107 & ~n1370 ;
  assign n1745 = x107 & n1373 ;
  assign n1746 = ( ~n1467 & n1744 ) | ( ~n1467 & n1745 ) | ( n1744 & n1745 ) ;
  assign n1747 = ( n1487 & n1744 ) | ( n1487 & n1745 ) | ( n1744 & n1745 ) ;
  assign n1748 = ( ~n1358 & n1746 ) | ( ~n1358 & n1747 ) | ( n1746 & n1747 ) ;
  assign n1749 = ( n1506 & n1746 ) | ( n1506 & n1747 ) | ( n1746 & n1747 ) ;
  assign n1750 = ( n1612 & n1748 ) | ( n1612 & n1749 ) | ( n1748 & n1749 ) ;
  assign n1751 = n1743 | n1750 ;
  assign n1752 = x491 & n812 ;
  assign n1753 = x491 & ~n815 ;
  assign n1754 = ( n909 & n1752 ) | ( n909 & n1753 ) | ( n1752 & n1753 ) ;
  assign n1755 = ( ~n929 & n1752 ) | ( ~n929 & n1753 ) | ( n1752 & n1753 ) ;
  assign n1756 = ( n800 & n1754 ) | ( n800 & n1755 ) | ( n1754 & n1755 ) ;
  assign n1757 = ( ~n948 & n1754 ) | ( ~n948 & n1755 ) | ( n1754 & n1755 ) ;
  assign n1758 = ( ~n1061 & n1756 ) | ( ~n1061 & n1757 ) | ( n1756 & n1757 ) ;
  assign n1759 = x363 & ~n812 ;
  assign n1760 = x363 & n815 ;
  assign n1761 = ( ~n909 & n1759 ) | ( ~n909 & n1760 ) | ( n1759 & n1760 ) ;
  assign n1762 = ( n929 & n1759 ) | ( n929 & n1760 ) | ( n1759 & n1760 ) ;
  assign n1763 = ( ~n800 & n1761 ) | ( ~n800 & n1762 ) | ( n1761 & n1762 ) ;
  assign n1764 = ( n948 & n1761 ) | ( n948 & n1762 ) | ( n1761 & n1762 ) ;
  assign n1765 = ( n1061 & n1763 ) | ( n1061 & n1764 ) | ( n1763 & n1764 ) ;
  assign n1766 = n1758 | n1765 ;
  assign n1767 = x490 & n812 ;
  assign n1768 = x490 & ~n815 ;
  assign n1769 = ( n909 & n1767 ) | ( n909 & n1768 ) | ( n1767 & n1768 ) ;
  assign n1770 = ( ~n929 & n1767 ) | ( ~n929 & n1768 ) | ( n1767 & n1768 ) ;
  assign n1771 = ( n800 & n1769 ) | ( n800 & n1770 ) | ( n1769 & n1770 ) ;
  assign n1772 = ( ~n948 & n1769 ) | ( ~n948 & n1770 ) | ( n1769 & n1770 ) ;
  assign n1773 = ( ~n1061 & n1771 ) | ( ~n1061 & n1772 ) | ( n1771 & n1772 ) ;
  assign n1774 = x362 & ~n812 ;
  assign n1775 = x362 & n815 ;
  assign n1776 = ( ~n909 & n1774 ) | ( ~n909 & n1775 ) | ( n1774 & n1775 ) ;
  assign n1777 = ( n929 & n1774 ) | ( n929 & n1775 ) | ( n1774 & n1775 ) ;
  assign n1778 = ( ~n800 & n1776 ) | ( ~n800 & n1777 ) | ( n1776 & n1777 ) ;
  assign n1779 = ( n948 & n1776 ) | ( n948 & n1777 ) | ( n1776 & n1777 ) ;
  assign n1780 = ( n1061 & n1778 ) | ( n1061 & n1779 ) | ( n1778 & n1779 ) ;
  assign n1781 = n1773 | n1780 ;
  assign n1782 = x234 & n1370 ;
  assign n1783 = x234 & ~n1373 ;
  assign n1784 = ( n1467 & n1782 ) | ( n1467 & n1783 ) | ( n1782 & n1783 ) ;
  assign n1785 = ( ~n1487 & n1782 ) | ( ~n1487 & n1783 ) | ( n1782 & n1783 ) ;
  assign n1786 = ( n1358 & n1784 ) | ( n1358 & n1785 ) | ( n1784 & n1785 ) ;
  assign n1787 = ( ~n1506 & n1784 ) | ( ~n1506 & n1785 ) | ( n1784 & n1785 ) ;
  assign n1788 = ( ~n1612 & n1786 ) | ( ~n1612 & n1787 ) | ( n1786 & n1787 ) ;
  assign n1789 = x106 & ~n1370 ;
  assign n1790 = x106 & n1373 ;
  assign n1791 = ( ~n1467 & n1789 ) | ( ~n1467 & n1790 ) | ( n1789 & n1790 ) ;
  assign n1792 = ( n1487 & n1789 ) | ( n1487 & n1790 ) | ( n1789 & n1790 ) ;
  assign n1793 = ( ~n1358 & n1791 ) | ( ~n1358 & n1792 ) | ( n1791 & n1792 ) ;
  assign n1794 = ( n1506 & n1791 ) | ( n1506 & n1792 ) | ( n1791 & n1792 ) ;
  assign n1795 = ( n1612 & n1793 ) | ( n1612 & n1794 ) | ( n1793 & n1794 ) ;
  assign n1796 = n1788 | n1795 ;
  assign n1797 = x233 & n1370 ;
  assign n1798 = x233 & ~n1373 ;
  assign n1799 = ( n1467 & n1797 ) | ( n1467 & n1798 ) | ( n1797 & n1798 ) ;
  assign n1800 = ( ~n1487 & n1797 ) | ( ~n1487 & n1798 ) | ( n1797 & n1798 ) ;
  assign n1801 = ( n1358 & n1799 ) | ( n1358 & n1800 ) | ( n1799 & n1800 ) ;
  assign n1802 = ( ~n1506 & n1799 ) | ( ~n1506 & n1800 ) | ( n1799 & n1800 ) ;
  assign n1803 = ( ~n1612 & n1801 ) | ( ~n1612 & n1802 ) | ( n1801 & n1802 ) ;
  assign n1804 = x105 & ~n1370 ;
  assign n1805 = x105 & n1373 ;
  assign n1806 = ( ~n1467 & n1804 ) | ( ~n1467 & n1805 ) | ( n1804 & n1805 ) ;
  assign n1807 = ( n1487 & n1804 ) | ( n1487 & n1805 ) | ( n1804 & n1805 ) ;
  assign n1808 = ( ~n1358 & n1806 ) | ( ~n1358 & n1807 ) | ( n1806 & n1807 ) ;
  assign n1809 = ( n1506 & n1806 ) | ( n1506 & n1807 ) | ( n1806 & n1807 ) ;
  assign n1810 = ( n1612 & n1808 ) | ( n1612 & n1809 ) | ( n1808 & n1809 ) ;
  assign n1811 = n1803 | n1810 ;
  assign n1812 = x489 & n812 ;
  assign n1813 = x489 & ~n815 ;
  assign n1814 = ( n909 & n1812 ) | ( n909 & n1813 ) | ( n1812 & n1813 ) ;
  assign n1815 = ( ~n929 & n1812 ) | ( ~n929 & n1813 ) | ( n1812 & n1813 ) ;
  assign n1816 = ( n800 & n1814 ) | ( n800 & n1815 ) | ( n1814 & n1815 ) ;
  assign n1817 = ( ~n948 & n1814 ) | ( ~n948 & n1815 ) | ( n1814 & n1815 ) ;
  assign n1818 = ( ~n1061 & n1816 ) | ( ~n1061 & n1817 ) | ( n1816 & n1817 ) ;
  assign n1819 = x361 & ~n812 ;
  assign n1820 = x361 & n815 ;
  assign n1821 = ( ~n909 & n1819 ) | ( ~n909 & n1820 ) | ( n1819 & n1820 ) ;
  assign n1822 = ( n929 & n1819 ) | ( n929 & n1820 ) | ( n1819 & n1820 ) ;
  assign n1823 = ( ~n800 & n1821 ) | ( ~n800 & n1822 ) | ( n1821 & n1822 ) ;
  assign n1824 = ( n948 & n1821 ) | ( n948 & n1822 ) | ( n1821 & n1822 ) ;
  assign n1825 = ( n1061 & n1823 ) | ( n1061 & n1824 ) | ( n1823 & n1824 ) ;
  assign n1826 = n1818 | n1825 ;
  assign n1827 = x488 & n812 ;
  assign n1828 = x488 & ~n815 ;
  assign n1829 = ( n909 & n1827 ) | ( n909 & n1828 ) | ( n1827 & n1828 ) ;
  assign n1830 = ( ~n929 & n1827 ) | ( ~n929 & n1828 ) | ( n1827 & n1828 ) ;
  assign n1831 = ( n800 & n1829 ) | ( n800 & n1830 ) | ( n1829 & n1830 ) ;
  assign n1832 = ( ~n948 & n1829 ) | ( ~n948 & n1830 ) | ( n1829 & n1830 ) ;
  assign n1833 = ( ~n1061 & n1831 ) | ( ~n1061 & n1832 ) | ( n1831 & n1832 ) ;
  assign n1834 = x360 & ~n812 ;
  assign n1835 = x360 & n815 ;
  assign n1836 = ( ~n909 & n1834 ) | ( ~n909 & n1835 ) | ( n1834 & n1835 ) ;
  assign n1837 = ( n929 & n1834 ) | ( n929 & n1835 ) | ( n1834 & n1835 ) ;
  assign n1838 = ( ~n800 & n1836 ) | ( ~n800 & n1837 ) | ( n1836 & n1837 ) ;
  assign n1839 = ( n948 & n1836 ) | ( n948 & n1837 ) | ( n1836 & n1837 ) ;
  assign n1840 = ( n1061 & n1838 ) | ( n1061 & n1839 ) | ( n1838 & n1839 ) ;
  assign n1841 = n1833 | n1840 ;
  assign n1842 = x232 & n1370 ;
  assign n1843 = x232 & ~n1373 ;
  assign n1844 = ( n1467 & n1842 ) | ( n1467 & n1843 ) | ( n1842 & n1843 ) ;
  assign n1845 = ( ~n1487 & n1842 ) | ( ~n1487 & n1843 ) | ( n1842 & n1843 ) ;
  assign n1846 = ( n1358 & n1844 ) | ( n1358 & n1845 ) | ( n1844 & n1845 ) ;
  assign n1847 = ( ~n1506 & n1844 ) | ( ~n1506 & n1845 ) | ( n1844 & n1845 ) ;
  assign n1848 = ( ~n1612 & n1846 ) | ( ~n1612 & n1847 ) | ( n1846 & n1847 ) ;
  assign n1849 = x104 & ~n1370 ;
  assign n1850 = x104 & n1373 ;
  assign n1851 = ( ~n1467 & n1849 ) | ( ~n1467 & n1850 ) | ( n1849 & n1850 ) ;
  assign n1852 = ( n1487 & n1849 ) | ( n1487 & n1850 ) | ( n1849 & n1850 ) ;
  assign n1853 = ( ~n1358 & n1851 ) | ( ~n1358 & n1852 ) | ( n1851 & n1852 ) ;
  assign n1854 = ( n1506 & n1851 ) | ( n1506 & n1852 ) | ( n1851 & n1852 ) ;
  assign n1855 = ( n1612 & n1853 ) | ( n1612 & n1854 ) | ( n1853 & n1854 ) ;
  assign n1856 = n1848 | n1855 ;
  assign n1857 = ~n1841 & n1856 ;
  assign n1858 = ( n1811 & ~n1826 ) | ( n1811 & n1857 ) | ( ~n1826 & n1857 ) ;
  assign n1859 = ( ~n1781 & n1796 ) | ( ~n1781 & n1858 ) | ( n1796 & n1858 ) ;
  assign n1860 = ( n1751 & ~n1766 ) | ( n1751 & n1859 ) | ( ~n1766 & n1859 ) ;
  assign n1861 = ( n1669 & ~n1736 ) | ( n1669 & n1860 ) | ( ~n1736 & n1860 ) ;
  assign n1862 = n1621 & ~n1636 ;
  assign n1863 = n1717 & ~n1732 ;
  assign n1864 = ( n1686 & ~n1701 ) | ( n1686 & n1863 ) | ( ~n1701 & n1863 ) ;
  assign n1865 = ~n1671 & n1864 ;
  assign n1866 = n1862 | n1865 ;
  assign n1867 = n1861 | n1866 ;
  assign n1868 = x251 & n1370 ;
  assign n1869 = x251 & ~n1373 ;
  assign n1870 = ( n1467 & n1868 ) | ( n1467 & n1869 ) | ( n1868 & n1869 ) ;
  assign n1871 = ( ~n1487 & n1868 ) | ( ~n1487 & n1869 ) | ( n1868 & n1869 ) ;
  assign n1872 = ( n1358 & n1870 ) | ( n1358 & n1871 ) | ( n1870 & n1871 ) ;
  assign n1873 = ( ~n1506 & n1870 ) | ( ~n1506 & n1871 ) | ( n1870 & n1871 ) ;
  assign n1874 = ( ~n1612 & n1872 ) | ( ~n1612 & n1873 ) | ( n1872 & n1873 ) ;
  assign n1875 = x123 & ~n1370 ;
  assign n1876 = x123 & n1373 ;
  assign n1877 = ( ~n1467 & n1875 ) | ( ~n1467 & n1876 ) | ( n1875 & n1876 ) ;
  assign n1878 = ( n1487 & n1875 ) | ( n1487 & n1876 ) | ( n1875 & n1876 ) ;
  assign n1879 = ( ~n1358 & n1877 ) | ( ~n1358 & n1878 ) | ( n1877 & n1878 ) ;
  assign n1880 = ( n1506 & n1877 ) | ( n1506 & n1878 ) | ( n1877 & n1878 ) ;
  assign n1881 = ( n1612 & n1879 ) | ( n1612 & n1880 ) | ( n1879 & n1880 ) ;
  assign n1882 = n1874 | n1881 ;
  assign n1883 = x507 & n812 ;
  assign n1884 = x507 & ~n815 ;
  assign n1885 = ( n909 & n1883 ) | ( n909 & n1884 ) | ( n1883 & n1884 ) ;
  assign n1886 = ( ~n929 & n1883 ) | ( ~n929 & n1884 ) | ( n1883 & n1884 ) ;
  assign n1887 = ( n800 & n1885 ) | ( n800 & n1886 ) | ( n1885 & n1886 ) ;
  assign n1888 = ( ~n948 & n1885 ) | ( ~n948 & n1886 ) | ( n1885 & n1886 ) ;
  assign n1889 = ( ~n1061 & n1887 ) | ( ~n1061 & n1888 ) | ( n1887 & n1888 ) ;
  assign n1890 = x379 & ~n812 ;
  assign n1891 = x379 & n815 ;
  assign n1892 = ( ~n909 & n1890 ) | ( ~n909 & n1891 ) | ( n1890 & n1891 ) ;
  assign n1893 = ( n929 & n1890 ) | ( n929 & n1891 ) | ( n1890 & n1891 ) ;
  assign n1894 = ( ~n800 & n1892 ) | ( ~n800 & n1893 ) | ( n1892 & n1893 ) ;
  assign n1895 = ( n948 & n1892 ) | ( n948 & n1893 ) | ( n1892 & n1893 ) ;
  assign n1896 = ( n1061 & n1894 ) | ( n1061 & n1895 ) | ( n1894 & n1895 ) ;
  assign n1897 = n1889 | n1896 ;
  assign n1898 = ~n1882 & n1897 ;
  assign n1899 = x506 & n812 ;
  assign n1900 = x506 & ~n815 ;
  assign n1901 = ( n909 & n1899 ) | ( n909 & n1900 ) | ( n1899 & n1900 ) ;
  assign n1902 = ( ~n929 & n1899 ) | ( ~n929 & n1900 ) | ( n1899 & n1900 ) ;
  assign n1903 = ( n800 & n1901 ) | ( n800 & n1902 ) | ( n1901 & n1902 ) ;
  assign n1904 = ( ~n948 & n1901 ) | ( ~n948 & n1902 ) | ( n1901 & n1902 ) ;
  assign n1905 = ( ~n1061 & n1903 ) | ( ~n1061 & n1904 ) | ( n1903 & n1904 ) ;
  assign n1906 = x378 & ~n812 ;
  assign n1907 = x378 & n815 ;
  assign n1908 = ( ~n909 & n1906 ) | ( ~n909 & n1907 ) | ( n1906 & n1907 ) ;
  assign n1909 = ( n929 & n1906 ) | ( n929 & n1907 ) | ( n1906 & n1907 ) ;
  assign n1910 = ( ~n800 & n1908 ) | ( ~n800 & n1909 ) | ( n1908 & n1909 ) ;
  assign n1911 = ( n948 & n1908 ) | ( n948 & n1909 ) | ( n1908 & n1909 ) ;
  assign n1912 = ( n1061 & n1910 ) | ( n1061 & n1911 ) | ( n1910 & n1911 ) ;
  assign n1913 = n1905 | n1912 ;
  assign n1914 = x250 & n1370 ;
  assign n1915 = x250 & ~n1373 ;
  assign n1916 = ( n1467 & n1914 ) | ( n1467 & n1915 ) | ( n1914 & n1915 ) ;
  assign n1917 = ( ~n1487 & n1914 ) | ( ~n1487 & n1915 ) | ( n1914 & n1915 ) ;
  assign n1918 = ( n1358 & n1916 ) | ( n1358 & n1917 ) | ( n1916 & n1917 ) ;
  assign n1919 = ( ~n1506 & n1916 ) | ( ~n1506 & n1917 ) | ( n1916 & n1917 ) ;
  assign n1920 = ( ~n1612 & n1918 ) | ( ~n1612 & n1919 ) | ( n1918 & n1919 ) ;
  assign n1921 = x122 & ~n1370 ;
  assign n1922 = x122 & n1373 ;
  assign n1923 = ( ~n1467 & n1921 ) | ( ~n1467 & n1922 ) | ( n1921 & n1922 ) ;
  assign n1924 = ( n1487 & n1921 ) | ( n1487 & n1922 ) | ( n1921 & n1922 ) ;
  assign n1925 = ( ~n1358 & n1923 ) | ( ~n1358 & n1924 ) | ( n1923 & n1924 ) ;
  assign n1926 = ( n1506 & n1923 ) | ( n1506 & n1924 ) | ( n1923 & n1924 ) ;
  assign n1927 = ( n1612 & n1925 ) | ( n1612 & n1926 ) | ( n1925 & n1926 ) ;
  assign n1928 = n1920 | n1927 ;
  assign n1929 = n1913 & ~n1928 ;
  assign n1930 = n1898 | n1929 ;
  assign n1931 = x249 & n1370 ;
  assign n1932 = x249 & ~n1373 ;
  assign n1933 = ( n1467 & n1931 ) | ( n1467 & n1932 ) | ( n1931 & n1932 ) ;
  assign n1934 = ( ~n1487 & n1931 ) | ( ~n1487 & n1932 ) | ( n1931 & n1932 ) ;
  assign n1935 = ( n1358 & n1933 ) | ( n1358 & n1934 ) | ( n1933 & n1934 ) ;
  assign n1936 = ( ~n1506 & n1933 ) | ( ~n1506 & n1934 ) | ( n1933 & n1934 ) ;
  assign n1937 = ( ~n1612 & n1935 ) | ( ~n1612 & n1936 ) | ( n1935 & n1936 ) ;
  assign n1938 = x121 & ~n1370 ;
  assign n1939 = x121 & n1373 ;
  assign n1940 = ( ~n1467 & n1938 ) | ( ~n1467 & n1939 ) | ( n1938 & n1939 ) ;
  assign n1941 = ( n1487 & n1938 ) | ( n1487 & n1939 ) | ( n1938 & n1939 ) ;
  assign n1942 = ( ~n1358 & n1940 ) | ( ~n1358 & n1941 ) | ( n1940 & n1941 ) ;
  assign n1943 = ( n1506 & n1940 ) | ( n1506 & n1941 ) | ( n1940 & n1941 ) ;
  assign n1944 = ( n1612 & n1942 ) | ( n1612 & n1943 ) | ( n1942 & n1943 ) ;
  assign n1945 = n1937 | n1944 ;
  assign n1946 = x505 & n812 ;
  assign n1947 = x505 & ~n815 ;
  assign n1948 = ( n909 & n1946 ) | ( n909 & n1947 ) | ( n1946 & n1947 ) ;
  assign n1949 = ( ~n929 & n1946 ) | ( ~n929 & n1947 ) | ( n1946 & n1947 ) ;
  assign n1950 = ( n800 & n1948 ) | ( n800 & n1949 ) | ( n1948 & n1949 ) ;
  assign n1951 = ( ~n948 & n1948 ) | ( ~n948 & n1949 ) | ( n1948 & n1949 ) ;
  assign n1952 = ( ~n1061 & n1950 ) | ( ~n1061 & n1951 ) | ( n1950 & n1951 ) ;
  assign n1953 = x377 & ~n812 ;
  assign n1954 = x377 & n815 ;
  assign n1955 = ( ~n909 & n1953 ) | ( ~n909 & n1954 ) | ( n1953 & n1954 ) ;
  assign n1956 = ( n929 & n1953 ) | ( n929 & n1954 ) | ( n1953 & n1954 ) ;
  assign n1957 = ( ~n800 & n1955 ) | ( ~n800 & n1956 ) | ( n1955 & n1956 ) ;
  assign n1958 = ( n948 & n1955 ) | ( n948 & n1956 ) | ( n1955 & n1956 ) ;
  assign n1959 = ( n1061 & n1957 ) | ( n1061 & n1958 ) | ( n1957 & n1958 ) ;
  assign n1960 = n1952 | n1959 ;
  assign n1961 = ~n1945 & n1960 ;
  assign n1962 = x504 & n812 ;
  assign n1963 = x504 & ~n815 ;
  assign n1964 = ( n909 & n1962 ) | ( n909 & n1963 ) | ( n1962 & n1963 ) ;
  assign n1965 = ( ~n929 & n1962 ) | ( ~n929 & n1963 ) | ( n1962 & n1963 ) ;
  assign n1966 = ( n800 & n1964 ) | ( n800 & n1965 ) | ( n1964 & n1965 ) ;
  assign n1967 = ( ~n948 & n1964 ) | ( ~n948 & n1965 ) | ( n1964 & n1965 ) ;
  assign n1968 = ( ~n1061 & n1966 ) | ( ~n1061 & n1967 ) | ( n1966 & n1967 ) ;
  assign n1969 = x376 & ~n812 ;
  assign n1970 = x376 & n815 ;
  assign n1971 = ( ~n909 & n1969 ) | ( ~n909 & n1970 ) | ( n1969 & n1970 ) ;
  assign n1972 = ( n929 & n1969 ) | ( n929 & n1970 ) | ( n1969 & n1970 ) ;
  assign n1973 = ( ~n800 & n1971 ) | ( ~n800 & n1972 ) | ( n1971 & n1972 ) ;
  assign n1974 = ( n948 & n1971 ) | ( n948 & n1972 ) | ( n1971 & n1972 ) ;
  assign n1975 = ( n1061 & n1973 ) | ( n1061 & n1974 ) | ( n1973 & n1974 ) ;
  assign n1976 = n1968 | n1975 ;
  assign n1977 = x248 & n1370 ;
  assign n1978 = x248 & ~n1373 ;
  assign n1979 = ( n1467 & n1977 ) | ( n1467 & n1978 ) | ( n1977 & n1978 ) ;
  assign n1980 = ( ~n1487 & n1977 ) | ( ~n1487 & n1978 ) | ( n1977 & n1978 ) ;
  assign n1981 = ( n1358 & n1979 ) | ( n1358 & n1980 ) | ( n1979 & n1980 ) ;
  assign n1982 = ( ~n1506 & n1979 ) | ( ~n1506 & n1980 ) | ( n1979 & n1980 ) ;
  assign n1983 = ( ~n1612 & n1981 ) | ( ~n1612 & n1982 ) | ( n1981 & n1982 ) ;
  assign n1984 = x120 & ~n1370 ;
  assign n1985 = x120 & n1373 ;
  assign n1986 = ( ~n1467 & n1984 ) | ( ~n1467 & n1985 ) | ( n1984 & n1985 ) ;
  assign n1987 = ( n1487 & n1984 ) | ( n1487 & n1985 ) | ( n1984 & n1985 ) ;
  assign n1988 = ( ~n1358 & n1986 ) | ( ~n1358 & n1987 ) | ( n1986 & n1987 ) ;
  assign n1989 = ( n1506 & n1986 ) | ( n1506 & n1987 ) | ( n1986 & n1987 ) ;
  assign n1990 = ( n1612 & n1988 ) | ( n1612 & n1989 ) | ( n1988 & n1989 ) ;
  assign n1991 = n1983 | n1990 ;
  assign n1992 = n1976 & ~n1991 ;
  assign n1993 = n1961 | n1992 ;
  assign n1994 = n1930 | n1993 ;
  assign n1995 = x247 & n1370 ;
  assign n1996 = x247 & ~n1373 ;
  assign n1997 = ( n1467 & n1995 ) | ( n1467 & n1996 ) | ( n1995 & n1996 ) ;
  assign n1998 = ( ~n1487 & n1995 ) | ( ~n1487 & n1996 ) | ( n1995 & n1996 ) ;
  assign n1999 = ( n1358 & n1997 ) | ( n1358 & n1998 ) | ( n1997 & n1998 ) ;
  assign n2000 = ( ~n1506 & n1997 ) | ( ~n1506 & n1998 ) | ( n1997 & n1998 ) ;
  assign n2001 = ( ~n1612 & n1999 ) | ( ~n1612 & n2000 ) | ( n1999 & n2000 ) ;
  assign n2002 = x119 & ~n1370 ;
  assign n2003 = x119 & n1373 ;
  assign n2004 = ( ~n1467 & n2002 ) | ( ~n1467 & n2003 ) | ( n2002 & n2003 ) ;
  assign n2005 = ( n1487 & n2002 ) | ( n1487 & n2003 ) | ( n2002 & n2003 ) ;
  assign n2006 = ( ~n1358 & n2004 ) | ( ~n1358 & n2005 ) | ( n2004 & n2005 ) ;
  assign n2007 = ( n1506 & n2004 ) | ( n1506 & n2005 ) | ( n2004 & n2005 ) ;
  assign n2008 = ( n1612 & n2006 ) | ( n1612 & n2007 ) | ( n2006 & n2007 ) ;
  assign n2009 = n2001 | n2008 ;
  assign n2010 = x503 & n812 ;
  assign n2011 = x503 & ~n815 ;
  assign n2012 = ( n909 & n2010 ) | ( n909 & n2011 ) | ( n2010 & n2011 ) ;
  assign n2013 = ( ~n929 & n2010 ) | ( ~n929 & n2011 ) | ( n2010 & n2011 ) ;
  assign n2014 = ( n800 & n2012 ) | ( n800 & n2013 ) | ( n2012 & n2013 ) ;
  assign n2015 = ( ~n948 & n2012 ) | ( ~n948 & n2013 ) | ( n2012 & n2013 ) ;
  assign n2016 = ( ~n1061 & n2014 ) | ( ~n1061 & n2015 ) | ( n2014 & n2015 ) ;
  assign n2017 = x375 & ~n812 ;
  assign n2018 = x375 & n815 ;
  assign n2019 = ( ~n909 & n2017 ) | ( ~n909 & n2018 ) | ( n2017 & n2018 ) ;
  assign n2020 = ( n929 & n2017 ) | ( n929 & n2018 ) | ( n2017 & n2018 ) ;
  assign n2021 = ( ~n800 & n2019 ) | ( ~n800 & n2020 ) | ( n2019 & n2020 ) ;
  assign n2022 = ( n948 & n2019 ) | ( n948 & n2020 ) | ( n2019 & n2020 ) ;
  assign n2023 = ( n1061 & n2021 ) | ( n1061 & n2022 ) | ( n2021 & n2022 ) ;
  assign n2024 = n2016 | n2023 ;
  assign n2025 = ~n2009 & n2024 ;
  assign n2026 = x502 & n812 ;
  assign n2027 = x502 & ~n815 ;
  assign n2028 = ( n909 & n2026 ) | ( n909 & n2027 ) | ( n2026 & n2027 ) ;
  assign n2029 = ( ~n929 & n2026 ) | ( ~n929 & n2027 ) | ( n2026 & n2027 ) ;
  assign n2030 = ( n800 & n2028 ) | ( n800 & n2029 ) | ( n2028 & n2029 ) ;
  assign n2031 = ( ~n948 & n2028 ) | ( ~n948 & n2029 ) | ( n2028 & n2029 ) ;
  assign n2032 = ( ~n1061 & n2030 ) | ( ~n1061 & n2031 ) | ( n2030 & n2031 ) ;
  assign n2033 = x374 & ~n812 ;
  assign n2034 = x374 & n815 ;
  assign n2035 = ( ~n909 & n2033 ) | ( ~n909 & n2034 ) | ( n2033 & n2034 ) ;
  assign n2036 = ( n929 & n2033 ) | ( n929 & n2034 ) | ( n2033 & n2034 ) ;
  assign n2037 = ( ~n800 & n2035 ) | ( ~n800 & n2036 ) | ( n2035 & n2036 ) ;
  assign n2038 = ( n948 & n2035 ) | ( n948 & n2036 ) | ( n2035 & n2036 ) ;
  assign n2039 = ( n1061 & n2037 ) | ( n1061 & n2038 ) | ( n2037 & n2038 ) ;
  assign n2040 = n2032 | n2039 ;
  assign n2041 = x246 & n1370 ;
  assign n2042 = x246 & ~n1373 ;
  assign n2043 = ( n1467 & n2041 ) | ( n1467 & n2042 ) | ( n2041 & n2042 ) ;
  assign n2044 = ( ~n1487 & n2041 ) | ( ~n1487 & n2042 ) | ( n2041 & n2042 ) ;
  assign n2045 = ( n1358 & n2043 ) | ( n1358 & n2044 ) | ( n2043 & n2044 ) ;
  assign n2046 = ( ~n1506 & n2043 ) | ( ~n1506 & n2044 ) | ( n2043 & n2044 ) ;
  assign n2047 = ( ~n1612 & n2045 ) | ( ~n1612 & n2046 ) | ( n2045 & n2046 ) ;
  assign n2048 = x118 & ~n1370 ;
  assign n2049 = x118 & n1373 ;
  assign n2050 = ( ~n1467 & n2048 ) | ( ~n1467 & n2049 ) | ( n2048 & n2049 ) ;
  assign n2051 = ( n1487 & n2048 ) | ( n1487 & n2049 ) | ( n2048 & n2049 ) ;
  assign n2052 = ( ~n1358 & n2050 ) | ( ~n1358 & n2051 ) | ( n2050 & n2051 ) ;
  assign n2053 = ( n1506 & n2050 ) | ( n1506 & n2051 ) | ( n2050 & n2051 ) ;
  assign n2054 = ( n1612 & n2052 ) | ( n1612 & n2053 ) | ( n2052 & n2053 ) ;
  assign n2055 = n2047 | n2054 ;
  assign n2056 = n2040 & ~n2055 ;
  assign n2057 = n2025 | n2056 ;
  assign n2058 = x245 & n1370 ;
  assign n2059 = x245 & ~n1373 ;
  assign n2060 = ( n1467 & n2058 ) | ( n1467 & n2059 ) | ( n2058 & n2059 ) ;
  assign n2061 = ( ~n1487 & n2058 ) | ( ~n1487 & n2059 ) | ( n2058 & n2059 ) ;
  assign n2062 = ( n1358 & n2060 ) | ( n1358 & n2061 ) | ( n2060 & n2061 ) ;
  assign n2063 = ( ~n1506 & n2060 ) | ( ~n1506 & n2061 ) | ( n2060 & n2061 ) ;
  assign n2064 = ( ~n1612 & n2062 ) | ( ~n1612 & n2063 ) | ( n2062 & n2063 ) ;
  assign n2065 = x117 & ~n1370 ;
  assign n2066 = x117 & n1373 ;
  assign n2067 = ( ~n1467 & n2065 ) | ( ~n1467 & n2066 ) | ( n2065 & n2066 ) ;
  assign n2068 = ( n1487 & n2065 ) | ( n1487 & n2066 ) | ( n2065 & n2066 ) ;
  assign n2069 = ( ~n1358 & n2067 ) | ( ~n1358 & n2068 ) | ( n2067 & n2068 ) ;
  assign n2070 = ( n1506 & n2067 ) | ( n1506 & n2068 ) | ( n2067 & n2068 ) ;
  assign n2071 = ( n1612 & n2069 ) | ( n1612 & n2070 ) | ( n2069 & n2070 ) ;
  assign n2072 = n2064 | n2071 ;
  assign n2073 = x501 & n812 ;
  assign n2074 = x501 & ~n815 ;
  assign n2075 = ( n909 & n2073 ) | ( n909 & n2074 ) | ( n2073 & n2074 ) ;
  assign n2076 = ( ~n929 & n2073 ) | ( ~n929 & n2074 ) | ( n2073 & n2074 ) ;
  assign n2077 = ( n800 & n2075 ) | ( n800 & n2076 ) | ( n2075 & n2076 ) ;
  assign n2078 = ( ~n948 & n2075 ) | ( ~n948 & n2076 ) | ( n2075 & n2076 ) ;
  assign n2079 = ( ~n1061 & n2077 ) | ( ~n1061 & n2078 ) | ( n2077 & n2078 ) ;
  assign n2080 = x373 & ~n812 ;
  assign n2081 = x373 & n815 ;
  assign n2082 = ( ~n909 & n2080 ) | ( ~n909 & n2081 ) | ( n2080 & n2081 ) ;
  assign n2083 = ( n929 & n2080 ) | ( n929 & n2081 ) | ( n2080 & n2081 ) ;
  assign n2084 = ( ~n800 & n2082 ) | ( ~n800 & n2083 ) | ( n2082 & n2083 ) ;
  assign n2085 = ( n948 & n2082 ) | ( n948 & n2083 ) | ( n2082 & n2083 ) ;
  assign n2086 = ( n1061 & n2084 ) | ( n1061 & n2085 ) | ( n2084 & n2085 ) ;
  assign n2087 = n2079 | n2086 ;
  assign n2088 = ~n2072 & n2087 ;
  assign n2089 = x244 & n1370 ;
  assign n2090 = x244 & ~n1373 ;
  assign n2091 = ( n1467 & n2089 ) | ( n1467 & n2090 ) | ( n2089 & n2090 ) ;
  assign n2092 = ( ~n1487 & n2089 ) | ( ~n1487 & n2090 ) | ( n2089 & n2090 ) ;
  assign n2093 = ( n1358 & n2091 ) | ( n1358 & n2092 ) | ( n2091 & n2092 ) ;
  assign n2094 = ( ~n1506 & n2091 ) | ( ~n1506 & n2092 ) | ( n2091 & n2092 ) ;
  assign n2095 = ( ~n1612 & n2093 ) | ( ~n1612 & n2094 ) | ( n2093 & n2094 ) ;
  assign n2096 = x116 & ~n1370 ;
  assign n2097 = x116 & n1373 ;
  assign n2098 = ( ~n1467 & n2096 ) | ( ~n1467 & n2097 ) | ( n2096 & n2097 ) ;
  assign n2099 = ( n1487 & n2096 ) | ( n1487 & n2097 ) | ( n2096 & n2097 ) ;
  assign n2100 = ( ~n1358 & n2098 ) | ( ~n1358 & n2099 ) | ( n2098 & n2099 ) ;
  assign n2101 = ( n1506 & n2098 ) | ( n1506 & n2099 ) | ( n2098 & n2099 ) ;
  assign n2102 = ( n1612 & n2100 ) | ( n1612 & n2101 ) | ( n2100 & n2101 ) ;
  assign n2103 = n2095 | n2102 ;
  assign n2104 = x500 & n812 ;
  assign n2105 = x500 & ~n815 ;
  assign n2106 = ( n909 & n2104 ) | ( n909 & n2105 ) | ( n2104 & n2105 ) ;
  assign n2107 = ( ~n929 & n2104 ) | ( ~n929 & n2105 ) | ( n2104 & n2105 ) ;
  assign n2108 = ( n800 & n2106 ) | ( n800 & n2107 ) | ( n2106 & n2107 ) ;
  assign n2109 = ( ~n948 & n2106 ) | ( ~n948 & n2107 ) | ( n2106 & n2107 ) ;
  assign n2110 = ( ~n1061 & n2108 ) | ( ~n1061 & n2109 ) | ( n2108 & n2109 ) ;
  assign n2111 = x372 & ~n812 ;
  assign n2112 = x372 & n815 ;
  assign n2113 = ( ~n909 & n2111 ) | ( ~n909 & n2112 ) | ( n2111 & n2112 ) ;
  assign n2114 = ( n929 & n2111 ) | ( n929 & n2112 ) | ( n2111 & n2112 ) ;
  assign n2115 = ( ~n800 & n2113 ) | ( ~n800 & n2114 ) | ( n2113 & n2114 ) ;
  assign n2116 = ( n948 & n2113 ) | ( n948 & n2114 ) | ( n2113 & n2114 ) ;
  assign n2117 = ( n1061 & n2115 ) | ( n1061 & n2116 ) | ( n2115 & n2116 ) ;
  assign n2118 = n2110 | n2117 ;
  assign n2119 = ~n2103 & n2118 ;
  assign n2120 = n2088 | n2119 ;
  assign n2121 = n2057 | n2120 ;
  assign n2122 = x243 & n1370 ;
  assign n2123 = x243 & ~n1373 ;
  assign n2124 = ( n1467 & n2122 ) | ( n1467 & n2123 ) | ( n2122 & n2123 ) ;
  assign n2125 = ( ~n1487 & n2122 ) | ( ~n1487 & n2123 ) | ( n2122 & n2123 ) ;
  assign n2126 = ( n1358 & n2124 ) | ( n1358 & n2125 ) | ( n2124 & n2125 ) ;
  assign n2127 = ( ~n1506 & n2124 ) | ( ~n1506 & n2125 ) | ( n2124 & n2125 ) ;
  assign n2128 = ( ~n1612 & n2126 ) | ( ~n1612 & n2127 ) | ( n2126 & n2127 ) ;
  assign n2129 = x115 & ~n1370 ;
  assign n2130 = x115 & n1373 ;
  assign n2131 = ( ~n1467 & n2129 ) | ( ~n1467 & n2130 ) | ( n2129 & n2130 ) ;
  assign n2132 = ( n1487 & n2129 ) | ( n1487 & n2130 ) | ( n2129 & n2130 ) ;
  assign n2133 = ( ~n1358 & n2131 ) | ( ~n1358 & n2132 ) | ( n2131 & n2132 ) ;
  assign n2134 = ( n1506 & n2131 ) | ( n1506 & n2132 ) | ( n2131 & n2132 ) ;
  assign n2135 = ( n1612 & n2133 ) | ( n1612 & n2134 ) | ( n2133 & n2134 ) ;
  assign n2136 = n2128 | n2135 ;
  assign n2137 = x499 & n812 ;
  assign n2138 = x499 & ~n815 ;
  assign n2139 = ( n909 & n2137 ) | ( n909 & n2138 ) | ( n2137 & n2138 ) ;
  assign n2140 = ( ~n929 & n2137 ) | ( ~n929 & n2138 ) | ( n2137 & n2138 ) ;
  assign n2141 = ( n800 & n2139 ) | ( n800 & n2140 ) | ( n2139 & n2140 ) ;
  assign n2142 = ( ~n948 & n2139 ) | ( ~n948 & n2140 ) | ( n2139 & n2140 ) ;
  assign n2143 = ( ~n1061 & n2141 ) | ( ~n1061 & n2142 ) | ( n2141 & n2142 ) ;
  assign n2144 = x371 & ~n812 ;
  assign n2145 = x371 & n815 ;
  assign n2146 = ( ~n909 & n2144 ) | ( ~n909 & n2145 ) | ( n2144 & n2145 ) ;
  assign n2147 = ( n929 & n2144 ) | ( n929 & n2145 ) | ( n2144 & n2145 ) ;
  assign n2148 = ( ~n800 & n2146 ) | ( ~n800 & n2147 ) | ( n2146 & n2147 ) ;
  assign n2149 = ( n948 & n2146 ) | ( n948 & n2147 ) | ( n2146 & n2147 ) ;
  assign n2150 = ( n1061 & n2148 ) | ( n1061 & n2149 ) | ( n2148 & n2149 ) ;
  assign n2151 = n2143 | n2150 ;
  assign n2152 = ~n2136 & n2151 ;
  assign n2153 = x498 & n812 ;
  assign n2154 = x498 & ~n815 ;
  assign n2155 = ( n909 & n2153 ) | ( n909 & n2154 ) | ( n2153 & n2154 ) ;
  assign n2156 = ( ~n929 & n2153 ) | ( ~n929 & n2154 ) | ( n2153 & n2154 ) ;
  assign n2157 = ( n800 & n2155 ) | ( n800 & n2156 ) | ( n2155 & n2156 ) ;
  assign n2158 = ( ~n948 & n2155 ) | ( ~n948 & n2156 ) | ( n2155 & n2156 ) ;
  assign n2159 = ( ~n1061 & n2157 ) | ( ~n1061 & n2158 ) | ( n2157 & n2158 ) ;
  assign n2160 = x370 & ~n812 ;
  assign n2161 = x370 & n815 ;
  assign n2162 = ( ~n909 & n2160 ) | ( ~n909 & n2161 ) | ( n2160 & n2161 ) ;
  assign n2163 = ( n929 & n2160 ) | ( n929 & n2161 ) | ( n2160 & n2161 ) ;
  assign n2164 = ( ~n800 & n2162 ) | ( ~n800 & n2163 ) | ( n2162 & n2163 ) ;
  assign n2165 = ( n948 & n2162 ) | ( n948 & n2163 ) | ( n2162 & n2163 ) ;
  assign n2166 = ( n1061 & n2164 ) | ( n1061 & n2165 ) | ( n2164 & n2165 ) ;
  assign n2167 = n2159 | n2166 ;
  assign n2168 = x242 & n1370 ;
  assign n2169 = x242 & ~n1373 ;
  assign n2170 = ( n1467 & n2168 ) | ( n1467 & n2169 ) | ( n2168 & n2169 ) ;
  assign n2171 = ( ~n1487 & n2168 ) | ( ~n1487 & n2169 ) | ( n2168 & n2169 ) ;
  assign n2172 = ( n1358 & n2170 ) | ( n1358 & n2171 ) | ( n2170 & n2171 ) ;
  assign n2173 = ( ~n1506 & n2170 ) | ( ~n1506 & n2171 ) | ( n2170 & n2171 ) ;
  assign n2174 = ( ~n1612 & n2172 ) | ( ~n1612 & n2173 ) | ( n2172 & n2173 ) ;
  assign n2175 = x114 & ~n1370 ;
  assign n2176 = x114 & n1373 ;
  assign n2177 = ( ~n1467 & n2175 ) | ( ~n1467 & n2176 ) | ( n2175 & n2176 ) ;
  assign n2178 = ( n1487 & n2175 ) | ( n1487 & n2176 ) | ( n2175 & n2176 ) ;
  assign n2179 = ( ~n1358 & n2177 ) | ( ~n1358 & n2178 ) | ( n2177 & n2178 ) ;
  assign n2180 = ( n1506 & n2177 ) | ( n1506 & n2178 ) | ( n2177 & n2178 ) ;
  assign n2181 = ( n1612 & n2179 ) | ( n1612 & n2180 ) | ( n2179 & n2180 ) ;
  assign n2182 = n2174 | n2181 ;
  assign n2183 = n2167 & ~n2182 ;
  assign n2184 = n2152 | n2183 ;
  assign n2185 = x241 & n1370 ;
  assign n2186 = x241 & ~n1373 ;
  assign n2187 = ( n1467 & n2185 ) | ( n1467 & n2186 ) | ( n2185 & n2186 ) ;
  assign n2188 = ( ~n1487 & n2185 ) | ( ~n1487 & n2186 ) | ( n2185 & n2186 ) ;
  assign n2189 = ( n1358 & n2187 ) | ( n1358 & n2188 ) | ( n2187 & n2188 ) ;
  assign n2190 = ( ~n1506 & n2187 ) | ( ~n1506 & n2188 ) | ( n2187 & n2188 ) ;
  assign n2191 = ( ~n1612 & n2189 ) | ( ~n1612 & n2190 ) | ( n2189 & n2190 ) ;
  assign n2192 = x113 & ~n1370 ;
  assign n2193 = x113 & n1373 ;
  assign n2194 = ( ~n1467 & n2192 ) | ( ~n1467 & n2193 ) | ( n2192 & n2193 ) ;
  assign n2195 = ( n1487 & n2192 ) | ( n1487 & n2193 ) | ( n2192 & n2193 ) ;
  assign n2196 = ( ~n1358 & n2194 ) | ( ~n1358 & n2195 ) | ( n2194 & n2195 ) ;
  assign n2197 = ( n1506 & n2194 ) | ( n1506 & n2195 ) | ( n2194 & n2195 ) ;
  assign n2198 = ( n1612 & n2196 ) | ( n1612 & n2197 ) | ( n2196 & n2197 ) ;
  assign n2199 = n2191 | n2198 ;
  assign n2200 = x497 & n812 ;
  assign n2201 = x497 & ~n815 ;
  assign n2202 = ( n909 & n2200 ) | ( n909 & n2201 ) | ( n2200 & n2201 ) ;
  assign n2203 = ( ~n929 & n2200 ) | ( ~n929 & n2201 ) | ( n2200 & n2201 ) ;
  assign n2204 = ( n800 & n2202 ) | ( n800 & n2203 ) | ( n2202 & n2203 ) ;
  assign n2205 = ( ~n948 & n2202 ) | ( ~n948 & n2203 ) | ( n2202 & n2203 ) ;
  assign n2206 = ( ~n1061 & n2204 ) | ( ~n1061 & n2205 ) | ( n2204 & n2205 ) ;
  assign n2207 = x369 & ~n812 ;
  assign n2208 = x369 & n815 ;
  assign n2209 = ( ~n909 & n2207 ) | ( ~n909 & n2208 ) | ( n2207 & n2208 ) ;
  assign n2210 = ( n929 & n2207 ) | ( n929 & n2208 ) | ( n2207 & n2208 ) ;
  assign n2211 = ( ~n800 & n2209 ) | ( ~n800 & n2210 ) | ( n2209 & n2210 ) ;
  assign n2212 = ( n948 & n2209 ) | ( n948 & n2210 ) | ( n2209 & n2210 ) ;
  assign n2213 = ( n1061 & n2211 ) | ( n1061 & n2212 ) | ( n2211 & n2212 ) ;
  assign n2214 = n2206 | n2213 ;
  assign n2215 = ~n2199 & n2214 ;
  assign n2216 = x496 & n812 ;
  assign n2217 = x496 & ~n815 ;
  assign n2218 = ( n909 & n2216 ) | ( n909 & n2217 ) | ( n2216 & n2217 ) ;
  assign n2219 = ( ~n929 & n2216 ) | ( ~n929 & n2217 ) | ( n2216 & n2217 ) ;
  assign n2220 = ( n800 & n2218 ) | ( n800 & n2219 ) | ( n2218 & n2219 ) ;
  assign n2221 = ( ~n948 & n2218 ) | ( ~n948 & n2219 ) | ( n2218 & n2219 ) ;
  assign n2222 = ( ~n1061 & n2220 ) | ( ~n1061 & n2221 ) | ( n2220 & n2221 ) ;
  assign n2223 = x368 & ~n812 ;
  assign n2224 = x368 & n815 ;
  assign n2225 = ( ~n909 & n2223 ) | ( ~n909 & n2224 ) | ( n2223 & n2224 ) ;
  assign n2226 = ( n929 & n2223 ) | ( n929 & n2224 ) | ( n2223 & n2224 ) ;
  assign n2227 = ( ~n800 & n2225 ) | ( ~n800 & n2226 ) | ( n2225 & n2226 ) ;
  assign n2228 = ( n948 & n2225 ) | ( n948 & n2226 ) | ( n2225 & n2226 ) ;
  assign n2229 = ( n1061 & n2227 ) | ( n1061 & n2228 ) | ( n2227 & n2228 ) ;
  assign n2230 = n2222 | n2229 ;
  assign n2231 = x240 & n1370 ;
  assign n2232 = x240 & ~n1373 ;
  assign n2233 = ( n1467 & n2231 ) | ( n1467 & n2232 ) | ( n2231 & n2232 ) ;
  assign n2234 = ( ~n1487 & n2231 ) | ( ~n1487 & n2232 ) | ( n2231 & n2232 ) ;
  assign n2235 = ( n1358 & n2233 ) | ( n1358 & n2234 ) | ( n2233 & n2234 ) ;
  assign n2236 = ( ~n1506 & n2233 ) | ( ~n1506 & n2234 ) | ( n2233 & n2234 ) ;
  assign n2237 = ( ~n1612 & n2235 ) | ( ~n1612 & n2236 ) | ( n2235 & n2236 ) ;
  assign n2238 = x112 & ~n1370 ;
  assign n2239 = x112 & n1373 ;
  assign n2240 = ( ~n1467 & n2238 ) | ( ~n1467 & n2239 ) | ( n2238 & n2239 ) ;
  assign n2241 = ( n1487 & n2238 ) | ( n1487 & n2239 ) | ( n2238 & n2239 ) ;
  assign n2242 = ( ~n1358 & n2240 ) | ( ~n1358 & n2241 ) | ( n2240 & n2241 ) ;
  assign n2243 = ( n1506 & n2240 ) | ( n1506 & n2241 ) | ( n2240 & n2241 ) ;
  assign n2244 = ( n1612 & n2242 ) | ( n1612 & n2243 ) | ( n2242 & n2243 ) ;
  assign n2245 = n2237 | n2244 ;
  assign n2246 = n2230 & ~n2245 ;
  assign n2247 = n2215 | n2246 ;
  assign n2248 = n2184 | n2247 ;
  assign n2249 = ~n2230 & n2245 ;
  assign n2250 = ( n2199 & ~n2214 ) | ( n2199 & n2249 ) | ( ~n2214 & n2249 ) ;
  assign n2251 = ( ~n2167 & n2182 ) | ( ~n2167 & n2250 ) | ( n2182 & n2250 ) ;
  assign n2252 = ( n2136 & ~n2151 ) | ( n2136 & n2251 ) | ( ~n2151 & n2251 ) ;
  assign n2253 = n2248 & ~n2252 ;
  assign n2254 = n2121 | n2253 ;
  assign n2255 = n2009 & ~n2024 ;
  assign n2256 = ~n2040 & n2055 ;
  assign n2257 = ~n2025 & n2256 ;
  assign n2258 = n2103 & ~n2118 ;
  assign n2259 = ( n2072 & ~n2087 ) | ( n2072 & n2258 ) | ( ~n2087 & n2258 ) ;
  assign n2260 = ~n2057 & n2259 ;
  assign n2261 = n2257 | n2260 ;
  assign n2262 = n2255 | n2261 ;
  assign n2263 = ~n1994 & n2262 ;
  assign n2264 = ( n1994 & n2254 ) | ( n1994 & ~n2263 ) | ( n2254 & ~n2263 ) ;
  assign n2265 = ~n2121 & n2252 ;
  assign n2266 = ( ~n1994 & n2263 ) | ( ~n1994 & n2265 ) | ( n2263 & n2265 ) ;
  assign n2267 = ( n1867 & ~n2264 ) | ( n1867 & n2266 ) | ( ~n2264 & n2266 ) ;
  assign n2268 = x254 & n1370 ;
  assign n2269 = x254 & ~n1373 ;
  assign n2270 = ( n1467 & n2268 ) | ( n1467 & n2269 ) | ( n2268 & n2269 ) ;
  assign n2271 = ( ~n1487 & n2268 ) | ( ~n1487 & n2269 ) | ( n2268 & n2269 ) ;
  assign n2272 = ( n1358 & n2270 ) | ( n1358 & n2271 ) | ( n2270 & n2271 ) ;
  assign n2273 = ( ~n1506 & n2270 ) | ( ~n1506 & n2271 ) | ( n2270 & n2271 ) ;
  assign n2274 = ( ~n1612 & n2272 ) | ( ~n1612 & n2273 ) | ( n2272 & n2273 ) ;
  assign n2275 = x126 & ~n1370 ;
  assign n2276 = x126 & n1373 ;
  assign n2277 = ( ~n1467 & n2275 ) | ( ~n1467 & n2276 ) | ( n2275 & n2276 ) ;
  assign n2278 = ( n1487 & n2275 ) | ( n1487 & n2276 ) | ( n2275 & n2276 ) ;
  assign n2279 = ( ~n1358 & n2277 ) | ( ~n1358 & n2278 ) | ( n2277 & n2278 ) ;
  assign n2280 = ( n1506 & n2277 ) | ( n1506 & n2278 ) | ( n2277 & n2278 ) ;
  assign n2281 = ( n1612 & n2279 ) | ( n1612 & n2280 ) | ( n2279 & n2280 ) ;
  assign n2282 = n2274 | n2281 ;
  assign n2283 = x510 & n812 ;
  assign n2284 = x510 & ~n815 ;
  assign n2285 = ( n909 & n2283 ) | ( n909 & n2284 ) | ( n2283 & n2284 ) ;
  assign n2286 = ( ~n929 & n2283 ) | ( ~n929 & n2284 ) | ( n2283 & n2284 ) ;
  assign n2287 = ( n800 & n2285 ) | ( n800 & n2286 ) | ( n2285 & n2286 ) ;
  assign n2288 = ( ~n948 & n2285 ) | ( ~n948 & n2286 ) | ( n2285 & n2286 ) ;
  assign n2289 = ( ~n1061 & n2287 ) | ( ~n1061 & n2288 ) | ( n2287 & n2288 ) ;
  assign n2290 = x382 & ~n812 ;
  assign n2291 = x382 & n815 ;
  assign n2292 = ( ~n909 & n2290 ) | ( ~n909 & n2291 ) | ( n2290 & n2291 ) ;
  assign n2293 = ( n929 & n2290 ) | ( n929 & n2291 ) | ( n2290 & n2291 ) ;
  assign n2294 = ( ~n800 & n2292 ) | ( ~n800 & n2293 ) | ( n2292 & n2293 ) ;
  assign n2295 = ( n948 & n2292 ) | ( n948 & n2293 ) | ( n2292 & n2293 ) ;
  assign n2296 = ( n1061 & n2294 ) | ( n1061 & n2295 ) | ( n2294 & n2295 ) ;
  assign n2297 = n2289 | n2296 ;
  assign n2298 = ~n2282 & n2297 ;
  assign n2299 = x253 & n1370 ;
  assign n2300 = x253 & ~n1373 ;
  assign n2301 = ( n1467 & n2299 ) | ( n1467 & n2300 ) | ( n2299 & n2300 ) ;
  assign n2302 = ( ~n1487 & n2299 ) | ( ~n1487 & n2300 ) | ( n2299 & n2300 ) ;
  assign n2303 = ( n1358 & n2301 ) | ( n1358 & n2302 ) | ( n2301 & n2302 ) ;
  assign n2304 = ( ~n1506 & n2301 ) | ( ~n1506 & n2302 ) | ( n2301 & n2302 ) ;
  assign n2305 = ( ~n1612 & n2303 ) | ( ~n1612 & n2304 ) | ( n2303 & n2304 ) ;
  assign n2306 = x125 & ~n1370 ;
  assign n2307 = x125 & n1373 ;
  assign n2308 = ( ~n1467 & n2306 ) | ( ~n1467 & n2307 ) | ( n2306 & n2307 ) ;
  assign n2309 = ( n1487 & n2306 ) | ( n1487 & n2307 ) | ( n2306 & n2307 ) ;
  assign n2310 = ( ~n1358 & n2308 ) | ( ~n1358 & n2309 ) | ( n2308 & n2309 ) ;
  assign n2311 = ( n1506 & n2308 ) | ( n1506 & n2309 ) | ( n2308 & n2309 ) ;
  assign n2312 = ( n1612 & n2310 ) | ( n1612 & n2311 ) | ( n2310 & n2311 ) ;
  assign n2313 = n2305 | n2312 ;
  assign n2314 = x509 & n812 ;
  assign n2315 = x509 & ~n815 ;
  assign n2316 = ( n909 & n2314 ) | ( n909 & n2315 ) | ( n2314 & n2315 ) ;
  assign n2317 = ( ~n929 & n2314 ) | ( ~n929 & n2315 ) | ( n2314 & n2315 ) ;
  assign n2318 = ( n800 & n2316 ) | ( n800 & n2317 ) | ( n2316 & n2317 ) ;
  assign n2319 = ( ~n948 & n2316 ) | ( ~n948 & n2317 ) | ( n2316 & n2317 ) ;
  assign n2320 = ( ~n1061 & n2318 ) | ( ~n1061 & n2319 ) | ( n2318 & n2319 ) ;
  assign n2321 = x381 & ~n812 ;
  assign n2322 = x381 & n815 ;
  assign n2323 = ( ~n909 & n2321 ) | ( ~n909 & n2322 ) | ( n2321 & n2322 ) ;
  assign n2324 = ( n929 & n2321 ) | ( n929 & n2322 ) | ( n2321 & n2322 ) ;
  assign n2325 = ( ~n800 & n2323 ) | ( ~n800 & n2324 ) | ( n2323 & n2324 ) ;
  assign n2326 = ( n948 & n2323 ) | ( n948 & n2324 ) | ( n2323 & n2324 ) ;
  assign n2327 = ( n1061 & n2325 ) | ( n1061 & n2326 ) | ( n2325 & n2326 ) ;
  assign n2328 = n2320 | n2327 ;
  assign n2329 = ~n2313 & n2328 ;
  assign n2330 = n2298 | n2329 ;
  assign n2331 = x252 & n1370 ;
  assign n2332 = x252 & ~n1373 ;
  assign n2333 = ( n1467 & n2331 ) | ( n1467 & n2332 ) | ( n2331 & n2332 ) ;
  assign n2334 = ( ~n1487 & n2331 ) | ( ~n1487 & n2332 ) | ( n2331 & n2332 ) ;
  assign n2335 = ( n1358 & n2333 ) | ( n1358 & n2334 ) | ( n2333 & n2334 ) ;
  assign n2336 = ( ~n1506 & n2333 ) | ( ~n1506 & n2334 ) | ( n2333 & n2334 ) ;
  assign n2337 = ( ~n1612 & n2335 ) | ( ~n1612 & n2336 ) | ( n2335 & n2336 ) ;
  assign n2338 = x124 & ~n1370 ;
  assign n2339 = x124 & n1373 ;
  assign n2340 = ( ~n1467 & n2338 ) | ( ~n1467 & n2339 ) | ( n2338 & n2339 ) ;
  assign n2341 = ( n1487 & n2338 ) | ( n1487 & n2339 ) | ( n2338 & n2339 ) ;
  assign n2342 = ( ~n1358 & n2340 ) | ( ~n1358 & n2341 ) | ( n2340 & n2341 ) ;
  assign n2343 = ( n1506 & n2340 ) | ( n1506 & n2341 ) | ( n2340 & n2341 ) ;
  assign n2344 = ( n1612 & n2342 ) | ( n1612 & n2343 ) | ( n2342 & n2343 ) ;
  assign n2345 = n2337 | n2344 ;
  assign n2346 = x508 & n812 ;
  assign n2347 = x508 & ~n815 ;
  assign n2348 = ( n909 & n2346 ) | ( n909 & n2347 ) | ( n2346 & n2347 ) ;
  assign n2349 = ( ~n929 & n2346 ) | ( ~n929 & n2347 ) | ( n2346 & n2347 ) ;
  assign n2350 = ( n800 & n2348 ) | ( n800 & n2349 ) | ( n2348 & n2349 ) ;
  assign n2351 = ( ~n948 & n2348 ) | ( ~n948 & n2349 ) | ( n2348 & n2349 ) ;
  assign n2352 = ( ~n1061 & n2350 ) | ( ~n1061 & n2351 ) | ( n2350 & n2351 ) ;
  assign n2353 = x380 & ~n812 ;
  assign n2354 = x380 & n815 ;
  assign n2355 = ( ~n909 & n2353 ) | ( ~n909 & n2354 ) | ( n2353 & n2354 ) ;
  assign n2356 = ( n929 & n2353 ) | ( n929 & n2354 ) | ( n2353 & n2354 ) ;
  assign n2357 = ( ~n800 & n2355 ) | ( ~n800 & n2356 ) | ( n2355 & n2356 ) ;
  assign n2358 = ( n948 & n2355 ) | ( n948 & n2356 ) | ( n2355 & n2356 ) ;
  assign n2359 = ( n1061 & n2357 ) | ( n1061 & n2358 ) | ( n2357 & n2358 ) ;
  assign n2360 = n2352 | n2359 ;
  assign n2361 = ~n2345 & n2360 ;
  assign n2362 = x383 & x511 ;
  assign n2363 = x127 & x255 ;
  assign n2364 = ~n2362 & n2363 ;
  assign n2365 = n2361 | n2364 ;
  assign n2366 = n2330 | n2365 ;
  assign n2367 = ~n1976 & n1991 ;
  assign n2368 = ( n1945 & ~n1960 ) | ( n1945 & n2367 ) | ( ~n1960 & n2367 ) ;
  assign n2369 = ( ~n1913 & n1928 ) | ( ~n1913 & n2368 ) | ( n1928 & n2368 ) ;
  assign n2370 = ( n1882 & ~n1897 ) | ( n1882 & n2369 ) | ( ~n1897 & n2369 ) ;
  assign n2371 = ~n2366 & n2370 ;
  assign n2372 = n2362 & ~n2363 ;
  assign n2373 = n2345 & ~n2360 ;
  assign n2374 = ( n2313 & ~n2328 ) | ( n2313 & n2373 ) | ( ~n2328 & n2373 ) ;
  assign n2375 = ( n2282 & ~n2297 ) | ( n2282 & n2374 ) | ( ~n2297 & n2374 ) ;
  assign n2376 = ~n2364 & n2375 ;
  assign n2377 = n2372 | n2376 ;
  assign n2378 = n2371 | n2377 ;
  assign n2379 = n2366 & ~n2377 ;
  assign n2380 = ( n2267 & n2378 ) | ( n2267 & ~n2379 ) | ( n2378 & ~n2379 ) ;
  assign n2381 = n1994 | n2366 ;
  assign n2382 = ( n2366 & ~n2370 ) | ( n2366 & n2381 ) | ( ~n2370 & n2381 ) ;
  assign n2383 = ~n2376 & n2382 ;
  assign n2384 = ~n2372 & n2383 ;
  assign n2385 = n1736 & ~n1865 ;
  assign n2386 = n1862 & ~n2215 ;
  assign n2387 = ~n2184 & n2386 ;
  assign n2388 = ~n2246 & n2387 ;
  assign n2389 = ( n2248 & n2385 ) | ( n2248 & ~n2388 ) | ( n2385 & ~n2388 ) ;
  assign n2390 = ~n2252 & n2389 ;
  assign n2391 = n2121 & ~n2261 ;
  assign n2392 = ( ~n2261 & n2390 ) | ( ~n2261 & n2391 ) | ( n2390 & n2391 ) ;
  assign n2393 = ~n2255 & n2392 ;
  assign n2394 = ( ~n2378 & n2384 ) | ( ~n2378 & n2393 ) | ( n2384 & n2393 ) ;
  assign n2395 = x183 & n1370 ;
  assign n2396 = x183 & ~n1373 ;
  assign n2397 = ( n1467 & n2395 ) | ( n1467 & n2396 ) | ( n2395 & n2396 ) ;
  assign n2398 = ( ~n1487 & n2395 ) | ( ~n1487 & n2396 ) | ( n2395 & n2396 ) ;
  assign n2399 = ( n1358 & n2397 ) | ( n1358 & n2398 ) | ( n2397 & n2398 ) ;
  assign n2400 = ( ~n1506 & n2397 ) | ( ~n1506 & n2398 ) | ( n2397 & n2398 ) ;
  assign n2401 = ( ~n1612 & n2399 ) | ( ~n1612 & n2400 ) | ( n2399 & n2400 ) ;
  assign n2402 = x55 & ~n1370 ;
  assign n2403 = x55 & n1373 ;
  assign n2404 = ( ~n1467 & n2402 ) | ( ~n1467 & n2403 ) | ( n2402 & n2403 ) ;
  assign n2405 = ( n1487 & n2402 ) | ( n1487 & n2403 ) | ( n2402 & n2403 ) ;
  assign n2406 = ( ~n1358 & n2404 ) | ( ~n1358 & n2405 ) | ( n2404 & n2405 ) ;
  assign n2407 = ( n1506 & n2404 ) | ( n1506 & n2405 ) | ( n2404 & n2405 ) ;
  assign n2408 = ( n1612 & n2406 ) | ( n1612 & n2407 ) | ( n2406 & n2407 ) ;
  assign n2409 = n2401 | n2408 ;
  assign n2410 = x439 & n812 ;
  assign n2411 = x439 & ~n815 ;
  assign n2412 = ( n909 & n2410 ) | ( n909 & n2411 ) | ( n2410 & n2411 ) ;
  assign n2413 = ( ~n929 & n2410 ) | ( ~n929 & n2411 ) | ( n2410 & n2411 ) ;
  assign n2414 = ( n800 & n2412 ) | ( n800 & n2413 ) | ( n2412 & n2413 ) ;
  assign n2415 = ( ~n948 & n2412 ) | ( ~n948 & n2413 ) | ( n2412 & n2413 ) ;
  assign n2416 = ( ~n1061 & n2414 ) | ( ~n1061 & n2415 ) | ( n2414 & n2415 ) ;
  assign n2417 = x311 & ~n812 ;
  assign n2418 = x311 & n815 ;
  assign n2419 = ( ~n909 & n2417 ) | ( ~n909 & n2418 ) | ( n2417 & n2418 ) ;
  assign n2420 = ( n929 & n2417 ) | ( n929 & n2418 ) | ( n2417 & n2418 ) ;
  assign n2421 = ( ~n800 & n2419 ) | ( ~n800 & n2420 ) | ( n2419 & n2420 ) ;
  assign n2422 = ( n948 & n2419 ) | ( n948 & n2420 ) | ( n2419 & n2420 ) ;
  assign n2423 = ( n1061 & n2421 ) | ( n1061 & n2422 ) | ( n2421 & n2422 ) ;
  assign n2424 = n2416 | n2423 ;
  assign n2425 = ~n2409 & n2424 ;
  assign n2426 = x438 & n812 ;
  assign n2427 = x438 & ~n815 ;
  assign n2428 = ( n909 & n2426 ) | ( n909 & n2427 ) | ( n2426 & n2427 ) ;
  assign n2429 = ( ~n929 & n2426 ) | ( ~n929 & n2427 ) | ( n2426 & n2427 ) ;
  assign n2430 = ( n800 & n2428 ) | ( n800 & n2429 ) | ( n2428 & n2429 ) ;
  assign n2431 = ( ~n948 & n2428 ) | ( ~n948 & n2429 ) | ( n2428 & n2429 ) ;
  assign n2432 = ( ~n1061 & n2430 ) | ( ~n1061 & n2431 ) | ( n2430 & n2431 ) ;
  assign n2433 = x310 & ~n812 ;
  assign n2434 = x310 & n815 ;
  assign n2435 = ( ~n909 & n2433 ) | ( ~n909 & n2434 ) | ( n2433 & n2434 ) ;
  assign n2436 = ( n929 & n2433 ) | ( n929 & n2434 ) | ( n2433 & n2434 ) ;
  assign n2437 = ( ~n800 & n2435 ) | ( ~n800 & n2436 ) | ( n2435 & n2436 ) ;
  assign n2438 = ( n948 & n2435 ) | ( n948 & n2436 ) | ( n2435 & n2436 ) ;
  assign n2439 = ( n1061 & n2437 ) | ( n1061 & n2438 ) | ( n2437 & n2438 ) ;
  assign n2440 = n2432 | n2439 ;
  assign n2441 = x182 & n1370 ;
  assign n2442 = x182 & ~n1373 ;
  assign n2443 = ( n1467 & n2441 ) | ( n1467 & n2442 ) | ( n2441 & n2442 ) ;
  assign n2444 = ( ~n1487 & n2441 ) | ( ~n1487 & n2442 ) | ( n2441 & n2442 ) ;
  assign n2445 = ( n1358 & n2443 ) | ( n1358 & n2444 ) | ( n2443 & n2444 ) ;
  assign n2446 = ( ~n1506 & n2443 ) | ( ~n1506 & n2444 ) | ( n2443 & n2444 ) ;
  assign n2447 = ( ~n1612 & n2445 ) | ( ~n1612 & n2446 ) | ( n2445 & n2446 ) ;
  assign n2448 = x54 & ~n1370 ;
  assign n2449 = x54 & n1373 ;
  assign n2450 = ( ~n1467 & n2448 ) | ( ~n1467 & n2449 ) | ( n2448 & n2449 ) ;
  assign n2451 = ( n1487 & n2448 ) | ( n1487 & n2449 ) | ( n2448 & n2449 ) ;
  assign n2452 = ( ~n1358 & n2450 ) | ( ~n1358 & n2451 ) | ( n2450 & n2451 ) ;
  assign n2453 = ( n1506 & n2450 ) | ( n1506 & n2451 ) | ( n2450 & n2451 ) ;
  assign n2454 = ( n1612 & n2452 ) | ( n1612 & n2453 ) | ( n2452 & n2453 ) ;
  assign n2455 = n2447 | n2454 ;
  assign n2456 = n2440 & ~n2455 ;
  assign n2457 = n2425 | n2456 ;
  assign n2458 = x181 & n1370 ;
  assign n2459 = x181 & ~n1373 ;
  assign n2460 = ( n1467 & n2458 ) | ( n1467 & n2459 ) | ( n2458 & n2459 ) ;
  assign n2461 = ( ~n1487 & n2458 ) | ( ~n1487 & n2459 ) | ( n2458 & n2459 ) ;
  assign n2462 = ( n1358 & n2460 ) | ( n1358 & n2461 ) | ( n2460 & n2461 ) ;
  assign n2463 = ( ~n1506 & n2460 ) | ( ~n1506 & n2461 ) | ( n2460 & n2461 ) ;
  assign n2464 = ( ~n1612 & n2462 ) | ( ~n1612 & n2463 ) | ( n2462 & n2463 ) ;
  assign n2465 = x53 & ~n1370 ;
  assign n2466 = x53 & n1373 ;
  assign n2467 = ( ~n1467 & n2465 ) | ( ~n1467 & n2466 ) | ( n2465 & n2466 ) ;
  assign n2468 = ( n1487 & n2465 ) | ( n1487 & n2466 ) | ( n2465 & n2466 ) ;
  assign n2469 = ( ~n1358 & n2467 ) | ( ~n1358 & n2468 ) | ( n2467 & n2468 ) ;
  assign n2470 = ( n1506 & n2467 ) | ( n1506 & n2468 ) | ( n2467 & n2468 ) ;
  assign n2471 = ( n1612 & n2469 ) | ( n1612 & n2470 ) | ( n2469 & n2470 ) ;
  assign n2472 = n2464 | n2471 ;
  assign n2473 = x437 & n812 ;
  assign n2474 = x437 & ~n815 ;
  assign n2475 = ( n909 & n2473 ) | ( n909 & n2474 ) | ( n2473 & n2474 ) ;
  assign n2476 = ( ~n929 & n2473 ) | ( ~n929 & n2474 ) | ( n2473 & n2474 ) ;
  assign n2477 = ( n800 & n2475 ) | ( n800 & n2476 ) | ( n2475 & n2476 ) ;
  assign n2478 = ( ~n948 & n2475 ) | ( ~n948 & n2476 ) | ( n2475 & n2476 ) ;
  assign n2479 = ( ~n1061 & n2477 ) | ( ~n1061 & n2478 ) | ( n2477 & n2478 ) ;
  assign n2480 = x309 & ~n812 ;
  assign n2481 = x309 & n815 ;
  assign n2482 = ( ~n909 & n2480 ) | ( ~n909 & n2481 ) | ( n2480 & n2481 ) ;
  assign n2483 = ( n929 & n2480 ) | ( n929 & n2481 ) | ( n2480 & n2481 ) ;
  assign n2484 = ( ~n800 & n2482 ) | ( ~n800 & n2483 ) | ( n2482 & n2483 ) ;
  assign n2485 = ( n948 & n2482 ) | ( n948 & n2483 ) | ( n2482 & n2483 ) ;
  assign n2486 = ( n1061 & n2484 ) | ( n1061 & n2485 ) | ( n2484 & n2485 ) ;
  assign n2487 = n2479 | n2486 ;
  assign n2488 = ~n2472 & n2487 ;
  assign n2489 = x436 & n812 ;
  assign n2490 = x436 & ~n815 ;
  assign n2491 = ( n909 & n2489 ) | ( n909 & n2490 ) | ( n2489 & n2490 ) ;
  assign n2492 = ( ~n929 & n2489 ) | ( ~n929 & n2490 ) | ( n2489 & n2490 ) ;
  assign n2493 = ( n800 & n2491 ) | ( n800 & n2492 ) | ( n2491 & n2492 ) ;
  assign n2494 = ( ~n948 & n2491 ) | ( ~n948 & n2492 ) | ( n2491 & n2492 ) ;
  assign n2495 = ( ~n1061 & n2493 ) | ( ~n1061 & n2494 ) | ( n2493 & n2494 ) ;
  assign n2496 = x308 & ~n812 ;
  assign n2497 = x308 & n815 ;
  assign n2498 = ( ~n909 & n2496 ) | ( ~n909 & n2497 ) | ( n2496 & n2497 ) ;
  assign n2499 = ( n929 & n2496 ) | ( n929 & n2497 ) | ( n2496 & n2497 ) ;
  assign n2500 = ( ~n800 & n2498 ) | ( ~n800 & n2499 ) | ( n2498 & n2499 ) ;
  assign n2501 = ( n948 & n2498 ) | ( n948 & n2499 ) | ( n2498 & n2499 ) ;
  assign n2502 = ( n1061 & n2500 ) | ( n1061 & n2501 ) | ( n2500 & n2501 ) ;
  assign n2503 = n2495 | n2502 ;
  assign n2504 = x180 & n1370 ;
  assign n2505 = x180 & ~n1373 ;
  assign n2506 = ( n1467 & n2504 ) | ( n1467 & n2505 ) | ( n2504 & n2505 ) ;
  assign n2507 = ( ~n1487 & n2504 ) | ( ~n1487 & n2505 ) | ( n2504 & n2505 ) ;
  assign n2508 = ( n1358 & n2506 ) | ( n1358 & n2507 ) | ( n2506 & n2507 ) ;
  assign n2509 = ( ~n1506 & n2506 ) | ( ~n1506 & n2507 ) | ( n2506 & n2507 ) ;
  assign n2510 = ( ~n1612 & n2508 ) | ( ~n1612 & n2509 ) | ( n2508 & n2509 ) ;
  assign n2511 = x52 & ~n1370 ;
  assign n2512 = x52 & n1373 ;
  assign n2513 = ( ~n1467 & n2511 ) | ( ~n1467 & n2512 ) | ( n2511 & n2512 ) ;
  assign n2514 = ( n1487 & n2511 ) | ( n1487 & n2512 ) | ( n2511 & n2512 ) ;
  assign n2515 = ( ~n1358 & n2513 ) | ( ~n1358 & n2514 ) | ( n2513 & n2514 ) ;
  assign n2516 = ( n1506 & n2513 ) | ( n1506 & n2514 ) | ( n2513 & n2514 ) ;
  assign n2517 = ( n1612 & n2515 ) | ( n1612 & n2516 ) | ( n2515 & n2516 ) ;
  assign n2518 = n2510 | n2517 ;
  assign n2519 = n2503 & ~n2518 ;
  assign n2520 = n2488 | n2519 ;
  assign n2521 = n2457 | n2520 ;
  assign n2522 = x177 & n1370 ;
  assign n2523 = x177 & ~n1373 ;
  assign n2524 = ( n1467 & n2522 ) | ( n1467 & n2523 ) | ( n2522 & n2523 ) ;
  assign n2525 = ( ~n1487 & n2522 ) | ( ~n1487 & n2523 ) | ( n2522 & n2523 ) ;
  assign n2526 = ( n1358 & n2524 ) | ( n1358 & n2525 ) | ( n2524 & n2525 ) ;
  assign n2527 = ( ~n1506 & n2524 ) | ( ~n1506 & n2525 ) | ( n2524 & n2525 ) ;
  assign n2528 = ( ~n1612 & n2526 ) | ( ~n1612 & n2527 ) | ( n2526 & n2527 ) ;
  assign n2529 = x49 & ~n1370 ;
  assign n2530 = x49 & n1373 ;
  assign n2531 = ( ~n1467 & n2529 ) | ( ~n1467 & n2530 ) | ( n2529 & n2530 ) ;
  assign n2532 = ( n1487 & n2529 ) | ( n1487 & n2530 ) | ( n2529 & n2530 ) ;
  assign n2533 = ( ~n1358 & n2531 ) | ( ~n1358 & n2532 ) | ( n2531 & n2532 ) ;
  assign n2534 = ( n1506 & n2531 ) | ( n1506 & n2532 ) | ( n2531 & n2532 ) ;
  assign n2535 = ( n1612 & n2533 ) | ( n1612 & n2534 ) | ( n2533 & n2534 ) ;
  assign n2536 = n2528 | n2535 ;
  assign n2537 = x433 & n812 ;
  assign n2538 = x433 & ~n815 ;
  assign n2539 = ( n909 & n2537 ) | ( n909 & n2538 ) | ( n2537 & n2538 ) ;
  assign n2540 = ( ~n929 & n2537 ) | ( ~n929 & n2538 ) | ( n2537 & n2538 ) ;
  assign n2541 = ( n800 & n2539 ) | ( n800 & n2540 ) | ( n2539 & n2540 ) ;
  assign n2542 = ( ~n948 & n2539 ) | ( ~n948 & n2540 ) | ( n2539 & n2540 ) ;
  assign n2543 = ( ~n1061 & n2541 ) | ( ~n1061 & n2542 ) | ( n2541 & n2542 ) ;
  assign n2544 = x305 & ~n812 ;
  assign n2545 = x305 & n815 ;
  assign n2546 = ( ~n909 & n2544 ) | ( ~n909 & n2545 ) | ( n2544 & n2545 ) ;
  assign n2547 = ( n929 & n2544 ) | ( n929 & n2545 ) | ( n2544 & n2545 ) ;
  assign n2548 = ( ~n800 & n2546 ) | ( ~n800 & n2547 ) | ( n2546 & n2547 ) ;
  assign n2549 = ( n948 & n2546 ) | ( n948 & n2547 ) | ( n2546 & n2547 ) ;
  assign n2550 = ( n1061 & n2548 ) | ( n1061 & n2549 ) | ( n2548 & n2549 ) ;
  assign n2551 = n2543 | n2550 ;
  assign n2552 = ~n2536 & n2551 ;
  assign n2553 = x179 & n1370 ;
  assign n2554 = x179 & ~n1373 ;
  assign n2555 = ( n1467 & n2553 ) | ( n1467 & n2554 ) | ( n2553 & n2554 ) ;
  assign n2556 = ( ~n1487 & n2553 ) | ( ~n1487 & n2554 ) | ( n2553 & n2554 ) ;
  assign n2557 = ( n1358 & n2555 ) | ( n1358 & n2556 ) | ( n2555 & n2556 ) ;
  assign n2558 = ( ~n1506 & n2555 ) | ( ~n1506 & n2556 ) | ( n2555 & n2556 ) ;
  assign n2559 = ( ~n1612 & n2557 ) | ( ~n1612 & n2558 ) | ( n2557 & n2558 ) ;
  assign n2560 = x51 & ~n1370 ;
  assign n2561 = x51 & n1373 ;
  assign n2562 = ( ~n1467 & n2560 ) | ( ~n1467 & n2561 ) | ( n2560 & n2561 ) ;
  assign n2563 = ( n1487 & n2560 ) | ( n1487 & n2561 ) | ( n2560 & n2561 ) ;
  assign n2564 = ( ~n1358 & n2562 ) | ( ~n1358 & n2563 ) | ( n2562 & n2563 ) ;
  assign n2565 = ( n1506 & n2562 ) | ( n1506 & n2563 ) | ( n2562 & n2563 ) ;
  assign n2566 = ( n1612 & n2564 ) | ( n1612 & n2565 ) | ( n2564 & n2565 ) ;
  assign n2567 = n2559 | n2566 ;
  assign n2568 = x435 & n812 ;
  assign n2569 = x435 & ~n815 ;
  assign n2570 = ( n909 & n2568 ) | ( n909 & n2569 ) | ( n2568 & n2569 ) ;
  assign n2571 = ( ~n929 & n2568 ) | ( ~n929 & n2569 ) | ( n2568 & n2569 ) ;
  assign n2572 = ( n800 & n2570 ) | ( n800 & n2571 ) | ( n2570 & n2571 ) ;
  assign n2573 = ( ~n948 & n2570 ) | ( ~n948 & n2571 ) | ( n2570 & n2571 ) ;
  assign n2574 = ( ~n1061 & n2572 ) | ( ~n1061 & n2573 ) | ( n2572 & n2573 ) ;
  assign n2575 = x307 & ~n812 ;
  assign n2576 = x307 & n815 ;
  assign n2577 = ( ~n909 & n2575 ) | ( ~n909 & n2576 ) | ( n2575 & n2576 ) ;
  assign n2578 = ( n929 & n2575 ) | ( n929 & n2576 ) | ( n2575 & n2576 ) ;
  assign n2579 = ( ~n800 & n2577 ) | ( ~n800 & n2578 ) | ( n2577 & n2578 ) ;
  assign n2580 = ( n948 & n2577 ) | ( n948 & n2578 ) | ( n2577 & n2578 ) ;
  assign n2581 = ( n1061 & n2579 ) | ( n1061 & n2580 ) | ( n2579 & n2580 ) ;
  assign n2582 = n2574 | n2581 ;
  assign n2583 = ~n2567 & n2582 ;
  assign n2584 = x434 & n812 ;
  assign n2585 = x434 & ~n815 ;
  assign n2586 = ( n909 & n2584 ) | ( n909 & n2585 ) | ( n2584 & n2585 ) ;
  assign n2587 = ( ~n929 & n2584 ) | ( ~n929 & n2585 ) | ( n2584 & n2585 ) ;
  assign n2588 = ( n800 & n2586 ) | ( n800 & n2587 ) | ( n2586 & n2587 ) ;
  assign n2589 = ( ~n948 & n2586 ) | ( ~n948 & n2587 ) | ( n2586 & n2587 ) ;
  assign n2590 = ( ~n1061 & n2588 ) | ( ~n1061 & n2589 ) | ( n2588 & n2589 ) ;
  assign n2591 = x306 & ~n812 ;
  assign n2592 = x306 & n815 ;
  assign n2593 = ( ~n909 & n2591 ) | ( ~n909 & n2592 ) | ( n2591 & n2592 ) ;
  assign n2594 = ( n929 & n2591 ) | ( n929 & n2592 ) | ( n2591 & n2592 ) ;
  assign n2595 = ( ~n800 & n2593 ) | ( ~n800 & n2594 ) | ( n2593 & n2594 ) ;
  assign n2596 = ( n948 & n2593 ) | ( n948 & n2594 ) | ( n2593 & n2594 ) ;
  assign n2597 = ( n1061 & n2595 ) | ( n1061 & n2596 ) | ( n2595 & n2596 ) ;
  assign n2598 = n2590 | n2597 ;
  assign n2599 = x178 & n1370 ;
  assign n2600 = x178 & ~n1373 ;
  assign n2601 = ( n1467 & n2599 ) | ( n1467 & n2600 ) | ( n2599 & n2600 ) ;
  assign n2602 = ( ~n1487 & n2599 ) | ( ~n1487 & n2600 ) | ( n2599 & n2600 ) ;
  assign n2603 = ( n1358 & n2601 ) | ( n1358 & n2602 ) | ( n2601 & n2602 ) ;
  assign n2604 = ( ~n1506 & n2601 ) | ( ~n1506 & n2602 ) | ( n2601 & n2602 ) ;
  assign n2605 = ( ~n1612 & n2603 ) | ( ~n1612 & n2604 ) | ( n2603 & n2604 ) ;
  assign n2606 = x50 & ~n1370 ;
  assign n2607 = x50 & n1373 ;
  assign n2608 = ( ~n1467 & n2606 ) | ( ~n1467 & n2607 ) | ( n2606 & n2607 ) ;
  assign n2609 = ( n1487 & n2606 ) | ( n1487 & n2607 ) | ( n2606 & n2607 ) ;
  assign n2610 = ( ~n1358 & n2608 ) | ( ~n1358 & n2609 ) | ( n2608 & n2609 ) ;
  assign n2611 = ( n1506 & n2608 ) | ( n1506 & n2609 ) | ( n2608 & n2609 ) ;
  assign n2612 = ( n1612 & n2610 ) | ( n1612 & n2611 ) | ( n2610 & n2611 ) ;
  assign n2613 = n2605 | n2612 ;
  assign n2614 = n2598 & ~n2613 ;
  assign n2615 = n2583 | n2614 ;
  assign n2616 = n2552 | n2615 ;
  assign n2617 = ~n2598 & n2613 ;
  assign n2618 = ~n2583 & n2617 ;
  assign n2619 = x432 & n812 ;
  assign n2620 = x432 & ~n815 ;
  assign n2621 = ( n909 & n2619 ) | ( n909 & n2620 ) | ( n2619 & n2620 ) ;
  assign n2622 = ( ~n929 & n2619 ) | ( ~n929 & n2620 ) | ( n2619 & n2620 ) ;
  assign n2623 = ( n800 & n2621 ) | ( n800 & n2622 ) | ( n2621 & n2622 ) ;
  assign n2624 = ( ~n948 & n2621 ) | ( ~n948 & n2622 ) | ( n2621 & n2622 ) ;
  assign n2625 = ( ~n1061 & n2623 ) | ( ~n1061 & n2624 ) | ( n2623 & n2624 ) ;
  assign n2626 = x304 & ~n812 ;
  assign n2627 = x304 & n815 ;
  assign n2628 = ( ~n909 & n2626 ) | ( ~n909 & n2627 ) | ( n2626 & n2627 ) ;
  assign n2629 = ( n929 & n2626 ) | ( n929 & n2627 ) | ( n2626 & n2627 ) ;
  assign n2630 = ( ~n800 & n2628 ) | ( ~n800 & n2629 ) | ( n2628 & n2629 ) ;
  assign n2631 = ( n948 & n2628 ) | ( n948 & n2629 ) | ( n2628 & n2629 ) ;
  assign n2632 = ( n1061 & n2630 ) | ( n1061 & n2631 ) | ( n2630 & n2631 ) ;
  assign n2633 = n2625 | n2632 ;
  assign n2634 = x176 & n1370 ;
  assign n2635 = x176 & ~n1373 ;
  assign n2636 = ( n1467 & n2634 ) | ( n1467 & n2635 ) | ( n2634 & n2635 ) ;
  assign n2637 = ( ~n1487 & n2634 ) | ( ~n1487 & n2635 ) | ( n2634 & n2635 ) ;
  assign n2638 = ( n1358 & n2636 ) | ( n1358 & n2637 ) | ( n2636 & n2637 ) ;
  assign n2639 = ( ~n1506 & n2636 ) | ( ~n1506 & n2637 ) | ( n2636 & n2637 ) ;
  assign n2640 = ( ~n1612 & n2638 ) | ( ~n1612 & n2639 ) | ( n2638 & n2639 ) ;
  assign n2641 = x48 & ~n1370 ;
  assign n2642 = x48 & n1373 ;
  assign n2643 = ( ~n1467 & n2641 ) | ( ~n1467 & n2642 ) | ( n2641 & n2642 ) ;
  assign n2644 = ( n1487 & n2641 ) | ( n1487 & n2642 ) | ( n2641 & n2642 ) ;
  assign n2645 = ( ~n1358 & n2643 ) | ( ~n1358 & n2644 ) | ( n2643 & n2644 ) ;
  assign n2646 = ( n1506 & n2643 ) | ( n1506 & n2644 ) | ( n2643 & n2644 ) ;
  assign n2647 = ( n1612 & n2645 ) | ( n1612 & n2646 ) | ( n2645 & n2646 ) ;
  assign n2648 = n2640 | n2647 ;
  assign n2649 = ~n2633 & n2648 ;
  assign n2650 = n2536 & ~n2551 ;
  assign n2651 = n2649 | n2650 ;
  assign n2652 = n2618 | n2651 ;
  assign n2653 = ( ~n2616 & n2618 ) | ( ~n2616 & n2652 ) | ( n2618 & n2652 ) ;
  assign n2654 = n2567 & ~n2582 ;
  assign n2655 = ~n2521 & n2654 ;
  assign n2656 = ( ~n2521 & n2653 ) | ( ~n2521 & n2655 ) | ( n2653 & n2655 ) ;
  assign n2657 = ~n2503 & n2518 ;
  assign n2658 = ( n2472 & ~n2487 ) | ( n2472 & n2657 ) | ( ~n2487 & n2657 ) ;
  assign n2659 = ( ~n2440 & n2455 ) | ( ~n2440 & n2658 ) | ( n2455 & n2658 ) ;
  assign n2660 = ( n2409 & ~n2424 ) | ( n2409 & n2659 ) | ( ~n2424 & n2659 ) ;
  assign n2661 = n2656 | n2660 ;
  assign n2662 = x175 & n1370 ;
  assign n2663 = x175 & ~n1373 ;
  assign n2664 = ( n1467 & n2662 ) | ( n1467 & n2663 ) | ( n2662 & n2663 ) ;
  assign n2665 = ( ~n1487 & n2662 ) | ( ~n1487 & n2663 ) | ( n2662 & n2663 ) ;
  assign n2666 = ( n1358 & n2664 ) | ( n1358 & n2665 ) | ( n2664 & n2665 ) ;
  assign n2667 = ( ~n1506 & n2664 ) | ( ~n1506 & n2665 ) | ( n2664 & n2665 ) ;
  assign n2668 = ( ~n1612 & n2666 ) | ( ~n1612 & n2667 ) | ( n2666 & n2667 ) ;
  assign n2669 = x47 & ~n1370 ;
  assign n2670 = x47 & n1373 ;
  assign n2671 = ( ~n1467 & n2669 ) | ( ~n1467 & n2670 ) | ( n2669 & n2670 ) ;
  assign n2672 = ( n1487 & n2669 ) | ( n1487 & n2670 ) | ( n2669 & n2670 ) ;
  assign n2673 = ( ~n1358 & n2671 ) | ( ~n1358 & n2672 ) | ( n2671 & n2672 ) ;
  assign n2674 = ( n1506 & n2671 ) | ( n1506 & n2672 ) | ( n2671 & n2672 ) ;
  assign n2675 = ( n1612 & n2673 ) | ( n1612 & n2674 ) | ( n2673 & n2674 ) ;
  assign n2676 = n2668 | n2675 ;
  assign n2677 = x431 & n812 ;
  assign n2678 = x431 & ~n815 ;
  assign n2679 = ( n909 & n2677 ) | ( n909 & n2678 ) | ( n2677 & n2678 ) ;
  assign n2680 = ( ~n929 & n2677 ) | ( ~n929 & n2678 ) | ( n2677 & n2678 ) ;
  assign n2681 = ( n800 & n2679 ) | ( n800 & n2680 ) | ( n2679 & n2680 ) ;
  assign n2682 = ( ~n948 & n2679 ) | ( ~n948 & n2680 ) | ( n2679 & n2680 ) ;
  assign n2683 = ( ~n1061 & n2681 ) | ( ~n1061 & n2682 ) | ( n2681 & n2682 ) ;
  assign n2684 = x303 & ~n812 ;
  assign n2685 = x303 & n815 ;
  assign n2686 = ( ~n909 & n2684 ) | ( ~n909 & n2685 ) | ( n2684 & n2685 ) ;
  assign n2687 = ( n929 & n2684 ) | ( n929 & n2685 ) | ( n2684 & n2685 ) ;
  assign n2688 = ( ~n800 & n2686 ) | ( ~n800 & n2687 ) | ( n2686 & n2687 ) ;
  assign n2689 = ( n948 & n2686 ) | ( n948 & n2687 ) | ( n2686 & n2687 ) ;
  assign n2690 = ( n1061 & n2688 ) | ( n1061 & n2689 ) | ( n2688 & n2689 ) ;
  assign n2691 = n2683 | n2690 ;
  assign n2692 = n2676 & ~n2691 ;
  assign n2693 = n2521 | n2616 ;
  assign n2694 = n2633 & ~n2648 ;
  assign n2695 = n2693 | n2694 ;
  assign n2696 = n2692 & ~n2695 ;
  assign n2697 = n2661 | n2696 ;
  assign n2698 = ~n2661 & n2695 ;
  assign n2699 = ~n2676 & n2691 ;
  assign n2700 = x430 & n812 ;
  assign n2701 = x430 & ~n815 ;
  assign n2702 = ( n909 & n2700 ) | ( n909 & n2701 ) | ( n2700 & n2701 ) ;
  assign n2703 = ( ~n929 & n2700 ) | ( ~n929 & n2701 ) | ( n2700 & n2701 ) ;
  assign n2704 = ( n800 & n2702 ) | ( n800 & n2703 ) | ( n2702 & n2703 ) ;
  assign n2705 = ( ~n948 & n2702 ) | ( ~n948 & n2703 ) | ( n2702 & n2703 ) ;
  assign n2706 = ( ~n1061 & n2704 ) | ( ~n1061 & n2705 ) | ( n2704 & n2705 ) ;
  assign n2707 = x302 & ~n812 ;
  assign n2708 = x302 & n815 ;
  assign n2709 = ( ~n909 & n2707 ) | ( ~n909 & n2708 ) | ( n2707 & n2708 ) ;
  assign n2710 = ( n929 & n2707 ) | ( n929 & n2708 ) | ( n2707 & n2708 ) ;
  assign n2711 = ( ~n800 & n2709 ) | ( ~n800 & n2710 ) | ( n2709 & n2710 ) ;
  assign n2712 = ( n948 & n2709 ) | ( n948 & n2710 ) | ( n2709 & n2710 ) ;
  assign n2713 = ( n1061 & n2711 ) | ( n1061 & n2712 ) | ( n2711 & n2712 ) ;
  assign n2714 = n2706 | n2713 ;
  assign n2715 = x174 & n1370 ;
  assign n2716 = x174 & ~n1373 ;
  assign n2717 = ( n1467 & n2715 ) | ( n1467 & n2716 ) | ( n2715 & n2716 ) ;
  assign n2718 = ( ~n1487 & n2715 ) | ( ~n1487 & n2716 ) | ( n2715 & n2716 ) ;
  assign n2719 = ( n1358 & n2717 ) | ( n1358 & n2718 ) | ( n2717 & n2718 ) ;
  assign n2720 = ( ~n1506 & n2717 ) | ( ~n1506 & n2718 ) | ( n2717 & n2718 ) ;
  assign n2721 = ( ~n1612 & n2719 ) | ( ~n1612 & n2720 ) | ( n2719 & n2720 ) ;
  assign n2722 = x46 & ~n1370 ;
  assign n2723 = x46 & n1373 ;
  assign n2724 = ( ~n1467 & n2722 ) | ( ~n1467 & n2723 ) | ( n2722 & n2723 ) ;
  assign n2725 = ( n1487 & n2722 ) | ( n1487 & n2723 ) | ( n2722 & n2723 ) ;
  assign n2726 = ( ~n1358 & n2724 ) | ( ~n1358 & n2725 ) | ( n2724 & n2725 ) ;
  assign n2727 = ( n1506 & n2724 ) | ( n1506 & n2725 ) | ( n2724 & n2725 ) ;
  assign n2728 = ( n1612 & n2726 ) | ( n1612 & n2727 ) | ( n2726 & n2727 ) ;
  assign n2729 = n2721 | n2728 ;
  assign n2730 = n2714 & ~n2729 ;
  assign n2731 = n2699 | n2730 ;
  assign n2732 = x172 & n1370 ;
  assign n2733 = x172 & ~n1373 ;
  assign n2734 = ( n1467 & n2732 ) | ( n1467 & n2733 ) | ( n2732 & n2733 ) ;
  assign n2735 = ( ~n1487 & n2732 ) | ( ~n1487 & n2733 ) | ( n2732 & n2733 ) ;
  assign n2736 = ( n1358 & n2734 ) | ( n1358 & n2735 ) | ( n2734 & n2735 ) ;
  assign n2737 = ( ~n1506 & n2734 ) | ( ~n1506 & n2735 ) | ( n2734 & n2735 ) ;
  assign n2738 = ( ~n1612 & n2736 ) | ( ~n1612 & n2737 ) | ( n2736 & n2737 ) ;
  assign n2739 = x44 & ~n1370 ;
  assign n2740 = x44 & n1373 ;
  assign n2741 = ( ~n1467 & n2739 ) | ( ~n1467 & n2740 ) | ( n2739 & n2740 ) ;
  assign n2742 = ( n1487 & n2739 ) | ( n1487 & n2740 ) | ( n2739 & n2740 ) ;
  assign n2743 = ( ~n1358 & n2741 ) | ( ~n1358 & n2742 ) | ( n2741 & n2742 ) ;
  assign n2744 = ( n1506 & n2741 ) | ( n1506 & n2742 ) | ( n2741 & n2742 ) ;
  assign n2745 = ( n1612 & n2743 ) | ( n1612 & n2744 ) | ( n2743 & n2744 ) ;
  assign n2746 = n2738 | n2745 ;
  assign n2747 = x428 & n812 ;
  assign n2748 = x428 & ~n815 ;
  assign n2749 = ( n909 & n2747 ) | ( n909 & n2748 ) | ( n2747 & n2748 ) ;
  assign n2750 = ( ~n929 & n2747 ) | ( ~n929 & n2748 ) | ( n2747 & n2748 ) ;
  assign n2751 = ( n800 & n2749 ) | ( n800 & n2750 ) | ( n2749 & n2750 ) ;
  assign n2752 = ( ~n948 & n2749 ) | ( ~n948 & n2750 ) | ( n2749 & n2750 ) ;
  assign n2753 = ( ~n1061 & n2751 ) | ( ~n1061 & n2752 ) | ( n2751 & n2752 ) ;
  assign n2754 = x300 & ~n812 ;
  assign n2755 = x300 & n815 ;
  assign n2756 = ( ~n909 & n2754 ) | ( ~n909 & n2755 ) | ( n2754 & n2755 ) ;
  assign n2757 = ( n929 & n2754 ) | ( n929 & n2755 ) | ( n2754 & n2755 ) ;
  assign n2758 = ( ~n800 & n2756 ) | ( ~n800 & n2757 ) | ( n2756 & n2757 ) ;
  assign n2759 = ( n948 & n2756 ) | ( n948 & n2757 ) | ( n2756 & n2757 ) ;
  assign n2760 = ( n1061 & n2758 ) | ( n1061 & n2759 ) | ( n2758 & n2759 ) ;
  assign n2761 = n2753 | n2760 ;
  assign n2762 = ~n2746 & n2761 ;
  assign n2763 = x173 & n1370 ;
  assign n2764 = x173 & ~n1373 ;
  assign n2765 = ( n1467 & n2763 ) | ( n1467 & n2764 ) | ( n2763 & n2764 ) ;
  assign n2766 = ( ~n1487 & n2763 ) | ( ~n1487 & n2764 ) | ( n2763 & n2764 ) ;
  assign n2767 = ( n1358 & n2765 ) | ( n1358 & n2766 ) | ( n2765 & n2766 ) ;
  assign n2768 = ( ~n1506 & n2765 ) | ( ~n1506 & n2766 ) | ( n2765 & n2766 ) ;
  assign n2769 = ( ~n1612 & n2767 ) | ( ~n1612 & n2768 ) | ( n2767 & n2768 ) ;
  assign n2770 = x45 & ~n1370 ;
  assign n2771 = x45 & n1373 ;
  assign n2772 = ( ~n1467 & n2770 ) | ( ~n1467 & n2771 ) | ( n2770 & n2771 ) ;
  assign n2773 = ( n1487 & n2770 ) | ( n1487 & n2771 ) | ( n2770 & n2771 ) ;
  assign n2774 = ( ~n1358 & n2772 ) | ( ~n1358 & n2773 ) | ( n2772 & n2773 ) ;
  assign n2775 = ( n1506 & n2772 ) | ( n1506 & n2773 ) | ( n2772 & n2773 ) ;
  assign n2776 = ( n1612 & n2774 ) | ( n1612 & n2775 ) | ( n2774 & n2775 ) ;
  assign n2777 = n2769 | n2776 ;
  assign n2778 = x429 & n812 ;
  assign n2779 = x429 & ~n815 ;
  assign n2780 = ( n909 & n2778 ) | ( n909 & n2779 ) | ( n2778 & n2779 ) ;
  assign n2781 = ( ~n929 & n2778 ) | ( ~n929 & n2779 ) | ( n2778 & n2779 ) ;
  assign n2782 = ( n800 & n2780 ) | ( n800 & n2781 ) | ( n2780 & n2781 ) ;
  assign n2783 = ( ~n948 & n2780 ) | ( ~n948 & n2781 ) | ( n2780 & n2781 ) ;
  assign n2784 = ( ~n1061 & n2782 ) | ( ~n1061 & n2783 ) | ( n2782 & n2783 ) ;
  assign n2785 = x301 & ~n812 ;
  assign n2786 = x301 & n815 ;
  assign n2787 = ( ~n909 & n2785 ) | ( ~n909 & n2786 ) | ( n2785 & n2786 ) ;
  assign n2788 = ( n929 & n2785 ) | ( n929 & n2786 ) | ( n2785 & n2786 ) ;
  assign n2789 = ( ~n800 & n2787 ) | ( ~n800 & n2788 ) | ( n2787 & n2788 ) ;
  assign n2790 = ( n948 & n2787 ) | ( n948 & n2788 ) | ( n2787 & n2788 ) ;
  assign n2791 = ( n1061 & n2789 ) | ( n1061 & n2790 ) | ( n2789 & n2790 ) ;
  assign n2792 = n2784 | n2791 ;
  assign n2793 = ~n2777 & n2792 ;
  assign n2794 = n2762 | n2793 ;
  assign n2795 = n2731 | n2794 ;
  assign n2796 = x171 & n1370 ;
  assign n2797 = x171 & ~n1373 ;
  assign n2798 = ( n1467 & n2796 ) | ( n1467 & n2797 ) | ( n2796 & n2797 ) ;
  assign n2799 = ( ~n1487 & n2796 ) | ( ~n1487 & n2797 ) | ( n2796 & n2797 ) ;
  assign n2800 = ( n1358 & n2798 ) | ( n1358 & n2799 ) | ( n2798 & n2799 ) ;
  assign n2801 = ( ~n1506 & n2798 ) | ( ~n1506 & n2799 ) | ( n2798 & n2799 ) ;
  assign n2802 = ( ~n1612 & n2800 ) | ( ~n1612 & n2801 ) | ( n2800 & n2801 ) ;
  assign n2803 = x43 & ~n1370 ;
  assign n2804 = x43 & n1373 ;
  assign n2805 = ( ~n1467 & n2803 ) | ( ~n1467 & n2804 ) | ( n2803 & n2804 ) ;
  assign n2806 = ( n1487 & n2803 ) | ( n1487 & n2804 ) | ( n2803 & n2804 ) ;
  assign n2807 = ( ~n1358 & n2805 ) | ( ~n1358 & n2806 ) | ( n2805 & n2806 ) ;
  assign n2808 = ( n1506 & n2805 ) | ( n1506 & n2806 ) | ( n2805 & n2806 ) ;
  assign n2809 = ( n1612 & n2807 ) | ( n1612 & n2808 ) | ( n2807 & n2808 ) ;
  assign n2810 = n2802 | n2809 ;
  assign n2811 = x427 & n812 ;
  assign n2812 = x427 & ~n815 ;
  assign n2813 = ( n909 & n2811 ) | ( n909 & n2812 ) | ( n2811 & n2812 ) ;
  assign n2814 = ( ~n929 & n2811 ) | ( ~n929 & n2812 ) | ( n2811 & n2812 ) ;
  assign n2815 = ( n800 & n2813 ) | ( n800 & n2814 ) | ( n2813 & n2814 ) ;
  assign n2816 = ( ~n948 & n2813 ) | ( ~n948 & n2814 ) | ( n2813 & n2814 ) ;
  assign n2817 = ( ~n1061 & n2815 ) | ( ~n1061 & n2816 ) | ( n2815 & n2816 ) ;
  assign n2818 = x299 & ~n812 ;
  assign n2819 = x299 & n815 ;
  assign n2820 = ( ~n909 & n2818 ) | ( ~n909 & n2819 ) | ( n2818 & n2819 ) ;
  assign n2821 = ( n929 & n2818 ) | ( n929 & n2819 ) | ( n2818 & n2819 ) ;
  assign n2822 = ( ~n800 & n2820 ) | ( ~n800 & n2821 ) | ( n2820 & n2821 ) ;
  assign n2823 = ( n948 & n2820 ) | ( n948 & n2821 ) | ( n2820 & n2821 ) ;
  assign n2824 = ( n1061 & n2822 ) | ( n1061 & n2823 ) | ( n2822 & n2823 ) ;
  assign n2825 = n2817 | n2824 ;
  assign n2826 = x170 & n1370 ;
  assign n2827 = x170 & ~n1373 ;
  assign n2828 = ( n1467 & n2826 ) | ( n1467 & n2827 ) | ( n2826 & n2827 ) ;
  assign n2829 = ( ~n1487 & n2826 ) | ( ~n1487 & n2827 ) | ( n2826 & n2827 ) ;
  assign n2830 = ( n1358 & n2828 ) | ( n1358 & n2829 ) | ( n2828 & n2829 ) ;
  assign n2831 = ( ~n1506 & n2828 ) | ( ~n1506 & n2829 ) | ( n2828 & n2829 ) ;
  assign n2832 = ( ~n1612 & n2830 ) | ( ~n1612 & n2831 ) | ( n2830 & n2831 ) ;
  assign n2833 = x42 & ~n1370 ;
  assign n2834 = x42 & n1373 ;
  assign n2835 = ( ~n1467 & n2833 ) | ( ~n1467 & n2834 ) | ( n2833 & n2834 ) ;
  assign n2836 = ( n1487 & n2833 ) | ( n1487 & n2834 ) | ( n2833 & n2834 ) ;
  assign n2837 = ( ~n1358 & n2835 ) | ( ~n1358 & n2836 ) | ( n2835 & n2836 ) ;
  assign n2838 = ( n1506 & n2835 ) | ( n1506 & n2836 ) | ( n2835 & n2836 ) ;
  assign n2839 = ( n1612 & n2837 ) | ( n1612 & n2838 ) | ( n2837 & n2838 ) ;
  assign n2840 = n2832 | n2839 ;
  assign n2841 = x426 & n812 ;
  assign n2842 = x426 & ~n815 ;
  assign n2843 = ( n909 & n2841 ) | ( n909 & n2842 ) | ( n2841 & n2842 ) ;
  assign n2844 = ( ~n929 & n2841 ) | ( ~n929 & n2842 ) | ( n2841 & n2842 ) ;
  assign n2845 = ( n800 & n2843 ) | ( n800 & n2844 ) | ( n2843 & n2844 ) ;
  assign n2846 = ( ~n948 & n2843 ) | ( ~n948 & n2844 ) | ( n2843 & n2844 ) ;
  assign n2847 = ( ~n1061 & n2845 ) | ( ~n1061 & n2846 ) | ( n2845 & n2846 ) ;
  assign n2848 = x298 & ~n812 ;
  assign n2849 = x298 & n815 ;
  assign n2850 = ( ~n909 & n2848 ) | ( ~n909 & n2849 ) | ( n2848 & n2849 ) ;
  assign n2851 = ( n929 & n2848 ) | ( n929 & n2849 ) | ( n2848 & n2849 ) ;
  assign n2852 = ( ~n800 & n2850 ) | ( ~n800 & n2851 ) | ( n2850 & n2851 ) ;
  assign n2853 = ( n948 & n2850 ) | ( n948 & n2851 ) | ( n2850 & n2851 ) ;
  assign n2854 = ( n1061 & n2852 ) | ( n1061 & n2853 ) | ( n2852 & n2853 ) ;
  assign n2855 = n2847 | n2854 ;
  assign n2856 = x169 & n1370 ;
  assign n2857 = x169 & ~n1373 ;
  assign n2858 = ( n1467 & n2856 ) | ( n1467 & n2857 ) | ( n2856 & n2857 ) ;
  assign n2859 = ( ~n1487 & n2856 ) | ( ~n1487 & n2857 ) | ( n2856 & n2857 ) ;
  assign n2860 = ( n1358 & n2858 ) | ( n1358 & n2859 ) | ( n2858 & n2859 ) ;
  assign n2861 = ( ~n1506 & n2858 ) | ( ~n1506 & n2859 ) | ( n2858 & n2859 ) ;
  assign n2862 = ( ~n1612 & n2860 ) | ( ~n1612 & n2861 ) | ( n2860 & n2861 ) ;
  assign n2863 = x41 & ~n1370 ;
  assign n2864 = x41 & n1373 ;
  assign n2865 = ( ~n1467 & n2863 ) | ( ~n1467 & n2864 ) | ( n2863 & n2864 ) ;
  assign n2866 = ( n1487 & n2863 ) | ( n1487 & n2864 ) | ( n2863 & n2864 ) ;
  assign n2867 = ( ~n1358 & n2865 ) | ( ~n1358 & n2866 ) | ( n2865 & n2866 ) ;
  assign n2868 = ( n1506 & n2865 ) | ( n1506 & n2866 ) | ( n2865 & n2866 ) ;
  assign n2869 = ( n1612 & n2867 ) | ( n1612 & n2868 ) | ( n2867 & n2868 ) ;
  assign n2870 = n2862 | n2869 ;
  assign n2871 = x425 & n812 ;
  assign n2872 = x425 & ~n815 ;
  assign n2873 = ( n909 & n2871 ) | ( n909 & n2872 ) | ( n2871 & n2872 ) ;
  assign n2874 = ( ~n929 & n2871 ) | ( ~n929 & n2872 ) | ( n2871 & n2872 ) ;
  assign n2875 = ( n800 & n2873 ) | ( n800 & n2874 ) | ( n2873 & n2874 ) ;
  assign n2876 = ( ~n948 & n2873 ) | ( ~n948 & n2874 ) | ( n2873 & n2874 ) ;
  assign n2877 = ( ~n1061 & n2875 ) | ( ~n1061 & n2876 ) | ( n2875 & n2876 ) ;
  assign n2878 = x297 & ~n812 ;
  assign n2879 = x297 & n815 ;
  assign n2880 = ( ~n909 & n2878 ) | ( ~n909 & n2879 ) | ( n2878 & n2879 ) ;
  assign n2881 = ( n929 & n2878 ) | ( n929 & n2879 ) | ( n2878 & n2879 ) ;
  assign n2882 = ( ~n800 & n2880 ) | ( ~n800 & n2881 ) | ( n2880 & n2881 ) ;
  assign n2883 = ( n948 & n2880 ) | ( n948 & n2881 ) | ( n2880 & n2881 ) ;
  assign n2884 = ( n1061 & n2882 ) | ( n1061 & n2883 ) | ( n2882 & n2883 ) ;
  assign n2885 = n2877 | n2884 ;
  assign n2886 = x168 & n1370 ;
  assign n2887 = x168 & ~n1373 ;
  assign n2888 = ( n1467 & n2886 ) | ( n1467 & n2887 ) | ( n2886 & n2887 ) ;
  assign n2889 = ( ~n1487 & n2886 ) | ( ~n1487 & n2887 ) | ( n2886 & n2887 ) ;
  assign n2890 = ( n1358 & n2888 ) | ( n1358 & n2889 ) | ( n2888 & n2889 ) ;
  assign n2891 = ( ~n1506 & n2888 ) | ( ~n1506 & n2889 ) | ( n2888 & n2889 ) ;
  assign n2892 = ( ~n1612 & n2890 ) | ( ~n1612 & n2891 ) | ( n2890 & n2891 ) ;
  assign n2893 = x40 & ~n1370 ;
  assign n2894 = x40 & n1373 ;
  assign n2895 = ( ~n1467 & n2893 ) | ( ~n1467 & n2894 ) | ( n2893 & n2894 ) ;
  assign n2896 = ( n1487 & n2893 ) | ( n1487 & n2894 ) | ( n2893 & n2894 ) ;
  assign n2897 = ( ~n1358 & n2895 ) | ( ~n1358 & n2896 ) | ( n2895 & n2896 ) ;
  assign n2898 = ( n1506 & n2895 ) | ( n1506 & n2896 ) | ( n2895 & n2896 ) ;
  assign n2899 = ( n1612 & n2897 ) | ( n1612 & n2898 ) | ( n2897 & n2898 ) ;
  assign n2900 = n2892 | n2899 ;
  assign n2901 = x424 & n812 ;
  assign n2902 = x424 & ~n815 ;
  assign n2903 = ( n909 & n2901 ) | ( n909 & n2902 ) | ( n2901 & n2902 ) ;
  assign n2904 = ( ~n929 & n2901 ) | ( ~n929 & n2902 ) | ( n2901 & n2902 ) ;
  assign n2905 = ( n800 & n2903 ) | ( n800 & n2904 ) | ( n2903 & n2904 ) ;
  assign n2906 = ( ~n948 & n2903 ) | ( ~n948 & n2904 ) | ( n2903 & n2904 ) ;
  assign n2907 = ( ~n1061 & n2905 ) | ( ~n1061 & n2906 ) | ( n2905 & n2906 ) ;
  assign n2908 = x296 & ~n812 ;
  assign n2909 = x296 & n815 ;
  assign n2910 = ( ~n909 & n2908 ) | ( ~n909 & n2909 ) | ( n2908 & n2909 ) ;
  assign n2911 = ( n929 & n2908 ) | ( n929 & n2909 ) | ( n2908 & n2909 ) ;
  assign n2912 = ( ~n800 & n2910 ) | ( ~n800 & n2911 ) | ( n2910 & n2911 ) ;
  assign n2913 = ( n948 & n2910 ) | ( n948 & n2911 ) | ( n2910 & n2911 ) ;
  assign n2914 = ( n1061 & n2912 ) | ( n1061 & n2913 ) | ( n2912 & n2913 ) ;
  assign n2915 = n2907 | n2914 ;
  assign n2916 = n2900 & ~n2915 ;
  assign n2917 = ( n2870 & ~n2885 ) | ( n2870 & n2916 ) | ( ~n2885 & n2916 ) ;
  assign n2918 = ( n2840 & ~n2855 ) | ( n2840 & n2917 ) | ( ~n2855 & n2917 ) ;
  assign n2919 = ( n2810 & ~n2825 ) | ( n2810 & n2918 ) | ( ~n2825 & n2918 ) ;
  assign n2920 = ~n2795 & n2919 ;
  assign n2921 = n2746 & ~n2761 ;
  assign n2922 = ( n2777 & ~n2792 ) | ( n2777 & n2921 ) | ( ~n2792 & n2921 ) ;
  assign n2923 = ~n2731 & n2922 ;
  assign n2924 = ~n2714 & n2729 ;
  assign n2925 = ~n2699 & n2924 ;
  assign n2926 = n2923 | n2925 ;
  assign n2927 = x416 & n812 ;
  assign n2928 = x416 & ~n815 ;
  assign n2929 = ( n909 & n2927 ) | ( n909 & n2928 ) | ( n2927 & n2928 ) ;
  assign n2930 = ( ~n929 & n2927 ) | ( ~n929 & n2928 ) | ( n2927 & n2928 ) ;
  assign n2931 = ( n800 & n2929 ) | ( n800 & n2930 ) | ( n2929 & n2930 ) ;
  assign n2932 = ( ~n948 & n2929 ) | ( ~n948 & n2930 ) | ( n2929 & n2930 ) ;
  assign n2933 = ( ~n1061 & n2931 ) | ( ~n1061 & n2932 ) | ( n2931 & n2932 ) ;
  assign n2934 = x288 & ~n812 ;
  assign n2935 = x288 & n815 ;
  assign n2936 = ( ~n909 & n2934 ) | ( ~n909 & n2935 ) | ( n2934 & n2935 ) ;
  assign n2937 = ( n929 & n2934 ) | ( n929 & n2935 ) | ( n2934 & n2935 ) ;
  assign n2938 = ( ~n800 & n2936 ) | ( ~n800 & n2937 ) | ( n2936 & n2937 ) ;
  assign n2939 = ( n948 & n2936 ) | ( n948 & n2937 ) | ( n2936 & n2937 ) ;
  assign n2940 = ( n1061 & n2938 ) | ( n1061 & n2939 ) | ( n2938 & n2939 ) ;
  assign n2941 = n2933 | n2940 ;
  assign n2942 = x160 & n1370 ;
  assign n2943 = x160 & ~n1373 ;
  assign n2944 = ( n1467 & n2942 ) | ( n1467 & n2943 ) | ( n2942 & n2943 ) ;
  assign n2945 = ( ~n1487 & n2942 ) | ( ~n1487 & n2943 ) | ( n2942 & n2943 ) ;
  assign n2946 = ( n1358 & n2944 ) | ( n1358 & n2945 ) | ( n2944 & n2945 ) ;
  assign n2947 = ( ~n1506 & n2944 ) | ( ~n1506 & n2945 ) | ( n2944 & n2945 ) ;
  assign n2948 = ( ~n1612 & n2946 ) | ( ~n1612 & n2947 ) | ( n2946 & n2947 ) ;
  assign n2949 = x32 & ~n1370 ;
  assign n2950 = x32 & n1373 ;
  assign n2951 = ( ~n1467 & n2949 ) | ( ~n1467 & n2950 ) | ( n2949 & n2950 ) ;
  assign n2952 = ( n1487 & n2949 ) | ( n1487 & n2950 ) | ( n2949 & n2950 ) ;
  assign n2953 = ( ~n1358 & n2951 ) | ( ~n1358 & n2952 ) | ( n2951 & n2952 ) ;
  assign n2954 = ( n1506 & n2951 ) | ( n1506 & n2952 ) | ( n2951 & n2952 ) ;
  assign n2955 = ( n1612 & n2953 ) | ( n1612 & n2954 ) | ( n2953 & n2954 ) ;
  assign n2956 = n2948 | n2955 ;
  assign n2957 = n2941 & ~n2956 ;
  assign n2958 = x167 & n1370 ;
  assign n2959 = x167 & ~n1373 ;
  assign n2960 = ( n1467 & n2958 ) | ( n1467 & n2959 ) | ( n2958 & n2959 ) ;
  assign n2961 = ( ~n1487 & n2958 ) | ( ~n1487 & n2959 ) | ( n2958 & n2959 ) ;
  assign n2962 = ( n1358 & n2960 ) | ( n1358 & n2961 ) | ( n2960 & n2961 ) ;
  assign n2963 = ( ~n1506 & n2960 ) | ( ~n1506 & n2961 ) | ( n2960 & n2961 ) ;
  assign n2964 = ( ~n1612 & n2962 ) | ( ~n1612 & n2963 ) | ( n2962 & n2963 ) ;
  assign n2965 = x39 & ~n1370 ;
  assign n2966 = x39 & n1373 ;
  assign n2967 = ( ~n1467 & n2965 ) | ( ~n1467 & n2966 ) | ( n2965 & n2966 ) ;
  assign n2968 = ( n1487 & n2965 ) | ( n1487 & n2966 ) | ( n2965 & n2966 ) ;
  assign n2969 = ( ~n1358 & n2967 ) | ( ~n1358 & n2968 ) | ( n2967 & n2968 ) ;
  assign n2970 = ( n1506 & n2967 ) | ( n1506 & n2968 ) | ( n2967 & n2968 ) ;
  assign n2971 = ( n1612 & n2969 ) | ( n1612 & n2970 ) | ( n2969 & n2970 ) ;
  assign n2972 = n2964 | n2971 ;
  assign n2973 = x423 & n812 ;
  assign n2974 = x423 & ~n815 ;
  assign n2975 = ( n909 & n2973 ) | ( n909 & n2974 ) | ( n2973 & n2974 ) ;
  assign n2976 = ( ~n929 & n2973 ) | ( ~n929 & n2974 ) | ( n2973 & n2974 ) ;
  assign n2977 = ( n800 & n2975 ) | ( n800 & n2976 ) | ( n2975 & n2976 ) ;
  assign n2978 = ( ~n948 & n2975 ) | ( ~n948 & n2976 ) | ( n2975 & n2976 ) ;
  assign n2979 = ( ~n1061 & n2977 ) | ( ~n1061 & n2978 ) | ( n2977 & n2978 ) ;
  assign n2980 = x295 & ~n812 ;
  assign n2981 = x295 & n815 ;
  assign n2982 = ( ~n909 & n2980 ) | ( ~n909 & n2981 ) | ( n2980 & n2981 ) ;
  assign n2983 = ( n929 & n2980 ) | ( n929 & n2981 ) | ( n2980 & n2981 ) ;
  assign n2984 = ( ~n800 & n2982 ) | ( ~n800 & n2983 ) | ( n2982 & n2983 ) ;
  assign n2985 = ( n948 & n2982 ) | ( n948 & n2983 ) | ( n2982 & n2983 ) ;
  assign n2986 = ( n1061 & n2984 ) | ( n1061 & n2985 ) | ( n2984 & n2985 ) ;
  assign n2987 = n2979 | n2986 ;
  assign n2988 = ~n2972 & n2987 ;
  assign n2989 = x422 & n812 ;
  assign n2990 = x422 & ~n815 ;
  assign n2991 = ( n909 & n2989 ) | ( n909 & n2990 ) | ( n2989 & n2990 ) ;
  assign n2992 = ( ~n929 & n2989 ) | ( ~n929 & n2990 ) | ( n2989 & n2990 ) ;
  assign n2993 = ( n800 & n2991 ) | ( n800 & n2992 ) | ( n2991 & n2992 ) ;
  assign n2994 = ( ~n948 & n2991 ) | ( ~n948 & n2992 ) | ( n2991 & n2992 ) ;
  assign n2995 = ( ~n1061 & n2993 ) | ( ~n1061 & n2994 ) | ( n2993 & n2994 ) ;
  assign n2996 = x294 & ~n812 ;
  assign n2997 = x294 & n815 ;
  assign n2998 = ( ~n909 & n2996 ) | ( ~n909 & n2997 ) | ( n2996 & n2997 ) ;
  assign n2999 = ( n929 & n2996 ) | ( n929 & n2997 ) | ( n2996 & n2997 ) ;
  assign n3000 = ( ~n800 & n2998 ) | ( ~n800 & n2999 ) | ( n2998 & n2999 ) ;
  assign n3001 = ( n948 & n2998 ) | ( n948 & n2999 ) | ( n2998 & n2999 ) ;
  assign n3002 = ( n1061 & n3000 ) | ( n1061 & n3001 ) | ( n3000 & n3001 ) ;
  assign n3003 = n2995 | n3002 ;
  assign n3004 = x166 & n1370 ;
  assign n3005 = x166 & ~n1373 ;
  assign n3006 = ( n1467 & n3004 ) | ( n1467 & n3005 ) | ( n3004 & n3005 ) ;
  assign n3007 = ( ~n1487 & n3004 ) | ( ~n1487 & n3005 ) | ( n3004 & n3005 ) ;
  assign n3008 = ( n1358 & n3006 ) | ( n1358 & n3007 ) | ( n3006 & n3007 ) ;
  assign n3009 = ( ~n1506 & n3006 ) | ( ~n1506 & n3007 ) | ( n3006 & n3007 ) ;
  assign n3010 = ( ~n1612 & n3008 ) | ( ~n1612 & n3009 ) | ( n3008 & n3009 ) ;
  assign n3011 = x38 & ~n1370 ;
  assign n3012 = x38 & n1373 ;
  assign n3013 = ( ~n1467 & n3011 ) | ( ~n1467 & n3012 ) | ( n3011 & n3012 ) ;
  assign n3014 = ( n1487 & n3011 ) | ( n1487 & n3012 ) | ( n3011 & n3012 ) ;
  assign n3015 = ( ~n1358 & n3013 ) | ( ~n1358 & n3014 ) | ( n3013 & n3014 ) ;
  assign n3016 = ( n1506 & n3013 ) | ( n1506 & n3014 ) | ( n3013 & n3014 ) ;
  assign n3017 = ( n1612 & n3015 ) | ( n1612 & n3016 ) | ( n3015 & n3016 ) ;
  assign n3018 = n3010 | n3017 ;
  assign n3019 = n3003 & ~n3018 ;
  assign n3020 = n2988 | n3019 ;
  assign n3021 = x164 & n1370 ;
  assign n3022 = x164 & ~n1373 ;
  assign n3023 = ( n1467 & n3021 ) | ( n1467 & n3022 ) | ( n3021 & n3022 ) ;
  assign n3024 = ( ~n1487 & n3021 ) | ( ~n1487 & n3022 ) | ( n3021 & n3022 ) ;
  assign n3025 = ( n1358 & n3023 ) | ( n1358 & n3024 ) | ( n3023 & n3024 ) ;
  assign n3026 = ( ~n1506 & n3023 ) | ( ~n1506 & n3024 ) | ( n3023 & n3024 ) ;
  assign n3027 = ( ~n1612 & n3025 ) | ( ~n1612 & n3026 ) | ( n3025 & n3026 ) ;
  assign n3028 = x36 & ~n1370 ;
  assign n3029 = x36 & n1373 ;
  assign n3030 = ( ~n1467 & n3028 ) | ( ~n1467 & n3029 ) | ( n3028 & n3029 ) ;
  assign n3031 = ( n1487 & n3028 ) | ( n1487 & n3029 ) | ( n3028 & n3029 ) ;
  assign n3032 = ( ~n1358 & n3030 ) | ( ~n1358 & n3031 ) | ( n3030 & n3031 ) ;
  assign n3033 = ( n1506 & n3030 ) | ( n1506 & n3031 ) | ( n3030 & n3031 ) ;
  assign n3034 = ( n1612 & n3032 ) | ( n1612 & n3033 ) | ( n3032 & n3033 ) ;
  assign n3035 = n3027 | n3034 ;
  assign n3036 = x420 & n812 ;
  assign n3037 = x420 & ~n815 ;
  assign n3038 = ( n909 & n3036 ) | ( n909 & n3037 ) | ( n3036 & n3037 ) ;
  assign n3039 = ( ~n929 & n3036 ) | ( ~n929 & n3037 ) | ( n3036 & n3037 ) ;
  assign n3040 = ( n800 & n3038 ) | ( n800 & n3039 ) | ( n3038 & n3039 ) ;
  assign n3041 = ( ~n948 & n3038 ) | ( ~n948 & n3039 ) | ( n3038 & n3039 ) ;
  assign n3042 = ( ~n1061 & n3040 ) | ( ~n1061 & n3041 ) | ( n3040 & n3041 ) ;
  assign n3043 = x292 & ~n812 ;
  assign n3044 = x292 & n815 ;
  assign n3045 = ( ~n909 & n3043 ) | ( ~n909 & n3044 ) | ( n3043 & n3044 ) ;
  assign n3046 = ( n929 & n3043 ) | ( n929 & n3044 ) | ( n3043 & n3044 ) ;
  assign n3047 = ( ~n800 & n3045 ) | ( ~n800 & n3046 ) | ( n3045 & n3046 ) ;
  assign n3048 = ( n948 & n3045 ) | ( n948 & n3046 ) | ( n3045 & n3046 ) ;
  assign n3049 = ( n1061 & n3047 ) | ( n1061 & n3048 ) | ( n3047 & n3048 ) ;
  assign n3050 = n3042 | n3049 ;
  assign n3051 = ~n3035 & n3050 ;
  assign n3052 = x165 & n1370 ;
  assign n3053 = x165 & ~n1373 ;
  assign n3054 = ( n1467 & n3052 ) | ( n1467 & n3053 ) | ( n3052 & n3053 ) ;
  assign n3055 = ( ~n1487 & n3052 ) | ( ~n1487 & n3053 ) | ( n3052 & n3053 ) ;
  assign n3056 = ( n1358 & n3054 ) | ( n1358 & n3055 ) | ( n3054 & n3055 ) ;
  assign n3057 = ( ~n1506 & n3054 ) | ( ~n1506 & n3055 ) | ( n3054 & n3055 ) ;
  assign n3058 = ( ~n1612 & n3056 ) | ( ~n1612 & n3057 ) | ( n3056 & n3057 ) ;
  assign n3059 = x37 & ~n1370 ;
  assign n3060 = x37 & n1373 ;
  assign n3061 = ( ~n1467 & n3059 ) | ( ~n1467 & n3060 ) | ( n3059 & n3060 ) ;
  assign n3062 = ( n1487 & n3059 ) | ( n1487 & n3060 ) | ( n3059 & n3060 ) ;
  assign n3063 = ( ~n1358 & n3061 ) | ( ~n1358 & n3062 ) | ( n3061 & n3062 ) ;
  assign n3064 = ( n1506 & n3061 ) | ( n1506 & n3062 ) | ( n3061 & n3062 ) ;
  assign n3065 = ( n1612 & n3063 ) | ( n1612 & n3064 ) | ( n3063 & n3064 ) ;
  assign n3066 = n3058 | n3065 ;
  assign n3067 = x421 & n812 ;
  assign n3068 = x421 & ~n815 ;
  assign n3069 = ( n909 & n3067 ) | ( n909 & n3068 ) | ( n3067 & n3068 ) ;
  assign n3070 = ( ~n929 & n3067 ) | ( ~n929 & n3068 ) | ( n3067 & n3068 ) ;
  assign n3071 = ( n800 & n3069 ) | ( n800 & n3070 ) | ( n3069 & n3070 ) ;
  assign n3072 = ( ~n948 & n3069 ) | ( ~n948 & n3070 ) | ( n3069 & n3070 ) ;
  assign n3073 = ( ~n1061 & n3071 ) | ( ~n1061 & n3072 ) | ( n3071 & n3072 ) ;
  assign n3074 = x293 & ~n812 ;
  assign n3075 = x293 & n815 ;
  assign n3076 = ( ~n909 & n3074 ) | ( ~n909 & n3075 ) | ( n3074 & n3075 ) ;
  assign n3077 = ( n929 & n3074 ) | ( n929 & n3075 ) | ( n3074 & n3075 ) ;
  assign n3078 = ( ~n800 & n3076 ) | ( ~n800 & n3077 ) | ( n3076 & n3077 ) ;
  assign n3079 = ( n948 & n3076 ) | ( n948 & n3077 ) | ( n3076 & n3077 ) ;
  assign n3080 = ( n1061 & n3078 ) | ( n1061 & n3079 ) | ( n3078 & n3079 ) ;
  assign n3081 = n3073 | n3080 ;
  assign n3082 = ~n3066 & n3081 ;
  assign n3083 = n3051 | n3082 ;
  assign n3084 = n3020 | n3083 ;
  assign n3085 = x161 & n1370 ;
  assign n3086 = x161 & ~n1373 ;
  assign n3087 = ( n1467 & n3085 ) | ( n1467 & n3086 ) | ( n3085 & n3086 ) ;
  assign n3088 = ( ~n1487 & n3085 ) | ( ~n1487 & n3086 ) | ( n3085 & n3086 ) ;
  assign n3089 = ( n1358 & n3087 ) | ( n1358 & n3088 ) | ( n3087 & n3088 ) ;
  assign n3090 = ( ~n1506 & n3087 ) | ( ~n1506 & n3088 ) | ( n3087 & n3088 ) ;
  assign n3091 = ( ~n1612 & n3089 ) | ( ~n1612 & n3090 ) | ( n3089 & n3090 ) ;
  assign n3092 = x33 & ~n1370 ;
  assign n3093 = x33 & n1373 ;
  assign n3094 = ( ~n1467 & n3092 ) | ( ~n1467 & n3093 ) | ( n3092 & n3093 ) ;
  assign n3095 = ( n1487 & n3092 ) | ( n1487 & n3093 ) | ( n3092 & n3093 ) ;
  assign n3096 = ( ~n1358 & n3094 ) | ( ~n1358 & n3095 ) | ( n3094 & n3095 ) ;
  assign n3097 = ( n1506 & n3094 ) | ( n1506 & n3095 ) | ( n3094 & n3095 ) ;
  assign n3098 = ( n1612 & n3096 ) | ( n1612 & n3097 ) | ( n3096 & n3097 ) ;
  assign n3099 = n3091 | n3098 ;
  assign n3100 = x417 & n812 ;
  assign n3101 = x417 & ~n815 ;
  assign n3102 = ( n909 & n3100 ) | ( n909 & n3101 ) | ( n3100 & n3101 ) ;
  assign n3103 = ( ~n929 & n3100 ) | ( ~n929 & n3101 ) | ( n3100 & n3101 ) ;
  assign n3104 = ( n800 & n3102 ) | ( n800 & n3103 ) | ( n3102 & n3103 ) ;
  assign n3105 = ( ~n948 & n3102 ) | ( ~n948 & n3103 ) | ( n3102 & n3103 ) ;
  assign n3106 = ( ~n1061 & n3104 ) | ( ~n1061 & n3105 ) | ( n3104 & n3105 ) ;
  assign n3107 = x289 & ~n812 ;
  assign n3108 = x289 & n815 ;
  assign n3109 = ( ~n909 & n3107 ) | ( ~n909 & n3108 ) | ( n3107 & n3108 ) ;
  assign n3110 = ( n929 & n3107 ) | ( n929 & n3108 ) | ( n3107 & n3108 ) ;
  assign n3111 = ( ~n800 & n3109 ) | ( ~n800 & n3110 ) | ( n3109 & n3110 ) ;
  assign n3112 = ( n948 & n3109 ) | ( n948 & n3110 ) | ( n3109 & n3110 ) ;
  assign n3113 = ( n1061 & n3111 ) | ( n1061 & n3112 ) | ( n3111 & n3112 ) ;
  assign n3114 = n3106 | n3113 ;
  assign n3115 = ~n3099 & n3114 ;
  assign n3116 = x163 & n1370 ;
  assign n3117 = x163 & ~n1373 ;
  assign n3118 = ( n1467 & n3116 ) | ( n1467 & n3117 ) | ( n3116 & n3117 ) ;
  assign n3119 = ( ~n1487 & n3116 ) | ( ~n1487 & n3117 ) | ( n3116 & n3117 ) ;
  assign n3120 = ( n1358 & n3118 ) | ( n1358 & n3119 ) | ( n3118 & n3119 ) ;
  assign n3121 = ( ~n1506 & n3118 ) | ( ~n1506 & n3119 ) | ( n3118 & n3119 ) ;
  assign n3122 = ( ~n1612 & n3120 ) | ( ~n1612 & n3121 ) | ( n3120 & n3121 ) ;
  assign n3123 = x35 & ~n1370 ;
  assign n3124 = x35 & n1373 ;
  assign n3125 = ( ~n1467 & n3123 ) | ( ~n1467 & n3124 ) | ( n3123 & n3124 ) ;
  assign n3126 = ( n1487 & n3123 ) | ( n1487 & n3124 ) | ( n3123 & n3124 ) ;
  assign n3127 = ( ~n1358 & n3125 ) | ( ~n1358 & n3126 ) | ( n3125 & n3126 ) ;
  assign n3128 = ( n1506 & n3125 ) | ( n1506 & n3126 ) | ( n3125 & n3126 ) ;
  assign n3129 = ( n1612 & n3127 ) | ( n1612 & n3128 ) | ( n3127 & n3128 ) ;
  assign n3130 = n3122 | n3129 ;
  assign n3131 = x419 & n812 ;
  assign n3132 = x419 & ~n815 ;
  assign n3133 = ( n909 & n3131 ) | ( n909 & n3132 ) | ( n3131 & n3132 ) ;
  assign n3134 = ( ~n929 & n3131 ) | ( ~n929 & n3132 ) | ( n3131 & n3132 ) ;
  assign n3135 = ( n800 & n3133 ) | ( n800 & n3134 ) | ( n3133 & n3134 ) ;
  assign n3136 = ( ~n948 & n3133 ) | ( ~n948 & n3134 ) | ( n3133 & n3134 ) ;
  assign n3137 = ( ~n1061 & n3135 ) | ( ~n1061 & n3136 ) | ( n3135 & n3136 ) ;
  assign n3138 = x291 & ~n812 ;
  assign n3139 = x291 & n815 ;
  assign n3140 = ( ~n909 & n3138 ) | ( ~n909 & n3139 ) | ( n3138 & n3139 ) ;
  assign n3141 = ( n929 & n3138 ) | ( n929 & n3139 ) | ( n3138 & n3139 ) ;
  assign n3142 = ( ~n800 & n3140 ) | ( ~n800 & n3141 ) | ( n3140 & n3141 ) ;
  assign n3143 = ( n948 & n3140 ) | ( n948 & n3141 ) | ( n3140 & n3141 ) ;
  assign n3144 = ( n1061 & n3142 ) | ( n1061 & n3143 ) | ( n3142 & n3143 ) ;
  assign n3145 = n3137 | n3144 ;
  assign n3146 = ~n3130 & n3145 ;
  assign n3147 = x418 & n812 ;
  assign n3148 = x418 & ~n815 ;
  assign n3149 = ( n909 & n3147 ) | ( n909 & n3148 ) | ( n3147 & n3148 ) ;
  assign n3150 = ( ~n929 & n3147 ) | ( ~n929 & n3148 ) | ( n3147 & n3148 ) ;
  assign n3151 = ( n800 & n3149 ) | ( n800 & n3150 ) | ( n3149 & n3150 ) ;
  assign n3152 = ( ~n948 & n3149 ) | ( ~n948 & n3150 ) | ( n3149 & n3150 ) ;
  assign n3153 = ( ~n1061 & n3151 ) | ( ~n1061 & n3152 ) | ( n3151 & n3152 ) ;
  assign n3154 = x290 & ~n812 ;
  assign n3155 = x290 & n815 ;
  assign n3156 = ( ~n909 & n3154 ) | ( ~n909 & n3155 ) | ( n3154 & n3155 ) ;
  assign n3157 = ( n929 & n3154 ) | ( n929 & n3155 ) | ( n3154 & n3155 ) ;
  assign n3158 = ( ~n800 & n3156 ) | ( ~n800 & n3157 ) | ( n3156 & n3157 ) ;
  assign n3159 = ( n948 & n3156 ) | ( n948 & n3157 ) | ( n3156 & n3157 ) ;
  assign n3160 = ( n1061 & n3158 ) | ( n1061 & n3159 ) | ( n3158 & n3159 ) ;
  assign n3161 = n3153 | n3160 ;
  assign n3162 = x162 & n1370 ;
  assign n3163 = x162 & ~n1373 ;
  assign n3164 = ( n1467 & n3162 ) | ( n1467 & n3163 ) | ( n3162 & n3163 ) ;
  assign n3165 = ( ~n1487 & n3162 ) | ( ~n1487 & n3163 ) | ( n3162 & n3163 ) ;
  assign n3166 = ( n1358 & n3164 ) | ( n1358 & n3165 ) | ( n3164 & n3165 ) ;
  assign n3167 = ( ~n1506 & n3164 ) | ( ~n1506 & n3165 ) | ( n3164 & n3165 ) ;
  assign n3168 = ( ~n1612 & n3166 ) | ( ~n1612 & n3167 ) | ( n3166 & n3167 ) ;
  assign n3169 = x34 & ~n1370 ;
  assign n3170 = x34 & n1373 ;
  assign n3171 = ( ~n1467 & n3169 ) | ( ~n1467 & n3170 ) | ( n3169 & n3170 ) ;
  assign n3172 = ( n1487 & n3169 ) | ( n1487 & n3170 ) | ( n3169 & n3170 ) ;
  assign n3173 = ( ~n1358 & n3171 ) | ( ~n1358 & n3172 ) | ( n3171 & n3172 ) ;
  assign n3174 = ( n1506 & n3171 ) | ( n1506 & n3172 ) | ( n3171 & n3172 ) ;
  assign n3175 = ( n1612 & n3173 ) | ( n1612 & n3174 ) | ( n3173 & n3174 ) ;
  assign n3176 = n3168 | n3175 ;
  assign n3177 = n3161 & ~n3176 ;
  assign n3178 = n3146 | n3177 ;
  assign n3179 = n3115 | n3178 ;
  assign n3180 = n3084 | n3179 ;
  assign n3181 = n2957 | n3180 ;
  assign n3182 = x159 & n1370 ;
  assign n3183 = x159 & ~n1373 ;
  assign n3184 = ( n1467 & n3182 ) | ( n1467 & n3183 ) | ( n3182 & n3183 ) ;
  assign n3185 = ( ~n1487 & n3182 ) | ( ~n1487 & n3183 ) | ( n3182 & n3183 ) ;
  assign n3186 = ( n1358 & n3184 ) | ( n1358 & n3185 ) | ( n3184 & n3185 ) ;
  assign n3187 = ( ~n1506 & n3184 ) | ( ~n1506 & n3185 ) | ( n3184 & n3185 ) ;
  assign n3188 = ( ~n1612 & n3186 ) | ( ~n1612 & n3187 ) | ( n3186 & n3187 ) ;
  assign n3189 = x31 & ~n1370 ;
  assign n3190 = x31 & n1373 ;
  assign n3191 = ( ~n1467 & n3189 ) | ( ~n1467 & n3190 ) | ( n3189 & n3190 ) ;
  assign n3192 = ( n1487 & n3189 ) | ( n1487 & n3190 ) | ( n3189 & n3190 ) ;
  assign n3193 = ( ~n1358 & n3191 ) | ( ~n1358 & n3192 ) | ( n3191 & n3192 ) ;
  assign n3194 = ( n1506 & n3191 ) | ( n1506 & n3192 ) | ( n3191 & n3192 ) ;
  assign n3195 = ( n1612 & n3193 ) | ( n1612 & n3194 ) | ( n3193 & n3194 ) ;
  assign n3196 = n3188 | n3195 ;
  assign n3197 = x415 & n812 ;
  assign n3198 = x415 & ~n815 ;
  assign n3199 = ( n909 & n3197 ) | ( n909 & n3198 ) | ( n3197 & n3198 ) ;
  assign n3200 = ( ~n929 & n3197 ) | ( ~n929 & n3198 ) | ( n3197 & n3198 ) ;
  assign n3201 = ( n800 & n3199 ) | ( n800 & n3200 ) | ( n3199 & n3200 ) ;
  assign n3202 = ( ~n948 & n3199 ) | ( ~n948 & n3200 ) | ( n3199 & n3200 ) ;
  assign n3203 = ( ~n1061 & n3201 ) | ( ~n1061 & n3202 ) | ( n3201 & n3202 ) ;
  assign n3204 = x287 & ~n812 ;
  assign n3205 = x287 & n815 ;
  assign n3206 = ( ~n909 & n3204 ) | ( ~n909 & n3205 ) | ( n3204 & n3205 ) ;
  assign n3207 = ( n929 & n3204 ) | ( n929 & n3205 ) | ( n3204 & n3205 ) ;
  assign n3208 = ( ~n800 & n3206 ) | ( ~n800 & n3207 ) | ( n3206 & n3207 ) ;
  assign n3209 = ( n948 & n3206 ) | ( n948 & n3207 ) | ( n3206 & n3207 ) ;
  assign n3210 = ( n1061 & n3208 ) | ( n1061 & n3209 ) | ( n3208 & n3209 ) ;
  assign n3211 = n3203 | n3210 ;
  assign n3212 = n3196 & ~n3211 ;
  assign n3213 = ~n3196 & n3211 ;
  assign n3214 = x158 & n1370 ;
  assign n3215 = x158 & ~n1373 ;
  assign n3216 = ( n1467 & n3214 ) | ( n1467 & n3215 ) | ( n3214 & n3215 ) ;
  assign n3217 = ( ~n1487 & n3214 ) | ( ~n1487 & n3215 ) | ( n3214 & n3215 ) ;
  assign n3218 = ( n1358 & n3216 ) | ( n1358 & n3217 ) | ( n3216 & n3217 ) ;
  assign n3219 = ( ~n1506 & n3216 ) | ( ~n1506 & n3217 ) | ( n3216 & n3217 ) ;
  assign n3220 = ( ~n1612 & n3218 ) | ( ~n1612 & n3219 ) | ( n3218 & n3219 ) ;
  assign n3221 = x30 & ~n1370 ;
  assign n3222 = x30 & n1373 ;
  assign n3223 = ( ~n1467 & n3221 ) | ( ~n1467 & n3222 ) | ( n3221 & n3222 ) ;
  assign n3224 = ( n1487 & n3221 ) | ( n1487 & n3222 ) | ( n3221 & n3222 ) ;
  assign n3225 = ( ~n1358 & n3223 ) | ( ~n1358 & n3224 ) | ( n3223 & n3224 ) ;
  assign n3226 = ( n1506 & n3223 ) | ( n1506 & n3224 ) | ( n3223 & n3224 ) ;
  assign n3227 = ( n1612 & n3225 ) | ( n1612 & n3226 ) | ( n3225 & n3226 ) ;
  assign n3228 = n3220 | n3227 ;
  assign n3229 = x414 & n812 ;
  assign n3230 = x414 & ~n815 ;
  assign n3231 = ( n909 & n3229 ) | ( n909 & n3230 ) | ( n3229 & n3230 ) ;
  assign n3232 = ( ~n929 & n3229 ) | ( ~n929 & n3230 ) | ( n3229 & n3230 ) ;
  assign n3233 = ( n800 & n3231 ) | ( n800 & n3232 ) | ( n3231 & n3232 ) ;
  assign n3234 = ( ~n948 & n3231 ) | ( ~n948 & n3232 ) | ( n3231 & n3232 ) ;
  assign n3235 = ( ~n1061 & n3233 ) | ( ~n1061 & n3234 ) | ( n3233 & n3234 ) ;
  assign n3236 = x286 & ~n812 ;
  assign n3237 = x286 & n815 ;
  assign n3238 = ( ~n909 & n3236 ) | ( ~n909 & n3237 ) | ( n3236 & n3237 ) ;
  assign n3239 = ( n929 & n3236 ) | ( n929 & n3237 ) | ( n3236 & n3237 ) ;
  assign n3240 = ( ~n800 & n3238 ) | ( ~n800 & n3239 ) | ( n3238 & n3239 ) ;
  assign n3241 = ( n948 & n3238 ) | ( n948 & n3239 ) | ( n3238 & n3239 ) ;
  assign n3242 = ( n1061 & n3240 ) | ( n1061 & n3241 ) | ( n3240 & n3241 ) ;
  assign n3243 = n3235 | n3242 ;
  assign n3244 = n3228 & ~n3243 ;
  assign n3245 = ~n3213 & n3244 ;
  assign n3246 = x156 & n1370 ;
  assign n3247 = x156 & ~n1373 ;
  assign n3248 = ( n1467 & n3246 ) | ( n1467 & n3247 ) | ( n3246 & n3247 ) ;
  assign n3249 = ( ~n1487 & n3246 ) | ( ~n1487 & n3247 ) | ( n3246 & n3247 ) ;
  assign n3250 = ( n1358 & n3248 ) | ( n1358 & n3249 ) | ( n3248 & n3249 ) ;
  assign n3251 = ( ~n1506 & n3248 ) | ( ~n1506 & n3249 ) | ( n3248 & n3249 ) ;
  assign n3252 = ( ~n1612 & n3250 ) | ( ~n1612 & n3251 ) | ( n3250 & n3251 ) ;
  assign n3253 = x28 & ~n1370 ;
  assign n3254 = x28 & n1373 ;
  assign n3255 = ( ~n1467 & n3253 ) | ( ~n1467 & n3254 ) | ( n3253 & n3254 ) ;
  assign n3256 = ( n1487 & n3253 ) | ( n1487 & n3254 ) | ( n3253 & n3254 ) ;
  assign n3257 = ( ~n1358 & n3255 ) | ( ~n1358 & n3256 ) | ( n3255 & n3256 ) ;
  assign n3258 = ( n1506 & n3255 ) | ( n1506 & n3256 ) | ( n3255 & n3256 ) ;
  assign n3259 = ( n1612 & n3257 ) | ( n1612 & n3258 ) | ( n3257 & n3258 ) ;
  assign n3260 = n3252 | n3259 ;
  assign n3261 = x412 & n812 ;
  assign n3262 = x412 & ~n815 ;
  assign n3263 = ( n909 & n3261 ) | ( n909 & n3262 ) | ( n3261 & n3262 ) ;
  assign n3264 = ( ~n929 & n3261 ) | ( ~n929 & n3262 ) | ( n3261 & n3262 ) ;
  assign n3265 = ( n800 & n3263 ) | ( n800 & n3264 ) | ( n3263 & n3264 ) ;
  assign n3266 = ( ~n948 & n3263 ) | ( ~n948 & n3264 ) | ( n3263 & n3264 ) ;
  assign n3267 = ( ~n1061 & n3265 ) | ( ~n1061 & n3266 ) | ( n3265 & n3266 ) ;
  assign n3268 = x284 & ~n812 ;
  assign n3269 = x284 & n815 ;
  assign n3270 = ( ~n909 & n3268 ) | ( ~n909 & n3269 ) | ( n3268 & n3269 ) ;
  assign n3271 = ( n929 & n3268 ) | ( n929 & n3269 ) | ( n3268 & n3269 ) ;
  assign n3272 = ( ~n800 & n3270 ) | ( ~n800 & n3271 ) | ( n3270 & n3271 ) ;
  assign n3273 = ( n948 & n3270 ) | ( n948 & n3271 ) | ( n3270 & n3271 ) ;
  assign n3274 = ( n1061 & n3272 ) | ( n1061 & n3273 ) | ( n3272 & n3273 ) ;
  assign n3275 = n3267 | n3274 ;
  assign n3276 = ~n3260 & n3275 ;
  assign n3277 = x155 & n1370 ;
  assign n3278 = x155 & ~n1373 ;
  assign n3279 = ( n1467 & n3277 ) | ( n1467 & n3278 ) | ( n3277 & n3278 ) ;
  assign n3280 = ( ~n1487 & n3277 ) | ( ~n1487 & n3278 ) | ( n3277 & n3278 ) ;
  assign n3281 = ( n1358 & n3279 ) | ( n1358 & n3280 ) | ( n3279 & n3280 ) ;
  assign n3282 = ( ~n1506 & n3279 ) | ( ~n1506 & n3280 ) | ( n3279 & n3280 ) ;
  assign n3283 = ( ~n1612 & n3281 ) | ( ~n1612 & n3282 ) | ( n3281 & n3282 ) ;
  assign n3284 = x27 & ~n1370 ;
  assign n3285 = x27 & n1373 ;
  assign n3286 = ( ~n1467 & n3284 ) | ( ~n1467 & n3285 ) | ( n3284 & n3285 ) ;
  assign n3287 = ( n1487 & n3284 ) | ( n1487 & n3285 ) | ( n3284 & n3285 ) ;
  assign n3288 = ( ~n1358 & n3286 ) | ( ~n1358 & n3287 ) | ( n3286 & n3287 ) ;
  assign n3289 = ( n1506 & n3286 ) | ( n1506 & n3287 ) | ( n3286 & n3287 ) ;
  assign n3290 = ( n1612 & n3288 ) | ( n1612 & n3289 ) | ( n3288 & n3289 ) ;
  assign n3291 = n3283 | n3290 ;
  assign n3292 = x411 & n812 ;
  assign n3293 = x411 & ~n815 ;
  assign n3294 = ( n909 & n3292 ) | ( n909 & n3293 ) | ( n3292 & n3293 ) ;
  assign n3295 = ( ~n929 & n3292 ) | ( ~n929 & n3293 ) | ( n3292 & n3293 ) ;
  assign n3296 = ( n800 & n3294 ) | ( n800 & n3295 ) | ( n3294 & n3295 ) ;
  assign n3297 = ( ~n948 & n3294 ) | ( ~n948 & n3295 ) | ( n3294 & n3295 ) ;
  assign n3298 = ( ~n1061 & n3296 ) | ( ~n1061 & n3297 ) | ( n3296 & n3297 ) ;
  assign n3299 = x283 & ~n812 ;
  assign n3300 = x283 & n815 ;
  assign n3301 = ( ~n909 & n3299 ) | ( ~n909 & n3300 ) | ( n3299 & n3300 ) ;
  assign n3302 = ( n929 & n3299 ) | ( n929 & n3300 ) | ( n3299 & n3300 ) ;
  assign n3303 = ( ~n800 & n3301 ) | ( ~n800 & n3302 ) | ( n3301 & n3302 ) ;
  assign n3304 = ( n948 & n3301 ) | ( n948 & n3302 ) | ( n3301 & n3302 ) ;
  assign n3305 = ( n1061 & n3303 ) | ( n1061 & n3304 ) | ( n3303 & n3304 ) ;
  assign n3306 = n3298 | n3305 ;
  assign n3307 = n3291 & ~n3306 ;
  assign n3308 = ~n3276 & n3307 ;
  assign n3309 = x154 & n1370 ;
  assign n3310 = x154 & ~n1373 ;
  assign n3311 = ( n1467 & n3309 ) | ( n1467 & n3310 ) | ( n3309 & n3310 ) ;
  assign n3312 = ( ~n1487 & n3309 ) | ( ~n1487 & n3310 ) | ( n3309 & n3310 ) ;
  assign n3313 = ( n1358 & n3311 ) | ( n1358 & n3312 ) | ( n3311 & n3312 ) ;
  assign n3314 = ( ~n1506 & n3311 ) | ( ~n1506 & n3312 ) | ( n3311 & n3312 ) ;
  assign n3315 = ( ~n1612 & n3313 ) | ( ~n1612 & n3314 ) | ( n3313 & n3314 ) ;
  assign n3316 = x26 & ~n1370 ;
  assign n3317 = x26 & n1373 ;
  assign n3318 = ( ~n1467 & n3316 ) | ( ~n1467 & n3317 ) | ( n3316 & n3317 ) ;
  assign n3319 = ( n1487 & n3316 ) | ( n1487 & n3317 ) | ( n3316 & n3317 ) ;
  assign n3320 = ( ~n1358 & n3318 ) | ( ~n1358 & n3319 ) | ( n3318 & n3319 ) ;
  assign n3321 = ( n1506 & n3318 ) | ( n1506 & n3319 ) | ( n3318 & n3319 ) ;
  assign n3322 = ( n1612 & n3320 ) | ( n1612 & n3321 ) | ( n3320 & n3321 ) ;
  assign n3323 = n3315 | n3322 ;
  assign n3324 = x410 & n812 ;
  assign n3325 = x410 & ~n815 ;
  assign n3326 = ( n909 & n3324 ) | ( n909 & n3325 ) | ( n3324 & n3325 ) ;
  assign n3327 = ( ~n929 & n3324 ) | ( ~n929 & n3325 ) | ( n3324 & n3325 ) ;
  assign n3328 = ( n800 & n3326 ) | ( n800 & n3327 ) | ( n3326 & n3327 ) ;
  assign n3329 = ( ~n948 & n3326 ) | ( ~n948 & n3327 ) | ( n3326 & n3327 ) ;
  assign n3330 = ( ~n1061 & n3328 ) | ( ~n1061 & n3329 ) | ( n3328 & n3329 ) ;
  assign n3331 = x282 & ~n812 ;
  assign n3332 = x282 & n815 ;
  assign n3333 = ( ~n909 & n3331 ) | ( ~n909 & n3332 ) | ( n3331 & n3332 ) ;
  assign n3334 = ( n929 & n3331 ) | ( n929 & n3332 ) | ( n3331 & n3332 ) ;
  assign n3335 = ( ~n800 & n3333 ) | ( ~n800 & n3334 ) | ( n3333 & n3334 ) ;
  assign n3336 = ( n948 & n3333 ) | ( n948 & n3334 ) | ( n3333 & n3334 ) ;
  assign n3337 = ( n1061 & n3335 ) | ( n1061 & n3336 ) | ( n3335 & n3336 ) ;
  assign n3338 = n3330 | n3337 ;
  assign n3339 = n3323 & ~n3338 ;
  assign n3340 = ~n3323 & n3338 ;
  assign n3341 = ( ~n3291 & n3306 ) | ( ~n3291 & n3340 ) | ( n3306 & n3340 ) ;
  assign n3342 = n3339 & ~n3341 ;
  assign n3343 = ( ~n3276 & n3308 ) | ( ~n3276 & n3342 ) | ( n3308 & n3342 ) ;
  assign n3344 = x157 & n1370 ;
  assign n3345 = x157 & ~n1373 ;
  assign n3346 = ( n1467 & n3344 ) | ( n1467 & n3345 ) | ( n3344 & n3345 ) ;
  assign n3347 = ( ~n1487 & n3344 ) | ( ~n1487 & n3345 ) | ( n3344 & n3345 ) ;
  assign n3348 = ( n1358 & n3346 ) | ( n1358 & n3347 ) | ( n3346 & n3347 ) ;
  assign n3349 = ( ~n1506 & n3346 ) | ( ~n1506 & n3347 ) | ( n3346 & n3347 ) ;
  assign n3350 = ( ~n1612 & n3348 ) | ( ~n1612 & n3349 ) | ( n3348 & n3349 ) ;
  assign n3351 = x29 & ~n1370 ;
  assign n3352 = x29 & n1373 ;
  assign n3353 = ( ~n1467 & n3351 ) | ( ~n1467 & n3352 ) | ( n3351 & n3352 ) ;
  assign n3354 = ( n1487 & n3351 ) | ( n1487 & n3352 ) | ( n3351 & n3352 ) ;
  assign n3355 = ( ~n1358 & n3353 ) | ( ~n1358 & n3354 ) | ( n3353 & n3354 ) ;
  assign n3356 = ( n1506 & n3353 ) | ( n1506 & n3354 ) | ( n3353 & n3354 ) ;
  assign n3357 = ( n1612 & n3355 ) | ( n1612 & n3356 ) | ( n3355 & n3356 ) ;
  assign n3358 = n3350 | n3357 ;
  assign n3359 = x413 & n812 ;
  assign n3360 = x413 & ~n815 ;
  assign n3361 = ( n909 & n3359 ) | ( n909 & n3360 ) | ( n3359 & n3360 ) ;
  assign n3362 = ( ~n929 & n3359 ) | ( ~n929 & n3360 ) | ( n3359 & n3360 ) ;
  assign n3363 = ( n800 & n3361 ) | ( n800 & n3362 ) | ( n3361 & n3362 ) ;
  assign n3364 = ( ~n948 & n3361 ) | ( ~n948 & n3362 ) | ( n3361 & n3362 ) ;
  assign n3365 = ( ~n1061 & n3363 ) | ( ~n1061 & n3364 ) | ( n3363 & n3364 ) ;
  assign n3366 = x285 & ~n812 ;
  assign n3367 = x285 & n815 ;
  assign n3368 = ( ~n909 & n3366 ) | ( ~n909 & n3367 ) | ( n3366 & n3367 ) ;
  assign n3369 = ( n929 & n3366 ) | ( n929 & n3367 ) | ( n3366 & n3367 ) ;
  assign n3370 = ( ~n800 & n3368 ) | ( ~n800 & n3369 ) | ( n3368 & n3369 ) ;
  assign n3371 = ( n948 & n3368 ) | ( n948 & n3369 ) | ( n3368 & n3369 ) ;
  assign n3372 = ( n1061 & n3370 ) | ( n1061 & n3371 ) | ( n3370 & n3371 ) ;
  assign n3373 = n3365 | n3372 ;
  assign n3374 = ~n3358 & n3373 ;
  assign n3375 = n3358 & ~n3373 ;
  assign n3376 = n3260 & ~n3275 ;
  assign n3377 = ~n3374 & n3376 ;
  assign n3378 = n3375 | n3377 ;
  assign n3379 = ( n3343 & ~n3374 ) | ( n3343 & n3378 ) | ( ~n3374 & n3378 ) ;
  assign n3380 = ~n3228 & n3243 ;
  assign n3381 = n3213 | n3380 ;
  assign n3382 = ( n3245 & n3379 ) | ( n3245 & ~n3381 ) | ( n3379 & ~n3381 ) ;
  assign n3383 = n3212 | n3382 ;
  assign n3384 = ~n3181 & n3383 ;
  assign n3385 = ~n3161 & n3176 ;
  assign n3386 = ~n3146 & n3385 ;
  assign n3387 = ~n2941 & n2956 ;
  assign n3388 = n3099 & ~n3114 ;
  assign n3389 = n3387 | n3388 ;
  assign n3390 = n3386 | n3389 ;
  assign n3391 = ( ~n3179 & n3386 ) | ( ~n3179 & n3390 ) | ( n3386 & n3390 ) ;
  assign n3392 = n3130 & ~n3145 ;
  assign n3393 = ~n3084 & n3392 ;
  assign n3394 = ( ~n3084 & n3391 ) | ( ~n3084 & n3393 ) | ( n3391 & n3393 ) ;
  assign n3395 = n3035 & ~n3050 ;
  assign n3396 = ( n3066 & ~n3081 ) | ( n3066 & n3395 ) | ( ~n3081 & n3395 ) ;
  assign n3397 = ( ~n3003 & n3018 ) | ( ~n3003 & n3396 ) | ( n3018 & n3396 ) ;
  assign n3398 = ( n2972 & ~n2987 ) | ( n2972 & n3397 ) | ( ~n2987 & n3397 ) ;
  assign n3399 = n3394 | n3398 ;
  assign n3400 = n3384 | n3399 ;
  assign n3401 = ~n2840 & n2855 ;
  assign n3402 = ~n2810 & n2825 ;
  assign n3403 = n3401 | n3402 ;
  assign n3404 = ~n2870 & n2885 ;
  assign n3405 = ~n2900 & n2915 ;
  assign n3406 = n3404 | n3405 ;
  assign n3407 = n3403 | n3406 ;
  assign n3408 = n2795 | n3407 ;
  assign n3409 = ( n2926 & n3400 ) | ( n2926 & ~n3408 ) | ( n3400 & ~n3408 ) ;
  assign n3410 = n2926 | n3409 ;
  assign n3411 = n2920 | n3410 ;
  assign n3412 = ( n2697 & ~n2698 ) | ( n2697 & n3411 ) | ( ~n2698 & n3411 ) ;
  assign n3413 = x209 & n1370 ;
  assign n3414 = x209 & ~n1373 ;
  assign n3415 = ( n1467 & n3413 ) | ( n1467 & n3414 ) | ( n3413 & n3414 ) ;
  assign n3416 = ( ~n1487 & n3413 ) | ( ~n1487 & n3414 ) | ( n3413 & n3414 ) ;
  assign n3417 = ( n1358 & n3415 ) | ( n1358 & n3416 ) | ( n3415 & n3416 ) ;
  assign n3418 = ( ~n1506 & n3415 ) | ( ~n1506 & n3416 ) | ( n3415 & n3416 ) ;
  assign n3419 = ( ~n1612 & n3417 ) | ( ~n1612 & n3418 ) | ( n3417 & n3418 ) ;
  assign n3420 = x81 & ~n1370 ;
  assign n3421 = x81 & n1373 ;
  assign n3422 = ( ~n1467 & n3420 ) | ( ~n1467 & n3421 ) | ( n3420 & n3421 ) ;
  assign n3423 = ( n1487 & n3420 ) | ( n1487 & n3421 ) | ( n3420 & n3421 ) ;
  assign n3424 = ( ~n1358 & n3422 ) | ( ~n1358 & n3423 ) | ( n3422 & n3423 ) ;
  assign n3425 = ( n1506 & n3422 ) | ( n1506 & n3423 ) | ( n3422 & n3423 ) ;
  assign n3426 = ( n1612 & n3424 ) | ( n1612 & n3425 ) | ( n3424 & n3425 ) ;
  assign n3427 = n3419 | n3426 ;
  assign n3428 = x465 & n812 ;
  assign n3429 = x465 & ~n815 ;
  assign n3430 = ( n909 & n3428 ) | ( n909 & n3429 ) | ( n3428 & n3429 ) ;
  assign n3431 = ( ~n929 & n3428 ) | ( ~n929 & n3429 ) | ( n3428 & n3429 ) ;
  assign n3432 = ( n800 & n3430 ) | ( n800 & n3431 ) | ( n3430 & n3431 ) ;
  assign n3433 = ( ~n948 & n3430 ) | ( ~n948 & n3431 ) | ( n3430 & n3431 ) ;
  assign n3434 = ( ~n1061 & n3432 ) | ( ~n1061 & n3433 ) | ( n3432 & n3433 ) ;
  assign n3435 = x337 & ~n812 ;
  assign n3436 = x337 & n815 ;
  assign n3437 = ( ~n909 & n3435 ) | ( ~n909 & n3436 ) | ( n3435 & n3436 ) ;
  assign n3438 = ( n929 & n3435 ) | ( n929 & n3436 ) | ( n3435 & n3436 ) ;
  assign n3439 = ( ~n800 & n3437 ) | ( ~n800 & n3438 ) | ( n3437 & n3438 ) ;
  assign n3440 = ( n948 & n3437 ) | ( n948 & n3438 ) | ( n3437 & n3438 ) ;
  assign n3441 = ( n1061 & n3439 ) | ( n1061 & n3440 ) | ( n3439 & n3440 ) ;
  assign n3442 = n3434 | n3441 ;
  assign n3443 = ~n3427 & n3442 ;
  assign n3444 = x199 & n1370 ;
  assign n3445 = x199 & ~n1373 ;
  assign n3446 = ( n1467 & n3444 ) | ( n1467 & n3445 ) | ( n3444 & n3445 ) ;
  assign n3447 = ( ~n1487 & n3444 ) | ( ~n1487 & n3445 ) | ( n3444 & n3445 ) ;
  assign n3448 = ( n1358 & n3446 ) | ( n1358 & n3447 ) | ( n3446 & n3447 ) ;
  assign n3449 = ( ~n1506 & n3446 ) | ( ~n1506 & n3447 ) | ( n3446 & n3447 ) ;
  assign n3450 = ( ~n1612 & n3448 ) | ( ~n1612 & n3449 ) | ( n3448 & n3449 ) ;
  assign n3451 = x71 & ~n1370 ;
  assign n3452 = x71 & n1373 ;
  assign n3453 = ( ~n1467 & n3451 ) | ( ~n1467 & n3452 ) | ( n3451 & n3452 ) ;
  assign n3454 = ( n1487 & n3451 ) | ( n1487 & n3452 ) | ( n3451 & n3452 ) ;
  assign n3455 = ( ~n1358 & n3453 ) | ( ~n1358 & n3454 ) | ( n3453 & n3454 ) ;
  assign n3456 = ( n1506 & n3453 ) | ( n1506 & n3454 ) | ( n3453 & n3454 ) ;
  assign n3457 = ( n1612 & n3455 ) | ( n1612 & n3456 ) | ( n3455 & n3456 ) ;
  assign n3458 = n3450 | n3457 ;
  assign n3459 = x455 & n812 ;
  assign n3460 = x455 & ~n815 ;
  assign n3461 = ( n909 & n3459 ) | ( n909 & n3460 ) | ( n3459 & n3460 ) ;
  assign n3462 = ( ~n929 & n3459 ) | ( ~n929 & n3460 ) | ( n3459 & n3460 ) ;
  assign n3463 = ( n800 & n3461 ) | ( n800 & n3462 ) | ( n3461 & n3462 ) ;
  assign n3464 = ( ~n948 & n3461 ) | ( ~n948 & n3462 ) | ( n3461 & n3462 ) ;
  assign n3465 = ( ~n1061 & n3463 ) | ( ~n1061 & n3464 ) | ( n3463 & n3464 ) ;
  assign n3466 = x327 & ~n812 ;
  assign n3467 = x327 & n815 ;
  assign n3468 = ( ~n909 & n3466 ) | ( ~n909 & n3467 ) | ( n3466 & n3467 ) ;
  assign n3469 = ( n929 & n3466 ) | ( n929 & n3467 ) | ( n3466 & n3467 ) ;
  assign n3470 = ( ~n800 & n3468 ) | ( ~n800 & n3469 ) | ( n3468 & n3469 ) ;
  assign n3471 = ( n948 & n3468 ) | ( n948 & n3469 ) | ( n3468 & n3469 ) ;
  assign n3472 = ( n1061 & n3470 ) | ( n1061 & n3471 ) | ( n3470 & n3471 ) ;
  assign n3473 = n3465 | n3472 ;
  assign n3474 = ~n3458 & n3473 ;
  assign n3475 = x454 & n812 ;
  assign n3476 = x454 & ~n815 ;
  assign n3477 = ( n909 & n3475 ) | ( n909 & n3476 ) | ( n3475 & n3476 ) ;
  assign n3478 = ( ~n929 & n3475 ) | ( ~n929 & n3476 ) | ( n3475 & n3476 ) ;
  assign n3479 = ( n800 & n3477 ) | ( n800 & n3478 ) | ( n3477 & n3478 ) ;
  assign n3480 = ( ~n948 & n3477 ) | ( ~n948 & n3478 ) | ( n3477 & n3478 ) ;
  assign n3481 = ( ~n1061 & n3479 ) | ( ~n1061 & n3480 ) | ( n3479 & n3480 ) ;
  assign n3482 = x326 & ~n812 ;
  assign n3483 = x326 & n815 ;
  assign n3484 = ( ~n909 & n3482 ) | ( ~n909 & n3483 ) | ( n3482 & n3483 ) ;
  assign n3485 = ( n929 & n3482 ) | ( n929 & n3483 ) | ( n3482 & n3483 ) ;
  assign n3486 = ( ~n800 & n3484 ) | ( ~n800 & n3485 ) | ( n3484 & n3485 ) ;
  assign n3487 = ( n948 & n3484 ) | ( n948 & n3485 ) | ( n3484 & n3485 ) ;
  assign n3488 = ( n1061 & n3486 ) | ( n1061 & n3487 ) | ( n3486 & n3487 ) ;
  assign n3489 = n3481 | n3488 ;
  assign n3490 = x198 & n1370 ;
  assign n3491 = x198 & ~n1373 ;
  assign n3492 = ( n1467 & n3490 ) | ( n1467 & n3491 ) | ( n3490 & n3491 ) ;
  assign n3493 = ( ~n1487 & n3490 ) | ( ~n1487 & n3491 ) | ( n3490 & n3491 ) ;
  assign n3494 = ( n1358 & n3492 ) | ( n1358 & n3493 ) | ( n3492 & n3493 ) ;
  assign n3495 = ( ~n1506 & n3492 ) | ( ~n1506 & n3493 ) | ( n3492 & n3493 ) ;
  assign n3496 = ( ~n1612 & n3494 ) | ( ~n1612 & n3495 ) | ( n3494 & n3495 ) ;
  assign n3497 = x70 & ~n1370 ;
  assign n3498 = x70 & n1373 ;
  assign n3499 = ( ~n1467 & n3497 ) | ( ~n1467 & n3498 ) | ( n3497 & n3498 ) ;
  assign n3500 = ( n1487 & n3497 ) | ( n1487 & n3498 ) | ( n3497 & n3498 ) ;
  assign n3501 = ( ~n1358 & n3499 ) | ( ~n1358 & n3500 ) | ( n3499 & n3500 ) ;
  assign n3502 = ( n1506 & n3499 ) | ( n1506 & n3500 ) | ( n3499 & n3500 ) ;
  assign n3503 = ( n1612 & n3501 ) | ( n1612 & n3502 ) | ( n3501 & n3502 ) ;
  assign n3504 = n3496 | n3503 ;
  assign n3505 = ~n3489 & n3504 ;
  assign n3506 = ~n3474 & n3505 ;
  assign n3507 = n3489 & ~n3504 ;
  assign n3508 = n3474 | n3507 ;
  assign n3509 = x197 & n1370 ;
  assign n3510 = x197 & ~n1373 ;
  assign n3511 = ( n1467 & n3509 ) | ( n1467 & n3510 ) | ( n3509 & n3510 ) ;
  assign n3512 = ( ~n1487 & n3509 ) | ( ~n1487 & n3510 ) | ( n3509 & n3510 ) ;
  assign n3513 = ( n1358 & n3511 ) | ( n1358 & n3512 ) | ( n3511 & n3512 ) ;
  assign n3514 = ( ~n1506 & n3511 ) | ( ~n1506 & n3512 ) | ( n3511 & n3512 ) ;
  assign n3515 = ( ~n1612 & n3513 ) | ( ~n1612 & n3514 ) | ( n3513 & n3514 ) ;
  assign n3516 = x69 & ~n1370 ;
  assign n3517 = x69 & n1373 ;
  assign n3518 = ( ~n1467 & n3516 ) | ( ~n1467 & n3517 ) | ( n3516 & n3517 ) ;
  assign n3519 = ( n1487 & n3516 ) | ( n1487 & n3517 ) | ( n3516 & n3517 ) ;
  assign n3520 = ( ~n1358 & n3518 ) | ( ~n1358 & n3519 ) | ( n3518 & n3519 ) ;
  assign n3521 = ( n1506 & n3518 ) | ( n1506 & n3519 ) | ( n3518 & n3519 ) ;
  assign n3522 = ( n1612 & n3520 ) | ( n1612 & n3521 ) | ( n3520 & n3521 ) ;
  assign n3523 = n3515 | n3522 ;
  assign n3524 = x453 & n812 ;
  assign n3525 = x453 & ~n815 ;
  assign n3526 = ( n909 & n3524 ) | ( n909 & n3525 ) | ( n3524 & n3525 ) ;
  assign n3527 = ( ~n929 & n3524 ) | ( ~n929 & n3525 ) | ( n3524 & n3525 ) ;
  assign n3528 = ( n800 & n3526 ) | ( n800 & n3527 ) | ( n3526 & n3527 ) ;
  assign n3529 = ( ~n948 & n3526 ) | ( ~n948 & n3527 ) | ( n3526 & n3527 ) ;
  assign n3530 = ( ~n1061 & n3528 ) | ( ~n1061 & n3529 ) | ( n3528 & n3529 ) ;
  assign n3531 = x325 & ~n812 ;
  assign n3532 = x325 & n815 ;
  assign n3533 = ( ~n909 & n3531 ) | ( ~n909 & n3532 ) | ( n3531 & n3532 ) ;
  assign n3534 = ( n929 & n3531 ) | ( n929 & n3532 ) | ( n3531 & n3532 ) ;
  assign n3535 = ( ~n800 & n3533 ) | ( ~n800 & n3534 ) | ( n3533 & n3534 ) ;
  assign n3536 = ( n948 & n3533 ) | ( n948 & n3534 ) | ( n3533 & n3534 ) ;
  assign n3537 = ( n1061 & n3535 ) | ( n1061 & n3536 ) | ( n3535 & n3536 ) ;
  assign n3538 = n3530 | n3537 ;
  assign n3539 = ~n3523 & n3538 ;
  assign n3540 = x196 & n1370 ;
  assign n3541 = x196 & ~n1373 ;
  assign n3542 = ( n1467 & n3540 ) | ( n1467 & n3541 ) | ( n3540 & n3541 ) ;
  assign n3543 = ( ~n1487 & n3540 ) | ( ~n1487 & n3541 ) | ( n3540 & n3541 ) ;
  assign n3544 = ( n1358 & n3542 ) | ( n1358 & n3543 ) | ( n3542 & n3543 ) ;
  assign n3545 = ( ~n1506 & n3542 ) | ( ~n1506 & n3543 ) | ( n3542 & n3543 ) ;
  assign n3546 = ( ~n1612 & n3544 ) | ( ~n1612 & n3545 ) | ( n3544 & n3545 ) ;
  assign n3547 = x68 & ~n1370 ;
  assign n3548 = x68 & n1373 ;
  assign n3549 = ( ~n1467 & n3547 ) | ( ~n1467 & n3548 ) | ( n3547 & n3548 ) ;
  assign n3550 = ( n1487 & n3547 ) | ( n1487 & n3548 ) | ( n3547 & n3548 ) ;
  assign n3551 = ( ~n1358 & n3549 ) | ( ~n1358 & n3550 ) | ( n3549 & n3550 ) ;
  assign n3552 = ( n1506 & n3549 ) | ( n1506 & n3550 ) | ( n3549 & n3550 ) ;
  assign n3553 = ( n1612 & n3551 ) | ( n1612 & n3552 ) | ( n3551 & n3552 ) ;
  assign n3554 = n3546 | n3553 ;
  assign n3555 = x452 & n812 ;
  assign n3556 = x452 & ~n815 ;
  assign n3557 = ( n909 & n3555 ) | ( n909 & n3556 ) | ( n3555 & n3556 ) ;
  assign n3558 = ( ~n929 & n3555 ) | ( ~n929 & n3556 ) | ( n3555 & n3556 ) ;
  assign n3559 = ( n800 & n3557 ) | ( n800 & n3558 ) | ( n3557 & n3558 ) ;
  assign n3560 = ( ~n948 & n3557 ) | ( ~n948 & n3558 ) | ( n3557 & n3558 ) ;
  assign n3561 = ( ~n1061 & n3559 ) | ( ~n1061 & n3560 ) | ( n3559 & n3560 ) ;
  assign n3562 = x324 & ~n812 ;
  assign n3563 = x324 & n815 ;
  assign n3564 = ( ~n909 & n3562 ) | ( ~n909 & n3563 ) | ( n3562 & n3563 ) ;
  assign n3565 = ( n929 & n3562 ) | ( n929 & n3563 ) | ( n3562 & n3563 ) ;
  assign n3566 = ( ~n800 & n3564 ) | ( ~n800 & n3565 ) | ( n3564 & n3565 ) ;
  assign n3567 = ( n948 & n3564 ) | ( n948 & n3565 ) | ( n3564 & n3565 ) ;
  assign n3568 = ( n1061 & n3566 ) | ( n1061 & n3567 ) | ( n3566 & n3567 ) ;
  assign n3569 = n3561 | n3568 ;
  assign n3570 = ~n3554 & n3569 ;
  assign n3571 = n3539 | n3570 ;
  assign n3572 = n3508 | n3571 ;
  assign n3573 = x195 & n1370 ;
  assign n3574 = x195 & ~n1373 ;
  assign n3575 = ( n1467 & n3573 ) | ( n1467 & n3574 ) | ( n3573 & n3574 ) ;
  assign n3576 = ( ~n1487 & n3573 ) | ( ~n1487 & n3574 ) | ( n3573 & n3574 ) ;
  assign n3577 = ( n1358 & n3575 ) | ( n1358 & n3576 ) | ( n3575 & n3576 ) ;
  assign n3578 = ( ~n1506 & n3575 ) | ( ~n1506 & n3576 ) | ( n3575 & n3576 ) ;
  assign n3579 = ( ~n1612 & n3577 ) | ( ~n1612 & n3578 ) | ( n3577 & n3578 ) ;
  assign n3580 = x67 & ~n1370 ;
  assign n3581 = x67 & n1373 ;
  assign n3582 = ( ~n1467 & n3580 ) | ( ~n1467 & n3581 ) | ( n3580 & n3581 ) ;
  assign n3583 = ( n1487 & n3580 ) | ( n1487 & n3581 ) | ( n3580 & n3581 ) ;
  assign n3584 = ( ~n1358 & n3582 ) | ( ~n1358 & n3583 ) | ( n3582 & n3583 ) ;
  assign n3585 = ( n1506 & n3582 ) | ( n1506 & n3583 ) | ( n3582 & n3583 ) ;
  assign n3586 = ( n1612 & n3584 ) | ( n1612 & n3585 ) | ( n3584 & n3585 ) ;
  assign n3587 = n3579 | n3586 ;
  assign n3588 = x451 & n812 ;
  assign n3589 = x451 & ~n815 ;
  assign n3590 = ( n909 & n3588 ) | ( n909 & n3589 ) | ( n3588 & n3589 ) ;
  assign n3591 = ( ~n929 & n3588 ) | ( ~n929 & n3589 ) | ( n3588 & n3589 ) ;
  assign n3592 = ( n800 & n3590 ) | ( n800 & n3591 ) | ( n3590 & n3591 ) ;
  assign n3593 = ( ~n948 & n3590 ) | ( ~n948 & n3591 ) | ( n3590 & n3591 ) ;
  assign n3594 = ( ~n1061 & n3592 ) | ( ~n1061 & n3593 ) | ( n3592 & n3593 ) ;
  assign n3595 = x323 & ~n812 ;
  assign n3596 = x323 & n815 ;
  assign n3597 = ( ~n909 & n3595 ) | ( ~n909 & n3596 ) | ( n3595 & n3596 ) ;
  assign n3598 = ( n929 & n3595 ) | ( n929 & n3596 ) | ( n3595 & n3596 ) ;
  assign n3599 = ( ~n800 & n3597 ) | ( ~n800 & n3598 ) | ( n3597 & n3598 ) ;
  assign n3600 = ( n948 & n3597 ) | ( n948 & n3598 ) | ( n3597 & n3598 ) ;
  assign n3601 = ( n1061 & n3599 ) | ( n1061 & n3600 ) | ( n3599 & n3600 ) ;
  assign n3602 = n3594 | n3601 ;
  assign n3603 = ~n3587 & n3602 ;
  assign n3604 = x450 & n812 ;
  assign n3605 = x450 & ~n815 ;
  assign n3606 = ( n909 & n3604 ) | ( n909 & n3605 ) | ( n3604 & n3605 ) ;
  assign n3607 = ( ~n929 & n3604 ) | ( ~n929 & n3605 ) | ( n3604 & n3605 ) ;
  assign n3608 = ( n800 & n3606 ) | ( n800 & n3607 ) | ( n3606 & n3607 ) ;
  assign n3609 = ( ~n948 & n3606 ) | ( ~n948 & n3607 ) | ( n3606 & n3607 ) ;
  assign n3610 = ( ~n1061 & n3608 ) | ( ~n1061 & n3609 ) | ( n3608 & n3609 ) ;
  assign n3611 = x322 & ~n812 ;
  assign n3612 = x322 & n815 ;
  assign n3613 = ( ~n909 & n3611 ) | ( ~n909 & n3612 ) | ( n3611 & n3612 ) ;
  assign n3614 = ( n929 & n3611 ) | ( n929 & n3612 ) | ( n3611 & n3612 ) ;
  assign n3615 = ( ~n800 & n3613 ) | ( ~n800 & n3614 ) | ( n3613 & n3614 ) ;
  assign n3616 = ( n948 & n3613 ) | ( n948 & n3614 ) | ( n3613 & n3614 ) ;
  assign n3617 = ( n1061 & n3615 ) | ( n1061 & n3616 ) | ( n3615 & n3616 ) ;
  assign n3618 = n3610 | n3617 ;
  assign n3619 = x194 & n1370 ;
  assign n3620 = x194 & ~n1373 ;
  assign n3621 = ( n1467 & n3619 ) | ( n1467 & n3620 ) | ( n3619 & n3620 ) ;
  assign n3622 = ( ~n1487 & n3619 ) | ( ~n1487 & n3620 ) | ( n3619 & n3620 ) ;
  assign n3623 = ( n1358 & n3621 ) | ( n1358 & n3622 ) | ( n3621 & n3622 ) ;
  assign n3624 = ( ~n1506 & n3621 ) | ( ~n1506 & n3622 ) | ( n3621 & n3622 ) ;
  assign n3625 = ( ~n1612 & n3623 ) | ( ~n1612 & n3624 ) | ( n3623 & n3624 ) ;
  assign n3626 = x66 & ~n1370 ;
  assign n3627 = x66 & n1373 ;
  assign n3628 = ( ~n1467 & n3626 ) | ( ~n1467 & n3627 ) | ( n3626 & n3627 ) ;
  assign n3629 = ( n1487 & n3626 ) | ( n1487 & n3627 ) | ( n3626 & n3627 ) ;
  assign n3630 = ( ~n1358 & n3628 ) | ( ~n1358 & n3629 ) | ( n3628 & n3629 ) ;
  assign n3631 = ( n1506 & n3628 ) | ( n1506 & n3629 ) | ( n3628 & n3629 ) ;
  assign n3632 = ( n1612 & n3630 ) | ( n1612 & n3631 ) | ( n3630 & n3631 ) ;
  assign n3633 = n3625 | n3632 ;
  assign n3634 = n3618 & ~n3633 ;
  assign n3635 = n3603 | n3634 ;
  assign n3636 = x193 & n1370 ;
  assign n3637 = x193 & ~n1373 ;
  assign n3638 = ( n1467 & n3636 ) | ( n1467 & n3637 ) | ( n3636 & n3637 ) ;
  assign n3639 = ( ~n1487 & n3636 ) | ( ~n1487 & n3637 ) | ( n3636 & n3637 ) ;
  assign n3640 = ( n1358 & n3638 ) | ( n1358 & n3639 ) | ( n3638 & n3639 ) ;
  assign n3641 = ( ~n1506 & n3638 ) | ( ~n1506 & n3639 ) | ( n3638 & n3639 ) ;
  assign n3642 = ( ~n1612 & n3640 ) | ( ~n1612 & n3641 ) | ( n3640 & n3641 ) ;
  assign n3643 = x65 & ~n1370 ;
  assign n3644 = x65 & n1373 ;
  assign n3645 = ( ~n1467 & n3643 ) | ( ~n1467 & n3644 ) | ( n3643 & n3644 ) ;
  assign n3646 = ( n1487 & n3643 ) | ( n1487 & n3644 ) | ( n3643 & n3644 ) ;
  assign n3647 = ( ~n1358 & n3645 ) | ( ~n1358 & n3646 ) | ( n3645 & n3646 ) ;
  assign n3648 = ( n1506 & n3645 ) | ( n1506 & n3646 ) | ( n3645 & n3646 ) ;
  assign n3649 = ( n1612 & n3647 ) | ( n1612 & n3648 ) | ( n3647 & n3648 ) ;
  assign n3650 = n3642 | n3649 ;
  assign n3651 = x449 & n812 ;
  assign n3652 = x449 & ~n815 ;
  assign n3653 = ( n909 & n3651 ) | ( n909 & n3652 ) | ( n3651 & n3652 ) ;
  assign n3654 = ( ~n929 & n3651 ) | ( ~n929 & n3652 ) | ( n3651 & n3652 ) ;
  assign n3655 = ( n800 & n3653 ) | ( n800 & n3654 ) | ( n3653 & n3654 ) ;
  assign n3656 = ( ~n948 & n3653 ) | ( ~n948 & n3654 ) | ( n3653 & n3654 ) ;
  assign n3657 = ( ~n1061 & n3655 ) | ( ~n1061 & n3656 ) | ( n3655 & n3656 ) ;
  assign n3658 = x321 & ~n812 ;
  assign n3659 = x321 & n815 ;
  assign n3660 = ( ~n909 & n3658 ) | ( ~n909 & n3659 ) | ( n3658 & n3659 ) ;
  assign n3661 = ( n929 & n3658 ) | ( n929 & n3659 ) | ( n3658 & n3659 ) ;
  assign n3662 = ( ~n800 & n3660 ) | ( ~n800 & n3661 ) | ( n3660 & n3661 ) ;
  assign n3663 = ( n948 & n3660 ) | ( n948 & n3661 ) | ( n3660 & n3661 ) ;
  assign n3664 = ( n1061 & n3662 ) | ( n1061 & n3663 ) | ( n3662 & n3663 ) ;
  assign n3665 = n3657 | n3664 ;
  assign n3666 = ~n3650 & n3665 ;
  assign n3667 = x448 & n812 ;
  assign n3668 = x448 & ~n815 ;
  assign n3669 = ( n909 & n3667 ) | ( n909 & n3668 ) | ( n3667 & n3668 ) ;
  assign n3670 = ( ~n929 & n3667 ) | ( ~n929 & n3668 ) | ( n3667 & n3668 ) ;
  assign n3671 = ( n800 & n3669 ) | ( n800 & n3670 ) | ( n3669 & n3670 ) ;
  assign n3672 = ( ~n948 & n3669 ) | ( ~n948 & n3670 ) | ( n3669 & n3670 ) ;
  assign n3673 = ( ~n1061 & n3671 ) | ( ~n1061 & n3672 ) | ( n3671 & n3672 ) ;
  assign n3674 = x320 & ~n812 ;
  assign n3675 = x320 & n815 ;
  assign n3676 = ( ~n909 & n3674 ) | ( ~n909 & n3675 ) | ( n3674 & n3675 ) ;
  assign n3677 = ( n929 & n3674 ) | ( n929 & n3675 ) | ( n3674 & n3675 ) ;
  assign n3678 = ( ~n800 & n3676 ) | ( ~n800 & n3677 ) | ( n3676 & n3677 ) ;
  assign n3679 = ( n948 & n3676 ) | ( n948 & n3677 ) | ( n3676 & n3677 ) ;
  assign n3680 = ( n1061 & n3678 ) | ( n1061 & n3679 ) | ( n3678 & n3679 ) ;
  assign n3681 = n3673 | n3680 ;
  assign n3682 = x192 & n1370 ;
  assign n3683 = x192 & ~n1373 ;
  assign n3684 = ( n1467 & n3682 ) | ( n1467 & n3683 ) | ( n3682 & n3683 ) ;
  assign n3685 = ( ~n1487 & n3682 ) | ( ~n1487 & n3683 ) | ( n3682 & n3683 ) ;
  assign n3686 = ( n1358 & n3684 ) | ( n1358 & n3685 ) | ( n3684 & n3685 ) ;
  assign n3687 = ( ~n1506 & n3684 ) | ( ~n1506 & n3685 ) | ( n3684 & n3685 ) ;
  assign n3688 = ( ~n1612 & n3686 ) | ( ~n1612 & n3687 ) | ( n3686 & n3687 ) ;
  assign n3689 = x64 & ~n1370 ;
  assign n3690 = x64 & n1373 ;
  assign n3691 = ( ~n1467 & n3689 ) | ( ~n1467 & n3690 ) | ( n3689 & n3690 ) ;
  assign n3692 = ( n1487 & n3689 ) | ( n1487 & n3690 ) | ( n3689 & n3690 ) ;
  assign n3693 = ( ~n1358 & n3691 ) | ( ~n1358 & n3692 ) | ( n3691 & n3692 ) ;
  assign n3694 = ( n1506 & n3691 ) | ( n1506 & n3692 ) | ( n3691 & n3692 ) ;
  assign n3695 = ( n1612 & n3693 ) | ( n1612 & n3694 ) | ( n3693 & n3694 ) ;
  assign n3696 = n3688 | n3695 ;
  assign n3697 = n3681 & ~n3696 ;
  assign n3698 = n3666 | n3697 ;
  assign n3699 = n3635 | n3698 ;
  assign n3700 = n3572 | n3699 ;
  assign n3701 = ~n3681 & n3696 ;
  assign n3702 = ( n3650 & ~n3665 ) | ( n3650 & n3701 ) | ( ~n3665 & n3701 ) ;
  assign n3703 = ( ~n3618 & n3633 ) | ( ~n3618 & n3702 ) | ( n3633 & n3702 ) ;
  assign n3704 = ( n3587 & ~n3602 ) | ( n3587 & n3703 ) | ( ~n3602 & n3703 ) ;
  assign n3705 = ( n3572 & n3700 ) | ( n3572 & ~n3704 ) | ( n3700 & ~n3704 ) ;
  assign n3706 = ~n3506 & n3705 ;
  assign n3707 = x207 & n1370 ;
  assign n3708 = x207 & ~n1373 ;
  assign n3709 = ( n1467 & n3707 ) | ( n1467 & n3708 ) | ( n3707 & n3708 ) ;
  assign n3710 = ( ~n1487 & n3707 ) | ( ~n1487 & n3708 ) | ( n3707 & n3708 ) ;
  assign n3711 = ( n1358 & n3709 ) | ( n1358 & n3710 ) | ( n3709 & n3710 ) ;
  assign n3712 = ( ~n1506 & n3709 ) | ( ~n1506 & n3710 ) | ( n3709 & n3710 ) ;
  assign n3713 = ( ~n1612 & n3711 ) | ( ~n1612 & n3712 ) | ( n3711 & n3712 ) ;
  assign n3714 = x79 & ~n1370 ;
  assign n3715 = x79 & n1373 ;
  assign n3716 = ( ~n1467 & n3714 ) | ( ~n1467 & n3715 ) | ( n3714 & n3715 ) ;
  assign n3717 = ( n1487 & n3714 ) | ( n1487 & n3715 ) | ( n3714 & n3715 ) ;
  assign n3718 = ( ~n1358 & n3716 ) | ( ~n1358 & n3717 ) | ( n3716 & n3717 ) ;
  assign n3719 = ( n1506 & n3716 ) | ( n1506 & n3717 ) | ( n3716 & n3717 ) ;
  assign n3720 = ( n1612 & n3718 ) | ( n1612 & n3719 ) | ( n3718 & n3719 ) ;
  assign n3721 = n3713 | n3720 ;
  assign n3722 = x463 & n812 ;
  assign n3723 = x463 & ~n815 ;
  assign n3724 = ( n909 & n3722 ) | ( n909 & n3723 ) | ( n3722 & n3723 ) ;
  assign n3725 = ( ~n929 & n3722 ) | ( ~n929 & n3723 ) | ( n3722 & n3723 ) ;
  assign n3726 = ( n800 & n3724 ) | ( n800 & n3725 ) | ( n3724 & n3725 ) ;
  assign n3727 = ( ~n948 & n3724 ) | ( ~n948 & n3725 ) | ( n3724 & n3725 ) ;
  assign n3728 = ( ~n1061 & n3726 ) | ( ~n1061 & n3727 ) | ( n3726 & n3727 ) ;
  assign n3729 = x335 & ~n812 ;
  assign n3730 = x335 & n815 ;
  assign n3731 = ( ~n909 & n3729 ) | ( ~n909 & n3730 ) | ( n3729 & n3730 ) ;
  assign n3732 = ( n929 & n3729 ) | ( n929 & n3730 ) | ( n3729 & n3730 ) ;
  assign n3733 = ( ~n800 & n3731 ) | ( ~n800 & n3732 ) | ( n3731 & n3732 ) ;
  assign n3734 = ( n948 & n3731 ) | ( n948 & n3732 ) | ( n3731 & n3732 ) ;
  assign n3735 = ( n1061 & n3733 ) | ( n1061 & n3734 ) | ( n3733 & n3734 ) ;
  assign n3736 = n3728 | n3735 ;
  assign n3737 = ~n3721 & n3736 ;
  assign n3738 = x462 & n812 ;
  assign n3739 = x462 & ~n815 ;
  assign n3740 = ( n909 & n3738 ) | ( n909 & n3739 ) | ( n3738 & n3739 ) ;
  assign n3741 = ( ~n929 & n3738 ) | ( ~n929 & n3739 ) | ( n3738 & n3739 ) ;
  assign n3742 = ( n800 & n3740 ) | ( n800 & n3741 ) | ( n3740 & n3741 ) ;
  assign n3743 = ( ~n948 & n3740 ) | ( ~n948 & n3741 ) | ( n3740 & n3741 ) ;
  assign n3744 = ( ~n1061 & n3742 ) | ( ~n1061 & n3743 ) | ( n3742 & n3743 ) ;
  assign n3745 = x334 & ~n812 ;
  assign n3746 = x334 & n815 ;
  assign n3747 = ( ~n909 & n3745 ) | ( ~n909 & n3746 ) | ( n3745 & n3746 ) ;
  assign n3748 = ( n929 & n3745 ) | ( n929 & n3746 ) | ( n3745 & n3746 ) ;
  assign n3749 = ( ~n800 & n3747 ) | ( ~n800 & n3748 ) | ( n3747 & n3748 ) ;
  assign n3750 = ( n948 & n3747 ) | ( n948 & n3748 ) | ( n3747 & n3748 ) ;
  assign n3751 = ( n1061 & n3749 ) | ( n1061 & n3750 ) | ( n3749 & n3750 ) ;
  assign n3752 = n3744 | n3751 ;
  assign n3753 = x206 & n1370 ;
  assign n3754 = x206 & ~n1373 ;
  assign n3755 = ( n1467 & n3753 ) | ( n1467 & n3754 ) | ( n3753 & n3754 ) ;
  assign n3756 = ( ~n1487 & n3753 ) | ( ~n1487 & n3754 ) | ( n3753 & n3754 ) ;
  assign n3757 = ( n1358 & n3755 ) | ( n1358 & n3756 ) | ( n3755 & n3756 ) ;
  assign n3758 = ( ~n1506 & n3755 ) | ( ~n1506 & n3756 ) | ( n3755 & n3756 ) ;
  assign n3759 = ( ~n1612 & n3757 ) | ( ~n1612 & n3758 ) | ( n3757 & n3758 ) ;
  assign n3760 = x78 & ~n1370 ;
  assign n3761 = x78 & n1373 ;
  assign n3762 = ( ~n1467 & n3760 ) | ( ~n1467 & n3761 ) | ( n3760 & n3761 ) ;
  assign n3763 = ( n1487 & n3760 ) | ( n1487 & n3761 ) | ( n3760 & n3761 ) ;
  assign n3764 = ( ~n1358 & n3762 ) | ( ~n1358 & n3763 ) | ( n3762 & n3763 ) ;
  assign n3765 = ( n1506 & n3762 ) | ( n1506 & n3763 ) | ( n3762 & n3763 ) ;
  assign n3766 = ( n1612 & n3764 ) | ( n1612 & n3765 ) | ( n3764 & n3765 ) ;
  assign n3767 = n3759 | n3766 ;
  assign n3768 = n3752 & ~n3767 ;
  assign n3769 = n3737 | n3768 ;
  assign n3770 = x205 & n1370 ;
  assign n3771 = x205 & ~n1373 ;
  assign n3772 = ( n1467 & n3770 ) | ( n1467 & n3771 ) | ( n3770 & n3771 ) ;
  assign n3773 = ( ~n1487 & n3770 ) | ( ~n1487 & n3771 ) | ( n3770 & n3771 ) ;
  assign n3774 = ( n1358 & n3772 ) | ( n1358 & n3773 ) | ( n3772 & n3773 ) ;
  assign n3775 = ( ~n1506 & n3772 ) | ( ~n1506 & n3773 ) | ( n3772 & n3773 ) ;
  assign n3776 = ( ~n1612 & n3774 ) | ( ~n1612 & n3775 ) | ( n3774 & n3775 ) ;
  assign n3777 = x77 & ~n1370 ;
  assign n3778 = x77 & n1373 ;
  assign n3779 = ( ~n1467 & n3777 ) | ( ~n1467 & n3778 ) | ( n3777 & n3778 ) ;
  assign n3780 = ( n1487 & n3777 ) | ( n1487 & n3778 ) | ( n3777 & n3778 ) ;
  assign n3781 = ( ~n1358 & n3779 ) | ( ~n1358 & n3780 ) | ( n3779 & n3780 ) ;
  assign n3782 = ( n1506 & n3779 ) | ( n1506 & n3780 ) | ( n3779 & n3780 ) ;
  assign n3783 = ( n1612 & n3781 ) | ( n1612 & n3782 ) | ( n3781 & n3782 ) ;
  assign n3784 = n3776 | n3783 ;
  assign n3785 = x461 & n812 ;
  assign n3786 = x461 & ~n815 ;
  assign n3787 = ( n909 & n3785 ) | ( n909 & n3786 ) | ( n3785 & n3786 ) ;
  assign n3788 = ( ~n929 & n3785 ) | ( ~n929 & n3786 ) | ( n3785 & n3786 ) ;
  assign n3789 = ( n800 & n3787 ) | ( n800 & n3788 ) | ( n3787 & n3788 ) ;
  assign n3790 = ( ~n948 & n3787 ) | ( ~n948 & n3788 ) | ( n3787 & n3788 ) ;
  assign n3791 = ( ~n1061 & n3789 ) | ( ~n1061 & n3790 ) | ( n3789 & n3790 ) ;
  assign n3792 = x333 & ~n812 ;
  assign n3793 = x333 & n815 ;
  assign n3794 = ( ~n909 & n3792 ) | ( ~n909 & n3793 ) | ( n3792 & n3793 ) ;
  assign n3795 = ( n929 & n3792 ) | ( n929 & n3793 ) | ( n3792 & n3793 ) ;
  assign n3796 = ( ~n800 & n3794 ) | ( ~n800 & n3795 ) | ( n3794 & n3795 ) ;
  assign n3797 = ( n948 & n3794 ) | ( n948 & n3795 ) | ( n3794 & n3795 ) ;
  assign n3798 = ( n1061 & n3796 ) | ( n1061 & n3797 ) | ( n3796 & n3797 ) ;
  assign n3799 = n3791 | n3798 ;
  assign n3800 = ~n3784 & n3799 ;
  assign n3801 = x204 & n1370 ;
  assign n3802 = x204 & ~n1373 ;
  assign n3803 = ( n1467 & n3801 ) | ( n1467 & n3802 ) | ( n3801 & n3802 ) ;
  assign n3804 = ( ~n1487 & n3801 ) | ( ~n1487 & n3802 ) | ( n3801 & n3802 ) ;
  assign n3805 = ( n1358 & n3803 ) | ( n1358 & n3804 ) | ( n3803 & n3804 ) ;
  assign n3806 = ( ~n1506 & n3803 ) | ( ~n1506 & n3804 ) | ( n3803 & n3804 ) ;
  assign n3807 = ( ~n1612 & n3805 ) | ( ~n1612 & n3806 ) | ( n3805 & n3806 ) ;
  assign n3808 = x76 & ~n1370 ;
  assign n3809 = x76 & n1373 ;
  assign n3810 = ( ~n1467 & n3808 ) | ( ~n1467 & n3809 ) | ( n3808 & n3809 ) ;
  assign n3811 = ( n1487 & n3808 ) | ( n1487 & n3809 ) | ( n3808 & n3809 ) ;
  assign n3812 = ( ~n1358 & n3810 ) | ( ~n1358 & n3811 ) | ( n3810 & n3811 ) ;
  assign n3813 = ( n1506 & n3810 ) | ( n1506 & n3811 ) | ( n3810 & n3811 ) ;
  assign n3814 = ( n1612 & n3812 ) | ( n1612 & n3813 ) | ( n3812 & n3813 ) ;
  assign n3815 = n3807 | n3814 ;
  assign n3816 = x460 & n812 ;
  assign n3817 = x460 & ~n815 ;
  assign n3818 = ( n909 & n3816 ) | ( n909 & n3817 ) | ( n3816 & n3817 ) ;
  assign n3819 = ( ~n929 & n3816 ) | ( ~n929 & n3817 ) | ( n3816 & n3817 ) ;
  assign n3820 = ( n800 & n3818 ) | ( n800 & n3819 ) | ( n3818 & n3819 ) ;
  assign n3821 = ( ~n948 & n3818 ) | ( ~n948 & n3819 ) | ( n3818 & n3819 ) ;
  assign n3822 = ( ~n1061 & n3820 ) | ( ~n1061 & n3821 ) | ( n3820 & n3821 ) ;
  assign n3823 = x332 & ~n812 ;
  assign n3824 = x332 & n815 ;
  assign n3825 = ( ~n909 & n3823 ) | ( ~n909 & n3824 ) | ( n3823 & n3824 ) ;
  assign n3826 = ( n929 & n3823 ) | ( n929 & n3824 ) | ( n3823 & n3824 ) ;
  assign n3827 = ( ~n800 & n3825 ) | ( ~n800 & n3826 ) | ( n3825 & n3826 ) ;
  assign n3828 = ( n948 & n3825 ) | ( n948 & n3826 ) | ( n3825 & n3826 ) ;
  assign n3829 = ( n1061 & n3827 ) | ( n1061 & n3828 ) | ( n3827 & n3828 ) ;
  assign n3830 = n3822 | n3829 ;
  assign n3831 = ~n3815 & n3830 ;
  assign n3832 = n3800 | n3831 ;
  assign n3833 = n3769 | n3832 ;
  assign n3834 = x203 & n1370 ;
  assign n3835 = x203 & ~n1373 ;
  assign n3836 = ( n1467 & n3834 ) | ( n1467 & n3835 ) | ( n3834 & n3835 ) ;
  assign n3837 = ( ~n1487 & n3834 ) | ( ~n1487 & n3835 ) | ( n3834 & n3835 ) ;
  assign n3838 = ( n1358 & n3836 ) | ( n1358 & n3837 ) | ( n3836 & n3837 ) ;
  assign n3839 = ( ~n1506 & n3836 ) | ( ~n1506 & n3837 ) | ( n3836 & n3837 ) ;
  assign n3840 = ( ~n1612 & n3838 ) | ( ~n1612 & n3839 ) | ( n3838 & n3839 ) ;
  assign n3841 = x75 & ~n1370 ;
  assign n3842 = x75 & n1373 ;
  assign n3843 = ( ~n1467 & n3841 ) | ( ~n1467 & n3842 ) | ( n3841 & n3842 ) ;
  assign n3844 = ( n1487 & n3841 ) | ( n1487 & n3842 ) | ( n3841 & n3842 ) ;
  assign n3845 = ( ~n1358 & n3843 ) | ( ~n1358 & n3844 ) | ( n3843 & n3844 ) ;
  assign n3846 = ( n1506 & n3843 ) | ( n1506 & n3844 ) | ( n3843 & n3844 ) ;
  assign n3847 = ( n1612 & n3845 ) | ( n1612 & n3846 ) | ( n3845 & n3846 ) ;
  assign n3848 = n3840 | n3847 ;
  assign n3849 = x459 & n812 ;
  assign n3850 = x459 & ~n815 ;
  assign n3851 = ( n909 & n3849 ) | ( n909 & n3850 ) | ( n3849 & n3850 ) ;
  assign n3852 = ( ~n929 & n3849 ) | ( ~n929 & n3850 ) | ( n3849 & n3850 ) ;
  assign n3853 = ( n800 & n3851 ) | ( n800 & n3852 ) | ( n3851 & n3852 ) ;
  assign n3854 = ( ~n948 & n3851 ) | ( ~n948 & n3852 ) | ( n3851 & n3852 ) ;
  assign n3855 = ( ~n1061 & n3853 ) | ( ~n1061 & n3854 ) | ( n3853 & n3854 ) ;
  assign n3856 = x331 & ~n812 ;
  assign n3857 = x331 & n815 ;
  assign n3858 = ( ~n909 & n3856 ) | ( ~n909 & n3857 ) | ( n3856 & n3857 ) ;
  assign n3859 = ( n929 & n3856 ) | ( n929 & n3857 ) | ( n3856 & n3857 ) ;
  assign n3860 = ( ~n800 & n3858 ) | ( ~n800 & n3859 ) | ( n3858 & n3859 ) ;
  assign n3861 = ( n948 & n3858 ) | ( n948 & n3859 ) | ( n3858 & n3859 ) ;
  assign n3862 = ( n1061 & n3860 ) | ( n1061 & n3861 ) | ( n3860 & n3861 ) ;
  assign n3863 = n3855 | n3862 ;
  assign n3864 = ~n3848 & n3863 ;
  assign n3865 = x458 & n812 ;
  assign n3866 = x458 & ~n815 ;
  assign n3867 = ( n909 & n3865 ) | ( n909 & n3866 ) | ( n3865 & n3866 ) ;
  assign n3868 = ( ~n929 & n3865 ) | ( ~n929 & n3866 ) | ( n3865 & n3866 ) ;
  assign n3869 = ( n800 & n3867 ) | ( n800 & n3868 ) | ( n3867 & n3868 ) ;
  assign n3870 = ( ~n948 & n3867 ) | ( ~n948 & n3868 ) | ( n3867 & n3868 ) ;
  assign n3871 = ( ~n1061 & n3869 ) | ( ~n1061 & n3870 ) | ( n3869 & n3870 ) ;
  assign n3872 = x330 & ~n812 ;
  assign n3873 = x330 & n815 ;
  assign n3874 = ( ~n909 & n3872 ) | ( ~n909 & n3873 ) | ( n3872 & n3873 ) ;
  assign n3875 = ( n929 & n3872 ) | ( n929 & n3873 ) | ( n3872 & n3873 ) ;
  assign n3876 = ( ~n800 & n3874 ) | ( ~n800 & n3875 ) | ( n3874 & n3875 ) ;
  assign n3877 = ( n948 & n3874 ) | ( n948 & n3875 ) | ( n3874 & n3875 ) ;
  assign n3878 = ( n1061 & n3876 ) | ( n1061 & n3877 ) | ( n3876 & n3877 ) ;
  assign n3879 = n3871 | n3878 ;
  assign n3880 = x202 & n1370 ;
  assign n3881 = x202 & ~n1373 ;
  assign n3882 = ( n1467 & n3880 ) | ( n1467 & n3881 ) | ( n3880 & n3881 ) ;
  assign n3883 = ( ~n1487 & n3880 ) | ( ~n1487 & n3881 ) | ( n3880 & n3881 ) ;
  assign n3884 = ( n1358 & n3882 ) | ( n1358 & n3883 ) | ( n3882 & n3883 ) ;
  assign n3885 = ( ~n1506 & n3882 ) | ( ~n1506 & n3883 ) | ( n3882 & n3883 ) ;
  assign n3886 = ( ~n1612 & n3884 ) | ( ~n1612 & n3885 ) | ( n3884 & n3885 ) ;
  assign n3887 = x74 & ~n1370 ;
  assign n3888 = x74 & n1373 ;
  assign n3889 = ( ~n1467 & n3887 ) | ( ~n1467 & n3888 ) | ( n3887 & n3888 ) ;
  assign n3890 = ( n1487 & n3887 ) | ( n1487 & n3888 ) | ( n3887 & n3888 ) ;
  assign n3891 = ( ~n1358 & n3889 ) | ( ~n1358 & n3890 ) | ( n3889 & n3890 ) ;
  assign n3892 = ( n1506 & n3889 ) | ( n1506 & n3890 ) | ( n3889 & n3890 ) ;
  assign n3893 = ( n1612 & n3891 ) | ( n1612 & n3892 ) | ( n3891 & n3892 ) ;
  assign n3894 = n3886 | n3893 ;
  assign n3895 = n3879 & ~n3894 ;
  assign n3896 = n3864 | n3895 ;
  assign n3897 = x201 & n1370 ;
  assign n3898 = x201 & ~n1373 ;
  assign n3899 = ( n1467 & n3897 ) | ( n1467 & n3898 ) | ( n3897 & n3898 ) ;
  assign n3900 = ( ~n1487 & n3897 ) | ( ~n1487 & n3898 ) | ( n3897 & n3898 ) ;
  assign n3901 = ( n1358 & n3899 ) | ( n1358 & n3900 ) | ( n3899 & n3900 ) ;
  assign n3902 = ( ~n1506 & n3899 ) | ( ~n1506 & n3900 ) | ( n3899 & n3900 ) ;
  assign n3903 = ( ~n1612 & n3901 ) | ( ~n1612 & n3902 ) | ( n3901 & n3902 ) ;
  assign n3904 = x73 & ~n1370 ;
  assign n3905 = x73 & n1373 ;
  assign n3906 = ( ~n1467 & n3904 ) | ( ~n1467 & n3905 ) | ( n3904 & n3905 ) ;
  assign n3907 = ( n1487 & n3904 ) | ( n1487 & n3905 ) | ( n3904 & n3905 ) ;
  assign n3908 = ( ~n1358 & n3906 ) | ( ~n1358 & n3907 ) | ( n3906 & n3907 ) ;
  assign n3909 = ( n1506 & n3906 ) | ( n1506 & n3907 ) | ( n3906 & n3907 ) ;
  assign n3910 = ( n1612 & n3908 ) | ( n1612 & n3909 ) | ( n3908 & n3909 ) ;
  assign n3911 = n3903 | n3910 ;
  assign n3912 = x457 & n812 ;
  assign n3913 = x457 & ~n815 ;
  assign n3914 = ( n909 & n3912 ) | ( n909 & n3913 ) | ( n3912 & n3913 ) ;
  assign n3915 = ( ~n929 & n3912 ) | ( ~n929 & n3913 ) | ( n3912 & n3913 ) ;
  assign n3916 = ( n800 & n3914 ) | ( n800 & n3915 ) | ( n3914 & n3915 ) ;
  assign n3917 = ( ~n948 & n3914 ) | ( ~n948 & n3915 ) | ( n3914 & n3915 ) ;
  assign n3918 = ( ~n1061 & n3916 ) | ( ~n1061 & n3917 ) | ( n3916 & n3917 ) ;
  assign n3919 = x329 & ~n812 ;
  assign n3920 = x329 & n815 ;
  assign n3921 = ( ~n909 & n3919 ) | ( ~n909 & n3920 ) | ( n3919 & n3920 ) ;
  assign n3922 = ( n929 & n3919 ) | ( n929 & n3920 ) | ( n3919 & n3920 ) ;
  assign n3923 = ( ~n800 & n3921 ) | ( ~n800 & n3922 ) | ( n3921 & n3922 ) ;
  assign n3924 = ( n948 & n3921 ) | ( n948 & n3922 ) | ( n3921 & n3922 ) ;
  assign n3925 = ( n1061 & n3923 ) | ( n1061 & n3924 ) | ( n3923 & n3924 ) ;
  assign n3926 = n3918 | n3925 ;
  assign n3927 = ~n3911 & n3926 ;
  assign n3928 = x456 & n812 ;
  assign n3929 = x456 & ~n815 ;
  assign n3930 = ( n909 & n3928 ) | ( n909 & n3929 ) | ( n3928 & n3929 ) ;
  assign n3931 = ( ~n929 & n3928 ) | ( ~n929 & n3929 ) | ( n3928 & n3929 ) ;
  assign n3932 = ( n800 & n3930 ) | ( n800 & n3931 ) | ( n3930 & n3931 ) ;
  assign n3933 = ( ~n948 & n3930 ) | ( ~n948 & n3931 ) | ( n3930 & n3931 ) ;
  assign n3934 = ( ~n1061 & n3932 ) | ( ~n1061 & n3933 ) | ( n3932 & n3933 ) ;
  assign n3935 = x328 & ~n812 ;
  assign n3936 = x328 & n815 ;
  assign n3937 = ( ~n909 & n3935 ) | ( ~n909 & n3936 ) | ( n3935 & n3936 ) ;
  assign n3938 = ( n929 & n3935 ) | ( n929 & n3936 ) | ( n3935 & n3936 ) ;
  assign n3939 = ( ~n800 & n3937 ) | ( ~n800 & n3938 ) | ( n3937 & n3938 ) ;
  assign n3940 = ( n948 & n3937 ) | ( n948 & n3938 ) | ( n3937 & n3938 ) ;
  assign n3941 = ( n1061 & n3939 ) | ( n1061 & n3940 ) | ( n3939 & n3940 ) ;
  assign n3942 = n3934 | n3941 ;
  assign n3943 = x200 & n1370 ;
  assign n3944 = x200 & ~n1373 ;
  assign n3945 = ( n1467 & n3943 ) | ( n1467 & n3944 ) | ( n3943 & n3944 ) ;
  assign n3946 = ( ~n1487 & n3943 ) | ( ~n1487 & n3944 ) | ( n3943 & n3944 ) ;
  assign n3947 = ( n1358 & n3945 ) | ( n1358 & n3946 ) | ( n3945 & n3946 ) ;
  assign n3948 = ( ~n1506 & n3945 ) | ( ~n1506 & n3946 ) | ( n3945 & n3946 ) ;
  assign n3949 = ( ~n1612 & n3947 ) | ( ~n1612 & n3948 ) | ( n3947 & n3948 ) ;
  assign n3950 = x72 & ~n1370 ;
  assign n3951 = x72 & n1373 ;
  assign n3952 = ( ~n1467 & n3950 ) | ( ~n1467 & n3951 ) | ( n3950 & n3951 ) ;
  assign n3953 = ( n1487 & n3950 ) | ( n1487 & n3951 ) | ( n3950 & n3951 ) ;
  assign n3954 = ( ~n1358 & n3952 ) | ( ~n1358 & n3953 ) | ( n3952 & n3953 ) ;
  assign n3955 = ( n1506 & n3952 ) | ( n1506 & n3953 ) | ( n3952 & n3953 ) ;
  assign n3956 = ( n1612 & n3954 ) | ( n1612 & n3955 ) | ( n3954 & n3955 ) ;
  assign n3957 = n3949 | n3956 ;
  assign n3958 = n3942 & ~n3957 ;
  assign n3959 = n3927 | n3958 ;
  assign n3960 = n3896 | n3959 ;
  assign n3961 = n3554 & ~n3569 ;
  assign n3962 = ( n3523 & ~n3538 ) | ( n3523 & n3961 ) | ( ~n3538 & n3961 ) ;
  assign n3963 = ~n3507 & n3962 ;
  assign n3964 = ( n3458 & ~n3473 ) | ( n3458 & n3963 ) | ( ~n3473 & n3963 ) ;
  assign n3965 = ~n3960 & n3964 ;
  assign n3966 = ~n3942 & n3957 ;
  assign n3967 = ( n3911 & ~n3926 ) | ( n3911 & n3966 ) | ( ~n3926 & n3966 ) ;
  assign n3968 = ( ~n3879 & n3894 ) | ( ~n3879 & n3967 ) | ( n3894 & n3967 ) ;
  assign n3969 = ( n3848 & ~n3863 ) | ( n3848 & n3968 ) | ( ~n3863 & n3968 ) ;
  assign n3970 = ~n3833 & n3969 ;
  assign n3971 = ( ~n3833 & n3965 ) | ( ~n3833 & n3970 ) | ( n3965 & n3970 ) ;
  assign n3972 = n3833 | n3960 ;
  assign n3973 = ( n3833 & ~n3969 ) | ( n3833 & n3972 ) | ( ~n3969 & n3972 ) ;
  assign n3974 = ( n3706 & ~n3971 ) | ( n3706 & n3973 ) | ( ~n3971 & n3973 ) ;
  assign n3975 = ~n3572 & n3704 ;
  assign n3976 = n3506 | n3975 ;
  assign n3977 = ( n3971 & ~n3973 ) | ( n3971 & n3976 ) | ( ~n3973 & n3976 ) ;
  assign n3978 = x191 & n1370 ;
  assign n3979 = x191 & ~n1373 ;
  assign n3980 = ( n1467 & n3978 ) | ( n1467 & n3979 ) | ( n3978 & n3979 ) ;
  assign n3981 = ( ~n1487 & n3978 ) | ( ~n1487 & n3979 ) | ( n3978 & n3979 ) ;
  assign n3982 = ( n1358 & n3980 ) | ( n1358 & n3981 ) | ( n3980 & n3981 ) ;
  assign n3983 = ( ~n1506 & n3980 ) | ( ~n1506 & n3981 ) | ( n3980 & n3981 ) ;
  assign n3984 = ( ~n1612 & n3982 ) | ( ~n1612 & n3983 ) | ( n3982 & n3983 ) ;
  assign n3985 = x63 & ~n1370 ;
  assign n3986 = x63 & n1373 ;
  assign n3987 = ( ~n1467 & n3985 ) | ( ~n1467 & n3986 ) | ( n3985 & n3986 ) ;
  assign n3988 = ( n1487 & n3985 ) | ( n1487 & n3986 ) | ( n3985 & n3986 ) ;
  assign n3989 = ( ~n1358 & n3987 ) | ( ~n1358 & n3988 ) | ( n3987 & n3988 ) ;
  assign n3990 = ( n1506 & n3987 ) | ( n1506 & n3988 ) | ( n3987 & n3988 ) ;
  assign n3991 = ( n1612 & n3989 ) | ( n1612 & n3990 ) | ( n3989 & n3990 ) ;
  assign n3992 = n3984 | n3991 ;
  assign n3993 = x447 & n812 ;
  assign n3994 = x447 & ~n815 ;
  assign n3995 = ( n909 & n3993 ) | ( n909 & n3994 ) | ( n3993 & n3994 ) ;
  assign n3996 = ( ~n929 & n3993 ) | ( ~n929 & n3994 ) | ( n3993 & n3994 ) ;
  assign n3997 = ( n800 & n3995 ) | ( n800 & n3996 ) | ( n3995 & n3996 ) ;
  assign n3998 = ( ~n948 & n3995 ) | ( ~n948 & n3996 ) | ( n3995 & n3996 ) ;
  assign n3999 = ( ~n1061 & n3997 ) | ( ~n1061 & n3998 ) | ( n3997 & n3998 ) ;
  assign n4000 = x319 & ~n812 ;
  assign n4001 = x319 & n815 ;
  assign n4002 = ( ~n909 & n4000 ) | ( ~n909 & n4001 ) | ( n4000 & n4001 ) ;
  assign n4003 = ( n929 & n4000 ) | ( n929 & n4001 ) | ( n4000 & n4001 ) ;
  assign n4004 = ( ~n800 & n4002 ) | ( ~n800 & n4003 ) | ( n4002 & n4003 ) ;
  assign n4005 = ( n948 & n4002 ) | ( n948 & n4003 ) | ( n4002 & n4003 ) ;
  assign n4006 = ( n1061 & n4004 ) | ( n1061 & n4005 ) | ( n4004 & n4005 ) ;
  assign n4007 = n3999 | n4006 ;
  assign n4008 = ~n3992 & n4007 ;
  assign n4009 = x446 & n812 ;
  assign n4010 = x446 & ~n815 ;
  assign n4011 = ( n909 & n4009 ) | ( n909 & n4010 ) | ( n4009 & n4010 ) ;
  assign n4012 = ( ~n929 & n4009 ) | ( ~n929 & n4010 ) | ( n4009 & n4010 ) ;
  assign n4013 = ( n800 & n4011 ) | ( n800 & n4012 ) | ( n4011 & n4012 ) ;
  assign n4014 = ( ~n948 & n4011 ) | ( ~n948 & n4012 ) | ( n4011 & n4012 ) ;
  assign n4015 = ( ~n1061 & n4013 ) | ( ~n1061 & n4014 ) | ( n4013 & n4014 ) ;
  assign n4016 = x318 & ~n812 ;
  assign n4017 = x318 & n815 ;
  assign n4018 = ( ~n909 & n4016 ) | ( ~n909 & n4017 ) | ( n4016 & n4017 ) ;
  assign n4019 = ( n929 & n4016 ) | ( n929 & n4017 ) | ( n4016 & n4017 ) ;
  assign n4020 = ( ~n800 & n4018 ) | ( ~n800 & n4019 ) | ( n4018 & n4019 ) ;
  assign n4021 = ( n948 & n4018 ) | ( n948 & n4019 ) | ( n4018 & n4019 ) ;
  assign n4022 = ( n1061 & n4020 ) | ( n1061 & n4021 ) | ( n4020 & n4021 ) ;
  assign n4023 = n4015 | n4022 ;
  assign n4024 = x190 & n1370 ;
  assign n4025 = x190 & ~n1373 ;
  assign n4026 = ( n1467 & n4024 ) | ( n1467 & n4025 ) | ( n4024 & n4025 ) ;
  assign n4027 = ( ~n1487 & n4024 ) | ( ~n1487 & n4025 ) | ( n4024 & n4025 ) ;
  assign n4028 = ( n1358 & n4026 ) | ( n1358 & n4027 ) | ( n4026 & n4027 ) ;
  assign n4029 = ( ~n1506 & n4026 ) | ( ~n1506 & n4027 ) | ( n4026 & n4027 ) ;
  assign n4030 = ( ~n1612 & n4028 ) | ( ~n1612 & n4029 ) | ( n4028 & n4029 ) ;
  assign n4031 = x62 & ~n1370 ;
  assign n4032 = x62 & n1373 ;
  assign n4033 = ( ~n1467 & n4031 ) | ( ~n1467 & n4032 ) | ( n4031 & n4032 ) ;
  assign n4034 = ( n1487 & n4031 ) | ( n1487 & n4032 ) | ( n4031 & n4032 ) ;
  assign n4035 = ( ~n1358 & n4033 ) | ( ~n1358 & n4034 ) | ( n4033 & n4034 ) ;
  assign n4036 = ( n1506 & n4033 ) | ( n1506 & n4034 ) | ( n4033 & n4034 ) ;
  assign n4037 = ( n1612 & n4035 ) | ( n1612 & n4036 ) | ( n4035 & n4036 ) ;
  assign n4038 = n4030 | n4037 ;
  assign n4039 = n4023 & ~n4038 ;
  assign n4040 = n4008 | n4039 ;
  assign n4041 = x189 & n1370 ;
  assign n4042 = x189 & ~n1373 ;
  assign n4043 = ( n1467 & n4041 ) | ( n1467 & n4042 ) | ( n4041 & n4042 ) ;
  assign n4044 = ( ~n1487 & n4041 ) | ( ~n1487 & n4042 ) | ( n4041 & n4042 ) ;
  assign n4045 = ( n1358 & n4043 ) | ( n1358 & n4044 ) | ( n4043 & n4044 ) ;
  assign n4046 = ( ~n1506 & n4043 ) | ( ~n1506 & n4044 ) | ( n4043 & n4044 ) ;
  assign n4047 = ( ~n1612 & n4045 ) | ( ~n1612 & n4046 ) | ( n4045 & n4046 ) ;
  assign n4048 = x61 & ~n1370 ;
  assign n4049 = x61 & n1373 ;
  assign n4050 = ( ~n1467 & n4048 ) | ( ~n1467 & n4049 ) | ( n4048 & n4049 ) ;
  assign n4051 = ( n1487 & n4048 ) | ( n1487 & n4049 ) | ( n4048 & n4049 ) ;
  assign n4052 = ( ~n1358 & n4050 ) | ( ~n1358 & n4051 ) | ( n4050 & n4051 ) ;
  assign n4053 = ( n1506 & n4050 ) | ( n1506 & n4051 ) | ( n4050 & n4051 ) ;
  assign n4054 = ( n1612 & n4052 ) | ( n1612 & n4053 ) | ( n4052 & n4053 ) ;
  assign n4055 = n4047 | n4054 ;
  assign n4056 = x445 & n812 ;
  assign n4057 = x445 & ~n815 ;
  assign n4058 = ( n909 & n4056 ) | ( n909 & n4057 ) | ( n4056 & n4057 ) ;
  assign n4059 = ( ~n929 & n4056 ) | ( ~n929 & n4057 ) | ( n4056 & n4057 ) ;
  assign n4060 = ( n800 & n4058 ) | ( n800 & n4059 ) | ( n4058 & n4059 ) ;
  assign n4061 = ( ~n948 & n4058 ) | ( ~n948 & n4059 ) | ( n4058 & n4059 ) ;
  assign n4062 = ( ~n1061 & n4060 ) | ( ~n1061 & n4061 ) | ( n4060 & n4061 ) ;
  assign n4063 = x317 & ~n812 ;
  assign n4064 = x317 & n815 ;
  assign n4065 = ( ~n909 & n4063 ) | ( ~n909 & n4064 ) | ( n4063 & n4064 ) ;
  assign n4066 = ( n929 & n4063 ) | ( n929 & n4064 ) | ( n4063 & n4064 ) ;
  assign n4067 = ( ~n800 & n4065 ) | ( ~n800 & n4066 ) | ( n4065 & n4066 ) ;
  assign n4068 = ( n948 & n4065 ) | ( n948 & n4066 ) | ( n4065 & n4066 ) ;
  assign n4069 = ( n1061 & n4067 ) | ( n1061 & n4068 ) | ( n4067 & n4068 ) ;
  assign n4070 = n4062 | n4069 ;
  assign n4071 = ~n4055 & n4070 ;
  assign n4072 = x188 & n1370 ;
  assign n4073 = x188 & ~n1373 ;
  assign n4074 = ( n1467 & n4072 ) | ( n1467 & n4073 ) | ( n4072 & n4073 ) ;
  assign n4075 = ( ~n1487 & n4072 ) | ( ~n1487 & n4073 ) | ( n4072 & n4073 ) ;
  assign n4076 = ( n1358 & n4074 ) | ( n1358 & n4075 ) | ( n4074 & n4075 ) ;
  assign n4077 = ( ~n1506 & n4074 ) | ( ~n1506 & n4075 ) | ( n4074 & n4075 ) ;
  assign n4078 = ( ~n1612 & n4076 ) | ( ~n1612 & n4077 ) | ( n4076 & n4077 ) ;
  assign n4079 = x60 & ~n1370 ;
  assign n4080 = x60 & n1373 ;
  assign n4081 = ( ~n1467 & n4079 ) | ( ~n1467 & n4080 ) | ( n4079 & n4080 ) ;
  assign n4082 = ( n1487 & n4079 ) | ( n1487 & n4080 ) | ( n4079 & n4080 ) ;
  assign n4083 = ( ~n1358 & n4081 ) | ( ~n1358 & n4082 ) | ( n4081 & n4082 ) ;
  assign n4084 = ( n1506 & n4081 ) | ( n1506 & n4082 ) | ( n4081 & n4082 ) ;
  assign n4085 = ( n1612 & n4083 ) | ( n1612 & n4084 ) | ( n4083 & n4084 ) ;
  assign n4086 = n4078 | n4085 ;
  assign n4087 = x444 & n812 ;
  assign n4088 = x444 & ~n815 ;
  assign n4089 = ( n909 & n4087 ) | ( n909 & n4088 ) | ( n4087 & n4088 ) ;
  assign n4090 = ( ~n929 & n4087 ) | ( ~n929 & n4088 ) | ( n4087 & n4088 ) ;
  assign n4091 = ( n800 & n4089 ) | ( n800 & n4090 ) | ( n4089 & n4090 ) ;
  assign n4092 = ( ~n948 & n4089 ) | ( ~n948 & n4090 ) | ( n4089 & n4090 ) ;
  assign n4093 = ( ~n1061 & n4091 ) | ( ~n1061 & n4092 ) | ( n4091 & n4092 ) ;
  assign n4094 = x316 & ~n812 ;
  assign n4095 = x316 & n815 ;
  assign n4096 = ( ~n909 & n4094 ) | ( ~n909 & n4095 ) | ( n4094 & n4095 ) ;
  assign n4097 = ( n929 & n4094 ) | ( n929 & n4095 ) | ( n4094 & n4095 ) ;
  assign n4098 = ( ~n800 & n4096 ) | ( ~n800 & n4097 ) | ( n4096 & n4097 ) ;
  assign n4099 = ( n948 & n4096 ) | ( n948 & n4097 ) | ( n4096 & n4097 ) ;
  assign n4100 = ( n1061 & n4098 ) | ( n1061 & n4099 ) | ( n4098 & n4099 ) ;
  assign n4101 = n4093 | n4100 ;
  assign n4102 = ~n4086 & n4101 ;
  assign n4103 = n4071 | n4102 ;
  assign n4104 = n4040 | n4103 ;
  assign n4105 = x187 & n1370 ;
  assign n4106 = x187 & ~n1373 ;
  assign n4107 = ( n1467 & n4105 ) | ( n1467 & n4106 ) | ( n4105 & n4106 ) ;
  assign n4108 = ( ~n1487 & n4105 ) | ( ~n1487 & n4106 ) | ( n4105 & n4106 ) ;
  assign n4109 = ( n1358 & n4107 ) | ( n1358 & n4108 ) | ( n4107 & n4108 ) ;
  assign n4110 = ( ~n1506 & n4107 ) | ( ~n1506 & n4108 ) | ( n4107 & n4108 ) ;
  assign n4111 = ( ~n1612 & n4109 ) | ( ~n1612 & n4110 ) | ( n4109 & n4110 ) ;
  assign n4112 = x59 & ~n1370 ;
  assign n4113 = x59 & n1373 ;
  assign n4114 = ( ~n1467 & n4112 ) | ( ~n1467 & n4113 ) | ( n4112 & n4113 ) ;
  assign n4115 = ( n1487 & n4112 ) | ( n1487 & n4113 ) | ( n4112 & n4113 ) ;
  assign n4116 = ( ~n1358 & n4114 ) | ( ~n1358 & n4115 ) | ( n4114 & n4115 ) ;
  assign n4117 = ( n1506 & n4114 ) | ( n1506 & n4115 ) | ( n4114 & n4115 ) ;
  assign n4118 = ( n1612 & n4116 ) | ( n1612 & n4117 ) | ( n4116 & n4117 ) ;
  assign n4119 = n4111 | n4118 ;
  assign n4120 = x443 & n812 ;
  assign n4121 = x443 & ~n815 ;
  assign n4122 = ( n909 & n4120 ) | ( n909 & n4121 ) | ( n4120 & n4121 ) ;
  assign n4123 = ( ~n929 & n4120 ) | ( ~n929 & n4121 ) | ( n4120 & n4121 ) ;
  assign n4124 = ( n800 & n4122 ) | ( n800 & n4123 ) | ( n4122 & n4123 ) ;
  assign n4125 = ( ~n948 & n4122 ) | ( ~n948 & n4123 ) | ( n4122 & n4123 ) ;
  assign n4126 = ( ~n1061 & n4124 ) | ( ~n1061 & n4125 ) | ( n4124 & n4125 ) ;
  assign n4127 = x315 & ~n812 ;
  assign n4128 = x315 & n815 ;
  assign n4129 = ( ~n909 & n4127 ) | ( ~n909 & n4128 ) | ( n4127 & n4128 ) ;
  assign n4130 = ( n929 & n4127 ) | ( n929 & n4128 ) | ( n4127 & n4128 ) ;
  assign n4131 = ( ~n800 & n4129 ) | ( ~n800 & n4130 ) | ( n4129 & n4130 ) ;
  assign n4132 = ( n948 & n4129 ) | ( n948 & n4130 ) | ( n4129 & n4130 ) ;
  assign n4133 = ( n1061 & n4131 ) | ( n1061 & n4132 ) | ( n4131 & n4132 ) ;
  assign n4134 = n4126 | n4133 ;
  assign n4135 = x186 & n1370 ;
  assign n4136 = x186 & ~n1373 ;
  assign n4137 = ( n1467 & n4135 ) | ( n1467 & n4136 ) | ( n4135 & n4136 ) ;
  assign n4138 = ( ~n1487 & n4135 ) | ( ~n1487 & n4136 ) | ( n4135 & n4136 ) ;
  assign n4139 = ( n1358 & n4137 ) | ( n1358 & n4138 ) | ( n4137 & n4138 ) ;
  assign n4140 = ( ~n1506 & n4137 ) | ( ~n1506 & n4138 ) | ( n4137 & n4138 ) ;
  assign n4141 = ( ~n1612 & n4139 ) | ( ~n1612 & n4140 ) | ( n4139 & n4140 ) ;
  assign n4142 = x58 & ~n1370 ;
  assign n4143 = x58 & n1373 ;
  assign n4144 = ( ~n1467 & n4142 ) | ( ~n1467 & n4143 ) | ( n4142 & n4143 ) ;
  assign n4145 = ( n1487 & n4142 ) | ( n1487 & n4143 ) | ( n4142 & n4143 ) ;
  assign n4146 = ( ~n1358 & n4144 ) | ( ~n1358 & n4145 ) | ( n4144 & n4145 ) ;
  assign n4147 = ( n1506 & n4144 ) | ( n1506 & n4145 ) | ( n4144 & n4145 ) ;
  assign n4148 = ( n1612 & n4146 ) | ( n1612 & n4147 ) | ( n4146 & n4147 ) ;
  assign n4149 = n4141 | n4148 ;
  assign n4150 = x442 & n812 ;
  assign n4151 = x442 & ~n815 ;
  assign n4152 = ( n909 & n4150 ) | ( n909 & n4151 ) | ( n4150 & n4151 ) ;
  assign n4153 = ( ~n929 & n4150 ) | ( ~n929 & n4151 ) | ( n4150 & n4151 ) ;
  assign n4154 = ( n800 & n4152 ) | ( n800 & n4153 ) | ( n4152 & n4153 ) ;
  assign n4155 = ( ~n948 & n4152 ) | ( ~n948 & n4153 ) | ( n4152 & n4153 ) ;
  assign n4156 = ( ~n1061 & n4154 ) | ( ~n1061 & n4155 ) | ( n4154 & n4155 ) ;
  assign n4157 = x314 & ~n812 ;
  assign n4158 = x314 & n815 ;
  assign n4159 = ( ~n909 & n4157 ) | ( ~n909 & n4158 ) | ( n4157 & n4158 ) ;
  assign n4160 = ( n929 & n4157 ) | ( n929 & n4158 ) | ( n4157 & n4158 ) ;
  assign n4161 = ( ~n800 & n4159 ) | ( ~n800 & n4160 ) | ( n4159 & n4160 ) ;
  assign n4162 = ( n948 & n4159 ) | ( n948 & n4160 ) | ( n4159 & n4160 ) ;
  assign n4163 = ( n1061 & n4161 ) | ( n1061 & n4162 ) | ( n4161 & n4162 ) ;
  assign n4164 = n4156 | n4163 ;
  assign n4165 = x185 & n1370 ;
  assign n4166 = x185 & ~n1373 ;
  assign n4167 = ( n1467 & n4165 ) | ( n1467 & n4166 ) | ( n4165 & n4166 ) ;
  assign n4168 = ( ~n1487 & n4165 ) | ( ~n1487 & n4166 ) | ( n4165 & n4166 ) ;
  assign n4169 = ( n1358 & n4167 ) | ( n1358 & n4168 ) | ( n4167 & n4168 ) ;
  assign n4170 = ( ~n1506 & n4167 ) | ( ~n1506 & n4168 ) | ( n4167 & n4168 ) ;
  assign n4171 = ( ~n1612 & n4169 ) | ( ~n1612 & n4170 ) | ( n4169 & n4170 ) ;
  assign n4172 = x57 & ~n1370 ;
  assign n4173 = x57 & n1373 ;
  assign n4174 = ( ~n1467 & n4172 ) | ( ~n1467 & n4173 ) | ( n4172 & n4173 ) ;
  assign n4175 = ( n1487 & n4172 ) | ( n1487 & n4173 ) | ( n4172 & n4173 ) ;
  assign n4176 = ( ~n1358 & n4174 ) | ( ~n1358 & n4175 ) | ( n4174 & n4175 ) ;
  assign n4177 = ( n1506 & n4174 ) | ( n1506 & n4175 ) | ( n4174 & n4175 ) ;
  assign n4178 = ( n1612 & n4176 ) | ( n1612 & n4177 ) | ( n4176 & n4177 ) ;
  assign n4179 = n4171 | n4178 ;
  assign n4180 = x441 & n812 ;
  assign n4181 = x441 & ~n815 ;
  assign n4182 = ( n909 & n4180 ) | ( n909 & n4181 ) | ( n4180 & n4181 ) ;
  assign n4183 = ( ~n929 & n4180 ) | ( ~n929 & n4181 ) | ( n4180 & n4181 ) ;
  assign n4184 = ( n800 & n4182 ) | ( n800 & n4183 ) | ( n4182 & n4183 ) ;
  assign n4185 = ( ~n948 & n4182 ) | ( ~n948 & n4183 ) | ( n4182 & n4183 ) ;
  assign n4186 = ( ~n1061 & n4184 ) | ( ~n1061 & n4185 ) | ( n4184 & n4185 ) ;
  assign n4187 = x313 & ~n812 ;
  assign n4188 = x313 & n815 ;
  assign n4189 = ( ~n909 & n4187 ) | ( ~n909 & n4188 ) | ( n4187 & n4188 ) ;
  assign n4190 = ( n929 & n4187 ) | ( n929 & n4188 ) | ( n4187 & n4188 ) ;
  assign n4191 = ( ~n800 & n4189 ) | ( ~n800 & n4190 ) | ( n4189 & n4190 ) ;
  assign n4192 = ( n948 & n4189 ) | ( n948 & n4190 ) | ( n4189 & n4190 ) ;
  assign n4193 = ( n1061 & n4191 ) | ( n1061 & n4192 ) | ( n4191 & n4192 ) ;
  assign n4194 = n4186 | n4193 ;
  assign n4195 = x184 & n1370 ;
  assign n4196 = x184 & ~n1373 ;
  assign n4197 = ( n1467 & n4195 ) | ( n1467 & n4196 ) | ( n4195 & n4196 ) ;
  assign n4198 = ( ~n1487 & n4195 ) | ( ~n1487 & n4196 ) | ( n4195 & n4196 ) ;
  assign n4199 = ( n1358 & n4197 ) | ( n1358 & n4198 ) | ( n4197 & n4198 ) ;
  assign n4200 = ( ~n1506 & n4197 ) | ( ~n1506 & n4198 ) | ( n4197 & n4198 ) ;
  assign n4201 = ( ~n1612 & n4199 ) | ( ~n1612 & n4200 ) | ( n4199 & n4200 ) ;
  assign n4202 = x56 & ~n1370 ;
  assign n4203 = x56 & n1373 ;
  assign n4204 = ( ~n1467 & n4202 ) | ( ~n1467 & n4203 ) | ( n4202 & n4203 ) ;
  assign n4205 = ( n1487 & n4202 ) | ( n1487 & n4203 ) | ( n4202 & n4203 ) ;
  assign n4206 = ( ~n1358 & n4204 ) | ( ~n1358 & n4205 ) | ( n4204 & n4205 ) ;
  assign n4207 = ( n1506 & n4204 ) | ( n1506 & n4205 ) | ( n4204 & n4205 ) ;
  assign n4208 = ( n1612 & n4206 ) | ( n1612 & n4207 ) | ( n4206 & n4207 ) ;
  assign n4209 = n4201 | n4208 ;
  assign n4210 = x440 & n812 ;
  assign n4211 = x440 & ~n815 ;
  assign n4212 = ( n909 & n4210 ) | ( n909 & n4211 ) | ( n4210 & n4211 ) ;
  assign n4213 = ( ~n929 & n4210 ) | ( ~n929 & n4211 ) | ( n4210 & n4211 ) ;
  assign n4214 = ( n800 & n4212 ) | ( n800 & n4213 ) | ( n4212 & n4213 ) ;
  assign n4215 = ( ~n948 & n4212 ) | ( ~n948 & n4213 ) | ( n4212 & n4213 ) ;
  assign n4216 = ( ~n1061 & n4214 ) | ( ~n1061 & n4215 ) | ( n4214 & n4215 ) ;
  assign n4217 = x312 & ~n812 ;
  assign n4218 = x312 & n815 ;
  assign n4219 = ( ~n909 & n4217 ) | ( ~n909 & n4218 ) | ( n4217 & n4218 ) ;
  assign n4220 = ( n929 & n4217 ) | ( n929 & n4218 ) | ( n4217 & n4218 ) ;
  assign n4221 = ( ~n800 & n4219 ) | ( ~n800 & n4220 ) | ( n4219 & n4220 ) ;
  assign n4222 = ( n948 & n4219 ) | ( n948 & n4220 ) | ( n4219 & n4220 ) ;
  assign n4223 = ( n1061 & n4221 ) | ( n1061 & n4222 ) | ( n4221 & n4222 ) ;
  assign n4224 = n4216 | n4223 ;
  assign n4225 = n4209 & ~n4224 ;
  assign n4226 = ( n4179 & ~n4194 ) | ( n4179 & n4225 ) | ( ~n4194 & n4225 ) ;
  assign n4227 = ( n4149 & ~n4164 ) | ( n4149 & n4226 ) | ( ~n4164 & n4226 ) ;
  assign n4228 = ( n4119 & ~n4134 ) | ( n4119 & n4227 ) | ( ~n4134 & n4227 ) ;
  assign n4229 = ~n4104 & n4228 ;
  assign n4230 = n4086 & ~n4101 ;
  assign n4231 = ( n4055 & ~n4070 ) | ( n4055 & n4230 ) | ( ~n4070 & n4230 ) ;
  assign n4232 = ~n4040 & n4231 ;
  assign n4233 = ~n4023 & n4038 ;
  assign n4234 = ( n3992 & ~n4007 ) | ( n3992 & n4233 ) | ( ~n4007 & n4233 ) ;
  assign n4235 = n4232 | n4234 ;
  assign n4236 = n4229 | n4235 ;
  assign n4237 = ~n4119 & n4134 ;
  assign n4238 = ~n4149 & n4164 ;
  assign n4239 = n4237 | n4238 ;
  assign n4240 = ~n4179 & n4194 ;
  assign n4241 = ~n4209 & n4224 ;
  assign n4242 = n4240 | n4241 ;
  assign n4243 = n4239 | n4242 ;
  assign n4244 = ( n4232 & n4233 ) | ( n4232 & n4235 ) | ( n4233 & n4235 ) ;
  assign n4245 = ( n4104 & n4243 ) | ( n4104 & ~n4244 ) | ( n4243 & ~n4244 ) ;
  assign n4246 = ~n4236 & n4245 ;
  assign n4247 = ( n3974 & ~n3977 ) | ( n3974 & n4246 ) | ( ~n3977 & n4246 ) ;
  assign n4248 = ~n3752 & n3767 ;
  assign n4249 = ~n3737 & n4248 ;
  assign n4250 = n3721 & ~n3736 ;
  assign n4251 = ~n3443 & n4250 ;
  assign n4252 = n3815 & ~n3830 ;
  assign n4253 = ( n3784 & ~n3799 ) | ( n3784 & n4252 ) | ( ~n3799 & n4252 ) ;
  assign n4254 = ~n3769 & n4253 ;
  assign n4255 = ( ~n3443 & n4251 ) | ( ~n3443 & n4254 ) | ( n4251 & n4254 ) ;
  assign n4256 = ( ~n3443 & n4249 ) | ( ~n3443 & n4255 ) | ( n4249 & n4255 ) ;
  assign n4257 = ( n3443 & n4247 ) | ( n3443 & ~n4256 ) | ( n4247 & ~n4256 ) ;
  assign n4258 = ( n3506 & ~n3508 ) | ( n3506 & n3962 ) | ( ~n3508 & n3962 ) ;
  assign n4259 = ( ~n3960 & n3965 ) | ( ~n3960 & n4258 ) | ( n3965 & n4258 ) ;
  assign n4260 = ( n3705 & n3960 ) | ( n3705 & ~n4259 ) | ( n3960 & ~n4259 ) ;
  assign n4261 = ( ~n3960 & n3975 ) | ( ~n3960 & n4259 ) | ( n3975 & n4259 ) ;
  assign n4262 = ( n4236 & ~n4260 ) | ( n4236 & n4261 ) | ( ~n4260 & n4261 ) ;
  assign n4263 = ( ~n3443 & n3970 ) | ( ~n3443 & n4256 ) | ( n3970 & n4256 ) ;
  assign n4264 = ( n3443 & n3833 ) | ( n3443 & ~n4256 ) | ( n3833 & ~n4256 ) ;
  assign n4265 = ( n4262 & n4263 ) | ( n4262 & ~n4264 ) | ( n4263 & ~n4264 ) ;
  assign n4266 = ( n3412 & ~n4257 ) | ( n3412 & n4265 ) | ( ~n4257 & n4265 ) ;
  assign n4267 = n1781 & ~n1796 ;
  assign n4268 = ~n1751 & n1766 ;
  assign n4269 = n4267 | n4268 ;
  assign n4270 = ~n1811 & n1826 ;
  assign n4271 = n1841 & ~n1856 ;
  assign n4272 = n4270 | n4271 ;
  assign n4273 = n4269 | n4272 ;
  assign n4274 = x231 & n1370 ;
  assign n4275 = x231 & ~n1373 ;
  assign n4276 = ( n1467 & n4274 ) | ( n1467 & n4275 ) | ( n4274 & n4275 ) ;
  assign n4277 = ( ~n1487 & n4274 ) | ( ~n1487 & n4275 ) | ( n4274 & n4275 ) ;
  assign n4278 = ( n1358 & n4276 ) | ( n1358 & n4277 ) | ( n4276 & n4277 ) ;
  assign n4279 = ( ~n1506 & n4276 ) | ( ~n1506 & n4277 ) | ( n4276 & n4277 ) ;
  assign n4280 = ( ~n1612 & n4278 ) | ( ~n1612 & n4279 ) | ( n4278 & n4279 ) ;
  assign n4281 = x103 & ~n1370 ;
  assign n4282 = x103 & n1373 ;
  assign n4283 = ( ~n1467 & n4281 ) | ( ~n1467 & n4282 ) | ( n4281 & n4282 ) ;
  assign n4284 = ( n1487 & n4281 ) | ( n1487 & n4282 ) | ( n4281 & n4282 ) ;
  assign n4285 = ( ~n1358 & n4283 ) | ( ~n1358 & n4284 ) | ( n4283 & n4284 ) ;
  assign n4286 = ( n1506 & n4283 ) | ( n1506 & n4284 ) | ( n4283 & n4284 ) ;
  assign n4287 = ( n1612 & n4285 ) | ( n1612 & n4286 ) | ( n4285 & n4286 ) ;
  assign n4288 = n4280 | n4287 ;
  assign n4289 = x487 & n812 ;
  assign n4290 = x487 & ~n815 ;
  assign n4291 = ( n909 & n4289 ) | ( n909 & n4290 ) | ( n4289 & n4290 ) ;
  assign n4292 = ( ~n929 & n4289 ) | ( ~n929 & n4290 ) | ( n4289 & n4290 ) ;
  assign n4293 = ( n800 & n4291 ) | ( n800 & n4292 ) | ( n4291 & n4292 ) ;
  assign n4294 = ( ~n948 & n4291 ) | ( ~n948 & n4292 ) | ( n4291 & n4292 ) ;
  assign n4295 = ( ~n1061 & n4293 ) | ( ~n1061 & n4294 ) | ( n4293 & n4294 ) ;
  assign n4296 = x359 & ~n812 ;
  assign n4297 = x359 & n815 ;
  assign n4298 = ( ~n909 & n4296 ) | ( ~n909 & n4297 ) | ( n4296 & n4297 ) ;
  assign n4299 = ( n929 & n4296 ) | ( n929 & n4297 ) | ( n4296 & n4297 ) ;
  assign n4300 = ( ~n800 & n4298 ) | ( ~n800 & n4299 ) | ( n4298 & n4299 ) ;
  assign n4301 = ( n948 & n4298 ) | ( n948 & n4299 ) | ( n4298 & n4299 ) ;
  assign n4302 = ( n1061 & n4300 ) | ( n1061 & n4301 ) | ( n4300 & n4301 ) ;
  assign n4303 = n4295 | n4302 ;
  assign n4304 = n4288 & ~n4303 ;
  assign n4305 = ~n4273 & n4304 ;
  assign n4306 = ~n4288 & n4303 ;
  assign n4307 = x486 & n812 ;
  assign n4308 = x486 & ~n815 ;
  assign n4309 = ( n909 & n4307 ) | ( n909 & n4308 ) | ( n4307 & n4308 ) ;
  assign n4310 = ( ~n929 & n4307 ) | ( ~n929 & n4308 ) | ( n4307 & n4308 ) ;
  assign n4311 = ( n800 & n4309 ) | ( n800 & n4310 ) | ( n4309 & n4310 ) ;
  assign n4312 = ( ~n948 & n4309 ) | ( ~n948 & n4310 ) | ( n4309 & n4310 ) ;
  assign n4313 = ( ~n1061 & n4311 ) | ( ~n1061 & n4312 ) | ( n4311 & n4312 ) ;
  assign n4314 = x358 & ~n812 ;
  assign n4315 = x358 & n815 ;
  assign n4316 = ( ~n909 & n4314 ) | ( ~n909 & n4315 ) | ( n4314 & n4315 ) ;
  assign n4317 = ( n929 & n4314 ) | ( n929 & n4315 ) | ( n4314 & n4315 ) ;
  assign n4318 = ( ~n800 & n4316 ) | ( ~n800 & n4317 ) | ( n4316 & n4317 ) ;
  assign n4319 = ( n948 & n4316 ) | ( n948 & n4317 ) | ( n4316 & n4317 ) ;
  assign n4320 = ( n1061 & n4318 ) | ( n1061 & n4319 ) | ( n4318 & n4319 ) ;
  assign n4321 = n4313 | n4320 ;
  assign n4322 = x230 & n1370 ;
  assign n4323 = x230 & ~n1373 ;
  assign n4324 = ( n1467 & n4322 ) | ( n1467 & n4323 ) | ( n4322 & n4323 ) ;
  assign n4325 = ( ~n1487 & n4322 ) | ( ~n1487 & n4323 ) | ( n4322 & n4323 ) ;
  assign n4326 = ( n1358 & n4324 ) | ( n1358 & n4325 ) | ( n4324 & n4325 ) ;
  assign n4327 = ( ~n1506 & n4324 ) | ( ~n1506 & n4325 ) | ( n4324 & n4325 ) ;
  assign n4328 = ( ~n1612 & n4326 ) | ( ~n1612 & n4327 ) | ( n4326 & n4327 ) ;
  assign n4329 = x102 & ~n1370 ;
  assign n4330 = x102 & n1373 ;
  assign n4331 = ( ~n1467 & n4329 ) | ( ~n1467 & n4330 ) | ( n4329 & n4330 ) ;
  assign n4332 = ( n1487 & n4329 ) | ( n1487 & n4330 ) | ( n4329 & n4330 ) ;
  assign n4333 = ( ~n1358 & n4331 ) | ( ~n1358 & n4332 ) | ( n4331 & n4332 ) ;
  assign n4334 = ( n1506 & n4331 ) | ( n1506 & n4332 ) | ( n4331 & n4332 ) ;
  assign n4335 = ( n1612 & n4333 ) | ( n1612 & n4334 ) | ( n4333 & n4334 ) ;
  assign n4336 = n4328 | n4335 ;
  assign n4337 = n4321 & ~n4336 ;
  assign n4338 = n4306 | n4337 ;
  assign n4339 = x229 & n1370 ;
  assign n4340 = x229 & ~n1373 ;
  assign n4341 = ( n1467 & n4339 ) | ( n1467 & n4340 ) | ( n4339 & n4340 ) ;
  assign n4342 = ( ~n1487 & n4339 ) | ( ~n1487 & n4340 ) | ( n4339 & n4340 ) ;
  assign n4343 = ( n1358 & n4341 ) | ( n1358 & n4342 ) | ( n4341 & n4342 ) ;
  assign n4344 = ( ~n1506 & n4341 ) | ( ~n1506 & n4342 ) | ( n4341 & n4342 ) ;
  assign n4345 = ( ~n1612 & n4343 ) | ( ~n1612 & n4344 ) | ( n4343 & n4344 ) ;
  assign n4346 = x101 & ~n1370 ;
  assign n4347 = x101 & n1373 ;
  assign n4348 = ( ~n1467 & n4346 ) | ( ~n1467 & n4347 ) | ( n4346 & n4347 ) ;
  assign n4349 = ( n1487 & n4346 ) | ( n1487 & n4347 ) | ( n4346 & n4347 ) ;
  assign n4350 = ( ~n1358 & n4348 ) | ( ~n1358 & n4349 ) | ( n4348 & n4349 ) ;
  assign n4351 = ( n1506 & n4348 ) | ( n1506 & n4349 ) | ( n4348 & n4349 ) ;
  assign n4352 = ( n1612 & n4350 ) | ( n1612 & n4351 ) | ( n4350 & n4351 ) ;
  assign n4353 = n4345 | n4352 ;
  assign n4354 = x485 & n812 ;
  assign n4355 = x485 & ~n815 ;
  assign n4356 = ( n909 & n4354 ) | ( n909 & n4355 ) | ( n4354 & n4355 ) ;
  assign n4357 = ( ~n929 & n4354 ) | ( ~n929 & n4355 ) | ( n4354 & n4355 ) ;
  assign n4358 = ( n800 & n4356 ) | ( n800 & n4357 ) | ( n4356 & n4357 ) ;
  assign n4359 = ( ~n948 & n4356 ) | ( ~n948 & n4357 ) | ( n4356 & n4357 ) ;
  assign n4360 = ( ~n1061 & n4358 ) | ( ~n1061 & n4359 ) | ( n4358 & n4359 ) ;
  assign n4361 = x357 & ~n812 ;
  assign n4362 = x357 & n815 ;
  assign n4363 = ( ~n909 & n4361 ) | ( ~n909 & n4362 ) | ( n4361 & n4362 ) ;
  assign n4364 = ( n929 & n4361 ) | ( n929 & n4362 ) | ( n4361 & n4362 ) ;
  assign n4365 = ( ~n800 & n4363 ) | ( ~n800 & n4364 ) | ( n4363 & n4364 ) ;
  assign n4366 = ( n948 & n4363 ) | ( n948 & n4364 ) | ( n4363 & n4364 ) ;
  assign n4367 = ( n1061 & n4365 ) | ( n1061 & n4366 ) | ( n4365 & n4366 ) ;
  assign n4368 = n4360 | n4367 ;
  assign n4369 = x228 & n1370 ;
  assign n4370 = x228 & ~n1373 ;
  assign n4371 = ( n1467 & n4369 ) | ( n1467 & n4370 ) | ( n4369 & n4370 ) ;
  assign n4372 = ( ~n1487 & n4369 ) | ( ~n1487 & n4370 ) | ( n4369 & n4370 ) ;
  assign n4373 = ( n1358 & n4371 ) | ( n1358 & n4372 ) | ( n4371 & n4372 ) ;
  assign n4374 = ( ~n1506 & n4371 ) | ( ~n1506 & n4372 ) | ( n4371 & n4372 ) ;
  assign n4375 = ( ~n1612 & n4373 ) | ( ~n1612 & n4374 ) | ( n4373 & n4374 ) ;
  assign n4376 = x100 & ~n1370 ;
  assign n4377 = x100 & n1373 ;
  assign n4378 = ( ~n1467 & n4376 ) | ( ~n1467 & n4377 ) | ( n4376 & n4377 ) ;
  assign n4379 = ( n1487 & n4376 ) | ( n1487 & n4377 ) | ( n4376 & n4377 ) ;
  assign n4380 = ( ~n1358 & n4378 ) | ( ~n1358 & n4379 ) | ( n4378 & n4379 ) ;
  assign n4381 = ( n1506 & n4378 ) | ( n1506 & n4379 ) | ( n4378 & n4379 ) ;
  assign n4382 = ( n1612 & n4380 ) | ( n1612 & n4381 ) | ( n4380 & n4381 ) ;
  assign n4383 = n4375 | n4382 ;
  assign n4384 = x484 & n812 ;
  assign n4385 = x484 & ~n815 ;
  assign n4386 = ( n909 & n4384 ) | ( n909 & n4385 ) | ( n4384 & n4385 ) ;
  assign n4387 = ( ~n929 & n4384 ) | ( ~n929 & n4385 ) | ( n4384 & n4385 ) ;
  assign n4388 = ( n800 & n4386 ) | ( n800 & n4387 ) | ( n4386 & n4387 ) ;
  assign n4389 = ( ~n948 & n4386 ) | ( ~n948 & n4387 ) | ( n4386 & n4387 ) ;
  assign n4390 = ( ~n1061 & n4388 ) | ( ~n1061 & n4389 ) | ( n4388 & n4389 ) ;
  assign n4391 = x356 & ~n812 ;
  assign n4392 = x356 & n815 ;
  assign n4393 = ( ~n909 & n4391 ) | ( ~n909 & n4392 ) | ( n4391 & n4392 ) ;
  assign n4394 = ( n929 & n4391 ) | ( n929 & n4392 ) | ( n4391 & n4392 ) ;
  assign n4395 = ( ~n800 & n4393 ) | ( ~n800 & n4394 ) | ( n4393 & n4394 ) ;
  assign n4396 = ( n948 & n4393 ) | ( n948 & n4394 ) | ( n4393 & n4394 ) ;
  assign n4397 = ( n1061 & n4395 ) | ( n1061 & n4396 ) | ( n4395 & n4396 ) ;
  assign n4398 = n4390 | n4397 ;
  assign n4399 = n4383 & ~n4398 ;
  assign n4400 = ( n4353 & ~n4368 ) | ( n4353 & n4399 ) | ( ~n4368 & n4399 ) ;
  assign n4401 = ~n4338 & n4400 ;
  assign n4402 = ~n4321 & n4336 ;
  assign n4403 = ~n4306 & n4402 ;
  assign n4404 = ~n4353 & n4368 ;
  assign n4405 = ~n4383 & n4398 ;
  assign n4406 = n4404 | n4405 ;
  assign n4407 = n4338 | n4406 ;
  assign n4408 = ~n4403 & n4407 ;
  assign n4409 = x227 & n1370 ;
  assign n4410 = x227 & ~n1373 ;
  assign n4411 = ( n1467 & n4409 ) | ( n1467 & n4410 ) | ( n4409 & n4410 ) ;
  assign n4412 = ( ~n1487 & n4409 ) | ( ~n1487 & n4410 ) | ( n4409 & n4410 ) ;
  assign n4413 = ( n1358 & n4411 ) | ( n1358 & n4412 ) | ( n4411 & n4412 ) ;
  assign n4414 = ( ~n1506 & n4411 ) | ( ~n1506 & n4412 ) | ( n4411 & n4412 ) ;
  assign n4415 = ( ~n1612 & n4413 ) | ( ~n1612 & n4414 ) | ( n4413 & n4414 ) ;
  assign n4416 = x99 & ~n1370 ;
  assign n4417 = x99 & n1373 ;
  assign n4418 = ( ~n1467 & n4416 ) | ( ~n1467 & n4417 ) | ( n4416 & n4417 ) ;
  assign n4419 = ( n1487 & n4416 ) | ( n1487 & n4417 ) | ( n4416 & n4417 ) ;
  assign n4420 = ( ~n1358 & n4418 ) | ( ~n1358 & n4419 ) | ( n4418 & n4419 ) ;
  assign n4421 = ( n1506 & n4418 ) | ( n1506 & n4419 ) | ( n4418 & n4419 ) ;
  assign n4422 = ( n1612 & n4420 ) | ( n1612 & n4421 ) | ( n4420 & n4421 ) ;
  assign n4423 = n4415 | n4422 ;
  assign n4424 = x483 & n812 ;
  assign n4425 = x483 & ~n815 ;
  assign n4426 = ( n909 & n4424 ) | ( n909 & n4425 ) | ( n4424 & n4425 ) ;
  assign n4427 = ( ~n929 & n4424 ) | ( ~n929 & n4425 ) | ( n4424 & n4425 ) ;
  assign n4428 = ( n800 & n4426 ) | ( n800 & n4427 ) | ( n4426 & n4427 ) ;
  assign n4429 = ( ~n948 & n4426 ) | ( ~n948 & n4427 ) | ( n4426 & n4427 ) ;
  assign n4430 = ( ~n1061 & n4428 ) | ( ~n1061 & n4429 ) | ( n4428 & n4429 ) ;
  assign n4431 = x355 & ~n812 ;
  assign n4432 = x355 & n815 ;
  assign n4433 = ( ~n909 & n4431 ) | ( ~n909 & n4432 ) | ( n4431 & n4432 ) ;
  assign n4434 = ( n929 & n4431 ) | ( n929 & n4432 ) | ( n4431 & n4432 ) ;
  assign n4435 = ( ~n800 & n4433 ) | ( ~n800 & n4434 ) | ( n4433 & n4434 ) ;
  assign n4436 = ( n948 & n4433 ) | ( n948 & n4434 ) | ( n4433 & n4434 ) ;
  assign n4437 = ( n1061 & n4435 ) | ( n1061 & n4436 ) | ( n4435 & n4436 ) ;
  assign n4438 = n4430 | n4437 ;
  assign n4439 = x482 & n812 ;
  assign n4440 = x482 & ~n815 ;
  assign n4441 = ( n909 & n4439 ) | ( n909 & n4440 ) | ( n4439 & n4440 ) ;
  assign n4442 = ( ~n929 & n4439 ) | ( ~n929 & n4440 ) | ( n4439 & n4440 ) ;
  assign n4443 = ( n800 & n4441 ) | ( n800 & n4442 ) | ( n4441 & n4442 ) ;
  assign n4444 = ( ~n948 & n4441 ) | ( ~n948 & n4442 ) | ( n4441 & n4442 ) ;
  assign n4445 = ( ~n1061 & n4443 ) | ( ~n1061 & n4444 ) | ( n4443 & n4444 ) ;
  assign n4446 = x354 & ~n812 ;
  assign n4447 = x354 & n815 ;
  assign n4448 = ( ~n909 & n4446 ) | ( ~n909 & n4447 ) | ( n4446 & n4447 ) ;
  assign n4449 = ( n929 & n4446 ) | ( n929 & n4447 ) | ( n4446 & n4447 ) ;
  assign n4450 = ( ~n800 & n4448 ) | ( ~n800 & n4449 ) | ( n4448 & n4449 ) ;
  assign n4451 = ( n948 & n4448 ) | ( n948 & n4449 ) | ( n4448 & n4449 ) ;
  assign n4452 = ( n1061 & n4450 ) | ( n1061 & n4451 ) | ( n4450 & n4451 ) ;
  assign n4453 = n4445 | n4452 ;
  assign n4454 = x226 & n1370 ;
  assign n4455 = x226 & ~n1373 ;
  assign n4456 = ( n1467 & n4454 ) | ( n1467 & n4455 ) | ( n4454 & n4455 ) ;
  assign n4457 = ( ~n1487 & n4454 ) | ( ~n1487 & n4455 ) | ( n4454 & n4455 ) ;
  assign n4458 = ( n1358 & n4456 ) | ( n1358 & n4457 ) | ( n4456 & n4457 ) ;
  assign n4459 = ( ~n1506 & n4456 ) | ( ~n1506 & n4457 ) | ( n4456 & n4457 ) ;
  assign n4460 = ( ~n1612 & n4458 ) | ( ~n1612 & n4459 ) | ( n4458 & n4459 ) ;
  assign n4461 = x98 & ~n1370 ;
  assign n4462 = x98 & n1373 ;
  assign n4463 = ( ~n1467 & n4461 ) | ( ~n1467 & n4462 ) | ( n4461 & n4462 ) ;
  assign n4464 = ( n1487 & n4461 ) | ( n1487 & n4462 ) | ( n4461 & n4462 ) ;
  assign n4465 = ( ~n1358 & n4463 ) | ( ~n1358 & n4464 ) | ( n4463 & n4464 ) ;
  assign n4466 = ( n1506 & n4463 ) | ( n1506 & n4464 ) | ( n4463 & n4464 ) ;
  assign n4467 = ( n1612 & n4465 ) | ( n1612 & n4466 ) | ( n4465 & n4466 ) ;
  assign n4468 = n4460 | n4467 ;
  assign n4469 = x225 & n1370 ;
  assign n4470 = x225 & ~n1373 ;
  assign n4471 = ( n1467 & n4469 ) | ( n1467 & n4470 ) | ( n4469 & n4470 ) ;
  assign n4472 = ( ~n1487 & n4469 ) | ( ~n1487 & n4470 ) | ( n4469 & n4470 ) ;
  assign n4473 = ( n1358 & n4471 ) | ( n1358 & n4472 ) | ( n4471 & n4472 ) ;
  assign n4474 = ( ~n1506 & n4471 ) | ( ~n1506 & n4472 ) | ( n4471 & n4472 ) ;
  assign n4475 = ( ~n1612 & n4473 ) | ( ~n1612 & n4474 ) | ( n4473 & n4474 ) ;
  assign n4476 = x97 & ~n1370 ;
  assign n4477 = x97 & n1373 ;
  assign n4478 = ( ~n1467 & n4476 ) | ( ~n1467 & n4477 ) | ( n4476 & n4477 ) ;
  assign n4479 = ( n1487 & n4476 ) | ( n1487 & n4477 ) | ( n4476 & n4477 ) ;
  assign n4480 = ( ~n1358 & n4478 ) | ( ~n1358 & n4479 ) | ( n4478 & n4479 ) ;
  assign n4481 = ( n1506 & n4478 ) | ( n1506 & n4479 ) | ( n4478 & n4479 ) ;
  assign n4482 = ( n1612 & n4480 ) | ( n1612 & n4481 ) | ( n4480 & n4481 ) ;
  assign n4483 = n4475 | n4482 ;
  assign n4484 = x481 & n812 ;
  assign n4485 = x481 & ~n815 ;
  assign n4486 = ( n909 & n4484 ) | ( n909 & n4485 ) | ( n4484 & n4485 ) ;
  assign n4487 = ( ~n929 & n4484 ) | ( ~n929 & n4485 ) | ( n4484 & n4485 ) ;
  assign n4488 = ( n800 & n4486 ) | ( n800 & n4487 ) | ( n4486 & n4487 ) ;
  assign n4489 = ( ~n948 & n4486 ) | ( ~n948 & n4487 ) | ( n4486 & n4487 ) ;
  assign n4490 = ( ~n1061 & n4488 ) | ( ~n1061 & n4489 ) | ( n4488 & n4489 ) ;
  assign n4491 = x353 & ~n812 ;
  assign n4492 = x353 & n815 ;
  assign n4493 = ( ~n909 & n4491 ) | ( ~n909 & n4492 ) | ( n4491 & n4492 ) ;
  assign n4494 = ( n929 & n4491 ) | ( n929 & n4492 ) | ( n4491 & n4492 ) ;
  assign n4495 = ( ~n800 & n4493 ) | ( ~n800 & n4494 ) | ( n4493 & n4494 ) ;
  assign n4496 = ( n948 & n4493 ) | ( n948 & n4494 ) | ( n4493 & n4494 ) ;
  assign n4497 = ( n1061 & n4495 ) | ( n1061 & n4496 ) | ( n4495 & n4496 ) ;
  assign n4498 = n4490 | n4497 ;
  assign n4499 = x480 & n812 ;
  assign n4500 = x480 & ~n815 ;
  assign n4501 = ( n909 & n4499 ) | ( n909 & n4500 ) | ( n4499 & n4500 ) ;
  assign n4502 = ( ~n929 & n4499 ) | ( ~n929 & n4500 ) | ( n4499 & n4500 ) ;
  assign n4503 = ( n800 & n4501 ) | ( n800 & n4502 ) | ( n4501 & n4502 ) ;
  assign n4504 = ( ~n948 & n4501 ) | ( ~n948 & n4502 ) | ( n4501 & n4502 ) ;
  assign n4505 = ( ~n1061 & n4503 ) | ( ~n1061 & n4504 ) | ( n4503 & n4504 ) ;
  assign n4506 = x352 & ~n812 ;
  assign n4507 = x352 & n815 ;
  assign n4508 = ( ~n909 & n4506 ) | ( ~n909 & n4507 ) | ( n4506 & n4507 ) ;
  assign n4509 = ( n929 & n4506 ) | ( n929 & n4507 ) | ( n4506 & n4507 ) ;
  assign n4510 = ( ~n800 & n4508 ) | ( ~n800 & n4509 ) | ( n4508 & n4509 ) ;
  assign n4511 = ( n948 & n4508 ) | ( n948 & n4509 ) | ( n4508 & n4509 ) ;
  assign n4512 = ( n1061 & n4510 ) | ( n1061 & n4511 ) | ( n4510 & n4511 ) ;
  assign n4513 = n4505 | n4512 ;
  assign n4514 = x224 & n1370 ;
  assign n4515 = x224 & ~n1373 ;
  assign n4516 = ( n1467 & n4514 ) | ( n1467 & n4515 ) | ( n4514 & n4515 ) ;
  assign n4517 = ( ~n1487 & n4514 ) | ( ~n1487 & n4515 ) | ( n4514 & n4515 ) ;
  assign n4518 = ( n1358 & n4516 ) | ( n1358 & n4517 ) | ( n4516 & n4517 ) ;
  assign n4519 = ( ~n1506 & n4516 ) | ( ~n1506 & n4517 ) | ( n4516 & n4517 ) ;
  assign n4520 = ( ~n1612 & n4518 ) | ( ~n1612 & n4519 ) | ( n4518 & n4519 ) ;
  assign n4521 = x96 & ~n1370 ;
  assign n4522 = x96 & n1373 ;
  assign n4523 = ( ~n1467 & n4521 ) | ( ~n1467 & n4522 ) | ( n4521 & n4522 ) ;
  assign n4524 = ( n1487 & n4521 ) | ( n1487 & n4522 ) | ( n4521 & n4522 ) ;
  assign n4525 = ( ~n1358 & n4523 ) | ( ~n1358 & n4524 ) | ( n4523 & n4524 ) ;
  assign n4526 = ( n1506 & n4523 ) | ( n1506 & n4524 ) | ( n4523 & n4524 ) ;
  assign n4527 = ( n1612 & n4525 ) | ( n1612 & n4526 ) | ( n4525 & n4526 ) ;
  assign n4528 = n4520 | n4527 ;
  assign n4529 = ~n4513 & n4528 ;
  assign n4530 = ( n4483 & ~n4498 ) | ( n4483 & n4529 ) | ( ~n4498 & n4529 ) ;
  assign n4531 = ( ~n4453 & n4468 ) | ( ~n4453 & n4530 ) | ( n4468 & n4530 ) ;
  assign n4532 = ( n4423 & ~n4438 ) | ( n4423 & n4531 ) | ( ~n4438 & n4531 ) ;
  assign n4533 = ( n4403 & ~n4408 ) | ( n4403 & n4532 ) | ( ~n4408 & n4532 ) ;
  assign n4534 = n4401 | n4533 ;
  assign n4535 = ~n4483 & n4498 ;
  assign n4536 = x223 & n1370 ;
  assign n4537 = x223 & ~n1373 ;
  assign n4538 = ( n1467 & n4536 ) | ( n1467 & n4537 ) | ( n4536 & n4537 ) ;
  assign n4539 = ( ~n1487 & n4536 ) | ( ~n1487 & n4537 ) | ( n4536 & n4537 ) ;
  assign n4540 = ( n1358 & n4538 ) | ( n1358 & n4539 ) | ( n4538 & n4539 ) ;
  assign n4541 = ( ~n1506 & n4538 ) | ( ~n1506 & n4539 ) | ( n4538 & n4539 ) ;
  assign n4542 = ( ~n1612 & n4540 ) | ( ~n1612 & n4541 ) | ( n4540 & n4541 ) ;
  assign n4543 = x95 & ~n1370 ;
  assign n4544 = x95 & n1373 ;
  assign n4545 = ( ~n1467 & n4543 ) | ( ~n1467 & n4544 ) | ( n4543 & n4544 ) ;
  assign n4546 = ( n1487 & n4543 ) | ( n1487 & n4544 ) | ( n4543 & n4544 ) ;
  assign n4547 = ( ~n1358 & n4545 ) | ( ~n1358 & n4546 ) | ( n4545 & n4546 ) ;
  assign n4548 = ( n1506 & n4545 ) | ( n1506 & n4546 ) | ( n4545 & n4546 ) ;
  assign n4549 = ( n1612 & n4547 ) | ( n1612 & n4548 ) | ( n4547 & n4548 ) ;
  assign n4550 = n4542 | n4549 ;
  assign n4551 = x479 & n812 ;
  assign n4552 = x479 & ~n815 ;
  assign n4553 = ( n909 & n4551 ) | ( n909 & n4552 ) | ( n4551 & n4552 ) ;
  assign n4554 = ( ~n929 & n4551 ) | ( ~n929 & n4552 ) | ( n4551 & n4552 ) ;
  assign n4555 = ( n800 & n4553 ) | ( n800 & n4554 ) | ( n4553 & n4554 ) ;
  assign n4556 = ( ~n948 & n4553 ) | ( ~n948 & n4554 ) | ( n4553 & n4554 ) ;
  assign n4557 = ( ~n1061 & n4555 ) | ( ~n1061 & n4556 ) | ( n4555 & n4556 ) ;
  assign n4558 = x351 & ~n812 ;
  assign n4559 = x351 & n815 ;
  assign n4560 = ( ~n909 & n4558 ) | ( ~n909 & n4559 ) | ( n4558 & n4559 ) ;
  assign n4561 = ( n929 & n4558 ) | ( n929 & n4559 ) | ( n4558 & n4559 ) ;
  assign n4562 = ( ~n800 & n4560 ) | ( ~n800 & n4561 ) | ( n4560 & n4561 ) ;
  assign n4563 = ( n948 & n4560 ) | ( n948 & n4561 ) | ( n4560 & n4561 ) ;
  assign n4564 = ( n1061 & n4562 ) | ( n1061 & n4563 ) | ( n4562 & n4563 ) ;
  assign n4565 = n4557 | n4564 ;
  assign n4566 = x478 & n812 ;
  assign n4567 = x478 & ~n815 ;
  assign n4568 = ( n909 & n4566 ) | ( n909 & n4567 ) | ( n4566 & n4567 ) ;
  assign n4569 = ( ~n929 & n4566 ) | ( ~n929 & n4567 ) | ( n4566 & n4567 ) ;
  assign n4570 = ( n800 & n4568 ) | ( n800 & n4569 ) | ( n4568 & n4569 ) ;
  assign n4571 = ( ~n948 & n4568 ) | ( ~n948 & n4569 ) | ( n4568 & n4569 ) ;
  assign n4572 = ( ~n1061 & n4570 ) | ( ~n1061 & n4571 ) | ( n4570 & n4571 ) ;
  assign n4573 = x350 & ~n812 ;
  assign n4574 = x350 & n815 ;
  assign n4575 = ( ~n909 & n4573 ) | ( ~n909 & n4574 ) | ( n4573 & n4574 ) ;
  assign n4576 = ( n929 & n4573 ) | ( n929 & n4574 ) | ( n4573 & n4574 ) ;
  assign n4577 = ( ~n800 & n4575 ) | ( ~n800 & n4576 ) | ( n4575 & n4576 ) ;
  assign n4578 = ( n948 & n4575 ) | ( n948 & n4576 ) | ( n4575 & n4576 ) ;
  assign n4579 = ( n1061 & n4577 ) | ( n1061 & n4578 ) | ( n4577 & n4578 ) ;
  assign n4580 = n4572 | n4579 ;
  assign n4581 = x222 & n1370 ;
  assign n4582 = x222 & ~n1373 ;
  assign n4583 = ( n1467 & n4581 ) | ( n1467 & n4582 ) | ( n4581 & n4582 ) ;
  assign n4584 = ( ~n1487 & n4581 ) | ( ~n1487 & n4582 ) | ( n4581 & n4582 ) ;
  assign n4585 = ( n1358 & n4583 ) | ( n1358 & n4584 ) | ( n4583 & n4584 ) ;
  assign n4586 = ( ~n1506 & n4583 ) | ( ~n1506 & n4584 ) | ( n4583 & n4584 ) ;
  assign n4587 = ( ~n1612 & n4585 ) | ( ~n1612 & n4586 ) | ( n4585 & n4586 ) ;
  assign n4588 = x94 & ~n1370 ;
  assign n4589 = x94 & n1373 ;
  assign n4590 = ( ~n1467 & n4588 ) | ( ~n1467 & n4589 ) | ( n4588 & n4589 ) ;
  assign n4591 = ( n1487 & n4588 ) | ( n1487 & n4589 ) | ( n4588 & n4589 ) ;
  assign n4592 = ( ~n1358 & n4590 ) | ( ~n1358 & n4591 ) | ( n4590 & n4591 ) ;
  assign n4593 = ( n1506 & n4590 ) | ( n1506 & n4591 ) | ( n4590 & n4591 ) ;
  assign n4594 = ( n1612 & n4592 ) | ( n1612 & n4593 ) | ( n4592 & n4593 ) ;
  assign n4595 = n4587 | n4594 ;
  assign n4596 = x221 & n1370 ;
  assign n4597 = x221 & ~n1373 ;
  assign n4598 = ( n1467 & n4596 ) | ( n1467 & n4597 ) | ( n4596 & n4597 ) ;
  assign n4599 = ( ~n1487 & n4596 ) | ( ~n1487 & n4597 ) | ( n4596 & n4597 ) ;
  assign n4600 = ( n1358 & n4598 ) | ( n1358 & n4599 ) | ( n4598 & n4599 ) ;
  assign n4601 = ( ~n1506 & n4598 ) | ( ~n1506 & n4599 ) | ( n4598 & n4599 ) ;
  assign n4602 = ( ~n1612 & n4600 ) | ( ~n1612 & n4601 ) | ( n4600 & n4601 ) ;
  assign n4603 = x93 & ~n1370 ;
  assign n4604 = x93 & n1373 ;
  assign n4605 = ( ~n1467 & n4603 ) | ( ~n1467 & n4604 ) | ( n4603 & n4604 ) ;
  assign n4606 = ( n1487 & n4603 ) | ( n1487 & n4604 ) | ( n4603 & n4604 ) ;
  assign n4607 = ( ~n1358 & n4605 ) | ( ~n1358 & n4606 ) | ( n4605 & n4606 ) ;
  assign n4608 = ( n1506 & n4605 ) | ( n1506 & n4606 ) | ( n4605 & n4606 ) ;
  assign n4609 = ( n1612 & n4607 ) | ( n1612 & n4608 ) | ( n4607 & n4608 ) ;
  assign n4610 = n4602 | n4609 ;
  assign n4611 = x477 & n812 ;
  assign n4612 = x477 & ~n815 ;
  assign n4613 = ( n909 & n4611 ) | ( n909 & n4612 ) | ( n4611 & n4612 ) ;
  assign n4614 = ( ~n929 & n4611 ) | ( ~n929 & n4612 ) | ( n4611 & n4612 ) ;
  assign n4615 = ( n800 & n4613 ) | ( n800 & n4614 ) | ( n4613 & n4614 ) ;
  assign n4616 = ( ~n948 & n4613 ) | ( ~n948 & n4614 ) | ( n4613 & n4614 ) ;
  assign n4617 = ( ~n1061 & n4615 ) | ( ~n1061 & n4616 ) | ( n4615 & n4616 ) ;
  assign n4618 = x349 & ~n812 ;
  assign n4619 = x349 & n815 ;
  assign n4620 = ( ~n909 & n4618 ) | ( ~n909 & n4619 ) | ( n4618 & n4619 ) ;
  assign n4621 = ( n929 & n4618 ) | ( n929 & n4619 ) | ( n4618 & n4619 ) ;
  assign n4622 = ( ~n800 & n4620 ) | ( ~n800 & n4621 ) | ( n4620 & n4621 ) ;
  assign n4623 = ( n948 & n4620 ) | ( n948 & n4621 ) | ( n4620 & n4621 ) ;
  assign n4624 = ( n1061 & n4622 ) | ( n1061 & n4623 ) | ( n4622 & n4623 ) ;
  assign n4625 = n4617 | n4624 ;
  assign n4626 = x220 & n1370 ;
  assign n4627 = x220 & ~n1373 ;
  assign n4628 = ( n1467 & n4626 ) | ( n1467 & n4627 ) | ( n4626 & n4627 ) ;
  assign n4629 = ( ~n1487 & n4626 ) | ( ~n1487 & n4627 ) | ( n4626 & n4627 ) ;
  assign n4630 = ( n1358 & n4628 ) | ( n1358 & n4629 ) | ( n4628 & n4629 ) ;
  assign n4631 = ( ~n1506 & n4628 ) | ( ~n1506 & n4629 ) | ( n4628 & n4629 ) ;
  assign n4632 = ( ~n1612 & n4630 ) | ( ~n1612 & n4631 ) | ( n4630 & n4631 ) ;
  assign n4633 = x92 & ~n1370 ;
  assign n4634 = x92 & n1373 ;
  assign n4635 = ( ~n1467 & n4633 ) | ( ~n1467 & n4634 ) | ( n4633 & n4634 ) ;
  assign n4636 = ( n1487 & n4633 ) | ( n1487 & n4634 ) | ( n4633 & n4634 ) ;
  assign n4637 = ( ~n1358 & n4635 ) | ( ~n1358 & n4636 ) | ( n4635 & n4636 ) ;
  assign n4638 = ( n1506 & n4635 ) | ( n1506 & n4636 ) | ( n4635 & n4636 ) ;
  assign n4639 = ( n1612 & n4637 ) | ( n1612 & n4638 ) | ( n4637 & n4638 ) ;
  assign n4640 = n4632 | n4639 ;
  assign n4641 = x476 & n812 ;
  assign n4642 = x476 & ~n815 ;
  assign n4643 = ( n909 & n4641 ) | ( n909 & n4642 ) | ( n4641 & n4642 ) ;
  assign n4644 = ( ~n929 & n4641 ) | ( ~n929 & n4642 ) | ( n4641 & n4642 ) ;
  assign n4645 = ( n800 & n4643 ) | ( n800 & n4644 ) | ( n4643 & n4644 ) ;
  assign n4646 = ( ~n948 & n4643 ) | ( ~n948 & n4644 ) | ( n4643 & n4644 ) ;
  assign n4647 = ( ~n1061 & n4645 ) | ( ~n1061 & n4646 ) | ( n4645 & n4646 ) ;
  assign n4648 = x348 & ~n812 ;
  assign n4649 = x348 & n815 ;
  assign n4650 = ( ~n909 & n4648 ) | ( ~n909 & n4649 ) | ( n4648 & n4649 ) ;
  assign n4651 = ( n929 & n4648 ) | ( n929 & n4649 ) | ( n4648 & n4649 ) ;
  assign n4652 = ( ~n800 & n4650 ) | ( ~n800 & n4651 ) | ( n4650 & n4651 ) ;
  assign n4653 = ( n948 & n4650 ) | ( n948 & n4651 ) | ( n4650 & n4651 ) ;
  assign n4654 = ( n1061 & n4652 ) | ( n1061 & n4653 ) | ( n4652 & n4653 ) ;
  assign n4655 = n4647 | n4654 ;
  assign n4656 = n4640 & ~n4655 ;
  assign n4657 = ( n4610 & ~n4625 ) | ( n4610 & n4656 ) | ( ~n4625 & n4656 ) ;
  assign n4658 = ( ~n4580 & n4595 ) | ( ~n4580 & n4657 ) | ( n4595 & n4657 ) ;
  assign n4659 = ( n4550 & ~n4565 ) | ( n4550 & n4658 ) | ( ~n4565 & n4658 ) ;
  assign n4660 = ~n4535 & n4659 ;
  assign n4661 = n4453 & ~n4468 ;
  assign n4662 = ~n4423 & n4438 ;
  assign n4663 = n4661 | n4662 ;
  assign n4664 = n4513 & ~n4528 ;
  assign n4665 = n4663 | n4664 ;
  assign n4666 = n4407 | n4665 ;
  assign n4667 = ~n4534 & n4666 ;
  assign n4668 = ( n4534 & n4660 ) | ( n4534 & ~n4667 ) | ( n4660 & ~n4667 ) ;
  assign n4669 = ( ~n4534 & n4535 ) | ( ~n4534 & n4667 ) | ( n4535 & n4667 ) ;
  assign n4670 = x215 & n1370 ;
  assign n4671 = x215 & ~n1373 ;
  assign n4672 = ( n1467 & n4670 ) | ( n1467 & n4671 ) | ( n4670 & n4671 ) ;
  assign n4673 = ( ~n1487 & n4670 ) | ( ~n1487 & n4671 ) | ( n4670 & n4671 ) ;
  assign n4674 = ( n1358 & n4672 ) | ( n1358 & n4673 ) | ( n4672 & n4673 ) ;
  assign n4675 = ( ~n1506 & n4672 ) | ( ~n1506 & n4673 ) | ( n4672 & n4673 ) ;
  assign n4676 = ( ~n1612 & n4674 ) | ( ~n1612 & n4675 ) | ( n4674 & n4675 ) ;
  assign n4677 = x87 & ~n1370 ;
  assign n4678 = x87 & n1373 ;
  assign n4679 = ( ~n1467 & n4677 ) | ( ~n1467 & n4678 ) | ( n4677 & n4678 ) ;
  assign n4680 = ( n1487 & n4677 ) | ( n1487 & n4678 ) | ( n4677 & n4678 ) ;
  assign n4681 = ( ~n1358 & n4679 ) | ( ~n1358 & n4680 ) | ( n4679 & n4680 ) ;
  assign n4682 = ( n1506 & n4679 ) | ( n1506 & n4680 ) | ( n4679 & n4680 ) ;
  assign n4683 = ( n1612 & n4681 ) | ( n1612 & n4682 ) | ( n4681 & n4682 ) ;
  assign n4684 = n4676 | n4683 ;
  assign n4685 = x471 & n812 ;
  assign n4686 = x471 & ~n815 ;
  assign n4687 = ( n909 & n4685 ) | ( n909 & n4686 ) | ( n4685 & n4686 ) ;
  assign n4688 = ( ~n929 & n4685 ) | ( ~n929 & n4686 ) | ( n4685 & n4686 ) ;
  assign n4689 = ( n800 & n4687 ) | ( n800 & n4688 ) | ( n4687 & n4688 ) ;
  assign n4690 = ( ~n948 & n4687 ) | ( ~n948 & n4688 ) | ( n4687 & n4688 ) ;
  assign n4691 = ( ~n1061 & n4689 ) | ( ~n1061 & n4690 ) | ( n4689 & n4690 ) ;
  assign n4692 = x343 & ~n812 ;
  assign n4693 = x343 & n815 ;
  assign n4694 = ( ~n909 & n4692 ) | ( ~n909 & n4693 ) | ( n4692 & n4693 ) ;
  assign n4695 = ( n929 & n4692 ) | ( n929 & n4693 ) | ( n4692 & n4693 ) ;
  assign n4696 = ( ~n800 & n4694 ) | ( ~n800 & n4695 ) | ( n4694 & n4695 ) ;
  assign n4697 = ( n948 & n4694 ) | ( n948 & n4695 ) | ( n4694 & n4695 ) ;
  assign n4698 = ( n1061 & n4696 ) | ( n1061 & n4697 ) | ( n4696 & n4697 ) ;
  assign n4699 = n4691 | n4698 ;
  assign n4700 = ~n4684 & n4699 ;
  assign n4701 = x470 & n812 ;
  assign n4702 = x470 & ~n815 ;
  assign n4703 = ( n909 & n4701 ) | ( n909 & n4702 ) | ( n4701 & n4702 ) ;
  assign n4704 = ( ~n929 & n4701 ) | ( ~n929 & n4702 ) | ( n4701 & n4702 ) ;
  assign n4705 = ( n800 & n4703 ) | ( n800 & n4704 ) | ( n4703 & n4704 ) ;
  assign n4706 = ( ~n948 & n4703 ) | ( ~n948 & n4704 ) | ( n4703 & n4704 ) ;
  assign n4707 = ( ~n1061 & n4705 ) | ( ~n1061 & n4706 ) | ( n4705 & n4706 ) ;
  assign n4708 = x342 & ~n812 ;
  assign n4709 = x342 & n815 ;
  assign n4710 = ( ~n909 & n4708 ) | ( ~n909 & n4709 ) | ( n4708 & n4709 ) ;
  assign n4711 = ( n929 & n4708 ) | ( n929 & n4709 ) | ( n4708 & n4709 ) ;
  assign n4712 = ( ~n800 & n4710 ) | ( ~n800 & n4711 ) | ( n4710 & n4711 ) ;
  assign n4713 = ( n948 & n4710 ) | ( n948 & n4711 ) | ( n4710 & n4711 ) ;
  assign n4714 = ( n1061 & n4712 ) | ( n1061 & n4713 ) | ( n4712 & n4713 ) ;
  assign n4715 = n4707 | n4714 ;
  assign n4716 = x214 & n1370 ;
  assign n4717 = x214 & ~n1373 ;
  assign n4718 = ( n1467 & n4716 ) | ( n1467 & n4717 ) | ( n4716 & n4717 ) ;
  assign n4719 = ( ~n1487 & n4716 ) | ( ~n1487 & n4717 ) | ( n4716 & n4717 ) ;
  assign n4720 = ( n1358 & n4718 ) | ( n1358 & n4719 ) | ( n4718 & n4719 ) ;
  assign n4721 = ( ~n1506 & n4718 ) | ( ~n1506 & n4719 ) | ( n4718 & n4719 ) ;
  assign n4722 = ( ~n1612 & n4720 ) | ( ~n1612 & n4721 ) | ( n4720 & n4721 ) ;
  assign n4723 = x86 & ~n1370 ;
  assign n4724 = x86 & n1373 ;
  assign n4725 = ( ~n1467 & n4723 ) | ( ~n1467 & n4724 ) | ( n4723 & n4724 ) ;
  assign n4726 = ( n1487 & n4723 ) | ( n1487 & n4724 ) | ( n4723 & n4724 ) ;
  assign n4727 = ( ~n1358 & n4725 ) | ( ~n1358 & n4726 ) | ( n4725 & n4726 ) ;
  assign n4728 = ( n1506 & n4725 ) | ( n1506 & n4726 ) | ( n4725 & n4726 ) ;
  assign n4729 = ( n1612 & n4727 ) | ( n1612 & n4728 ) | ( n4727 & n4728 ) ;
  assign n4730 = n4722 | n4729 ;
  assign n4731 = n4715 & ~n4730 ;
  assign n4732 = n4700 | n4731 ;
  assign n4733 = x213 & n1370 ;
  assign n4734 = x213 & ~n1373 ;
  assign n4735 = ( n1467 & n4733 ) | ( n1467 & n4734 ) | ( n4733 & n4734 ) ;
  assign n4736 = ( ~n1487 & n4733 ) | ( ~n1487 & n4734 ) | ( n4733 & n4734 ) ;
  assign n4737 = ( n1358 & n4735 ) | ( n1358 & n4736 ) | ( n4735 & n4736 ) ;
  assign n4738 = ( ~n1506 & n4735 ) | ( ~n1506 & n4736 ) | ( n4735 & n4736 ) ;
  assign n4739 = ( ~n1612 & n4737 ) | ( ~n1612 & n4738 ) | ( n4737 & n4738 ) ;
  assign n4740 = x85 & ~n1370 ;
  assign n4741 = x85 & n1373 ;
  assign n4742 = ( ~n1467 & n4740 ) | ( ~n1467 & n4741 ) | ( n4740 & n4741 ) ;
  assign n4743 = ( n1487 & n4740 ) | ( n1487 & n4741 ) | ( n4740 & n4741 ) ;
  assign n4744 = ( ~n1358 & n4742 ) | ( ~n1358 & n4743 ) | ( n4742 & n4743 ) ;
  assign n4745 = ( n1506 & n4742 ) | ( n1506 & n4743 ) | ( n4742 & n4743 ) ;
  assign n4746 = ( n1612 & n4744 ) | ( n1612 & n4745 ) | ( n4744 & n4745 ) ;
  assign n4747 = n4739 | n4746 ;
  assign n4748 = x469 & n812 ;
  assign n4749 = x469 & ~n815 ;
  assign n4750 = ( n909 & n4748 ) | ( n909 & n4749 ) | ( n4748 & n4749 ) ;
  assign n4751 = ( ~n929 & n4748 ) | ( ~n929 & n4749 ) | ( n4748 & n4749 ) ;
  assign n4752 = ( n800 & n4750 ) | ( n800 & n4751 ) | ( n4750 & n4751 ) ;
  assign n4753 = ( ~n948 & n4750 ) | ( ~n948 & n4751 ) | ( n4750 & n4751 ) ;
  assign n4754 = ( ~n1061 & n4752 ) | ( ~n1061 & n4753 ) | ( n4752 & n4753 ) ;
  assign n4755 = x341 & ~n812 ;
  assign n4756 = x341 & n815 ;
  assign n4757 = ( ~n909 & n4755 ) | ( ~n909 & n4756 ) | ( n4755 & n4756 ) ;
  assign n4758 = ( n929 & n4755 ) | ( n929 & n4756 ) | ( n4755 & n4756 ) ;
  assign n4759 = ( ~n800 & n4757 ) | ( ~n800 & n4758 ) | ( n4757 & n4758 ) ;
  assign n4760 = ( n948 & n4757 ) | ( n948 & n4758 ) | ( n4757 & n4758 ) ;
  assign n4761 = ( n1061 & n4759 ) | ( n1061 & n4760 ) | ( n4759 & n4760 ) ;
  assign n4762 = n4754 | n4761 ;
  assign n4763 = ~n4747 & n4762 ;
  assign n4764 = x212 & n1370 ;
  assign n4765 = x212 & ~n1373 ;
  assign n4766 = ( n1467 & n4764 ) | ( n1467 & n4765 ) | ( n4764 & n4765 ) ;
  assign n4767 = ( ~n1487 & n4764 ) | ( ~n1487 & n4765 ) | ( n4764 & n4765 ) ;
  assign n4768 = ( n1358 & n4766 ) | ( n1358 & n4767 ) | ( n4766 & n4767 ) ;
  assign n4769 = ( ~n1506 & n4766 ) | ( ~n1506 & n4767 ) | ( n4766 & n4767 ) ;
  assign n4770 = ( ~n1612 & n4768 ) | ( ~n1612 & n4769 ) | ( n4768 & n4769 ) ;
  assign n4771 = x84 & ~n1370 ;
  assign n4772 = x84 & n1373 ;
  assign n4773 = ( ~n1467 & n4771 ) | ( ~n1467 & n4772 ) | ( n4771 & n4772 ) ;
  assign n4774 = ( n1487 & n4771 ) | ( n1487 & n4772 ) | ( n4771 & n4772 ) ;
  assign n4775 = ( ~n1358 & n4773 ) | ( ~n1358 & n4774 ) | ( n4773 & n4774 ) ;
  assign n4776 = ( n1506 & n4773 ) | ( n1506 & n4774 ) | ( n4773 & n4774 ) ;
  assign n4777 = ( n1612 & n4775 ) | ( n1612 & n4776 ) | ( n4775 & n4776 ) ;
  assign n4778 = n4770 | n4777 ;
  assign n4779 = x468 & n812 ;
  assign n4780 = x468 & ~n815 ;
  assign n4781 = ( n909 & n4779 ) | ( n909 & n4780 ) | ( n4779 & n4780 ) ;
  assign n4782 = ( ~n929 & n4779 ) | ( ~n929 & n4780 ) | ( n4779 & n4780 ) ;
  assign n4783 = ( n800 & n4781 ) | ( n800 & n4782 ) | ( n4781 & n4782 ) ;
  assign n4784 = ( ~n948 & n4781 ) | ( ~n948 & n4782 ) | ( n4781 & n4782 ) ;
  assign n4785 = ( ~n1061 & n4783 ) | ( ~n1061 & n4784 ) | ( n4783 & n4784 ) ;
  assign n4786 = x340 & ~n812 ;
  assign n4787 = x340 & n815 ;
  assign n4788 = ( ~n909 & n4786 ) | ( ~n909 & n4787 ) | ( n4786 & n4787 ) ;
  assign n4789 = ( n929 & n4786 ) | ( n929 & n4787 ) | ( n4786 & n4787 ) ;
  assign n4790 = ( ~n800 & n4788 ) | ( ~n800 & n4789 ) | ( n4788 & n4789 ) ;
  assign n4791 = ( n948 & n4788 ) | ( n948 & n4789 ) | ( n4788 & n4789 ) ;
  assign n4792 = ( n1061 & n4790 ) | ( n1061 & n4791 ) | ( n4790 & n4791 ) ;
  assign n4793 = n4785 | n4792 ;
  assign n4794 = ~n4778 & n4793 ;
  assign n4795 = n4763 | n4794 ;
  assign n4796 = n4732 | n4795 ;
  assign n4797 = x211 & n1370 ;
  assign n4798 = x211 & ~n1373 ;
  assign n4799 = ( n1467 & n4797 ) | ( n1467 & n4798 ) | ( n4797 & n4798 ) ;
  assign n4800 = ( ~n1487 & n4797 ) | ( ~n1487 & n4798 ) | ( n4797 & n4798 ) ;
  assign n4801 = ( n1358 & n4799 ) | ( n1358 & n4800 ) | ( n4799 & n4800 ) ;
  assign n4802 = ( ~n1506 & n4799 ) | ( ~n1506 & n4800 ) | ( n4799 & n4800 ) ;
  assign n4803 = ( ~n1612 & n4801 ) | ( ~n1612 & n4802 ) | ( n4801 & n4802 ) ;
  assign n4804 = x83 & ~n1370 ;
  assign n4805 = x83 & n1373 ;
  assign n4806 = ( ~n1467 & n4804 ) | ( ~n1467 & n4805 ) | ( n4804 & n4805 ) ;
  assign n4807 = ( n1487 & n4804 ) | ( n1487 & n4805 ) | ( n4804 & n4805 ) ;
  assign n4808 = ( ~n1358 & n4806 ) | ( ~n1358 & n4807 ) | ( n4806 & n4807 ) ;
  assign n4809 = ( n1506 & n4806 ) | ( n1506 & n4807 ) | ( n4806 & n4807 ) ;
  assign n4810 = ( n1612 & n4808 ) | ( n1612 & n4809 ) | ( n4808 & n4809 ) ;
  assign n4811 = n4803 | n4810 ;
  assign n4812 = x467 & n812 ;
  assign n4813 = x467 & ~n815 ;
  assign n4814 = ( n909 & n4812 ) | ( n909 & n4813 ) | ( n4812 & n4813 ) ;
  assign n4815 = ( ~n929 & n4812 ) | ( ~n929 & n4813 ) | ( n4812 & n4813 ) ;
  assign n4816 = ( n800 & n4814 ) | ( n800 & n4815 ) | ( n4814 & n4815 ) ;
  assign n4817 = ( ~n948 & n4814 ) | ( ~n948 & n4815 ) | ( n4814 & n4815 ) ;
  assign n4818 = ( ~n1061 & n4816 ) | ( ~n1061 & n4817 ) | ( n4816 & n4817 ) ;
  assign n4819 = x339 & ~n812 ;
  assign n4820 = x339 & n815 ;
  assign n4821 = ( ~n909 & n4819 ) | ( ~n909 & n4820 ) | ( n4819 & n4820 ) ;
  assign n4822 = ( n929 & n4819 ) | ( n929 & n4820 ) | ( n4819 & n4820 ) ;
  assign n4823 = ( ~n800 & n4821 ) | ( ~n800 & n4822 ) | ( n4821 & n4822 ) ;
  assign n4824 = ( n948 & n4821 ) | ( n948 & n4822 ) | ( n4821 & n4822 ) ;
  assign n4825 = ( n1061 & n4823 ) | ( n1061 & n4824 ) | ( n4823 & n4824 ) ;
  assign n4826 = n4818 | n4825 ;
  assign n4827 = ~n4811 & n4826 ;
  assign n4828 = x466 & n812 ;
  assign n4829 = x466 & ~n815 ;
  assign n4830 = ( n909 & n4828 ) | ( n909 & n4829 ) | ( n4828 & n4829 ) ;
  assign n4831 = ( ~n929 & n4828 ) | ( ~n929 & n4829 ) | ( n4828 & n4829 ) ;
  assign n4832 = ( n800 & n4830 ) | ( n800 & n4831 ) | ( n4830 & n4831 ) ;
  assign n4833 = ( ~n948 & n4830 ) | ( ~n948 & n4831 ) | ( n4830 & n4831 ) ;
  assign n4834 = ( ~n1061 & n4832 ) | ( ~n1061 & n4833 ) | ( n4832 & n4833 ) ;
  assign n4835 = x338 & ~n812 ;
  assign n4836 = x338 & n815 ;
  assign n4837 = ( ~n909 & n4835 ) | ( ~n909 & n4836 ) | ( n4835 & n4836 ) ;
  assign n4838 = ( n929 & n4835 ) | ( n929 & n4836 ) | ( n4835 & n4836 ) ;
  assign n4839 = ( ~n800 & n4837 ) | ( ~n800 & n4838 ) | ( n4837 & n4838 ) ;
  assign n4840 = ( n948 & n4837 ) | ( n948 & n4838 ) | ( n4837 & n4838 ) ;
  assign n4841 = ( n1061 & n4839 ) | ( n1061 & n4840 ) | ( n4839 & n4840 ) ;
  assign n4842 = n4834 | n4841 ;
  assign n4843 = x210 & n1370 ;
  assign n4844 = x210 & ~n1373 ;
  assign n4845 = ( n1467 & n4843 ) | ( n1467 & n4844 ) | ( n4843 & n4844 ) ;
  assign n4846 = ( ~n1487 & n4843 ) | ( ~n1487 & n4844 ) | ( n4843 & n4844 ) ;
  assign n4847 = ( n1358 & n4845 ) | ( n1358 & n4846 ) | ( n4845 & n4846 ) ;
  assign n4848 = ( ~n1506 & n4845 ) | ( ~n1506 & n4846 ) | ( n4845 & n4846 ) ;
  assign n4849 = ( ~n1612 & n4847 ) | ( ~n1612 & n4848 ) | ( n4847 & n4848 ) ;
  assign n4850 = x82 & ~n1370 ;
  assign n4851 = x82 & n1373 ;
  assign n4852 = ( ~n1467 & n4850 ) | ( ~n1467 & n4851 ) | ( n4850 & n4851 ) ;
  assign n4853 = ( n1487 & n4850 ) | ( n1487 & n4851 ) | ( n4850 & n4851 ) ;
  assign n4854 = ( ~n1358 & n4852 ) | ( ~n1358 & n4853 ) | ( n4852 & n4853 ) ;
  assign n4855 = ( n1506 & n4852 ) | ( n1506 & n4853 ) | ( n4852 & n4853 ) ;
  assign n4856 = ( n1612 & n4854 ) | ( n1612 & n4855 ) | ( n4854 & n4855 ) ;
  assign n4857 = n4849 | n4856 ;
  assign n4858 = n4842 & ~n4857 ;
  assign n4859 = n4827 | n4858 ;
  assign n4860 = x464 & n812 ;
  assign n4861 = x464 & ~n815 ;
  assign n4862 = ( n909 & n4860 ) | ( n909 & n4861 ) | ( n4860 & n4861 ) ;
  assign n4863 = ( ~n929 & n4860 ) | ( ~n929 & n4861 ) | ( n4860 & n4861 ) ;
  assign n4864 = ( n800 & n4862 ) | ( n800 & n4863 ) | ( n4862 & n4863 ) ;
  assign n4865 = ( ~n948 & n4862 ) | ( ~n948 & n4863 ) | ( n4862 & n4863 ) ;
  assign n4866 = ( ~n1061 & n4864 ) | ( ~n1061 & n4865 ) | ( n4864 & n4865 ) ;
  assign n4867 = x336 & ~n812 ;
  assign n4868 = x336 & n815 ;
  assign n4869 = ( ~n909 & n4867 ) | ( ~n909 & n4868 ) | ( n4867 & n4868 ) ;
  assign n4870 = ( n929 & n4867 ) | ( n929 & n4868 ) | ( n4867 & n4868 ) ;
  assign n4871 = ( ~n800 & n4869 ) | ( ~n800 & n4870 ) | ( n4869 & n4870 ) ;
  assign n4872 = ( n948 & n4869 ) | ( n948 & n4870 ) | ( n4869 & n4870 ) ;
  assign n4873 = ( n1061 & n4871 ) | ( n1061 & n4872 ) | ( n4871 & n4872 ) ;
  assign n4874 = n4866 | n4873 ;
  assign n4875 = x208 & n1370 ;
  assign n4876 = x208 & ~n1373 ;
  assign n4877 = ( n1467 & n4875 ) | ( n1467 & n4876 ) | ( n4875 & n4876 ) ;
  assign n4878 = ( ~n1487 & n4875 ) | ( ~n1487 & n4876 ) | ( n4875 & n4876 ) ;
  assign n4879 = ( n1358 & n4877 ) | ( n1358 & n4878 ) | ( n4877 & n4878 ) ;
  assign n4880 = ( ~n1506 & n4877 ) | ( ~n1506 & n4878 ) | ( n4877 & n4878 ) ;
  assign n4881 = ( ~n1612 & n4879 ) | ( ~n1612 & n4880 ) | ( n4879 & n4880 ) ;
  assign n4882 = x80 & ~n1370 ;
  assign n4883 = x80 & n1373 ;
  assign n4884 = ( ~n1467 & n4882 ) | ( ~n1467 & n4883 ) | ( n4882 & n4883 ) ;
  assign n4885 = ( n1487 & n4882 ) | ( n1487 & n4883 ) | ( n4882 & n4883 ) ;
  assign n4886 = ( ~n1358 & n4884 ) | ( ~n1358 & n4885 ) | ( n4884 & n4885 ) ;
  assign n4887 = ( n1506 & n4884 ) | ( n1506 & n4885 ) | ( n4884 & n4885 ) ;
  assign n4888 = ( n1612 & n4886 ) | ( n1612 & n4887 ) | ( n4886 & n4887 ) ;
  assign n4889 = n4881 | n4888 ;
  assign n4890 = n4874 & ~n4889 ;
  assign n4891 = n4859 | n4890 ;
  assign n4892 = n4796 | n4891 ;
  assign n4893 = ~n4874 & n4889 ;
  assign n4894 = ( n3427 & ~n3442 ) | ( n3427 & n4893 ) | ( ~n3442 & n4893 ) ;
  assign n4895 = ( ~n4842 & n4857 ) | ( ~n4842 & n4894 ) | ( n4857 & n4894 ) ;
  assign n4896 = ( n4811 & ~n4826 ) | ( n4811 & n4895 ) | ( ~n4826 & n4895 ) ;
  assign n4897 = ( n4796 & n4892 ) | ( n4796 & ~n4896 ) | ( n4892 & ~n4896 ) ;
  assign n4898 = ~n4715 & n4730 ;
  assign n4899 = ~n4700 & n4898 ;
  assign n4900 = n4778 & ~n4793 ;
  assign n4901 = ( n4747 & ~n4762 ) | ( n4747 & n4900 ) | ( ~n4762 & n4900 ) ;
  assign n4902 = ( ~n4732 & n4899 ) | ( ~n4732 & n4901 ) | ( n4899 & n4901 ) ;
  assign n4903 = n4897 & ~n4902 ;
  assign n4904 = ~n4550 & n4565 ;
  assign n4905 = n4580 & ~n4595 ;
  assign n4906 = n4904 | n4905 ;
  assign n4907 = ~n4610 & n4625 ;
  assign n4908 = ~n4640 & n4655 ;
  assign n4909 = n4907 | n4908 ;
  assign n4910 = n4906 | n4909 ;
  assign n4911 = x219 & n1370 ;
  assign n4912 = x219 & ~n1373 ;
  assign n4913 = ( n1467 & n4911 ) | ( n1467 & n4912 ) | ( n4911 & n4912 ) ;
  assign n4914 = ( ~n1487 & n4911 ) | ( ~n1487 & n4912 ) | ( n4911 & n4912 ) ;
  assign n4915 = ( n1358 & n4913 ) | ( n1358 & n4914 ) | ( n4913 & n4914 ) ;
  assign n4916 = ( ~n1506 & n4913 ) | ( ~n1506 & n4914 ) | ( n4913 & n4914 ) ;
  assign n4917 = ( ~n1612 & n4915 ) | ( ~n1612 & n4916 ) | ( n4915 & n4916 ) ;
  assign n4918 = x91 & ~n1370 ;
  assign n4919 = x91 & n1373 ;
  assign n4920 = ( ~n1467 & n4918 ) | ( ~n1467 & n4919 ) | ( n4918 & n4919 ) ;
  assign n4921 = ( n1487 & n4918 ) | ( n1487 & n4919 ) | ( n4918 & n4919 ) ;
  assign n4922 = ( ~n1358 & n4920 ) | ( ~n1358 & n4921 ) | ( n4920 & n4921 ) ;
  assign n4923 = ( n1506 & n4920 ) | ( n1506 & n4921 ) | ( n4920 & n4921 ) ;
  assign n4924 = ( n1612 & n4922 ) | ( n1612 & n4923 ) | ( n4922 & n4923 ) ;
  assign n4925 = n4917 | n4924 ;
  assign n4926 = x475 & n812 ;
  assign n4927 = x475 & ~n815 ;
  assign n4928 = ( n909 & n4926 ) | ( n909 & n4927 ) | ( n4926 & n4927 ) ;
  assign n4929 = ( ~n929 & n4926 ) | ( ~n929 & n4927 ) | ( n4926 & n4927 ) ;
  assign n4930 = ( n800 & n4928 ) | ( n800 & n4929 ) | ( n4928 & n4929 ) ;
  assign n4931 = ( ~n948 & n4928 ) | ( ~n948 & n4929 ) | ( n4928 & n4929 ) ;
  assign n4932 = ( ~n1061 & n4930 ) | ( ~n1061 & n4931 ) | ( n4930 & n4931 ) ;
  assign n4933 = x347 & ~n812 ;
  assign n4934 = x347 & n815 ;
  assign n4935 = ( ~n909 & n4933 ) | ( ~n909 & n4934 ) | ( n4933 & n4934 ) ;
  assign n4936 = ( n929 & n4933 ) | ( n929 & n4934 ) | ( n4933 & n4934 ) ;
  assign n4937 = ( ~n800 & n4935 ) | ( ~n800 & n4936 ) | ( n4935 & n4936 ) ;
  assign n4938 = ( n948 & n4935 ) | ( n948 & n4936 ) | ( n4935 & n4936 ) ;
  assign n4939 = ( n1061 & n4937 ) | ( n1061 & n4938 ) | ( n4937 & n4938 ) ;
  assign n4940 = n4932 | n4939 ;
  assign n4941 = x474 & n812 ;
  assign n4942 = x474 & ~n815 ;
  assign n4943 = ( n909 & n4941 ) | ( n909 & n4942 ) | ( n4941 & n4942 ) ;
  assign n4944 = ( ~n929 & n4941 ) | ( ~n929 & n4942 ) | ( n4941 & n4942 ) ;
  assign n4945 = ( n800 & n4943 ) | ( n800 & n4944 ) | ( n4943 & n4944 ) ;
  assign n4946 = ( ~n948 & n4943 ) | ( ~n948 & n4944 ) | ( n4943 & n4944 ) ;
  assign n4947 = ( ~n1061 & n4945 ) | ( ~n1061 & n4946 ) | ( n4945 & n4946 ) ;
  assign n4948 = x346 & ~n812 ;
  assign n4949 = x346 & n815 ;
  assign n4950 = ( ~n909 & n4948 ) | ( ~n909 & n4949 ) | ( n4948 & n4949 ) ;
  assign n4951 = ( n929 & n4948 ) | ( n929 & n4949 ) | ( n4948 & n4949 ) ;
  assign n4952 = ( ~n800 & n4950 ) | ( ~n800 & n4951 ) | ( n4950 & n4951 ) ;
  assign n4953 = ( n948 & n4950 ) | ( n948 & n4951 ) | ( n4950 & n4951 ) ;
  assign n4954 = ( n1061 & n4952 ) | ( n1061 & n4953 ) | ( n4952 & n4953 ) ;
  assign n4955 = n4947 | n4954 ;
  assign n4956 = x218 & n1370 ;
  assign n4957 = x218 & ~n1373 ;
  assign n4958 = ( n1467 & n4956 ) | ( n1467 & n4957 ) | ( n4956 & n4957 ) ;
  assign n4959 = ( ~n1487 & n4956 ) | ( ~n1487 & n4957 ) | ( n4956 & n4957 ) ;
  assign n4960 = ( n1358 & n4958 ) | ( n1358 & n4959 ) | ( n4958 & n4959 ) ;
  assign n4961 = ( ~n1506 & n4958 ) | ( ~n1506 & n4959 ) | ( n4958 & n4959 ) ;
  assign n4962 = ( ~n1612 & n4960 ) | ( ~n1612 & n4961 ) | ( n4960 & n4961 ) ;
  assign n4963 = x90 & ~n1370 ;
  assign n4964 = x90 & n1373 ;
  assign n4965 = ( ~n1467 & n4963 ) | ( ~n1467 & n4964 ) | ( n4963 & n4964 ) ;
  assign n4966 = ( n1487 & n4963 ) | ( n1487 & n4964 ) | ( n4963 & n4964 ) ;
  assign n4967 = ( ~n1358 & n4965 ) | ( ~n1358 & n4966 ) | ( n4965 & n4966 ) ;
  assign n4968 = ( n1506 & n4965 ) | ( n1506 & n4966 ) | ( n4965 & n4966 ) ;
  assign n4969 = ( n1612 & n4967 ) | ( n1612 & n4968 ) | ( n4967 & n4968 ) ;
  assign n4970 = n4962 | n4969 ;
  assign n4971 = x217 & n1370 ;
  assign n4972 = x217 & ~n1373 ;
  assign n4973 = ( n1467 & n4971 ) | ( n1467 & n4972 ) | ( n4971 & n4972 ) ;
  assign n4974 = ( ~n1487 & n4971 ) | ( ~n1487 & n4972 ) | ( n4971 & n4972 ) ;
  assign n4975 = ( n1358 & n4973 ) | ( n1358 & n4974 ) | ( n4973 & n4974 ) ;
  assign n4976 = ( ~n1506 & n4973 ) | ( ~n1506 & n4974 ) | ( n4973 & n4974 ) ;
  assign n4977 = ( ~n1612 & n4975 ) | ( ~n1612 & n4976 ) | ( n4975 & n4976 ) ;
  assign n4978 = x89 & ~n1370 ;
  assign n4979 = x89 & n1373 ;
  assign n4980 = ( ~n1467 & n4978 ) | ( ~n1467 & n4979 ) | ( n4978 & n4979 ) ;
  assign n4981 = ( n1487 & n4978 ) | ( n1487 & n4979 ) | ( n4978 & n4979 ) ;
  assign n4982 = ( ~n1358 & n4980 ) | ( ~n1358 & n4981 ) | ( n4980 & n4981 ) ;
  assign n4983 = ( n1506 & n4980 ) | ( n1506 & n4981 ) | ( n4980 & n4981 ) ;
  assign n4984 = ( n1612 & n4982 ) | ( n1612 & n4983 ) | ( n4982 & n4983 ) ;
  assign n4985 = n4977 | n4984 ;
  assign n4986 = x473 & n812 ;
  assign n4987 = x473 & ~n815 ;
  assign n4988 = ( n909 & n4986 ) | ( n909 & n4987 ) | ( n4986 & n4987 ) ;
  assign n4989 = ( ~n929 & n4986 ) | ( ~n929 & n4987 ) | ( n4986 & n4987 ) ;
  assign n4990 = ( n800 & n4988 ) | ( n800 & n4989 ) | ( n4988 & n4989 ) ;
  assign n4991 = ( ~n948 & n4988 ) | ( ~n948 & n4989 ) | ( n4988 & n4989 ) ;
  assign n4992 = ( ~n1061 & n4990 ) | ( ~n1061 & n4991 ) | ( n4990 & n4991 ) ;
  assign n4993 = x345 & ~n812 ;
  assign n4994 = x345 & n815 ;
  assign n4995 = ( ~n909 & n4993 ) | ( ~n909 & n4994 ) | ( n4993 & n4994 ) ;
  assign n4996 = ( n929 & n4993 ) | ( n929 & n4994 ) | ( n4993 & n4994 ) ;
  assign n4997 = ( ~n800 & n4995 ) | ( ~n800 & n4996 ) | ( n4995 & n4996 ) ;
  assign n4998 = ( n948 & n4995 ) | ( n948 & n4996 ) | ( n4995 & n4996 ) ;
  assign n4999 = ( n1061 & n4997 ) | ( n1061 & n4998 ) | ( n4997 & n4998 ) ;
  assign n5000 = n4992 | n4999 ;
  assign n5001 = x472 & n812 ;
  assign n5002 = x472 & ~n815 ;
  assign n5003 = ( n909 & n5001 ) | ( n909 & n5002 ) | ( n5001 & n5002 ) ;
  assign n5004 = ( ~n929 & n5001 ) | ( ~n929 & n5002 ) | ( n5001 & n5002 ) ;
  assign n5005 = ( n800 & n5003 ) | ( n800 & n5004 ) | ( n5003 & n5004 ) ;
  assign n5006 = ( ~n948 & n5003 ) | ( ~n948 & n5004 ) | ( n5003 & n5004 ) ;
  assign n5007 = ( ~n1061 & n5005 ) | ( ~n1061 & n5006 ) | ( n5005 & n5006 ) ;
  assign n5008 = x344 & ~n812 ;
  assign n5009 = x344 & n815 ;
  assign n5010 = ( ~n909 & n5008 ) | ( ~n909 & n5009 ) | ( n5008 & n5009 ) ;
  assign n5011 = ( n929 & n5008 ) | ( n929 & n5009 ) | ( n5008 & n5009 ) ;
  assign n5012 = ( ~n800 & n5010 ) | ( ~n800 & n5011 ) | ( n5010 & n5011 ) ;
  assign n5013 = ( n948 & n5010 ) | ( n948 & n5011 ) | ( n5010 & n5011 ) ;
  assign n5014 = ( n1061 & n5012 ) | ( n1061 & n5013 ) | ( n5012 & n5013 ) ;
  assign n5015 = n5007 | n5014 ;
  assign n5016 = x216 & n1370 ;
  assign n5017 = x216 & ~n1373 ;
  assign n5018 = ( n1467 & n5016 ) | ( n1467 & n5017 ) | ( n5016 & n5017 ) ;
  assign n5019 = ( ~n1487 & n5016 ) | ( ~n1487 & n5017 ) | ( n5016 & n5017 ) ;
  assign n5020 = ( n1358 & n5018 ) | ( n1358 & n5019 ) | ( n5018 & n5019 ) ;
  assign n5021 = ( ~n1506 & n5018 ) | ( ~n1506 & n5019 ) | ( n5018 & n5019 ) ;
  assign n5022 = ( ~n1612 & n5020 ) | ( ~n1612 & n5021 ) | ( n5020 & n5021 ) ;
  assign n5023 = x88 & ~n1370 ;
  assign n5024 = x88 & n1373 ;
  assign n5025 = ( ~n1467 & n5023 ) | ( ~n1467 & n5024 ) | ( n5023 & n5024 ) ;
  assign n5026 = ( n1487 & n5023 ) | ( n1487 & n5024 ) | ( n5023 & n5024 ) ;
  assign n5027 = ( ~n1358 & n5025 ) | ( ~n1358 & n5026 ) | ( n5025 & n5026 ) ;
  assign n5028 = ( n1506 & n5025 ) | ( n1506 & n5026 ) | ( n5025 & n5026 ) ;
  assign n5029 = ( n1612 & n5027 ) | ( n1612 & n5028 ) | ( n5027 & n5028 ) ;
  assign n5030 = n5022 | n5029 ;
  assign n5031 = ~n5015 & n5030 ;
  assign n5032 = ( n4985 & ~n5000 ) | ( n4985 & n5031 ) | ( ~n5000 & n5031 ) ;
  assign n5033 = ( ~n4955 & n4970 ) | ( ~n4955 & n5032 ) | ( n4970 & n5032 ) ;
  assign n5034 = ( n4925 & ~n4940 ) | ( n4925 & n5033 ) | ( ~n4940 & n5033 ) ;
  assign n5035 = ~n4925 & n4940 ;
  assign n5036 = n4955 & ~n4970 ;
  assign n5037 = n5035 | n5036 ;
  assign n5038 = ~n4985 & n5000 ;
  assign n5039 = n5015 & ~n5030 ;
  assign n5040 = n5038 | n5039 ;
  assign n5041 = n5037 | n5040 ;
  assign n5042 = n4910 | n5041 ;
  assign n5043 = ( n4910 & ~n5034 ) | ( n4910 & n5042 ) | ( ~n5034 & n5042 ) ;
  assign n5044 = n4684 & ~n4699 ;
  assign n5045 = ~n4910 & n5034 ;
  assign n5046 = ( ~n5043 & n5044 ) | ( ~n5043 & n5045 ) | ( n5044 & n5045 ) ;
  assign n5047 = ( n4903 & n5043 ) | ( n4903 & ~n5046 ) | ( n5043 & ~n5046 ) ;
  assign n5048 = ( ~n4668 & n4669 ) | ( ~n4668 & n5047 ) | ( n4669 & n5047 ) ;
  assign n5049 = ( n4273 & ~n4305 ) | ( n4273 & n5048 ) | ( ~n4305 & n5048 ) ;
  assign n5050 = n4796 & ~n4899 ;
  assign n5051 = ( n4896 & n4899 ) | ( n4896 & ~n5050 ) | ( n4899 & ~n5050 ) ;
  assign n5052 = n4732 & ~n5044 ;
  assign n5053 = ( n4901 & n5044 ) | ( n4901 & ~n5052 ) | ( n5044 & ~n5052 ) ;
  assign n5054 = n5051 | n5053 ;
  assign n5055 = ( n4535 & ~n4660 ) | ( n4535 & n5043 ) | ( ~n4660 & n5043 ) ;
  assign n5056 = ( ~n4535 & n4660 ) | ( ~n4535 & n5045 ) | ( n4660 & n5045 ) ;
  assign n5057 = ( n5054 & ~n5055 ) | ( n5054 & n5056 ) | ( ~n5055 & n5056 ) ;
  assign n5058 = ( n4273 & ~n4305 ) | ( n4273 & n4667 ) | ( ~n4305 & n4667 ) ;
  assign n5059 = ( ~n4273 & n4305 ) | ( ~n4273 & n4534 ) | ( n4305 & n4534 ) ;
  assign n5060 = ( n5057 & ~n5058 ) | ( n5057 & n5059 ) | ( ~n5058 & n5059 ) ;
  assign n5061 = ( n4266 & ~n5049 ) | ( n4266 & n5060 ) | ( ~n5049 & n5060 ) ;
  assign n5062 = n3399 & ~n3408 ;
  assign n5063 = n3276 | n3374 ;
  assign n5064 = ( n3341 & ~n3377 ) | ( n3341 & n5063 ) | ( ~n3377 & n5063 ) ;
  assign n5065 = n3375 & ~n3380 ;
  assign n5066 = ( ~n3213 & n3245 ) | ( ~n3213 & n5065 ) | ( n3245 & n5065 ) ;
  assign n5067 = ( n3381 & n5064 ) | ( n3381 & ~n5066 ) | ( n5064 & ~n5066 ) ;
  assign n5068 = ( n3181 & ~n3212 ) | ( n3181 & n5067 ) | ( ~n3212 & n5067 ) ;
  assign n5069 = n3181 | n5068 ;
  assign n5070 = ( n3408 & ~n5062 ) | ( n3408 & n5069 ) | ( ~n5062 & n5069 ) ;
  assign n5071 = n2920 | n2926 ;
  assign n5072 = ( ~n2695 & n2696 ) | ( ~n2695 & n5071 ) | ( n2696 & n5071 ) ;
  assign n5073 = n2661 | n5072 ;
  assign n5074 = ( n2698 & n5070 ) | ( n2698 & ~n5073 ) | ( n5070 & ~n5073 ) ;
  assign n5075 = ( n4257 & ~n4265 ) | ( n4257 & n5074 ) | ( ~n4265 & n5074 ) ;
  assign n5076 = ( n5049 & ~n5060 ) | ( n5049 & n5075 ) | ( ~n5060 & n5075 ) ;
  assign n5077 = x149 & n1370 ;
  assign n5078 = x149 & ~n1373 ;
  assign n5079 = ( n1467 & n5077 ) | ( n1467 & n5078 ) | ( n5077 & n5078 ) ;
  assign n5080 = ( ~n1487 & n5077 ) | ( ~n1487 & n5078 ) | ( n5077 & n5078 ) ;
  assign n5081 = ( n1358 & n5079 ) | ( n1358 & n5080 ) | ( n5079 & n5080 ) ;
  assign n5082 = ( ~n1506 & n5079 ) | ( ~n1506 & n5080 ) | ( n5079 & n5080 ) ;
  assign n5083 = ( ~n1612 & n5081 ) | ( ~n1612 & n5082 ) | ( n5081 & n5082 ) ;
  assign n5084 = x21 & ~n1370 ;
  assign n5085 = x21 & n1373 ;
  assign n5086 = ( ~n1467 & n5084 ) | ( ~n1467 & n5085 ) | ( n5084 & n5085 ) ;
  assign n5087 = ( n1487 & n5084 ) | ( n1487 & n5085 ) | ( n5084 & n5085 ) ;
  assign n5088 = ( ~n1358 & n5086 ) | ( ~n1358 & n5087 ) | ( n5086 & n5087 ) ;
  assign n5089 = ( n1506 & n5086 ) | ( n1506 & n5087 ) | ( n5086 & n5087 ) ;
  assign n5090 = ( n1612 & n5088 ) | ( n1612 & n5089 ) | ( n5088 & n5089 ) ;
  assign n5091 = n5083 | n5090 ;
  assign n5092 = x405 & n812 ;
  assign n5093 = x405 & ~n815 ;
  assign n5094 = ( n909 & n5092 ) | ( n909 & n5093 ) | ( n5092 & n5093 ) ;
  assign n5095 = ( ~n929 & n5092 ) | ( ~n929 & n5093 ) | ( n5092 & n5093 ) ;
  assign n5096 = ( n800 & n5094 ) | ( n800 & n5095 ) | ( n5094 & n5095 ) ;
  assign n5097 = ( ~n948 & n5094 ) | ( ~n948 & n5095 ) | ( n5094 & n5095 ) ;
  assign n5098 = ( ~n1061 & n5096 ) | ( ~n1061 & n5097 ) | ( n5096 & n5097 ) ;
  assign n5099 = x277 & ~n812 ;
  assign n5100 = x277 & n815 ;
  assign n5101 = ( ~n909 & n5099 ) | ( ~n909 & n5100 ) | ( n5099 & n5100 ) ;
  assign n5102 = ( n929 & n5099 ) | ( n929 & n5100 ) | ( n5099 & n5100 ) ;
  assign n5103 = ( ~n800 & n5101 ) | ( ~n800 & n5102 ) | ( n5101 & n5102 ) ;
  assign n5104 = ( n948 & n5101 ) | ( n948 & n5102 ) | ( n5101 & n5102 ) ;
  assign n5105 = ( n1061 & n5103 ) | ( n1061 & n5104 ) | ( n5103 & n5104 ) ;
  assign n5106 = n5098 | n5105 ;
  assign n5107 = ~n5091 & n5106 ;
  assign n5108 = x148 & n1370 ;
  assign n5109 = x148 & ~n1373 ;
  assign n5110 = ( n1467 & n5108 ) | ( n1467 & n5109 ) | ( n5108 & n5109 ) ;
  assign n5111 = ( ~n1487 & n5108 ) | ( ~n1487 & n5109 ) | ( n5108 & n5109 ) ;
  assign n5112 = ( n1358 & n5110 ) | ( n1358 & n5111 ) | ( n5110 & n5111 ) ;
  assign n5113 = ( ~n1506 & n5110 ) | ( ~n1506 & n5111 ) | ( n5110 & n5111 ) ;
  assign n5114 = ( ~n1612 & n5112 ) | ( ~n1612 & n5113 ) | ( n5112 & n5113 ) ;
  assign n5115 = x20 & ~n1370 ;
  assign n5116 = x20 & n1373 ;
  assign n5117 = ( ~n1467 & n5115 ) | ( ~n1467 & n5116 ) | ( n5115 & n5116 ) ;
  assign n5118 = ( n1487 & n5115 ) | ( n1487 & n5116 ) | ( n5115 & n5116 ) ;
  assign n5119 = ( ~n1358 & n5117 ) | ( ~n1358 & n5118 ) | ( n5117 & n5118 ) ;
  assign n5120 = ( n1506 & n5117 ) | ( n1506 & n5118 ) | ( n5117 & n5118 ) ;
  assign n5121 = ( n1612 & n5119 ) | ( n1612 & n5120 ) | ( n5119 & n5120 ) ;
  assign n5122 = n5114 | n5121 ;
  assign n5123 = x404 & n812 ;
  assign n5124 = x404 & ~n815 ;
  assign n5125 = ( n909 & n5123 ) | ( n909 & n5124 ) | ( n5123 & n5124 ) ;
  assign n5126 = ( ~n929 & n5123 ) | ( ~n929 & n5124 ) | ( n5123 & n5124 ) ;
  assign n5127 = ( n800 & n5125 ) | ( n800 & n5126 ) | ( n5125 & n5126 ) ;
  assign n5128 = ( ~n948 & n5125 ) | ( ~n948 & n5126 ) | ( n5125 & n5126 ) ;
  assign n5129 = ( ~n1061 & n5127 ) | ( ~n1061 & n5128 ) | ( n5127 & n5128 ) ;
  assign n5130 = x276 & ~n812 ;
  assign n5131 = x276 & n815 ;
  assign n5132 = ( ~n909 & n5130 ) | ( ~n909 & n5131 ) | ( n5130 & n5131 ) ;
  assign n5133 = ( n929 & n5130 ) | ( n929 & n5131 ) | ( n5130 & n5131 ) ;
  assign n5134 = ( ~n800 & n5132 ) | ( ~n800 & n5133 ) | ( n5132 & n5133 ) ;
  assign n5135 = ( n948 & n5132 ) | ( n948 & n5133 ) | ( n5132 & n5133 ) ;
  assign n5136 = ( n1061 & n5134 ) | ( n1061 & n5135 ) | ( n5134 & n5135 ) ;
  assign n5137 = n5129 | n5136 ;
  assign n5138 = n5122 & ~n5137 ;
  assign n5139 = ~n5107 & n5138 ;
  assign n5140 = x147 & n1370 ;
  assign n5141 = x147 & ~n1373 ;
  assign n5142 = ( n1467 & n5140 ) | ( n1467 & n5141 ) | ( n5140 & n5141 ) ;
  assign n5143 = ( ~n1487 & n5140 ) | ( ~n1487 & n5141 ) | ( n5140 & n5141 ) ;
  assign n5144 = ( n1358 & n5142 ) | ( n1358 & n5143 ) | ( n5142 & n5143 ) ;
  assign n5145 = ( ~n1506 & n5142 ) | ( ~n1506 & n5143 ) | ( n5142 & n5143 ) ;
  assign n5146 = ( ~n1612 & n5144 ) | ( ~n1612 & n5145 ) | ( n5144 & n5145 ) ;
  assign n5147 = x19 & ~n1370 ;
  assign n5148 = x19 & n1373 ;
  assign n5149 = ( ~n1467 & n5147 ) | ( ~n1467 & n5148 ) | ( n5147 & n5148 ) ;
  assign n5150 = ( n1487 & n5147 ) | ( n1487 & n5148 ) | ( n5147 & n5148 ) ;
  assign n5151 = ( ~n1358 & n5149 ) | ( ~n1358 & n5150 ) | ( n5149 & n5150 ) ;
  assign n5152 = ( n1506 & n5149 ) | ( n1506 & n5150 ) | ( n5149 & n5150 ) ;
  assign n5153 = ( n1612 & n5151 ) | ( n1612 & n5152 ) | ( n5151 & n5152 ) ;
  assign n5154 = n5146 | n5153 ;
  assign n5155 = x403 & n812 ;
  assign n5156 = x403 & ~n815 ;
  assign n5157 = ( n909 & n5155 ) | ( n909 & n5156 ) | ( n5155 & n5156 ) ;
  assign n5158 = ( ~n929 & n5155 ) | ( ~n929 & n5156 ) | ( n5155 & n5156 ) ;
  assign n5159 = ( n800 & n5157 ) | ( n800 & n5158 ) | ( n5157 & n5158 ) ;
  assign n5160 = ( ~n948 & n5157 ) | ( ~n948 & n5158 ) | ( n5157 & n5158 ) ;
  assign n5161 = ( ~n1061 & n5159 ) | ( ~n1061 & n5160 ) | ( n5159 & n5160 ) ;
  assign n5162 = x275 & ~n812 ;
  assign n5163 = x275 & n815 ;
  assign n5164 = ( ~n909 & n5162 ) | ( ~n909 & n5163 ) | ( n5162 & n5163 ) ;
  assign n5165 = ( n929 & n5162 ) | ( n929 & n5163 ) | ( n5162 & n5163 ) ;
  assign n5166 = ( ~n800 & n5164 ) | ( ~n800 & n5165 ) | ( n5164 & n5165 ) ;
  assign n5167 = ( n948 & n5164 ) | ( n948 & n5165 ) | ( n5164 & n5165 ) ;
  assign n5168 = ( n1061 & n5166 ) | ( n1061 & n5167 ) | ( n5166 & n5167 ) ;
  assign n5169 = n5161 | n5168 ;
  assign n5170 = x146 & n1370 ;
  assign n5171 = x146 & ~n1373 ;
  assign n5172 = ( n1467 & n5170 ) | ( n1467 & n5171 ) | ( n5170 & n5171 ) ;
  assign n5173 = ( ~n1487 & n5170 ) | ( ~n1487 & n5171 ) | ( n5170 & n5171 ) ;
  assign n5174 = ( n1358 & n5172 ) | ( n1358 & n5173 ) | ( n5172 & n5173 ) ;
  assign n5175 = ( ~n1506 & n5172 ) | ( ~n1506 & n5173 ) | ( n5172 & n5173 ) ;
  assign n5176 = ( ~n1612 & n5174 ) | ( ~n1612 & n5175 ) | ( n5174 & n5175 ) ;
  assign n5177 = x18 & ~n1370 ;
  assign n5178 = x18 & n1373 ;
  assign n5179 = ( ~n1467 & n5177 ) | ( ~n1467 & n5178 ) | ( n5177 & n5178 ) ;
  assign n5180 = ( n1487 & n5177 ) | ( n1487 & n5178 ) | ( n5177 & n5178 ) ;
  assign n5181 = ( ~n1358 & n5179 ) | ( ~n1358 & n5180 ) | ( n5179 & n5180 ) ;
  assign n5182 = ( n1506 & n5179 ) | ( n1506 & n5180 ) | ( n5179 & n5180 ) ;
  assign n5183 = ( n1612 & n5181 ) | ( n1612 & n5182 ) | ( n5181 & n5182 ) ;
  assign n5184 = n5176 | n5183 ;
  assign n5185 = x402 & n812 ;
  assign n5186 = x402 & ~n815 ;
  assign n5187 = ( n909 & n5185 ) | ( n909 & n5186 ) | ( n5185 & n5186 ) ;
  assign n5188 = ( ~n929 & n5185 ) | ( ~n929 & n5186 ) | ( n5185 & n5186 ) ;
  assign n5189 = ( n800 & n5187 ) | ( n800 & n5188 ) | ( n5187 & n5188 ) ;
  assign n5190 = ( ~n948 & n5187 ) | ( ~n948 & n5188 ) | ( n5187 & n5188 ) ;
  assign n5191 = ( ~n1061 & n5189 ) | ( ~n1061 & n5190 ) | ( n5189 & n5190 ) ;
  assign n5192 = x274 & ~n812 ;
  assign n5193 = x274 & n815 ;
  assign n5194 = ( ~n909 & n5192 ) | ( ~n909 & n5193 ) | ( n5192 & n5193 ) ;
  assign n5195 = ( n929 & n5192 ) | ( n929 & n5193 ) | ( n5192 & n5193 ) ;
  assign n5196 = ( ~n800 & n5194 ) | ( ~n800 & n5195 ) | ( n5194 & n5195 ) ;
  assign n5197 = ( n948 & n5194 ) | ( n948 & n5195 ) | ( n5194 & n5195 ) ;
  assign n5198 = ( n1061 & n5196 ) | ( n1061 & n5197 ) | ( n5196 & n5197 ) ;
  assign n5199 = n5191 | n5198 ;
  assign n5200 = ~n5184 & n5199 ;
  assign n5201 = ( ~n5154 & n5169 ) | ( ~n5154 & n5200 ) | ( n5169 & n5200 ) ;
  assign n5202 = ~n5122 & n5137 ;
  assign n5203 = n5107 | n5202 ;
  assign n5204 = ( ~n5139 & n5201 ) | ( ~n5139 & n5203 ) | ( n5201 & n5203 ) ;
  assign n5205 = x408 & n812 ;
  assign n5206 = x408 & ~n815 ;
  assign n5207 = ( n909 & n5205 ) | ( n909 & n5206 ) | ( n5205 & n5206 ) ;
  assign n5208 = ( ~n929 & n5205 ) | ( ~n929 & n5206 ) | ( n5205 & n5206 ) ;
  assign n5209 = ( n800 & n5207 ) | ( n800 & n5208 ) | ( n5207 & n5208 ) ;
  assign n5210 = ( ~n948 & n5207 ) | ( ~n948 & n5208 ) | ( n5207 & n5208 ) ;
  assign n5211 = ( ~n1061 & n5209 ) | ( ~n1061 & n5210 ) | ( n5209 & n5210 ) ;
  assign n5212 = x280 & ~n812 ;
  assign n5213 = x280 & n815 ;
  assign n5214 = ( ~n909 & n5212 ) | ( ~n909 & n5213 ) | ( n5212 & n5213 ) ;
  assign n5215 = ( n929 & n5212 ) | ( n929 & n5213 ) | ( n5212 & n5213 ) ;
  assign n5216 = ( ~n800 & n5214 ) | ( ~n800 & n5215 ) | ( n5214 & n5215 ) ;
  assign n5217 = ( n948 & n5214 ) | ( n948 & n5215 ) | ( n5214 & n5215 ) ;
  assign n5218 = ( n1061 & n5216 ) | ( n1061 & n5217 ) | ( n5216 & n5217 ) ;
  assign n5219 = n5211 | n5218 ;
  assign n5220 = x151 & n1370 ;
  assign n5221 = x151 & ~n1373 ;
  assign n5222 = ( n1467 & n5220 ) | ( n1467 & n5221 ) | ( n5220 & n5221 ) ;
  assign n5223 = ( ~n1487 & n5220 ) | ( ~n1487 & n5221 ) | ( n5220 & n5221 ) ;
  assign n5224 = ( n1358 & n5222 ) | ( n1358 & n5223 ) | ( n5222 & n5223 ) ;
  assign n5225 = ( ~n1506 & n5222 ) | ( ~n1506 & n5223 ) | ( n5222 & n5223 ) ;
  assign n5226 = ( ~n1612 & n5224 ) | ( ~n1612 & n5225 ) | ( n5224 & n5225 ) ;
  assign n5227 = x23 & ~n1370 ;
  assign n5228 = x23 & n1373 ;
  assign n5229 = ( ~n1467 & n5227 ) | ( ~n1467 & n5228 ) | ( n5227 & n5228 ) ;
  assign n5230 = ( n1487 & n5227 ) | ( n1487 & n5228 ) | ( n5227 & n5228 ) ;
  assign n5231 = ( ~n1358 & n5229 ) | ( ~n1358 & n5230 ) | ( n5229 & n5230 ) ;
  assign n5232 = ( n1506 & n5229 ) | ( n1506 & n5230 ) | ( n5229 & n5230 ) ;
  assign n5233 = ( n1612 & n5231 ) | ( n1612 & n5232 ) | ( n5231 & n5232 ) ;
  assign n5234 = n5226 | n5233 ;
  assign n5235 = x407 & n812 ;
  assign n5236 = x407 & ~n815 ;
  assign n5237 = ( n909 & n5235 ) | ( n909 & n5236 ) | ( n5235 & n5236 ) ;
  assign n5238 = ( ~n929 & n5235 ) | ( ~n929 & n5236 ) | ( n5235 & n5236 ) ;
  assign n5239 = ( n800 & n5237 ) | ( n800 & n5238 ) | ( n5237 & n5238 ) ;
  assign n5240 = ( ~n948 & n5237 ) | ( ~n948 & n5238 ) | ( n5237 & n5238 ) ;
  assign n5241 = ( ~n1061 & n5239 ) | ( ~n1061 & n5240 ) | ( n5239 & n5240 ) ;
  assign n5242 = x279 & ~n812 ;
  assign n5243 = x279 & n815 ;
  assign n5244 = ( ~n909 & n5242 ) | ( ~n909 & n5243 ) | ( n5242 & n5243 ) ;
  assign n5245 = ( n929 & n5242 ) | ( n929 & n5243 ) | ( n5242 & n5243 ) ;
  assign n5246 = ( ~n800 & n5244 ) | ( ~n800 & n5245 ) | ( n5244 & n5245 ) ;
  assign n5247 = ( n948 & n5244 ) | ( n948 & n5245 ) | ( n5244 & n5245 ) ;
  assign n5248 = ( n1061 & n5246 ) | ( n1061 & n5247 ) | ( n5246 & n5247 ) ;
  assign n5249 = n5241 | n5248 ;
  assign n5250 = ~n5234 & n5249 ;
  assign n5251 = x150 & n1370 ;
  assign n5252 = x150 & ~n1373 ;
  assign n5253 = ( n1467 & n5251 ) | ( n1467 & n5252 ) | ( n5251 & n5252 ) ;
  assign n5254 = ( ~n1487 & n5251 ) | ( ~n1487 & n5252 ) | ( n5251 & n5252 ) ;
  assign n5255 = ( n1358 & n5253 ) | ( n1358 & n5254 ) | ( n5253 & n5254 ) ;
  assign n5256 = ( ~n1506 & n5253 ) | ( ~n1506 & n5254 ) | ( n5253 & n5254 ) ;
  assign n5257 = ( ~n1612 & n5255 ) | ( ~n1612 & n5256 ) | ( n5255 & n5256 ) ;
  assign n5258 = x22 & ~n1370 ;
  assign n5259 = x22 & n1373 ;
  assign n5260 = ( ~n1467 & n5258 ) | ( ~n1467 & n5259 ) | ( n5258 & n5259 ) ;
  assign n5261 = ( n1487 & n5258 ) | ( n1487 & n5259 ) | ( n5258 & n5259 ) ;
  assign n5262 = ( ~n1358 & n5260 ) | ( ~n1358 & n5261 ) | ( n5260 & n5261 ) ;
  assign n5263 = ( n1506 & n5260 ) | ( n1506 & n5261 ) | ( n5260 & n5261 ) ;
  assign n5264 = ( n1612 & n5262 ) | ( n1612 & n5263 ) | ( n5262 & n5263 ) ;
  assign n5265 = n5257 | n5264 ;
  assign n5266 = x406 & n812 ;
  assign n5267 = x406 & ~n815 ;
  assign n5268 = ( n909 & n5266 ) | ( n909 & n5267 ) | ( n5266 & n5267 ) ;
  assign n5269 = ( ~n929 & n5266 ) | ( ~n929 & n5267 ) | ( n5266 & n5267 ) ;
  assign n5270 = ( n800 & n5268 ) | ( n800 & n5269 ) | ( n5268 & n5269 ) ;
  assign n5271 = ( ~n948 & n5268 ) | ( ~n948 & n5269 ) | ( n5268 & n5269 ) ;
  assign n5272 = ( ~n1061 & n5270 ) | ( ~n1061 & n5271 ) | ( n5270 & n5271 ) ;
  assign n5273 = x278 & ~n812 ;
  assign n5274 = x278 & n815 ;
  assign n5275 = ( ~n909 & n5273 ) | ( ~n909 & n5274 ) | ( n5273 & n5274 ) ;
  assign n5276 = ( n929 & n5273 ) | ( n929 & n5274 ) | ( n5273 & n5274 ) ;
  assign n5277 = ( ~n800 & n5275 ) | ( ~n800 & n5276 ) | ( n5275 & n5276 ) ;
  assign n5278 = ( n948 & n5275 ) | ( n948 & n5276 ) | ( n5275 & n5276 ) ;
  assign n5279 = ( n1061 & n5277 ) | ( n1061 & n5278 ) | ( n5277 & n5278 ) ;
  assign n5280 = n5272 | n5279 ;
  assign n5281 = ~n5265 & n5280 ;
  assign n5282 = n5091 & ~n5106 ;
  assign n5283 = ~n5281 & n5282 ;
  assign n5284 = n5265 & ~n5280 ;
  assign n5285 = ~n5250 & n5284 ;
  assign n5286 = ( ~n5250 & n5283 ) | ( ~n5250 & n5285 ) | ( n5283 & n5285 ) ;
  assign n5287 = n5234 & ~n5249 ;
  assign n5288 = x152 & n1370 ;
  assign n5289 = x152 & ~n1373 ;
  assign n5290 = ( n1467 & n5288 ) | ( n1467 & n5289 ) | ( n5288 & n5289 ) ;
  assign n5291 = ( ~n1487 & n5288 ) | ( ~n1487 & n5289 ) | ( n5288 & n5289 ) ;
  assign n5292 = ( n1358 & n5290 ) | ( n1358 & n5291 ) | ( n5290 & n5291 ) ;
  assign n5293 = ( ~n1506 & n5290 ) | ( ~n1506 & n5291 ) | ( n5290 & n5291 ) ;
  assign n5294 = ( ~n1612 & n5292 ) | ( ~n1612 & n5293 ) | ( n5292 & n5293 ) ;
  assign n5295 = x24 & ~n1370 ;
  assign n5296 = x24 & n1373 ;
  assign n5297 = ( ~n1467 & n5295 ) | ( ~n1467 & n5296 ) | ( n5295 & n5296 ) ;
  assign n5298 = ( n1487 & n5295 ) | ( n1487 & n5296 ) | ( n5295 & n5296 ) ;
  assign n5299 = ( ~n1358 & n5297 ) | ( ~n1358 & n5298 ) | ( n5297 & n5298 ) ;
  assign n5300 = ( n1506 & n5297 ) | ( n1506 & n5298 ) | ( n5297 & n5298 ) ;
  assign n5301 = ( n1612 & n5299 ) | ( n1612 & n5300 ) | ( n5299 & n5300 ) ;
  assign n5302 = n5294 | n5301 ;
  assign n5303 = ~n5219 & n5302 ;
  assign n5304 = ( ~n5219 & n5287 ) | ( ~n5219 & n5303 ) | ( n5287 & n5303 ) ;
  assign n5305 = ( ~n5219 & n5286 ) | ( ~n5219 & n5304 ) | ( n5286 & n5304 ) ;
  assign n5306 = n5250 | n5281 ;
  assign n5307 = ~n5287 & n5306 ;
  assign n5308 = ( n5219 & ~n5303 ) | ( n5219 & n5307 ) | ( ~n5303 & n5307 ) ;
  assign n5309 = ( n5204 & ~n5305 ) | ( n5204 & n5308 ) | ( ~n5305 & n5308 ) ;
  assign n5310 = ( ~n5219 & n5285 ) | ( ~n5219 & n5304 ) | ( n5285 & n5304 ) ;
  assign n5311 = n5154 & ~n5169 ;
  assign n5312 = ~n5202 & n5311 ;
  assign n5313 = n5184 & ~n5199 ;
  assign n5314 = ~n5201 & n5313 ;
  assign n5315 = ( ~n5202 & n5312 ) | ( ~n5202 & n5314 ) | ( n5312 & n5314 ) ;
  assign n5316 = ( ~n5107 & n5139 ) | ( ~n5107 & n5315 ) | ( n5139 & n5315 ) ;
  assign n5317 = n5282 | n5316 ;
  assign n5318 = ( ~n5308 & n5310 ) | ( ~n5308 & n5317 ) | ( n5310 & n5317 ) ;
  assign n5319 = x141 & n1370 ;
  assign n5320 = x141 & ~n1373 ;
  assign n5321 = ( n1467 & n5319 ) | ( n1467 & n5320 ) | ( n5319 & n5320 ) ;
  assign n5322 = ( ~n1487 & n5319 ) | ( ~n1487 & n5320 ) | ( n5319 & n5320 ) ;
  assign n5323 = ( n1358 & n5321 ) | ( n1358 & n5322 ) | ( n5321 & n5322 ) ;
  assign n5324 = ( ~n1506 & n5321 ) | ( ~n1506 & n5322 ) | ( n5321 & n5322 ) ;
  assign n5325 = ( ~n1612 & n5323 ) | ( ~n1612 & n5324 ) | ( n5323 & n5324 ) ;
  assign n5326 = x13 & ~n1370 ;
  assign n5327 = x13 & n1373 ;
  assign n5328 = ( ~n1467 & n5326 ) | ( ~n1467 & n5327 ) | ( n5326 & n5327 ) ;
  assign n5329 = ( n1487 & n5326 ) | ( n1487 & n5327 ) | ( n5326 & n5327 ) ;
  assign n5330 = ( ~n1358 & n5328 ) | ( ~n1358 & n5329 ) | ( n5328 & n5329 ) ;
  assign n5331 = ( n1506 & n5328 ) | ( n1506 & n5329 ) | ( n5328 & n5329 ) ;
  assign n5332 = ( n1612 & n5330 ) | ( n1612 & n5331 ) | ( n5330 & n5331 ) ;
  assign n5333 = n5325 | n5332 ;
  assign n5334 = x397 & n812 ;
  assign n5335 = x397 & ~n815 ;
  assign n5336 = ( n909 & n5334 ) | ( n909 & n5335 ) | ( n5334 & n5335 ) ;
  assign n5337 = ( ~n929 & n5334 ) | ( ~n929 & n5335 ) | ( n5334 & n5335 ) ;
  assign n5338 = ( n800 & n5336 ) | ( n800 & n5337 ) | ( n5336 & n5337 ) ;
  assign n5339 = ( ~n948 & n5336 ) | ( ~n948 & n5337 ) | ( n5336 & n5337 ) ;
  assign n5340 = ( ~n1061 & n5338 ) | ( ~n1061 & n5339 ) | ( n5338 & n5339 ) ;
  assign n5341 = x269 & ~n812 ;
  assign n5342 = x269 & n815 ;
  assign n5343 = ( ~n909 & n5341 ) | ( ~n909 & n5342 ) | ( n5341 & n5342 ) ;
  assign n5344 = ( n929 & n5341 ) | ( n929 & n5342 ) | ( n5341 & n5342 ) ;
  assign n5345 = ( ~n800 & n5343 ) | ( ~n800 & n5344 ) | ( n5343 & n5344 ) ;
  assign n5346 = ( n948 & n5343 ) | ( n948 & n5344 ) | ( n5343 & n5344 ) ;
  assign n5347 = ( n1061 & n5345 ) | ( n1061 & n5346 ) | ( n5345 & n5346 ) ;
  assign n5348 = n5340 | n5347 ;
  assign n5349 = ~n5333 & n5348 ;
  assign n5350 = x140 & n1370 ;
  assign n5351 = x140 & ~n1373 ;
  assign n5352 = ( n1467 & n5350 ) | ( n1467 & n5351 ) | ( n5350 & n5351 ) ;
  assign n5353 = ( ~n1487 & n5350 ) | ( ~n1487 & n5351 ) | ( n5350 & n5351 ) ;
  assign n5354 = ( n1358 & n5352 ) | ( n1358 & n5353 ) | ( n5352 & n5353 ) ;
  assign n5355 = ( ~n1506 & n5352 ) | ( ~n1506 & n5353 ) | ( n5352 & n5353 ) ;
  assign n5356 = ( ~n1612 & n5354 ) | ( ~n1612 & n5355 ) | ( n5354 & n5355 ) ;
  assign n5357 = x12 & ~n1370 ;
  assign n5358 = x12 & n1373 ;
  assign n5359 = ( ~n1467 & n5357 ) | ( ~n1467 & n5358 ) | ( n5357 & n5358 ) ;
  assign n5360 = ( n1487 & n5357 ) | ( n1487 & n5358 ) | ( n5357 & n5358 ) ;
  assign n5361 = ( ~n1358 & n5359 ) | ( ~n1358 & n5360 ) | ( n5359 & n5360 ) ;
  assign n5362 = ( n1506 & n5359 ) | ( n1506 & n5360 ) | ( n5359 & n5360 ) ;
  assign n5363 = ( n1612 & n5361 ) | ( n1612 & n5362 ) | ( n5361 & n5362 ) ;
  assign n5364 = n5356 | n5363 ;
  assign n5365 = x396 & n812 ;
  assign n5366 = x396 & ~n815 ;
  assign n5367 = ( n909 & n5365 ) | ( n909 & n5366 ) | ( n5365 & n5366 ) ;
  assign n5368 = ( ~n929 & n5365 ) | ( ~n929 & n5366 ) | ( n5365 & n5366 ) ;
  assign n5369 = ( n800 & n5367 ) | ( n800 & n5368 ) | ( n5367 & n5368 ) ;
  assign n5370 = ( ~n948 & n5367 ) | ( ~n948 & n5368 ) | ( n5367 & n5368 ) ;
  assign n5371 = ( ~n1061 & n5369 ) | ( ~n1061 & n5370 ) | ( n5369 & n5370 ) ;
  assign n5372 = x268 & ~n812 ;
  assign n5373 = x268 & n815 ;
  assign n5374 = ( ~n909 & n5372 ) | ( ~n909 & n5373 ) | ( n5372 & n5373 ) ;
  assign n5375 = ( n929 & n5372 ) | ( n929 & n5373 ) | ( n5372 & n5373 ) ;
  assign n5376 = ( ~n800 & n5374 ) | ( ~n800 & n5375 ) | ( n5374 & n5375 ) ;
  assign n5377 = ( n948 & n5374 ) | ( n948 & n5375 ) | ( n5374 & n5375 ) ;
  assign n5378 = ( n1061 & n5376 ) | ( n1061 & n5377 ) | ( n5376 & n5377 ) ;
  assign n5379 = n5371 | n5378 ;
  assign n5380 = n5364 & ~n5379 ;
  assign n5381 = ~n5349 & n5380 ;
  assign n5382 = x139 & n1370 ;
  assign n5383 = x139 & ~n1373 ;
  assign n5384 = ( n1467 & n5382 ) | ( n1467 & n5383 ) | ( n5382 & n5383 ) ;
  assign n5385 = ( ~n1487 & n5382 ) | ( ~n1487 & n5383 ) | ( n5382 & n5383 ) ;
  assign n5386 = ( n1358 & n5384 ) | ( n1358 & n5385 ) | ( n5384 & n5385 ) ;
  assign n5387 = ( ~n1506 & n5384 ) | ( ~n1506 & n5385 ) | ( n5384 & n5385 ) ;
  assign n5388 = ( ~n1612 & n5386 ) | ( ~n1612 & n5387 ) | ( n5386 & n5387 ) ;
  assign n5389 = x11 & ~n1370 ;
  assign n5390 = x11 & n1373 ;
  assign n5391 = ( ~n1467 & n5389 ) | ( ~n1467 & n5390 ) | ( n5389 & n5390 ) ;
  assign n5392 = ( n1487 & n5389 ) | ( n1487 & n5390 ) | ( n5389 & n5390 ) ;
  assign n5393 = ( ~n1358 & n5391 ) | ( ~n1358 & n5392 ) | ( n5391 & n5392 ) ;
  assign n5394 = ( n1506 & n5391 ) | ( n1506 & n5392 ) | ( n5391 & n5392 ) ;
  assign n5395 = ( n1612 & n5393 ) | ( n1612 & n5394 ) | ( n5393 & n5394 ) ;
  assign n5396 = n5388 | n5395 ;
  assign n5397 = x395 & n812 ;
  assign n5398 = x395 & ~n815 ;
  assign n5399 = ( n909 & n5397 ) | ( n909 & n5398 ) | ( n5397 & n5398 ) ;
  assign n5400 = ( ~n929 & n5397 ) | ( ~n929 & n5398 ) | ( n5397 & n5398 ) ;
  assign n5401 = ( n800 & n5399 ) | ( n800 & n5400 ) | ( n5399 & n5400 ) ;
  assign n5402 = ( ~n948 & n5399 ) | ( ~n948 & n5400 ) | ( n5399 & n5400 ) ;
  assign n5403 = ( ~n1061 & n5401 ) | ( ~n1061 & n5402 ) | ( n5401 & n5402 ) ;
  assign n5404 = x267 & ~n812 ;
  assign n5405 = x267 & n815 ;
  assign n5406 = ( ~n909 & n5404 ) | ( ~n909 & n5405 ) | ( n5404 & n5405 ) ;
  assign n5407 = ( n929 & n5404 ) | ( n929 & n5405 ) | ( n5404 & n5405 ) ;
  assign n5408 = ( ~n800 & n5406 ) | ( ~n800 & n5407 ) | ( n5406 & n5407 ) ;
  assign n5409 = ( n948 & n5406 ) | ( n948 & n5407 ) | ( n5406 & n5407 ) ;
  assign n5410 = ( n1061 & n5408 ) | ( n1061 & n5409 ) | ( n5408 & n5409 ) ;
  assign n5411 = n5403 | n5410 ;
  assign n5412 = x138 & n1370 ;
  assign n5413 = x138 & ~n1373 ;
  assign n5414 = ( n1467 & n5412 ) | ( n1467 & n5413 ) | ( n5412 & n5413 ) ;
  assign n5415 = ( ~n1487 & n5412 ) | ( ~n1487 & n5413 ) | ( n5412 & n5413 ) ;
  assign n5416 = ( n1358 & n5414 ) | ( n1358 & n5415 ) | ( n5414 & n5415 ) ;
  assign n5417 = ( ~n1506 & n5414 ) | ( ~n1506 & n5415 ) | ( n5414 & n5415 ) ;
  assign n5418 = ( ~n1612 & n5416 ) | ( ~n1612 & n5417 ) | ( n5416 & n5417 ) ;
  assign n5419 = x10 & ~n1370 ;
  assign n5420 = x10 & n1373 ;
  assign n5421 = ( ~n1467 & n5419 ) | ( ~n1467 & n5420 ) | ( n5419 & n5420 ) ;
  assign n5422 = ( n1487 & n5419 ) | ( n1487 & n5420 ) | ( n5419 & n5420 ) ;
  assign n5423 = ( ~n1358 & n5421 ) | ( ~n1358 & n5422 ) | ( n5421 & n5422 ) ;
  assign n5424 = ( n1506 & n5421 ) | ( n1506 & n5422 ) | ( n5421 & n5422 ) ;
  assign n5425 = ( n1612 & n5423 ) | ( n1612 & n5424 ) | ( n5423 & n5424 ) ;
  assign n5426 = n5418 | n5425 ;
  assign n5427 = x394 & n812 ;
  assign n5428 = x394 & ~n815 ;
  assign n5429 = ( n909 & n5427 ) | ( n909 & n5428 ) | ( n5427 & n5428 ) ;
  assign n5430 = ( ~n929 & n5427 ) | ( ~n929 & n5428 ) | ( n5427 & n5428 ) ;
  assign n5431 = ( n800 & n5429 ) | ( n800 & n5430 ) | ( n5429 & n5430 ) ;
  assign n5432 = ( ~n948 & n5429 ) | ( ~n948 & n5430 ) | ( n5429 & n5430 ) ;
  assign n5433 = ( ~n1061 & n5431 ) | ( ~n1061 & n5432 ) | ( n5431 & n5432 ) ;
  assign n5434 = x266 & ~n812 ;
  assign n5435 = x266 & n815 ;
  assign n5436 = ( ~n909 & n5434 ) | ( ~n909 & n5435 ) | ( n5434 & n5435 ) ;
  assign n5437 = ( n929 & n5434 ) | ( n929 & n5435 ) | ( n5434 & n5435 ) ;
  assign n5438 = ( ~n800 & n5436 ) | ( ~n800 & n5437 ) | ( n5436 & n5437 ) ;
  assign n5439 = ( n948 & n5436 ) | ( n948 & n5437 ) | ( n5436 & n5437 ) ;
  assign n5440 = ( n1061 & n5438 ) | ( n1061 & n5439 ) | ( n5438 & n5439 ) ;
  assign n5441 = n5433 | n5440 ;
  assign n5442 = ~n5426 & n5441 ;
  assign n5443 = ( ~n5396 & n5411 ) | ( ~n5396 & n5442 ) | ( n5411 & n5442 ) ;
  assign n5444 = ~n5364 & n5379 ;
  assign n5445 = n5349 | n5444 ;
  assign n5446 = ( ~n5381 & n5443 ) | ( ~n5381 & n5445 ) | ( n5443 & n5445 ) ;
  assign n5447 = x400 & n812 ;
  assign n5448 = x400 & ~n815 ;
  assign n5449 = ( n909 & n5447 ) | ( n909 & n5448 ) | ( n5447 & n5448 ) ;
  assign n5450 = ( ~n929 & n5447 ) | ( ~n929 & n5448 ) | ( n5447 & n5448 ) ;
  assign n5451 = ( n800 & n5449 ) | ( n800 & n5450 ) | ( n5449 & n5450 ) ;
  assign n5452 = ( ~n948 & n5449 ) | ( ~n948 & n5450 ) | ( n5449 & n5450 ) ;
  assign n5453 = ( ~n1061 & n5451 ) | ( ~n1061 & n5452 ) | ( n5451 & n5452 ) ;
  assign n5454 = x272 & ~n812 ;
  assign n5455 = x272 & n815 ;
  assign n5456 = ( ~n909 & n5454 ) | ( ~n909 & n5455 ) | ( n5454 & n5455 ) ;
  assign n5457 = ( n929 & n5454 ) | ( n929 & n5455 ) | ( n5454 & n5455 ) ;
  assign n5458 = ( ~n800 & n5456 ) | ( ~n800 & n5457 ) | ( n5456 & n5457 ) ;
  assign n5459 = ( n948 & n5456 ) | ( n948 & n5457 ) | ( n5456 & n5457 ) ;
  assign n5460 = ( n1061 & n5458 ) | ( n1061 & n5459 ) | ( n5458 & n5459 ) ;
  assign n5461 = n5453 | n5460 ;
  assign n5462 = x143 & n1370 ;
  assign n5463 = x143 & ~n1373 ;
  assign n5464 = ( n1467 & n5462 ) | ( n1467 & n5463 ) | ( n5462 & n5463 ) ;
  assign n5465 = ( ~n1487 & n5462 ) | ( ~n1487 & n5463 ) | ( n5462 & n5463 ) ;
  assign n5466 = ( n1358 & n5464 ) | ( n1358 & n5465 ) | ( n5464 & n5465 ) ;
  assign n5467 = ( ~n1506 & n5464 ) | ( ~n1506 & n5465 ) | ( n5464 & n5465 ) ;
  assign n5468 = ( ~n1612 & n5466 ) | ( ~n1612 & n5467 ) | ( n5466 & n5467 ) ;
  assign n5469 = x15 & ~n1370 ;
  assign n5470 = x15 & n1373 ;
  assign n5471 = ( ~n1467 & n5469 ) | ( ~n1467 & n5470 ) | ( n5469 & n5470 ) ;
  assign n5472 = ( n1487 & n5469 ) | ( n1487 & n5470 ) | ( n5469 & n5470 ) ;
  assign n5473 = ( ~n1358 & n5471 ) | ( ~n1358 & n5472 ) | ( n5471 & n5472 ) ;
  assign n5474 = ( n1506 & n5471 ) | ( n1506 & n5472 ) | ( n5471 & n5472 ) ;
  assign n5475 = ( n1612 & n5473 ) | ( n1612 & n5474 ) | ( n5473 & n5474 ) ;
  assign n5476 = n5468 | n5475 ;
  assign n5477 = x399 & n812 ;
  assign n5478 = x399 & ~n815 ;
  assign n5479 = ( n909 & n5477 ) | ( n909 & n5478 ) | ( n5477 & n5478 ) ;
  assign n5480 = ( ~n929 & n5477 ) | ( ~n929 & n5478 ) | ( n5477 & n5478 ) ;
  assign n5481 = ( n800 & n5479 ) | ( n800 & n5480 ) | ( n5479 & n5480 ) ;
  assign n5482 = ( ~n948 & n5479 ) | ( ~n948 & n5480 ) | ( n5479 & n5480 ) ;
  assign n5483 = ( ~n1061 & n5481 ) | ( ~n1061 & n5482 ) | ( n5481 & n5482 ) ;
  assign n5484 = x271 & ~n812 ;
  assign n5485 = x271 & n815 ;
  assign n5486 = ( ~n909 & n5484 ) | ( ~n909 & n5485 ) | ( n5484 & n5485 ) ;
  assign n5487 = ( n929 & n5484 ) | ( n929 & n5485 ) | ( n5484 & n5485 ) ;
  assign n5488 = ( ~n800 & n5486 ) | ( ~n800 & n5487 ) | ( n5486 & n5487 ) ;
  assign n5489 = ( n948 & n5486 ) | ( n948 & n5487 ) | ( n5486 & n5487 ) ;
  assign n5490 = ( n1061 & n5488 ) | ( n1061 & n5489 ) | ( n5488 & n5489 ) ;
  assign n5491 = n5483 | n5490 ;
  assign n5492 = ~n5476 & n5491 ;
  assign n5493 = x142 & n1370 ;
  assign n5494 = x142 & ~n1373 ;
  assign n5495 = ( n1467 & n5493 ) | ( n1467 & n5494 ) | ( n5493 & n5494 ) ;
  assign n5496 = ( ~n1487 & n5493 ) | ( ~n1487 & n5494 ) | ( n5493 & n5494 ) ;
  assign n5497 = ( n1358 & n5495 ) | ( n1358 & n5496 ) | ( n5495 & n5496 ) ;
  assign n5498 = ( ~n1506 & n5495 ) | ( ~n1506 & n5496 ) | ( n5495 & n5496 ) ;
  assign n5499 = ( ~n1612 & n5497 ) | ( ~n1612 & n5498 ) | ( n5497 & n5498 ) ;
  assign n5500 = x14 & ~n1370 ;
  assign n5501 = x14 & n1373 ;
  assign n5502 = ( ~n1467 & n5500 ) | ( ~n1467 & n5501 ) | ( n5500 & n5501 ) ;
  assign n5503 = ( n1487 & n5500 ) | ( n1487 & n5501 ) | ( n5500 & n5501 ) ;
  assign n5504 = ( ~n1358 & n5502 ) | ( ~n1358 & n5503 ) | ( n5502 & n5503 ) ;
  assign n5505 = ( n1506 & n5502 ) | ( n1506 & n5503 ) | ( n5502 & n5503 ) ;
  assign n5506 = ( n1612 & n5504 ) | ( n1612 & n5505 ) | ( n5504 & n5505 ) ;
  assign n5507 = n5499 | n5506 ;
  assign n5508 = x398 & n812 ;
  assign n5509 = x398 & ~n815 ;
  assign n5510 = ( n909 & n5508 ) | ( n909 & n5509 ) | ( n5508 & n5509 ) ;
  assign n5511 = ( ~n929 & n5508 ) | ( ~n929 & n5509 ) | ( n5508 & n5509 ) ;
  assign n5512 = ( n800 & n5510 ) | ( n800 & n5511 ) | ( n5510 & n5511 ) ;
  assign n5513 = ( ~n948 & n5510 ) | ( ~n948 & n5511 ) | ( n5510 & n5511 ) ;
  assign n5514 = ( ~n1061 & n5512 ) | ( ~n1061 & n5513 ) | ( n5512 & n5513 ) ;
  assign n5515 = x270 & ~n812 ;
  assign n5516 = x270 & n815 ;
  assign n5517 = ( ~n909 & n5515 ) | ( ~n909 & n5516 ) | ( n5515 & n5516 ) ;
  assign n5518 = ( n929 & n5515 ) | ( n929 & n5516 ) | ( n5515 & n5516 ) ;
  assign n5519 = ( ~n800 & n5517 ) | ( ~n800 & n5518 ) | ( n5517 & n5518 ) ;
  assign n5520 = ( n948 & n5517 ) | ( n948 & n5518 ) | ( n5517 & n5518 ) ;
  assign n5521 = ( n1061 & n5519 ) | ( n1061 & n5520 ) | ( n5519 & n5520 ) ;
  assign n5522 = n5514 | n5521 ;
  assign n5523 = ~n5507 & n5522 ;
  assign n5524 = n5333 & ~n5348 ;
  assign n5525 = ~n5523 & n5524 ;
  assign n5526 = n5507 & ~n5522 ;
  assign n5527 = ~n5492 & n5526 ;
  assign n5528 = ( ~n5492 & n5525 ) | ( ~n5492 & n5527 ) | ( n5525 & n5527 ) ;
  assign n5529 = n5476 & ~n5491 ;
  assign n5530 = x144 & n1370 ;
  assign n5531 = x144 & ~n1373 ;
  assign n5532 = ( n1467 & n5530 ) | ( n1467 & n5531 ) | ( n5530 & n5531 ) ;
  assign n5533 = ( ~n1487 & n5530 ) | ( ~n1487 & n5531 ) | ( n5530 & n5531 ) ;
  assign n5534 = ( n1358 & n5532 ) | ( n1358 & n5533 ) | ( n5532 & n5533 ) ;
  assign n5535 = ( ~n1506 & n5532 ) | ( ~n1506 & n5533 ) | ( n5532 & n5533 ) ;
  assign n5536 = ( ~n1612 & n5534 ) | ( ~n1612 & n5535 ) | ( n5534 & n5535 ) ;
  assign n5537 = x16 & ~n1370 ;
  assign n5538 = x16 & n1373 ;
  assign n5539 = ( ~n1467 & n5537 ) | ( ~n1467 & n5538 ) | ( n5537 & n5538 ) ;
  assign n5540 = ( n1487 & n5537 ) | ( n1487 & n5538 ) | ( n5537 & n5538 ) ;
  assign n5541 = ( ~n1358 & n5539 ) | ( ~n1358 & n5540 ) | ( n5539 & n5540 ) ;
  assign n5542 = ( n1506 & n5539 ) | ( n1506 & n5540 ) | ( n5539 & n5540 ) ;
  assign n5543 = ( n1612 & n5541 ) | ( n1612 & n5542 ) | ( n5541 & n5542 ) ;
  assign n5544 = n5536 | n5543 ;
  assign n5545 = ~n5461 & n5544 ;
  assign n5546 = ( ~n5461 & n5529 ) | ( ~n5461 & n5545 ) | ( n5529 & n5545 ) ;
  assign n5547 = ( ~n5461 & n5528 ) | ( ~n5461 & n5546 ) | ( n5528 & n5546 ) ;
  assign n5548 = n5492 | n5523 ;
  assign n5549 = ~n5529 & n5548 ;
  assign n5550 = ( n5461 & ~n5545 ) | ( n5461 & n5549 ) | ( ~n5545 & n5549 ) ;
  assign n5551 = ( n5446 & ~n5547 ) | ( n5446 & n5550 ) | ( ~n5547 & n5550 ) ;
  assign n5552 = ( ~n5461 & n5527 ) | ( ~n5461 & n5546 ) | ( n5527 & n5546 ) ;
  assign n5553 = n5396 & ~n5411 ;
  assign n5554 = ~n5444 & n5553 ;
  assign n5555 = n5426 & ~n5441 ;
  assign n5556 = ~n5443 & n5555 ;
  assign n5557 = ( ~n5444 & n5554 ) | ( ~n5444 & n5556 ) | ( n5554 & n5556 ) ;
  assign n5558 = ( ~n5349 & n5381 ) | ( ~n5349 & n5557 ) | ( n5381 & n5557 ) ;
  assign n5559 = n5524 | n5558 ;
  assign n5560 = ( ~n5550 & n5552 ) | ( ~n5550 & n5559 ) | ( n5552 & n5559 ) ;
  assign n5561 = x392 & n812 ;
  assign n5562 = x392 & ~n815 ;
  assign n5563 = ( n909 & n5561 ) | ( n909 & n5562 ) | ( n5561 & n5562 ) ;
  assign n5564 = ( ~n929 & n5561 ) | ( ~n929 & n5562 ) | ( n5561 & n5562 ) ;
  assign n5565 = ( n800 & n5563 ) | ( n800 & n5564 ) | ( n5563 & n5564 ) ;
  assign n5566 = ( ~n948 & n5563 ) | ( ~n948 & n5564 ) | ( n5563 & n5564 ) ;
  assign n5567 = ( ~n1061 & n5565 ) | ( ~n1061 & n5566 ) | ( n5565 & n5566 ) ;
  assign n5568 = x264 & ~n812 ;
  assign n5569 = x264 & n815 ;
  assign n5570 = ( ~n909 & n5568 ) | ( ~n909 & n5569 ) | ( n5568 & n5569 ) ;
  assign n5571 = ( n929 & n5568 ) | ( n929 & n5569 ) | ( n5568 & n5569 ) ;
  assign n5572 = ( ~n800 & n5570 ) | ( ~n800 & n5571 ) | ( n5570 & n5571 ) ;
  assign n5573 = ( n948 & n5570 ) | ( n948 & n5571 ) | ( n5570 & n5571 ) ;
  assign n5574 = ( n1061 & n5572 ) | ( n1061 & n5573 ) | ( n5572 & n5573 ) ;
  assign n5575 = n5567 | n5574 ;
  assign n5576 = x135 & n1370 ;
  assign n5577 = x135 & ~n1373 ;
  assign n5578 = ( n1467 & n5576 ) | ( n1467 & n5577 ) | ( n5576 & n5577 ) ;
  assign n5579 = ( ~n1487 & n5576 ) | ( ~n1487 & n5577 ) | ( n5576 & n5577 ) ;
  assign n5580 = ( n1358 & n5578 ) | ( n1358 & n5579 ) | ( n5578 & n5579 ) ;
  assign n5581 = ( ~n1506 & n5578 ) | ( ~n1506 & n5579 ) | ( n5578 & n5579 ) ;
  assign n5582 = ( ~n1612 & n5580 ) | ( ~n1612 & n5581 ) | ( n5580 & n5581 ) ;
  assign n5583 = x7 & ~n1370 ;
  assign n5584 = x7 & n1373 ;
  assign n5585 = ( ~n1467 & n5583 ) | ( ~n1467 & n5584 ) | ( n5583 & n5584 ) ;
  assign n5586 = ( n1487 & n5583 ) | ( n1487 & n5584 ) | ( n5583 & n5584 ) ;
  assign n5587 = ( ~n1358 & n5585 ) | ( ~n1358 & n5586 ) | ( n5585 & n5586 ) ;
  assign n5588 = ( n1506 & n5585 ) | ( n1506 & n5586 ) | ( n5585 & n5586 ) ;
  assign n5589 = ( n1612 & n5587 ) | ( n1612 & n5588 ) | ( n5587 & n5588 ) ;
  assign n5590 = n5582 | n5589 ;
  assign n5591 = x391 & n812 ;
  assign n5592 = x391 & ~n815 ;
  assign n5593 = ( n909 & n5591 ) | ( n909 & n5592 ) | ( n5591 & n5592 ) ;
  assign n5594 = ( ~n929 & n5591 ) | ( ~n929 & n5592 ) | ( n5591 & n5592 ) ;
  assign n5595 = ( n800 & n5593 ) | ( n800 & n5594 ) | ( n5593 & n5594 ) ;
  assign n5596 = ( ~n948 & n5593 ) | ( ~n948 & n5594 ) | ( n5593 & n5594 ) ;
  assign n5597 = ( ~n1061 & n5595 ) | ( ~n1061 & n5596 ) | ( n5595 & n5596 ) ;
  assign n5598 = x263 & ~n812 ;
  assign n5599 = x263 & n815 ;
  assign n5600 = ( ~n909 & n5598 ) | ( ~n909 & n5599 ) | ( n5598 & n5599 ) ;
  assign n5601 = ( n929 & n5598 ) | ( n929 & n5599 ) | ( n5598 & n5599 ) ;
  assign n5602 = ( ~n800 & n5600 ) | ( ~n800 & n5601 ) | ( n5600 & n5601 ) ;
  assign n5603 = ( n948 & n5600 ) | ( n948 & n5601 ) | ( n5600 & n5601 ) ;
  assign n5604 = ( n1061 & n5602 ) | ( n1061 & n5603 ) | ( n5602 & n5603 ) ;
  assign n5605 = n5597 | n5604 ;
  assign n5606 = ~n5590 & n5605 ;
  assign n5607 = x136 & n1370 ;
  assign n5608 = x136 & ~n1373 ;
  assign n5609 = ( n1467 & n5607 ) | ( n1467 & n5608 ) | ( n5607 & n5608 ) ;
  assign n5610 = ( ~n1487 & n5607 ) | ( ~n1487 & n5608 ) | ( n5607 & n5608 ) ;
  assign n5611 = ( n1358 & n5609 ) | ( n1358 & n5610 ) | ( n5609 & n5610 ) ;
  assign n5612 = ( ~n1506 & n5609 ) | ( ~n1506 & n5610 ) | ( n5609 & n5610 ) ;
  assign n5613 = ( ~n1612 & n5611 ) | ( ~n1612 & n5612 ) | ( n5611 & n5612 ) ;
  assign n5614 = x8 & ~n1370 ;
  assign n5615 = x8 & n1373 ;
  assign n5616 = ( ~n1467 & n5614 ) | ( ~n1467 & n5615 ) | ( n5614 & n5615 ) ;
  assign n5617 = ( n1487 & n5614 ) | ( n1487 & n5615 ) | ( n5614 & n5615 ) ;
  assign n5618 = ( ~n1358 & n5616 ) | ( ~n1358 & n5617 ) | ( n5616 & n5617 ) ;
  assign n5619 = ( n1506 & n5616 ) | ( n1506 & n5617 ) | ( n5616 & n5617 ) ;
  assign n5620 = ( n1612 & n5618 ) | ( n1612 & n5619 ) | ( n5618 & n5619 ) ;
  assign n5621 = n5613 | n5620 ;
  assign n5622 = ~n5575 & n5621 ;
  assign n5623 = ( n5575 & n5606 ) | ( n5575 & ~n5622 ) | ( n5606 & ~n5622 ) ;
  assign n5624 = n5590 & ~n5605 ;
  assign n5625 = ( ~n5575 & n5622 ) | ( ~n5575 & n5624 ) | ( n5622 & n5624 ) ;
  assign n5626 = x134 & n1370 ;
  assign n5627 = x134 & ~n1373 ;
  assign n5628 = ( n1467 & n5626 ) | ( n1467 & n5627 ) | ( n5626 & n5627 ) ;
  assign n5629 = ( ~n1487 & n5626 ) | ( ~n1487 & n5627 ) | ( n5626 & n5627 ) ;
  assign n5630 = ( n1358 & n5628 ) | ( n1358 & n5629 ) | ( n5628 & n5629 ) ;
  assign n5631 = ( ~n1506 & n5628 ) | ( ~n1506 & n5629 ) | ( n5628 & n5629 ) ;
  assign n5632 = ( ~n1612 & n5630 ) | ( ~n1612 & n5631 ) | ( n5630 & n5631 ) ;
  assign n5633 = x6 & ~n1370 ;
  assign n5634 = x6 & n1373 ;
  assign n5635 = ( ~n1467 & n5633 ) | ( ~n1467 & n5634 ) | ( n5633 & n5634 ) ;
  assign n5636 = ( n1487 & n5633 ) | ( n1487 & n5634 ) | ( n5633 & n5634 ) ;
  assign n5637 = ( ~n1358 & n5635 ) | ( ~n1358 & n5636 ) | ( n5635 & n5636 ) ;
  assign n5638 = ( n1506 & n5635 ) | ( n1506 & n5636 ) | ( n5635 & n5636 ) ;
  assign n5639 = ( n1612 & n5637 ) | ( n1612 & n5638 ) | ( n5637 & n5638 ) ;
  assign n5640 = n5632 | n5639 ;
  assign n5641 = x390 & n812 ;
  assign n5642 = x390 & ~n815 ;
  assign n5643 = ( n909 & n5641 ) | ( n909 & n5642 ) | ( n5641 & n5642 ) ;
  assign n5644 = ( ~n929 & n5641 ) | ( ~n929 & n5642 ) | ( n5641 & n5642 ) ;
  assign n5645 = ( n800 & n5643 ) | ( n800 & n5644 ) | ( n5643 & n5644 ) ;
  assign n5646 = ( ~n948 & n5643 ) | ( ~n948 & n5644 ) | ( n5643 & n5644 ) ;
  assign n5647 = ( ~n1061 & n5645 ) | ( ~n1061 & n5646 ) | ( n5645 & n5646 ) ;
  assign n5648 = x262 & ~n812 ;
  assign n5649 = x262 & n815 ;
  assign n5650 = ( ~n909 & n5648 ) | ( ~n909 & n5649 ) | ( n5648 & n5649 ) ;
  assign n5651 = ( n929 & n5648 ) | ( n929 & n5649 ) | ( n5648 & n5649 ) ;
  assign n5652 = ( ~n800 & n5650 ) | ( ~n800 & n5651 ) | ( n5650 & n5651 ) ;
  assign n5653 = ( n948 & n5650 ) | ( n948 & n5651 ) | ( n5650 & n5651 ) ;
  assign n5654 = ( n1061 & n5652 ) | ( n1061 & n5653 ) | ( n5652 & n5653 ) ;
  assign n5655 = n5647 | n5654 ;
  assign n5656 = x133 & n1370 ;
  assign n5657 = x133 & ~n1373 ;
  assign n5658 = ( n1467 & n5656 ) | ( n1467 & n5657 ) | ( n5656 & n5657 ) ;
  assign n5659 = ( ~n1487 & n5656 ) | ( ~n1487 & n5657 ) | ( n5656 & n5657 ) ;
  assign n5660 = ( n1358 & n5658 ) | ( n1358 & n5659 ) | ( n5658 & n5659 ) ;
  assign n5661 = ( ~n1506 & n5658 ) | ( ~n1506 & n5659 ) | ( n5658 & n5659 ) ;
  assign n5662 = ( ~n1612 & n5660 ) | ( ~n1612 & n5661 ) | ( n5660 & n5661 ) ;
  assign n5663 = x5 & ~n1370 ;
  assign n5664 = x5 & n1373 ;
  assign n5665 = ( ~n1467 & n5663 ) | ( ~n1467 & n5664 ) | ( n5663 & n5664 ) ;
  assign n5666 = ( n1487 & n5663 ) | ( n1487 & n5664 ) | ( n5663 & n5664 ) ;
  assign n5667 = ( ~n1358 & n5665 ) | ( ~n1358 & n5666 ) | ( n5665 & n5666 ) ;
  assign n5668 = ( n1506 & n5665 ) | ( n1506 & n5666 ) | ( n5665 & n5666 ) ;
  assign n5669 = ( n1612 & n5667 ) | ( n1612 & n5668 ) | ( n5667 & n5668 ) ;
  assign n5670 = n5662 | n5669 ;
  assign n5671 = x389 & n812 ;
  assign n5672 = x389 & ~n815 ;
  assign n5673 = ( n909 & n5671 ) | ( n909 & n5672 ) | ( n5671 & n5672 ) ;
  assign n5674 = ( ~n929 & n5671 ) | ( ~n929 & n5672 ) | ( n5671 & n5672 ) ;
  assign n5675 = ( n800 & n5673 ) | ( n800 & n5674 ) | ( n5673 & n5674 ) ;
  assign n5676 = ( ~n948 & n5673 ) | ( ~n948 & n5674 ) | ( n5673 & n5674 ) ;
  assign n5677 = ( ~n1061 & n5675 ) | ( ~n1061 & n5676 ) | ( n5675 & n5676 ) ;
  assign n5678 = x261 & ~n812 ;
  assign n5679 = x261 & n815 ;
  assign n5680 = ( ~n909 & n5678 ) | ( ~n909 & n5679 ) | ( n5678 & n5679 ) ;
  assign n5681 = ( n929 & n5678 ) | ( n929 & n5679 ) | ( n5678 & n5679 ) ;
  assign n5682 = ( ~n800 & n5680 ) | ( ~n800 & n5681 ) | ( n5680 & n5681 ) ;
  assign n5683 = ( n948 & n5680 ) | ( n948 & n5681 ) | ( n5680 & n5681 ) ;
  assign n5684 = ( n1061 & n5682 ) | ( n1061 & n5683 ) | ( n5682 & n5683 ) ;
  assign n5685 = n5677 | n5684 ;
  assign n5686 = x132 & n1370 ;
  assign n5687 = x132 & ~n1373 ;
  assign n5688 = ( n1467 & n5686 ) | ( n1467 & n5687 ) | ( n5686 & n5687 ) ;
  assign n5689 = ( ~n1487 & n5686 ) | ( ~n1487 & n5687 ) | ( n5686 & n5687 ) ;
  assign n5690 = ( n1358 & n5688 ) | ( n1358 & n5689 ) | ( n5688 & n5689 ) ;
  assign n5691 = ( ~n1506 & n5688 ) | ( ~n1506 & n5689 ) | ( n5688 & n5689 ) ;
  assign n5692 = ( ~n1612 & n5690 ) | ( ~n1612 & n5691 ) | ( n5690 & n5691 ) ;
  assign n5693 = x4 & ~n1370 ;
  assign n5694 = x4 & n1373 ;
  assign n5695 = ( ~n1467 & n5693 ) | ( ~n1467 & n5694 ) | ( n5693 & n5694 ) ;
  assign n5696 = ( n1487 & n5693 ) | ( n1487 & n5694 ) | ( n5693 & n5694 ) ;
  assign n5697 = ( ~n1358 & n5695 ) | ( ~n1358 & n5696 ) | ( n5695 & n5696 ) ;
  assign n5698 = ( n1506 & n5695 ) | ( n1506 & n5696 ) | ( n5695 & n5696 ) ;
  assign n5699 = ( n1612 & n5697 ) | ( n1612 & n5698 ) | ( n5697 & n5698 ) ;
  assign n5700 = n5692 | n5699 ;
  assign n5701 = x388 & n812 ;
  assign n5702 = x388 & ~n815 ;
  assign n5703 = ( n909 & n5701 ) | ( n909 & n5702 ) | ( n5701 & n5702 ) ;
  assign n5704 = ( ~n929 & n5701 ) | ( ~n929 & n5702 ) | ( n5701 & n5702 ) ;
  assign n5705 = ( n800 & n5703 ) | ( n800 & n5704 ) | ( n5703 & n5704 ) ;
  assign n5706 = ( ~n948 & n5703 ) | ( ~n948 & n5704 ) | ( n5703 & n5704 ) ;
  assign n5707 = ( ~n1061 & n5705 ) | ( ~n1061 & n5706 ) | ( n5705 & n5706 ) ;
  assign n5708 = x260 & ~n812 ;
  assign n5709 = x260 & n815 ;
  assign n5710 = ( ~n909 & n5708 ) | ( ~n909 & n5709 ) | ( n5708 & n5709 ) ;
  assign n5711 = ( n929 & n5708 ) | ( n929 & n5709 ) | ( n5708 & n5709 ) ;
  assign n5712 = ( ~n800 & n5710 ) | ( ~n800 & n5711 ) | ( n5710 & n5711 ) ;
  assign n5713 = ( n948 & n5710 ) | ( n948 & n5711 ) | ( n5710 & n5711 ) ;
  assign n5714 = ( n1061 & n5712 ) | ( n1061 & n5713 ) | ( n5712 & n5713 ) ;
  assign n5715 = n5707 | n5714 ;
  assign n5716 = x131 & n1370 ;
  assign n5717 = x131 & ~n1373 ;
  assign n5718 = ( n1467 & n5716 ) | ( n1467 & n5717 ) | ( n5716 & n5717 ) ;
  assign n5719 = ( ~n1487 & n5716 ) | ( ~n1487 & n5717 ) | ( n5716 & n5717 ) ;
  assign n5720 = ( n1358 & n5718 ) | ( n1358 & n5719 ) | ( n5718 & n5719 ) ;
  assign n5721 = ( ~n1506 & n5718 ) | ( ~n1506 & n5719 ) | ( n5718 & n5719 ) ;
  assign n5722 = ( ~n1612 & n5720 ) | ( ~n1612 & n5721 ) | ( n5720 & n5721 ) ;
  assign n5723 = x3 & ~n1370 ;
  assign n5724 = x3 & n1373 ;
  assign n5725 = ( ~n1467 & n5723 ) | ( ~n1467 & n5724 ) | ( n5723 & n5724 ) ;
  assign n5726 = ( n1487 & n5723 ) | ( n1487 & n5724 ) | ( n5723 & n5724 ) ;
  assign n5727 = ( ~n1358 & n5725 ) | ( ~n1358 & n5726 ) | ( n5725 & n5726 ) ;
  assign n5728 = ( n1506 & n5725 ) | ( n1506 & n5726 ) | ( n5725 & n5726 ) ;
  assign n5729 = ( n1612 & n5727 ) | ( n1612 & n5728 ) | ( n5727 & n5728 ) ;
  assign n5730 = n5722 | n5729 ;
  assign n5731 = x387 & n812 ;
  assign n5732 = x387 & ~n815 ;
  assign n5733 = ( n909 & n5731 ) | ( n909 & n5732 ) | ( n5731 & n5732 ) ;
  assign n5734 = ( ~n929 & n5731 ) | ( ~n929 & n5732 ) | ( n5731 & n5732 ) ;
  assign n5735 = ( n800 & n5733 ) | ( n800 & n5734 ) | ( n5733 & n5734 ) ;
  assign n5736 = ( ~n948 & n5733 ) | ( ~n948 & n5734 ) | ( n5733 & n5734 ) ;
  assign n5737 = ( ~n1061 & n5735 ) | ( ~n1061 & n5736 ) | ( n5735 & n5736 ) ;
  assign n5738 = x259 & ~n812 ;
  assign n5739 = x259 & n815 ;
  assign n5740 = ( ~n909 & n5738 ) | ( ~n909 & n5739 ) | ( n5738 & n5739 ) ;
  assign n5741 = ( n929 & n5738 ) | ( n929 & n5739 ) | ( n5738 & n5739 ) ;
  assign n5742 = ( ~n800 & n5740 ) | ( ~n800 & n5741 ) | ( n5740 & n5741 ) ;
  assign n5743 = ( n948 & n5740 ) | ( n948 & n5741 ) | ( n5740 & n5741 ) ;
  assign n5744 = ( n1061 & n5742 ) | ( n1061 & n5743 ) | ( n5742 & n5743 ) ;
  assign n5745 = n5737 | n5744 ;
  assign n5746 = x130 & n1370 ;
  assign n5747 = x130 & ~n1373 ;
  assign n5748 = ( n1467 & n5746 ) | ( n1467 & n5747 ) | ( n5746 & n5747 ) ;
  assign n5749 = ( ~n1487 & n5746 ) | ( ~n1487 & n5747 ) | ( n5746 & n5747 ) ;
  assign n5750 = ( n1358 & n5748 ) | ( n1358 & n5749 ) | ( n5748 & n5749 ) ;
  assign n5751 = ( ~n1506 & n5748 ) | ( ~n1506 & n5749 ) | ( n5748 & n5749 ) ;
  assign n5752 = ( ~n1612 & n5750 ) | ( ~n1612 & n5751 ) | ( n5750 & n5751 ) ;
  assign n5753 = x2 & ~n1370 ;
  assign n5754 = x2 & n1373 ;
  assign n5755 = ( ~n1467 & n5753 ) | ( ~n1467 & n5754 ) | ( n5753 & n5754 ) ;
  assign n5756 = ( n1487 & n5753 ) | ( n1487 & n5754 ) | ( n5753 & n5754 ) ;
  assign n5757 = ( ~n1358 & n5755 ) | ( ~n1358 & n5756 ) | ( n5755 & n5756 ) ;
  assign n5758 = ( n1506 & n5755 ) | ( n1506 & n5756 ) | ( n5755 & n5756 ) ;
  assign n5759 = ( n1612 & n5757 ) | ( n1612 & n5758 ) | ( n5757 & n5758 ) ;
  assign n5760 = n5752 | n5759 ;
  assign n5761 = x386 & n812 ;
  assign n5762 = x386 & ~n815 ;
  assign n5763 = ( n909 & n5761 ) | ( n909 & n5762 ) | ( n5761 & n5762 ) ;
  assign n5764 = ( ~n929 & n5761 ) | ( ~n929 & n5762 ) | ( n5761 & n5762 ) ;
  assign n5765 = ( n800 & n5763 ) | ( n800 & n5764 ) | ( n5763 & n5764 ) ;
  assign n5766 = ( ~n948 & n5763 ) | ( ~n948 & n5764 ) | ( n5763 & n5764 ) ;
  assign n5767 = ( ~n1061 & n5765 ) | ( ~n1061 & n5766 ) | ( n5765 & n5766 ) ;
  assign n5768 = x258 & ~n812 ;
  assign n5769 = x258 & n815 ;
  assign n5770 = ( ~n909 & n5768 ) | ( ~n909 & n5769 ) | ( n5768 & n5769 ) ;
  assign n5771 = ( n929 & n5768 ) | ( n929 & n5769 ) | ( n5768 & n5769 ) ;
  assign n5772 = ( ~n800 & n5770 ) | ( ~n800 & n5771 ) | ( n5770 & n5771 ) ;
  assign n5773 = ( n948 & n5770 ) | ( n948 & n5771 ) | ( n5770 & n5771 ) ;
  assign n5774 = ( n1061 & n5772 ) | ( n1061 & n5773 ) | ( n5772 & n5773 ) ;
  assign n5775 = n5767 | n5774 ;
  assign n5776 = x385 & n812 ;
  assign n5777 = x385 & ~n815 ;
  assign n5778 = ( n909 & n5776 ) | ( n909 & n5777 ) | ( n5776 & n5777 ) ;
  assign n5779 = ( ~n929 & n5776 ) | ( ~n929 & n5777 ) | ( n5776 & n5777 ) ;
  assign n5780 = ( n800 & n5778 ) | ( n800 & n5779 ) | ( n5778 & n5779 ) ;
  assign n5781 = ( ~n948 & n5778 ) | ( ~n948 & n5779 ) | ( n5778 & n5779 ) ;
  assign n5782 = ( ~n1061 & n5780 ) | ( ~n1061 & n5781 ) | ( n5780 & n5781 ) ;
  assign n5783 = x257 & ~n812 ;
  assign n5784 = x257 & n815 ;
  assign n5785 = ( ~n909 & n5783 ) | ( ~n909 & n5784 ) | ( n5783 & n5784 ) ;
  assign n5786 = ( n929 & n5783 ) | ( n929 & n5784 ) | ( n5783 & n5784 ) ;
  assign n5787 = ( ~n800 & n5785 ) | ( ~n800 & n5786 ) | ( n5785 & n5786 ) ;
  assign n5788 = ( n948 & n5785 ) | ( n948 & n5786 ) | ( n5785 & n5786 ) ;
  assign n5789 = ( n1061 & n5787 ) | ( n1061 & n5788 ) | ( n5787 & n5788 ) ;
  assign n5790 = n5782 | n5789 ;
  assign n5791 = x128 & n1370 ;
  assign n5792 = x128 & ~n1373 ;
  assign n5793 = ( n1467 & n5791 ) | ( n1467 & n5792 ) | ( n5791 & n5792 ) ;
  assign n5794 = ( ~n1487 & n5791 ) | ( ~n1487 & n5792 ) | ( n5791 & n5792 ) ;
  assign n5795 = ( n1358 & n5793 ) | ( n1358 & n5794 ) | ( n5793 & n5794 ) ;
  assign n5796 = ( ~n1506 & n5793 ) | ( ~n1506 & n5794 ) | ( n5793 & n5794 ) ;
  assign n5797 = ( ~n1612 & n5795 ) | ( ~n1612 & n5796 ) | ( n5795 & n5796 ) ;
  assign n5798 = x0 & ~n1370 ;
  assign n5799 = x0 & n1373 ;
  assign n5800 = ( ~n1467 & n5798 ) | ( ~n1467 & n5799 ) | ( n5798 & n5799 ) ;
  assign n5801 = ( n1487 & n5798 ) | ( n1487 & n5799 ) | ( n5798 & n5799 ) ;
  assign n5802 = ( ~n1358 & n5800 ) | ( ~n1358 & n5801 ) | ( n5800 & n5801 ) ;
  assign n5803 = ( n1506 & n5800 ) | ( n1506 & n5801 ) | ( n5800 & n5801 ) ;
  assign n5804 = ( n1612 & n5802 ) | ( n1612 & n5803 ) | ( n5802 & n5803 ) ;
  assign n5805 = n5797 | n5804 ;
  assign n5806 = ~n1070 & n5805 ;
  assign n5807 = x129 & n1370 ;
  assign n5808 = x129 & ~n1373 ;
  assign n5809 = ( n1467 & n5807 ) | ( n1467 & n5808 ) | ( n5807 & n5808 ) ;
  assign n5810 = ( ~n1487 & n5807 ) | ( ~n1487 & n5808 ) | ( n5807 & n5808 ) ;
  assign n5811 = ( n1358 & n5809 ) | ( n1358 & n5810 ) | ( n5809 & n5810 ) ;
  assign n5812 = ( ~n1506 & n5809 ) | ( ~n1506 & n5810 ) | ( n5809 & n5810 ) ;
  assign n5813 = ( ~n1612 & n5811 ) | ( ~n1612 & n5812 ) | ( n5811 & n5812 ) ;
  assign n5814 = x1 & ~n1370 ;
  assign n5815 = x1 & n1373 ;
  assign n5816 = ( ~n1467 & n5814 ) | ( ~n1467 & n5815 ) | ( n5814 & n5815 ) ;
  assign n5817 = ( n1487 & n5814 ) | ( n1487 & n5815 ) | ( n5814 & n5815 ) ;
  assign n5818 = ( ~n1358 & n5816 ) | ( ~n1358 & n5817 ) | ( n5816 & n5817 ) ;
  assign n5819 = ( n1506 & n5816 ) | ( n1506 & n5817 ) | ( n5816 & n5817 ) ;
  assign n5820 = ( n1612 & n5818 ) | ( n1612 & n5819 ) | ( n5818 & n5819 ) ;
  assign n5821 = n5813 | n5820 ;
  assign n5822 = ( ~n5790 & n5806 ) | ( ~n5790 & n5821 ) | ( n5806 & n5821 ) ;
  assign n5823 = ( n5760 & ~n5775 ) | ( n5760 & n5822 ) | ( ~n5775 & n5822 ) ;
  assign n5824 = ( n5730 & ~n5745 ) | ( n5730 & n5823 ) | ( ~n5745 & n5823 ) ;
  assign n5825 = ( n5700 & ~n5715 ) | ( n5700 & n5824 ) | ( ~n5715 & n5824 ) ;
  assign n5826 = ( n5670 & ~n5685 ) | ( n5670 & n5825 ) | ( ~n5685 & n5825 ) ;
  assign n5827 = ( n5640 & ~n5655 ) | ( n5640 & n5826 ) | ( ~n5655 & n5826 ) ;
  assign n5828 = ( ~n5623 & n5625 ) | ( ~n5623 & n5827 ) | ( n5625 & n5827 ) ;
  assign n5829 = ( ~n5606 & n5624 ) | ( ~n5606 & n5827 ) | ( n5624 & n5827 ) ;
  assign n5830 = n5621 & n5829 ;
  assign n5831 = n5828 | n5830 ;
  assign n5832 = x137 & n1370 ;
  assign n5833 = x137 & ~n1373 ;
  assign n5834 = ( n1467 & n5832 ) | ( n1467 & n5833 ) | ( n5832 & n5833 ) ;
  assign n5835 = ( ~n1487 & n5832 ) | ( ~n1487 & n5833 ) | ( n5832 & n5833 ) ;
  assign n5836 = ( n1358 & n5834 ) | ( n1358 & n5835 ) | ( n5834 & n5835 ) ;
  assign n5837 = ( ~n1506 & n5834 ) | ( ~n1506 & n5835 ) | ( n5834 & n5835 ) ;
  assign n5838 = ( ~n1612 & n5836 ) | ( ~n1612 & n5837 ) | ( n5836 & n5837 ) ;
  assign n5839 = x9 & ~n1370 ;
  assign n5840 = x9 & n1373 ;
  assign n5841 = ( ~n1467 & n5839 ) | ( ~n1467 & n5840 ) | ( n5839 & n5840 ) ;
  assign n5842 = ( n1487 & n5839 ) | ( n1487 & n5840 ) | ( n5839 & n5840 ) ;
  assign n5843 = ( ~n1358 & n5841 ) | ( ~n1358 & n5842 ) | ( n5841 & n5842 ) ;
  assign n5844 = ( n1506 & n5841 ) | ( n1506 & n5842 ) | ( n5841 & n5842 ) ;
  assign n5845 = ( n1612 & n5843 ) | ( n1612 & n5844 ) | ( n5843 & n5844 ) ;
  assign n5846 = n5838 | n5845 ;
  assign n5847 = x393 & n812 ;
  assign n5848 = x393 & ~n815 ;
  assign n5849 = ( n909 & n5847 ) | ( n909 & n5848 ) | ( n5847 & n5848 ) ;
  assign n5850 = ( ~n929 & n5847 ) | ( ~n929 & n5848 ) | ( n5847 & n5848 ) ;
  assign n5851 = ( n800 & n5849 ) | ( n800 & n5850 ) | ( n5849 & n5850 ) ;
  assign n5852 = ( ~n948 & n5849 ) | ( ~n948 & n5850 ) | ( n5849 & n5850 ) ;
  assign n5853 = ( ~n1061 & n5851 ) | ( ~n1061 & n5852 ) | ( n5851 & n5852 ) ;
  assign n5854 = x265 & ~n812 ;
  assign n5855 = x265 & n815 ;
  assign n5856 = ( ~n909 & n5854 ) | ( ~n909 & n5855 ) | ( n5854 & n5855 ) ;
  assign n5857 = ( n929 & n5854 ) | ( n929 & n5855 ) | ( n5854 & n5855 ) ;
  assign n5858 = ( ~n800 & n5856 ) | ( ~n800 & n5857 ) | ( n5856 & n5857 ) ;
  assign n5859 = ( n948 & n5856 ) | ( n948 & n5857 ) | ( n5856 & n5857 ) ;
  assign n5860 = ( n1061 & n5858 ) | ( n1061 & n5859 ) | ( n5858 & n5859 ) ;
  assign n5861 = n5853 | n5860 ;
  assign n5862 = ( n5831 & n5846 ) | ( n5831 & ~n5861 ) | ( n5846 & ~n5861 ) ;
  assign n5863 = ( ~n5551 & n5560 ) | ( ~n5551 & n5862 ) | ( n5560 & n5862 ) ;
  assign n5864 = n5529 & n5544 ;
  assign n5865 = ( n5527 & n5544 ) | ( n5527 & n5864 ) | ( n5544 & n5864 ) ;
  assign n5866 = ( n5544 & ~n5548 ) | ( n5544 & n5864 ) | ( ~n5548 & n5864 ) ;
  assign n5867 = ( n5559 & n5865 ) | ( n5559 & n5866 ) | ( n5865 & n5866 ) ;
  assign n5868 = ( n5528 & n5544 ) | ( n5528 & n5864 ) | ( n5544 & n5864 ) ;
  assign n5869 = ( ~n5446 & n5866 ) | ( ~n5446 & n5868 ) | ( n5866 & n5868 ) ;
  assign n5870 = ( n5862 & n5867 ) | ( n5862 & n5869 ) | ( n5867 & n5869 ) ;
  assign n5871 = n5863 | n5870 ;
  assign n5872 = x145 & n1370 ;
  assign n5873 = x145 & ~n1373 ;
  assign n5874 = ( n1467 & n5872 ) | ( n1467 & n5873 ) | ( n5872 & n5873 ) ;
  assign n5875 = ( ~n1487 & n5872 ) | ( ~n1487 & n5873 ) | ( n5872 & n5873 ) ;
  assign n5876 = ( n1358 & n5874 ) | ( n1358 & n5875 ) | ( n5874 & n5875 ) ;
  assign n5877 = ( ~n1506 & n5874 ) | ( ~n1506 & n5875 ) | ( n5874 & n5875 ) ;
  assign n5878 = ( ~n1612 & n5876 ) | ( ~n1612 & n5877 ) | ( n5876 & n5877 ) ;
  assign n5879 = x17 & ~n1370 ;
  assign n5880 = x17 & n1373 ;
  assign n5881 = ( ~n1467 & n5879 ) | ( ~n1467 & n5880 ) | ( n5879 & n5880 ) ;
  assign n5882 = ( n1487 & n5879 ) | ( n1487 & n5880 ) | ( n5879 & n5880 ) ;
  assign n5883 = ( ~n1358 & n5881 ) | ( ~n1358 & n5882 ) | ( n5881 & n5882 ) ;
  assign n5884 = ( n1506 & n5881 ) | ( n1506 & n5882 ) | ( n5881 & n5882 ) ;
  assign n5885 = ( n1612 & n5883 ) | ( n1612 & n5884 ) | ( n5883 & n5884 ) ;
  assign n5886 = n5878 | n5885 ;
  assign n5887 = x401 & n812 ;
  assign n5888 = x401 & ~n815 ;
  assign n5889 = ( n909 & n5887 ) | ( n909 & n5888 ) | ( n5887 & n5888 ) ;
  assign n5890 = ( ~n929 & n5887 ) | ( ~n929 & n5888 ) | ( n5887 & n5888 ) ;
  assign n5891 = ( n800 & n5889 ) | ( n800 & n5890 ) | ( n5889 & n5890 ) ;
  assign n5892 = ( ~n948 & n5889 ) | ( ~n948 & n5890 ) | ( n5889 & n5890 ) ;
  assign n5893 = ( ~n1061 & n5891 ) | ( ~n1061 & n5892 ) | ( n5891 & n5892 ) ;
  assign n5894 = x273 & ~n812 ;
  assign n5895 = x273 & n815 ;
  assign n5896 = ( ~n909 & n5894 ) | ( ~n909 & n5895 ) | ( n5894 & n5895 ) ;
  assign n5897 = ( n929 & n5894 ) | ( n929 & n5895 ) | ( n5894 & n5895 ) ;
  assign n5898 = ( ~n800 & n5896 ) | ( ~n800 & n5897 ) | ( n5896 & n5897 ) ;
  assign n5899 = ( n948 & n5896 ) | ( n948 & n5897 ) | ( n5896 & n5897 ) ;
  assign n5900 = ( n1061 & n5898 ) | ( n1061 & n5899 ) | ( n5898 & n5899 ) ;
  assign n5901 = n5893 | n5900 ;
  assign n5902 = ( n5871 & n5886 ) | ( n5871 & ~n5901 ) | ( n5886 & ~n5901 ) ;
  assign n5903 = ( ~n5309 & n5318 ) | ( ~n5309 & n5902 ) | ( n5318 & n5902 ) ;
  assign n5904 = n5287 & n5302 ;
  assign n5905 = ( n5285 & n5302 ) | ( n5285 & n5904 ) | ( n5302 & n5904 ) ;
  assign n5906 = ( n5302 & ~n5306 ) | ( n5302 & n5904 ) | ( ~n5306 & n5904 ) ;
  assign n5907 = ( n5317 & n5905 ) | ( n5317 & n5906 ) | ( n5905 & n5906 ) ;
  assign n5908 = ( n5286 & n5302 ) | ( n5286 & n5904 ) | ( n5302 & n5904 ) ;
  assign n5909 = ( ~n5204 & n5906 ) | ( ~n5204 & n5908 ) | ( n5906 & n5908 ) ;
  assign n5910 = ( n5902 & n5907 ) | ( n5902 & n5909 ) | ( n5907 & n5909 ) ;
  assign n5911 = n5903 | n5910 ;
  assign n5912 = x153 & n1370 ;
  assign n5913 = x153 & ~n1373 ;
  assign n5914 = ( n1467 & n5912 ) | ( n1467 & n5913 ) | ( n5912 & n5913 ) ;
  assign n5915 = ( ~n1487 & n5912 ) | ( ~n1487 & n5913 ) | ( n5912 & n5913 ) ;
  assign n5916 = ( n1358 & n5914 ) | ( n1358 & n5915 ) | ( n5914 & n5915 ) ;
  assign n5917 = ( ~n1506 & n5914 ) | ( ~n1506 & n5915 ) | ( n5914 & n5915 ) ;
  assign n5918 = ( ~n1612 & n5916 ) | ( ~n1612 & n5917 ) | ( n5916 & n5917 ) ;
  assign n5919 = x25 & ~n1370 ;
  assign n5920 = x25 & n1373 ;
  assign n5921 = ( ~n1467 & n5919 ) | ( ~n1467 & n5920 ) | ( n5919 & n5920 ) ;
  assign n5922 = ( n1487 & n5919 ) | ( n1487 & n5920 ) | ( n5919 & n5920 ) ;
  assign n5923 = ( ~n1358 & n5921 ) | ( ~n1358 & n5922 ) | ( n5921 & n5922 ) ;
  assign n5924 = ( n1506 & n5921 ) | ( n1506 & n5922 ) | ( n5921 & n5922 ) ;
  assign n5925 = ( n1612 & n5923 ) | ( n1612 & n5924 ) | ( n5923 & n5924 ) ;
  assign n5926 = n5918 | n5925 ;
  assign n5927 = x409 & n812 ;
  assign n5928 = x409 & ~n815 ;
  assign n5929 = ( n909 & n5927 ) | ( n909 & n5928 ) | ( n5927 & n5928 ) ;
  assign n5930 = ( ~n929 & n5927 ) | ( ~n929 & n5928 ) | ( n5927 & n5928 ) ;
  assign n5931 = ( n800 & n5929 ) | ( n800 & n5930 ) | ( n5929 & n5930 ) ;
  assign n5932 = ( ~n948 & n5929 ) | ( ~n948 & n5930 ) | ( n5929 & n5930 ) ;
  assign n5933 = ( ~n1061 & n5931 ) | ( ~n1061 & n5932 ) | ( n5931 & n5932 ) ;
  assign n5934 = x281 & ~n812 ;
  assign n5935 = x281 & n815 ;
  assign n5936 = ( ~n909 & n5934 ) | ( ~n909 & n5935 ) | ( n5934 & n5935 ) ;
  assign n5937 = ( n929 & n5934 ) | ( n929 & n5935 ) | ( n5934 & n5935 ) ;
  assign n5938 = ( ~n800 & n5936 ) | ( ~n800 & n5937 ) | ( n5936 & n5937 ) ;
  assign n5939 = ( n948 & n5936 ) | ( n948 & n5937 ) | ( n5936 & n5937 ) ;
  assign n5940 = ( n1061 & n5938 ) | ( n1061 & n5939 ) | ( n5938 & n5939 ) ;
  assign n5941 = n5933 | n5940 ;
  assign n5942 = ( n5911 & n5926 ) | ( n5911 & ~n5941 ) | ( n5926 & ~n5941 ) ;
  assign n5943 = ( n5061 & ~n5076 ) | ( n5061 & n5942 ) | ( ~n5076 & n5942 ) ;
  assign n5944 = ( n2380 & ~n2394 ) | ( n2380 & n5943 ) | ( ~n2394 & n5943 ) ;
  assign n5945 = n1070 & ~n5944 ;
  assign n5946 = n5805 & n5944 ;
  assign n5947 = n5945 | n5946 ;
  assign n5948 = ( ~n2380 & n2394 ) | ( ~n2380 & n5049 ) | ( n2394 & n5049 ) ;
  assign n5949 = ( n2380 & ~n2394 ) | ( n2380 & n5060 ) | ( ~n2394 & n5060 ) ;
  assign n5950 = ( n4266 & ~n5948 ) | ( n4266 & n5949 ) | ( ~n5948 & n5949 ) ;
  assign n5951 = ( n5075 & n5948 ) | ( n5075 & ~n5949 ) | ( n5948 & ~n5949 ) ;
  assign n5952 = ( n5942 & n5950 ) | ( n5942 & ~n5951 ) | ( n5950 & ~n5951 ) ;
  assign n5953 = n5790 & ~n5952 ;
  assign n5954 = n5821 & n5952 ;
  assign n5955 = n5953 | n5954 ;
  assign n5956 = n5775 & ~n5952 ;
  assign n5957 = n5760 & n5952 ;
  assign n5958 = n5956 | n5957 ;
  assign n5959 = n5745 & ~n5952 ;
  assign n5960 = n5730 & n5952 ;
  assign n5961 = n5959 | n5960 ;
  assign n5962 = n5715 & ~n5952 ;
  assign n5963 = n5700 & n5952 ;
  assign n5964 = n5962 | n5963 ;
  assign n5965 = n5685 & ~n5952 ;
  assign n5966 = n5670 & n5952 ;
  assign n5967 = n5965 | n5966 ;
  assign n5968 = n5655 & ~n5952 ;
  assign n5969 = n5640 & n5952 ;
  assign n5970 = n5968 | n5969 ;
  assign n5971 = n5605 & ~n5952 ;
  assign n5972 = n5590 & n5952 ;
  assign n5973 = n5971 | n5972 ;
  assign n5974 = n5575 & ~n5952 ;
  assign n5975 = n5621 & n5952 ;
  assign n5976 = n5974 | n5975 ;
  assign n5977 = n5861 & ~n5952 ;
  assign n5978 = n5846 & n5952 ;
  assign n5979 = n5977 | n5978 ;
  assign n5980 = n5441 & ~n5952 ;
  assign n5981 = n5426 & n5952 ;
  assign n5982 = n5980 | n5981 ;
  assign n5983 = n5411 & ~n5952 ;
  assign n5984 = n5396 & n5952 ;
  assign n5985 = n5983 | n5984 ;
  assign n5986 = n5379 & ~n5952 ;
  assign n5987 = n5364 & n5952 ;
  assign n5988 = n5986 | n5987 ;
  assign n5989 = n5348 & ~n5952 ;
  assign n5990 = n5333 & n5952 ;
  assign n5991 = n5989 | n5990 ;
  assign n5992 = n5522 & ~n5952 ;
  assign n5993 = n5507 & n5952 ;
  assign n5994 = n5992 | n5993 ;
  assign n5995 = n5491 & ~n5952 ;
  assign n5996 = n5476 & n5952 ;
  assign n5997 = n5995 | n5996 ;
  assign n5998 = n5461 & ~n5952 ;
  assign n5999 = n5544 & n5952 ;
  assign n6000 = n5998 | n5999 ;
  assign n6001 = n5901 & ~n5952 ;
  assign n6002 = n5886 & n5952 ;
  assign n6003 = n6001 | n6002 ;
  assign n6004 = n5199 & ~n5952 ;
  assign n6005 = n5184 & n5952 ;
  assign n6006 = n6004 | n6005 ;
  assign n6007 = n5169 & ~n5952 ;
  assign n6008 = n5154 & n5952 ;
  assign n6009 = n6007 | n6008 ;
  assign n6010 = n5137 & ~n5952 ;
  assign n6011 = n5122 & n5952 ;
  assign n6012 = n6010 | n6011 ;
  assign n6013 = n5106 & ~n5952 ;
  assign n6014 = n5091 & n5952 ;
  assign n6015 = n6013 | n6014 ;
  assign n6016 = n5280 & ~n5952 ;
  assign n6017 = n5265 & n5952 ;
  assign n6018 = n6016 | n6017 ;
  assign n6019 = n5249 & ~n5952 ;
  assign n6020 = n5234 & n5952 ;
  assign n6021 = n6019 | n6020 ;
  assign n6022 = n5219 & ~n5952 ;
  assign n6023 = n5302 & n5952 ;
  assign n6024 = n6022 | n6023 ;
  assign n6025 = n5941 & ~n5952 ;
  assign n6026 = n5926 & n5952 ;
  assign n6027 = n6025 | n6026 ;
  assign n6028 = n3338 & ~n5952 ;
  assign n6029 = n3323 & n5952 ;
  assign n6030 = n6028 | n6029 ;
  assign n6031 = n3306 & ~n5952 ;
  assign n6032 = n3291 & n5952 ;
  assign n6033 = n6031 | n6032 ;
  assign n6034 = n3275 & ~n5952 ;
  assign n6035 = n3260 & n5952 ;
  assign n6036 = n6034 | n6035 ;
  assign n6037 = n3373 & ~n5952 ;
  assign n6038 = n3358 & n5952 ;
  assign n6039 = n6037 | n6038 ;
  assign n6040 = n3243 & ~n5952 ;
  assign n6041 = n3228 & n5952 ;
  assign n6042 = n6040 | n6041 ;
  assign n6043 = n3211 & ~n5952 ;
  assign n6044 = n3196 & n5952 ;
  assign n6045 = n6043 | n6044 ;
  assign n6046 = n2941 & ~n5952 ;
  assign n6047 = n2956 & n5952 ;
  assign n6048 = n6046 | n6047 ;
  assign n6049 = n3114 & ~n5952 ;
  assign n6050 = n3099 & n5952 ;
  assign n6051 = n6049 | n6050 ;
  assign n6052 = n3161 & ~n5952 ;
  assign n6053 = n3176 & n5952 ;
  assign n6054 = n6052 | n6053 ;
  assign n6055 = n3145 & ~n5952 ;
  assign n6056 = n3130 & n5952 ;
  assign n6057 = n6055 | n6056 ;
  assign n6058 = n3050 & ~n5952 ;
  assign n6059 = n3035 & n5952 ;
  assign n6060 = n6058 | n6059 ;
  assign n6061 = n3081 & ~n5952 ;
  assign n6062 = n3066 & n5952 ;
  assign n6063 = n6061 | n6062 ;
  assign n6064 = n3003 & ~n5952 ;
  assign n6065 = n3018 & n5952 ;
  assign n6066 = n6064 | n6065 ;
  assign n6067 = n2987 & ~n5952 ;
  assign n6068 = n2972 & n5952 ;
  assign n6069 = n6067 | n6068 ;
  assign n6070 = n2915 & ~n5952 ;
  assign n6071 = n2900 & n5952 ;
  assign n6072 = n6070 | n6071 ;
  assign n6073 = n2885 & ~n5952 ;
  assign n6074 = n2870 & n5952 ;
  assign n6075 = n6073 | n6074 ;
  assign n6076 = n2855 & ~n5952 ;
  assign n6077 = n2840 & n5952 ;
  assign n6078 = n6076 | n6077 ;
  assign n6079 = n2825 & ~n5952 ;
  assign n6080 = n2810 & n5952 ;
  assign n6081 = n6079 | n6080 ;
  assign n6082 = n2761 & ~n5952 ;
  assign n6083 = n2746 & n5952 ;
  assign n6084 = n6082 | n6083 ;
  assign n6085 = n2792 & ~n5952 ;
  assign n6086 = n2777 & n5952 ;
  assign n6087 = n6085 | n6086 ;
  assign n6088 = n2714 & ~n5952 ;
  assign n6089 = n2729 & n5952 ;
  assign n6090 = n6088 | n6089 ;
  assign n6091 = n2691 & ~n5952 ;
  assign n6092 = n2676 & n5952 ;
  assign n6093 = n6091 | n6092 ;
  assign n6094 = n2633 & ~n5952 ;
  assign n6095 = n2648 & n5952 ;
  assign n6096 = n6094 | n6095 ;
  assign n6097 = n2551 & ~n5952 ;
  assign n6098 = n2536 & n5952 ;
  assign n6099 = n6097 | n6098 ;
  assign n6100 = n2598 & ~n5952 ;
  assign n6101 = n2613 & n5952 ;
  assign n6102 = n6100 | n6101 ;
  assign n6103 = n2582 & ~n5952 ;
  assign n6104 = n2567 & n5952 ;
  assign n6105 = n6103 | n6104 ;
  assign n6106 = n2503 & ~n5952 ;
  assign n6107 = n2518 & n5952 ;
  assign n6108 = n6106 | n6107 ;
  assign n6109 = n2487 & ~n5952 ;
  assign n6110 = n2472 & n5952 ;
  assign n6111 = n6109 | n6110 ;
  assign n6112 = n2440 & ~n5952 ;
  assign n6113 = n2455 & n5952 ;
  assign n6114 = n6112 | n6113 ;
  assign n6115 = n2424 & ~n5952 ;
  assign n6116 = n2409 & n5952 ;
  assign n6117 = n6115 | n6116 ;
  assign n6118 = n4224 & ~n5952 ;
  assign n6119 = n4209 & n5952 ;
  assign n6120 = n6118 | n6119 ;
  assign n6121 = n4194 & ~n5952 ;
  assign n6122 = n4179 & n5952 ;
  assign n6123 = n6121 | n6122 ;
  assign n6124 = n4164 & ~n5952 ;
  assign n6125 = n4149 & n5952 ;
  assign n6126 = n6124 | n6125 ;
  assign n6127 = n4134 & ~n5952 ;
  assign n6128 = n4119 & n5952 ;
  assign n6129 = n6127 | n6128 ;
  assign n6130 = n4101 & ~n5952 ;
  assign n6131 = n4086 & n5952 ;
  assign n6132 = n6130 | n6131 ;
  assign n6133 = n4070 & ~n5952 ;
  assign n6134 = n4055 & n5952 ;
  assign n6135 = n6133 | n6134 ;
  assign n6136 = n4023 & ~n5952 ;
  assign n6137 = n4038 & n5952 ;
  assign n6138 = n6136 | n6137 ;
  assign n6139 = n4007 & ~n5952 ;
  assign n6140 = n3992 & n5952 ;
  assign n6141 = n6139 | n6140 ;
  assign n6142 = n3681 & ~n5952 ;
  assign n6143 = n3696 & n5952 ;
  assign n6144 = n6142 | n6143 ;
  assign n6145 = n3665 & ~n5952 ;
  assign n6146 = n3650 & n5952 ;
  assign n6147 = n6145 | n6146 ;
  assign n6148 = n3618 & ~n5952 ;
  assign n6149 = n3633 & n5952 ;
  assign n6150 = n6148 | n6149 ;
  assign n6151 = n3602 & ~n5952 ;
  assign n6152 = n3587 & n5952 ;
  assign n6153 = n6151 | n6152 ;
  assign n6154 = n3569 & ~n5952 ;
  assign n6155 = n3554 & n5952 ;
  assign n6156 = n6154 | n6155 ;
  assign n6157 = n3538 & ~n5952 ;
  assign n6158 = n3523 & n5952 ;
  assign n6159 = n6157 | n6158 ;
  assign n6160 = n3489 & ~n5952 ;
  assign n6161 = n3504 & n5952 ;
  assign n6162 = n6160 | n6161 ;
  assign n6163 = n3473 & ~n5952 ;
  assign n6164 = n3458 & n5952 ;
  assign n6165 = n6163 | n6164 ;
  assign n6166 = n3942 & ~n5952 ;
  assign n6167 = n3957 & n5952 ;
  assign n6168 = n6166 | n6167 ;
  assign n6169 = n3926 & ~n5952 ;
  assign n6170 = n3911 & n5952 ;
  assign n6171 = n6169 | n6170 ;
  assign n6172 = n3879 & ~n5952 ;
  assign n6173 = n3894 & n5952 ;
  assign n6174 = n6172 | n6173 ;
  assign n6175 = n3863 & ~n5952 ;
  assign n6176 = n3848 & n5952 ;
  assign n6177 = n6175 | n6176 ;
  assign n6178 = n3830 & ~n5952 ;
  assign n6179 = n3815 & n5952 ;
  assign n6180 = n6178 | n6179 ;
  assign n6181 = n3799 & ~n5952 ;
  assign n6182 = n3784 & n5952 ;
  assign n6183 = n6181 | n6182 ;
  assign n6184 = n3752 & ~n5952 ;
  assign n6185 = n3767 & n5952 ;
  assign n6186 = n6184 | n6185 ;
  assign n6187 = n3736 & ~n5952 ;
  assign n6188 = n3721 & n5952 ;
  assign n6189 = n6187 | n6188 ;
  assign n6190 = n4874 & ~n5952 ;
  assign n6191 = n4889 & n5952 ;
  assign n6192 = n6190 | n6191 ;
  assign n6193 = n3442 & ~n5952 ;
  assign n6194 = n3427 & n5952 ;
  assign n6195 = n6193 | n6194 ;
  assign n6196 = n4842 & ~n5952 ;
  assign n6197 = n4857 & n5952 ;
  assign n6198 = n6196 | n6197 ;
  assign n6199 = n4826 & ~n5952 ;
  assign n6200 = n4811 & n5952 ;
  assign n6201 = n6199 | n6200 ;
  assign n6202 = n4793 & ~n5952 ;
  assign n6203 = n4778 & n5952 ;
  assign n6204 = n6202 | n6203 ;
  assign n6205 = n4762 & ~n5952 ;
  assign n6206 = n4747 & n5952 ;
  assign n6207 = n6205 | n6206 ;
  assign n6208 = n4715 & ~n5952 ;
  assign n6209 = n4730 & n5952 ;
  assign n6210 = n6208 | n6209 ;
  assign n6211 = n4699 & ~n5952 ;
  assign n6212 = n4684 & n5952 ;
  assign n6213 = n6211 | n6212 ;
  assign n6214 = n5015 & ~n5952 ;
  assign n6215 = n5030 & n5952 ;
  assign n6216 = n6214 | n6215 ;
  assign n6217 = n5000 & ~n5952 ;
  assign n6218 = n4985 & n5952 ;
  assign n6219 = n6217 | n6218 ;
  assign n6220 = n4955 & ~n5952 ;
  assign n6221 = n4970 & n5952 ;
  assign n6222 = n6220 | n6221 ;
  assign n6223 = n4940 & ~n5952 ;
  assign n6224 = n4925 & n5952 ;
  assign n6225 = n6223 | n6224 ;
  assign n6226 = n4655 & ~n5952 ;
  assign n6227 = n4640 & n5952 ;
  assign n6228 = n6226 | n6227 ;
  assign n6229 = n4625 & ~n5952 ;
  assign n6230 = n4610 & n5952 ;
  assign n6231 = n6229 | n6230 ;
  assign n6232 = n4580 & ~n5952 ;
  assign n6233 = n4595 & n5952 ;
  assign n6234 = n6232 | n6233 ;
  assign n6235 = n4565 & ~n5952 ;
  assign n6236 = n4550 & n5952 ;
  assign n6237 = n6235 | n6236 ;
  assign n6238 = n4513 & ~n5952 ;
  assign n6239 = n4528 & n5952 ;
  assign n6240 = n6238 | n6239 ;
  assign n6241 = n4498 & ~n5952 ;
  assign n6242 = n4483 & n5952 ;
  assign n6243 = n6241 | n6242 ;
  assign n6244 = n4453 & ~n5952 ;
  assign n6245 = n4468 & n5952 ;
  assign n6246 = n6244 | n6245 ;
  assign n6247 = n4438 & ~n5952 ;
  assign n6248 = n4423 & n5952 ;
  assign n6249 = n6247 | n6248 ;
  assign n6250 = n4398 & ~n5952 ;
  assign n6251 = n4383 & n5952 ;
  assign n6252 = n6250 | n6251 ;
  assign n6253 = n4368 & ~n5952 ;
  assign n6254 = n4353 & n5952 ;
  assign n6255 = n6253 | n6254 ;
  assign n6256 = n4321 & ~n5952 ;
  assign n6257 = n4336 & n5952 ;
  assign n6258 = n6256 | n6257 ;
  assign n6259 = n4303 & ~n5952 ;
  assign n6260 = n4288 & n5952 ;
  assign n6261 = n6259 | n6260 ;
  assign n6262 = n1841 & ~n5952 ;
  assign n6263 = n1856 & n5952 ;
  assign n6264 = n6262 | n6263 ;
  assign n6265 = n1826 & ~n5952 ;
  assign n6266 = n1811 & n5952 ;
  assign n6267 = n6265 | n6266 ;
  assign n6268 = n1781 & ~n5952 ;
  assign n6269 = n1796 & n5952 ;
  assign n6270 = n6268 | n6269 ;
  assign n6271 = n1766 & ~n5952 ;
  assign n6272 = n1751 & n5952 ;
  assign n6273 = n6271 | n6272 ;
  assign n6274 = n1732 & ~n5952 ;
  assign n6275 = n1717 & n5952 ;
  assign n6276 = n6274 | n6275 ;
  assign n6277 = n1701 & ~n5952 ;
  assign n6278 = n1686 & n5952 ;
  assign n6279 = n6277 | n6278 ;
  assign n6280 = n1652 & ~n5952 ;
  assign n6281 = n1667 & n5952 ;
  assign n6282 = n6280 | n6281 ;
  assign n6283 = n1636 & ~n5952 ;
  assign n6284 = n1621 & n5952 ;
  assign n6285 = n6283 | n6284 ;
  assign n6286 = n2230 & ~n5952 ;
  assign n6287 = n2245 & n5952 ;
  assign n6288 = n6286 | n6287 ;
  assign n6289 = n2214 & ~n5952 ;
  assign n6290 = n2199 & n5952 ;
  assign n6291 = n6289 | n6290 ;
  assign n6292 = n2167 & ~n5952 ;
  assign n6293 = n2182 & n5952 ;
  assign n6294 = n6292 | n6293 ;
  assign n6295 = n2151 & ~n5952 ;
  assign n6296 = n2136 & n5952 ;
  assign n6297 = n6295 | n6296 ;
  assign n6298 = n2118 & ~n5952 ;
  assign n6299 = n2103 & n5952 ;
  assign n6300 = n6298 | n6299 ;
  assign n6301 = n2087 & ~n5952 ;
  assign n6302 = n2072 & n5952 ;
  assign n6303 = n6301 | n6302 ;
  assign n6304 = n2040 & ~n5952 ;
  assign n6305 = n2055 & n5952 ;
  assign n6306 = n6304 | n6305 ;
  assign n6307 = n2024 & ~n5952 ;
  assign n6308 = n2009 & n5952 ;
  assign n6309 = n6307 | n6308 ;
  assign n6310 = n1976 & ~n5952 ;
  assign n6311 = n1991 & n5952 ;
  assign n6312 = n6310 | n6311 ;
  assign n6313 = n1960 & ~n5952 ;
  assign n6314 = n1945 & n5952 ;
  assign n6315 = n6313 | n6314 ;
  assign n6316 = n1913 & ~n5952 ;
  assign n6317 = n1928 & n5952 ;
  assign n6318 = n6316 | n6317 ;
  assign n6319 = n1897 & ~n5952 ;
  assign n6320 = n1882 & n5952 ;
  assign n6321 = n6319 | n6320 ;
  assign n6322 = n2360 & ~n5952 ;
  assign n6323 = n2345 & n5952 ;
  assign n6324 = n6322 | n6323 ;
  assign n6325 = n2328 & ~n5952 ;
  assign n6326 = n2313 & n5952 ;
  assign n6327 = n6325 | n6326 ;
  assign n6328 = n2297 & ~n5952 ;
  assign n6329 = n2282 & n5952 ;
  assign n6330 = n6328 | n6329 ;
  assign n6331 = n2371 | n2376 ;
  assign n6332 = n2366 & ~n2376 ;
  assign n6333 = ( n2267 & n6331 ) | ( n2267 & ~n6332 ) | ( n6331 & ~n6332 ) ;
  assign n6334 = ( n2383 & n2393 ) | ( n2383 & ~n6331 ) | ( n2393 & ~n6331 ) ;
  assign n6335 = ( n5076 & ~n6333 ) | ( n5076 & n6334 ) | ( ~n6333 & n6334 ) ;
  assign n6336 = ( n5061 & n6333 ) | ( n5061 & ~n6334 ) | ( n6333 & ~n6334 ) ;
  assign n6337 = ( n5942 & ~n6335 ) | ( n5942 & n6336 ) | ( ~n6335 & n6336 ) ;
  assign n6338 = n2362 | n6337 ;
  assign n6339 = n2363 & n6338 ;
  assign n6340 = ( n800 & n909 ) | ( n800 & ~n929 ) | ( n909 & ~n929 ) ;
  assign n6341 = ( n812 & ~n815 ) | ( n812 & n6340 ) | ( ~n815 & n6340 ) ;
  assign n6342 = ( ~n909 & n929 ) | ( ~n909 & n948 ) | ( n929 & n948 ) ;
  assign n6343 = ( ~n812 & n815 ) | ( ~n812 & n6342 ) | ( n815 & n6342 ) ;
  assign n6344 = ( n1061 & ~n6341 ) | ( n1061 & n6343 ) | ( ~n6341 & n6343 ) ;
  assign n6345 = n5952 | n6344 ;
  assign n6346 = ( n1358 & n1467 ) | ( n1358 & ~n1487 ) | ( n1467 & ~n1487 ) ;
  assign n6347 = ( n1370 & ~n1373 ) | ( n1370 & n6346 ) | ( ~n1373 & n6346 ) ;
  assign n6348 = ( ~n1467 & n1487 ) | ( ~n1467 & n1506 ) | ( n1487 & n1506 ) ;
  assign n6349 = ( ~n1370 & n1373 ) | ( ~n1370 & n6348 ) | ( n1373 & n6348 ) ;
  assign n6350 = ( n1612 & ~n6347 ) | ( n1612 & n6349 ) | ( ~n6347 & n6349 ) ;
  assign n6351 = n5952 & ~n6350 ;
  assign n6352 = n6345 & ~n6351 ;
  assign y0 = n5947 ;
  assign y1 = n5955 ;
  assign y2 = n5958 ;
  assign y3 = n5961 ;
  assign y4 = n5964 ;
  assign y5 = n5967 ;
  assign y6 = n5970 ;
  assign y7 = n5973 ;
  assign y8 = n5976 ;
  assign y9 = n5979 ;
  assign y10 = n5982 ;
  assign y11 = n5985 ;
  assign y12 = n5988 ;
  assign y13 = n5991 ;
  assign y14 = n5994 ;
  assign y15 = n5997 ;
  assign y16 = n6000 ;
  assign y17 = n6003 ;
  assign y18 = n6006 ;
  assign y19 = n6009 ;
  assign y20 = n6012 ;
  assign y21 = n6015 ;
  assign y22 = n6018 ;
  assign y23 = n6021 ;
  assign y24 = n6024 ;
  assign y25 = n6027 ;
  assign y26 = n6030 ;
  assign y27 = n6033 ;
  assign y28 = n6036 ;
  assign y29 = n6039 ;
  assign y30 = n6042 ;
  assign y31 = n6045 ;
  assign y32 = n6048 ;
  assign y33 = n6051 ;
  assign y34 = n6054 ;
  assign y35 = n6057 ;
  assign y36 = n6060 ;
  assign y37 = n6063 ;
  assign y38 = n6066 ;
  assign y39 = n6069 ;
  assign y40 = n6072 ;
  assign y41 = n6075 ;
  assign y42 = n6078 ;
  assign y43 = n6081 ;
  assign y44 = n6084 ;
  assign y45 = n6087 ;
  assign y46 = n6090 ;
  assign y47 = n6093 ;
  assign y48 = n6096 ;
  assign y49 = n6099 ;
  assign y50 = n6102 ;
  assign y51 = n6105 ;
  assign y52 = n6108 ;
  assign y53 = n6111 ;
  assign y54 = n6114 ;
  assign y55 = n6117 ;
  assign y56 = n6120 ;
  assign y57 = n6123 ;
  assign y58 = n6126 ;
  assign y59 = n6129 ;
  assign y60 = n6132 ;
  assign y61 = n6135 ;
  assign y62 = n6138 ;
  assign y63 = n6141 ;
  assign y64 = n6144 ;
  assign y65 = n6147 ;
  assign y66 = n6150 ;
  assign y67 = n6153 ;
  assign y68 = n6156 ;
  assign y69 = n6159 ;
  assign y70 = n6162 ;
  assign y71 = n6165 ;
  assign y72 = n6168 ;
  assign y73 = n6171 ;
  assign y74 = n6174 ;
  assign y75 = n6177 ;
  assign y76 = n6180 ;
  assign y77 = n6183 ;
  assign y78 = n6186 ;
  assign y79 = n6189 ;
  assign y80 = n6192 ;
  assign y81 = n6195 ;
  assign y82 = n6198 ;
  assign y83 = n6201 ;
  assign y84 = n6204 ;
  assign y85 = n6207 ;
  assign y86 = n6210 ;
  assign y87 = n6213 ;
  assign y88 = n6216 ;
  assign y89 = n6219 ;
  assign y90 = n6222 ;
  assign y91 = n6225 ;
  assign y92 = n6228 ;
  assign y93 = n6231 ;
  assign y94 = n6234 ;
  assign y95 = n6237 ;
  assign y96 = n6240 ;
  assign y97 = n6243 ;
  assign y98 = n6246 ;
  assign y99 = n6249 ;
  assign y100 = n6252 ;
  assign y101 = n6255 ;
  assign y102 = n6258 ;
  assign y103 = n6261 ;
  assign y104 = n6264 ;
  assign y105 = n6267 ;
  assign y106 = n6270 ;
  assign y107 = n6273 ;
  assign y108 = n6276 ;
  assign y109 = n6279 ;
  assign y110 = n6282 ;
  assign y111 = n6285 ;
  assign y112 = n6288 ;
  assign y113 = n6291 ;
  assign y114 = n6294 ;
  assign y115 = n6297 ;
  assign y116 = n6300 ;
  assign y117 = n6303 ;
  assign y118 = n6306 ;
  assign y119 = n6309 ;
  assign y120 = n6312 ;
  assign y121 = n6315 ;
  assign y122 = n6318 ;
  assign y123 = n6321 ;
  assign y124 = n6324 ;
  assign y125 = n6327 ;
  assign y126 = n6330 ;
  assign y127 = n6339 ;
  assign y128 = ~n6352 ;
  assign y129 = ~n5952 ;
endmodule
