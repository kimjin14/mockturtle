module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 ;
  assign n33 = x29 | x30 ;
  assign n34 = ~x27 & x28 ;
  assign n35 = ~n33 & n34 ;
  assign n36 = x24 | x25 ;
  assign n37 = x23 | x26 ;
  assign n38 = n36 | n37 ;
  assign n39 = n35 & ~n38 ;
  assign n40 = ~x24 & x25 ;
  assign n41 = ~x23 & x26 ;
  assign n42 = n40 & n41 ;
  assign n43 = x27 | x28 ;
  assign n44 = x29 & x30 ;
  assign n45 = ~n43 & n44 ;
  assign n46 = n42 & n45 ;
  assign n47 = ~x29 & x30 ;
  assign n48 = x27 & x28 ;
  assign n49 = n47 & n48 ;
  assign n50 = x24 & ~x25 ;
  assign n51 = x23 & x26 ;
  assign n52 = n50 & n51 ;
  assign n53 = n49 & n52 ;
  assign n54 = n46 | n53 ;
  assign n55 = n39 | n54 ;
  assign n56 = x23 & ~x26 ;
  assign n57 = n50 & n56 ;
  assign n58 = n33 | n43 ;
  assign n59 = n57 & ~n58 ;
  assign n60 = x27 & ~x28 ;
  assign n61 = n44 & n60 ;
  assign n62 = x24 & x25 ;
  assign n63 = n51 & n62 ;
  assign n64 = n61 & n63 ;
  assign n65 = n34 & n44 ;
  assign n66 = ~n36 & n56 ;
  assign n67 = n65 & n66 ;
  assign n68 = n64 | n67 ;
  assign n69 = n59 | n68 ;
  assign n70 = n55 | n69 ;
  assign n71 = n52 & ~n58 ;
  assign n72 = x29 & ~x30 ;
  assign n73 = ~n43 & n72 ;
  assign n74 = n40 & n51 ;
  assign n75 = n73 & n74 ;
  assign n76 = n71 | n75 ;
  assign n77 = n45 & n63 ;
  assign n78 = n56 & n62 ;
  assign n79 = n45 & n78 ;
  assign n80 = n77 | n79 ;
  assign n81 = n76 | n80 ;
  assign n82 = n70 | n81 ;
  assign n83 = n65 & n78 ;
  assign n84 = ~n43 & n47 ;
  assign n85 = ~n38 & n84 ;
  assign n86 = ~n37 & n50 ;
  assign n87 = n47 & n60 ;
  assign n88 = n86 & n87 ;
  assign n89 = n85 | n88 ;
  assign n90 = n83 | n89 ;
  assign n91 = ~n37 & n40 ;
  assign n92 = n45 & n91 ;
  assign n93 = n41 & n62 ;
  assign n94 = n87 & n93 ;
  assign n95 = n92 | n94 ;
  assign n96 = n35 & n86 ;
  assign n97 = n40 & n56 ;
  assign n98 = ~n33 & n48 ;
  assign n99 = n97 & n98 ;
  assign n100 = n96 | n99 ;
  assign n101 = n95 | n100 ;
  assign n102 = n60 & n72 ;
  assign n103 = n97 & n102 ;
  assign n104 = n42 & n102 ;
  assign n105 = n103 | n104 ;
  assign n106 = n101 | n105 ;
  assign n107 = n90 | n106 ;
  assign n108 = n82 | n107 ;
  assign n109 = n48 & n72 ;
  assign n110 = n86 & n109 ;
  assign n111 = ~n37 & n62 ;
  assign n112 = n49 & n111 ;
  assign n113 = n34 & n47 ;
  assign n114 = n93 & n113 ;
  assign n115 = n112 | n114 ;
  assign n116 = n41 & n50 ;
  assign n117 = n84 & n116 ;
  assign n118 = n35 & n57 ;
  assign n119 = n117 | n118 ;
  assign n120 = n115 | n119 ;
  assign n121 = n110 | n120 ;
  assign n122 = ~n33 & n60 ;
  assign n123 = n86 & n122 ;
  assign n124 = n49 & n78 ;
  assign n125 = n123 | n124 ;
  assign n126 = ~n38 & n73 ;
  assign n127 = ~n36 & n41 ;
  assign n128 = n45 & n127 ;
  assign n129 = n126 | n128 ;
  assign n130 = n125 | n129 ;
  assign n131 = n98 & n127 ;
  assign n132 = n44 & n48 ;
  assign n133 = n111 & n132 ;
  assign n134 = n52 & n132 ;
  assign n135 = n133 | n134 ;
  assign n136 = n131 | n135 ;
  assign n137 = n130 | n136 ;
  assign n138 = n97 & n113 ;
  assign n139 = n66 & n98 ;
  assign n140 = n138 | n139 ;
  assign n141 = n35 & n78 ;
  assign n142 = n98 & n116 ;
  assign n143 = n38 | n58 ;
  assign n144 = ~n142 & n143 ;
  assign n145 = ~n141 & n144 ;
  assign n146 = ~n140 & n145 ;
  assign n147 = ~n137 & n146 ;
  assign n148 = ~n121 & n147 ;
  assign n149 = ~n108 & n148 ;
  assign n150 = n34 & n72 ;
  assign n151 = n57 & n150 ;
  assign n152 = n65 & n91 ;
  assign n153 = n151 | n152 ;
  assign n154 = n91 & n109 ;
  assign n155 = n93 & n102 ;
  assign n156 = n154 | n155 ;
  assign n157 = n153 | n156 ;
  assign n158 = ~n36 & n51 ;
  assign n159 = n150 & n158 ;
  assign n160 = n63 & n122 ;
  assign n161 = n159 | n160 ;
  assign n162 = n87 & n97 ;
  assign n163 = n65 & n111 ;
  assign n164 = n162 | n163 ;
  assign n165 = n161 | n164 ;
  assign n166 = n157 | n165 ;
  assign n167 = n84 & n127 ;
  assign n168 = n49 & n97 ;
  assign n169 = n167 | n168 ;
  assign n170 = ~n38 & n87 ;
  assign n171 = n63 & n65 ;
  assign n172 = n170 | n171 ;
  assign n173 = n169 | n172 ;
  assign n174 = n166 | n173 ;
  assign n175 = n78 & n84 ;
  assign n176 = n87 & n91 ;
  assign n177 = n175 | n176 ;
  assign n178 = n84 & n86 ;
  assign n179 = n52 & n84 ;
  assign n180 = n178 | n179 ;
  assign n181 = n177 | n180 ;
  assign n182 = n74 & n109 ;
  assign n183 = n63 & n132 ;
  assign n184 = n73 & n91 ;
  assign n185 = n183 | n184 ;
  assign n186 = n182 | n185 ;
  assign n187 = n181 | n186 ;
  assign n188 = n174 | n187 ;
  assign n189 = n45 & n52 ;
  assign n190 = n61 & n111 ;
  assign n191 = n189 | n190 ;
  assign n192 = n98 & n111 ;
  assign n193 = n116 & n132 ;
  assign n194 = n192 | n193 ;
  assign n195 = n191 | n194 ;
  assign n196 = n74 & n150 ;
  assign n197 = n57 & n102 ;
  assign n198 = n97 & n150 ;
  assign n199 = n197 | n198 ;
  assign n200 = n196 | n199 ;
  assign n201 = n195 | n200 ;
  assign n202 = n49 & n158 ;
  assign n203 = n35 & n63 ;
  assign n204 = n202 | n203 ;
  assign n205 = n87 & n127 ;
  assign n206 = n111 & n122 ;
  assign n207 = n205 | n206 ;
  assign n208 = n63 & n98 ;
  assign n209 = n49 & n74 ;
  assign n210 = n208 | n209 ;
  assign n211 = n207 | n210 ;
  assign n212 = n86 & n150 ;
  assign n213 = n45 & n158 ;
  assign n214 = n61 & n66 ;
  assign n215 = n213 | n214 ;
  assign n216 = n212 | n215 ;
  assign n217 = n211 | n216 ;
  assign n218 = n204 | n217 ;
  assign n219 = n201 | n218 ;
  assign n220 = n188 | n219 ;
  assign n221 = n149 & ~n220 ;
  assign n222 = n45 & n66 ;
  assign n223 = ~n58 & n111 ;
  assign n224 = n222 | n223 ;
  assign n225 = n73 & n86 ;
  assign n226 = n74 & n122 ;
  assign n227 = n225 | n226 ;
  assign n228 = n63 & n113 ;
  assign n229 = n97 & n109 ;
  assign n230 = n228 | n229 ;
  assign n231 = n227 | n230 ;
  assign n232 = n224 | n231 ;
  assign n233 = n84 & n93 ;
  assign n234 = n91 & n102 ;
  assign n235 = n233 | n234 ;
  assign n236 = n65 & n158 ;
  assign n237 = n74 & n132 ;
  assign n238 = n236 | n237 ;
  assign n239 = n78 & n132 ;
  assign n240 = n35 & n91 ;
  assign n241 = n239 | n240 ;
  assign n242 = n238 | n241 ;
  assign n243 = n235 | n242 ;
  assign n244 = n232 | n243 ;
  assign n245 = ~n38 & n109 ;
  assign n246 = n78 & n113 ;
  assign n247 = n57 & n65 ;
  assign n248 = n246 | n247 ;
  assign n249 = ~n38 & n45 ;
  assign n250 = n66 & n150 ;
  assign n251 = n249 | n250 ;
  assign n252 = n248 | n251 ;
  assign n253 = n245 | n252 ;
  assign n254 = n73 & n111 ;
  assign n255 = n122 & n158 ;
  assign n256 = n254 | n255 ;
  assign n257 = n42 & n65 ;
  assign n258 = n66 & n84 ;
  assign n259 = n257 | n258 ;
  assign n260 = n256 | n259 ;
  assign n261 = n42 & n113 ;
  assign n262 = n97 & n122 ;
  assign n263 = n73 & n93 ;
  assign n264 = n262 | n263 ;
  assign n265 = n261 | n264 ;
  assign n266 = n260 | n265 ;
  assign n267 = n253 | n266 ;
  assign n268 = n244 | n267 ;
  assign n269 = n42 & n122 ;
  assign n270 = n116 & n122 ;
  assign n271 = n269 | n270 ;
  assign n272 = n93 & n98 ;
  assign n273 = n66 & n73 ;
  assign n274 = n272 | n273 ;
  assign n275 = n271 | n274 ;
  assign n276 = n268 | n275 ;
  assign n277 = n35 & n111 ;
  assign n278 = n78 & n98 ;
  assign n279 = n277 | n278 ;
  assign n280 = n52 & n102 ;
  assign n281 = n102 & n111 ;
  assign n282 = n280 | n281 ;
  assign n283 = n74 & n102 ;
  assign n284 = n65 & n93 ;
  assign n285 = n283 | n284 ;
  assign n286 = n282 | n285 ;
  assign n287 = n279 | n286 ;
  assign n288 = n57 & n84 ;
  assign n289 = n52 & n113 ;
  assign n290 = n288 | n289 ;
  assign n291 = n57 & n61 ;
  assign n292 = n49 & n116 ;
  assign n293 = n291 | n292 ;
  assign n294 = n290 | n293 ;
  assign n295 = n35 & n93 ;
  assign n296 = n42 & n84 ;
  assign n297 = n57 & n122 ;
  assign n298 = n296 | n297 ;
  assign n299 = n295 | n298 ;
  assign n300 = n294 | n299 ;
  assign n301 = n287 | n300 ;
  assign n302 = n35 & n74 ;
  assign n303 = ~n58 & n97 ;
  assign n304 = n302 | n303 ;
  assign n305 = n78 & n102 ;
  assign n306 = n57 & n98 ;
  assign n307 = n305 | n306 ;
  assign n308 = n304 | n307 ;
  assign n309 = ~n58 & n63 ;
  assign n310 = n91 & n122 ;
  assign n311 = n309 | n310 ;
  assign n312 = n102 & n158 ;
  assign n313 = n61 & n158 ;
  assign n314 = n312 | n313 ;
  assign n315 = n311 | n314 ;
  assign n316 = n308 | n315 ;
  assign n317 = n113 & n158 ;
  assign n318 = n74 & n84 ;
  assign n319 = n317 | n318 ;
  assign n320 = n61 & n78 ;
  assign n321 = n61 & n127 ;
  assign n322 = n320 | n321 ;
  assign n323 = n319 | n322 ;
  assign n324 = n63 & n150 ;
  assign n325 = ~n58 & n66 ;
  assign n326 = n324 | n325 ;
  assign n327 = n323 | n326 ;
  assign n328 = n316 | n327 ;
  assign n329 = n301 | n328 ;
  assign n330 = n45 & n93 ;
  assign n331 = n74 & n87 ;
  assign n332 = n57 & n109 ;
  assign n333 = n73 & n116 ;
  assign n334 = n332 | n333 ;
  assign n335 = n331 | n334 ;
  assign n336 = n330 | n335 ;
  assign n337 = n329 | n336 ;
  assign n338 = n276 | n337 ;
  assign n339 = n221 & ~n338 ;
  assign n340 = n61 & n97 ;
  assign n341 = n45 & n86 ;
  assign n342 = n340 | n341 ;
  assign n343 = ~n38 & n122 ;
  assign n344 = n93 & n122 ;
  assign n345 = n343 | n344 ;
  assign n346 = n342 | n345 ;
  assign n347 = n63 & n73 ;
  assign n348 = n42 & n150 ;
  assign n349 = ~n58 & n74 ;
  assign n350 = n348 | n349 ;
  assign n351 = n347 | n350 ;
  assign n352 = n346 | n351 ;
  assign n353 = n339 & ~n352 ;
  assign n354 = n109 & n116 ;
  assign n355 = n97 & n132 ;
  assign n356 = n66 & n122 ;
  assign n357 = n355 | n356 ;
  assign n358 = n110 | n357 ;
  assign n359 = n120 | n358 ;
  assign n360 = n354 | n359 ;
  assign n361 = n147 & ~n360 ;
  assign n362 = ~n108 & n361 ;
  assign n363 = n102 & n127 ;
  assign n364 = n111 & n113 ;
  assign n365 = n363 | n364 ;
  assign n366 = n255 | n349 ;
  assign n367 = n365 | n366 ;
  assign n368 = n197 | n367 ;
  assign n369 = n61 & n116 ;
  assign n370 = n42 & n61 ;
  assign n371 = n369 | n370 ;
  assign n372 = n35 & n52 ;
  assign n373 = n214 | n372 ;
  assign n374 = n73 & n127 ;
  assign n375 = n109 & n111 ;
  assign n376 = n374 | n375 ;
  assign n377 = n373 | n376 ;
  assign n378 = n371 | n377 ;
  assign n379 = n368 | n378 ;
  assign n380 = n362 & ~n379 ;
  assign n381 = ~n58 & n158 ;
  assign n382 = n325 | n381 ;
  assign n383 = n61 & n86 ;
  assign n384 = n57 & n87 ;
  assign n385 = n313 | n384 ;
  assign n386 = n383 | n385 ;
  assign n387 = n63 & n87 ;
  assign n388 = n45 & n116 ;
  assign n389 = n387 | n388 ;
  assign n390 = n93 & n109 ;
  assign n391 = n343 | n390 ;
  assign n392 = n389 | n391 ;
  assign n393 = n386 | n392 ;
  assign n394 = n193 | n228 ;
  assign n395 = ~n58 & n116 ;
  assign n396 = n305 | n395 ;
  assign n397 = n394 | n396 ;
  assign n398 = n393 | n397 ;
  assign n399 = n49 & n93 ;
  assign n400 = n331 | n399 ;
  assign n401 = n74 & n98 ;
  assign n402 = n57 & n132 ;
  assign n403 = n401 | n402 ;
  assign n404 = n400 | n403 ;
  assign n405 = n73 & n97 ;
  assign n406 = n91 & n113 ;
  assign n407 = n405 | n406 ;
  assign n408 = n295 | n407 ;
  assign n409 = n404 | n408 ;
  assign n410 = n398 | n409 ;
  assign n411 = n203 | n297 ;
  assign n412 = ~n38 & n49 ;
  assign n413 = n57 & n73 ;
  assign n414 = n412 | n413 ;
  assign n415 = n411 | n414 ;
  assign n416 = ~n38 & n132 ;
  assign n417 = n292 | n416 ;
  assign n418 = n42 & n87 ;
  assign n419 = n283 | n418 ;
  assign n420 = n417 | n419 ;
  assign n421 = n415 | n420 ;
  assign n422 = n257 | n421 ;
  assign n423 = n302 | n310 ;
  assign n424 = n111 & n150 ;
  assign n425 = n225 | n424 ;
  assign n426 = n423 | n425 ;
  assign n427 = n422 | n426 ;
  assign n428 = n410 | n427 ;
  assign n429 = n382 | n428 ;
  assign n430 = n380 & ~n429 ;
  assign n431 = n52 & n150 ;
  assign n432 = n91 & n98 ;
  assign n433 = n306 | n432 ;
  assign n434 = ~n58 & n93 ;
  assign n435 = n42 & n98 ;
  assign n436 = n434 | n435 ;
  assign n437 = n91 & n150 ;
  assign n438 = n167 | n437 ;
  assign n439 = n436 | n438 ;
  assign n440 = n433 | n439 ;
  assign n441 = n84 & n158 ;
  assign n442 = n296 | n441 ;
  assign n443 = n73 & n158 ;
  assign n444 = n132 & n158 ;
  assign n445 = n443 | n444 ;
  assign n446 = n442 | n445 ;
  assign n447 = ~n38 & n98 ;
  assign n448 = n127 & n150 ;
  assign n449 = n447 | n448 ;
  assign n450 = n65 & n86 ;
  assign n451 = n84 & n111 ;
  assign n452 = n450 | n451 ;
  assign n453 = n449 | n452 ;
  assign n454 = n446 | n453 ;
  assign n455 = n440 | n454 ;
  assign n456 = n45 & n97 ;
  assign n457 = n42 & n49 ;
  assign n458 = n66 & n87 ;
  assign n459 = n457 | n458 ;
  assign n460 = n86 & n113 ;
  assign n461 = n87 & n158 ;
  assign n462 = n460 | n461 ;
  assign n463 = n459 | n462 ;
  assign n464 = n456 | n463 ;
  assign n465 = n93 & n132 ;
  assign n466 = n320 | n341 ;
  assign n467 = n465 | n466 ;
  assign n468 = n66 & n102 ;
  assign n469 = ~n58 & n86 ;
  assign n470 = n281 | n469 ;
  assign n471 = n468 | n470 ;
  assign n472 = n467 | n471 ;
  assign n473 = n464 | n472 ;
  assign n474 = n455 | n473 ;
  assign n475 = n431 | n474 ;
  assign n476 = ~n58 & n127 ;
  assign n477 = n65 & n97 ;
  assign n478 = n476 | n477 ;
  assign n479 = n49 & n86 ;
  assign n480 = n84 & n91 ;
  assign n481 = n479 | n480 ;
  assign n482 = n478 | n481 ;
  assign n483 = n57 & n113 ;
  assign n484 = n237 | n483 ;
  assign n485 = n179 | n484 ;
  assign n486 = n482 | n485 ;
  assign n487 = n52 & n109 ;
  assign n488 = n154 | n487 ;
  assign n489 = n122 & n127 ;
  assign n490 = n247 | n489 ;
  assign n491 = n86 & n98 ;
  assign n492 = n223 | n491 ;
  assign n493 = n490 | n492 ;
  assign n494 = n488 | n493 ;
  assign n495 = n486 | n494 ;
  assign n496 = n240 | n277 ;
  assign n497 = ~n58 & n78 ;
  assign n498 = n312 | n497 ;
  assign n499 = n496 | n498 ;
  assign n500 = n66 & n109 ;
  assign n501 = n35 & n66 ;
  assign n502 = n500 | n501 ;
  assign n503 = n49 & n66 ;
  assign n504 = n171 | n503 ;
  assign n505 = n502 | n504 ;
  assign n506 = n499 | n505 ;
  assign n507 = n495 | n506 ;
  assign n508 = n178 | n507 ;
  assign n509 = n475 | n508 ;
  assign n510 = n61 & n93 ;
  assign n511 = n65 & n127 ;
  assign n512 = n510 | n511 ;
  assign n513 = n63 & n102 ;
  assign n514 = n35 & n97 ;
  assign n515 = n513 | n514 ;
  assign n516 = n512 | n515 ;
  assign n517 = n73 & n78 ;
  assign n518 = n116 & n150 ;
  assign n519 = n155 | n518 ;
  assign n520 = n517 | n519 ;
  assign n521 = n516 | n520 ;
  assign n522 = n509 | n521 ;
  assign n523 = n430 & ~n522 ;
  assign n524 = n353 | n523 ;
  assign n525 = n353 & n523 ;
  assign n526 = n524 & ~n525 ;
  assign n527 = n98 & n158 ;
  assign n528 = n432 | n527 ;
  assign n529 = n162 | n257 ;
  assign n530 = n343 | n529 ;
  assign n531 = n208 | n510 ;
  assign n532 = n530 | n531 ;
  assign n533 = n99 | n189 ;
  assign n534 = n399 | n469 ;
  assign n535 = n324 | n534 ;
  assign n536 = n533 | n535 ;
  assign n537 = n532 | n536 ;
  assign n538 = n371 | n537 ;
  assign n539 = n71 | n205 ;
  assign n540 = n302 | n503 ;
  assign n541 = n539 | n540 ;
  assign n542 = n65 & n74 ;
  assign n543 = n412 | n542 ;
  assign n544 = n77 | n543 ;
  assign n545 = n541 | n544 ;
  assign n546 = n123 | n151 ;
  assign n547 = n431 | n546 ;
  assign n548 = n545 | n547 ;
  assign n549 = n538 | n548 ;
  assign n550 = n197 | n288 ;
  assign n551 = n178 | n491 ;
  assign n552 = n550 | n551 ;
  assign n553 = n405 | n552 ;
  assign n554 = n141 | n202 ;
  assign n555 = n42 & ~n58 ;
  assign n556 = n142 | n555 ;
  assign n557 = n96 | n556 ;
  assign n558 = n554 | n557 ;
  assign n559 = n553 | n558 ;
  assign n560 = n35 & n42 ;
  assign n561 = n354 | n560 ;
  assign n562 = n249 | n476 ;
  assign n563 = n561 | n562 ;
  assign n564 = n236 | n384 ;
  assign n565 = n563 | n564 ;
  assign n566 = ~n38 & n102 ;
  assign n567 = n213 | n566 ;
  assign n568 = n109 & n127 ;
  assign n569 = n518 | n568 ;
  assign n570 = n567 | n569 ;
  assign n571 = n565 | n570 ;
  assign n572 = n559 | n571 ;
  assign n573 = n198 | n296 ;
  assign n574 = n49 & n91 ;
  assign n575 = n513 | n574 ;
  assign n576 = n573 | n575 ;
  assign n577 = n78 & n109 ;
  assign n578 = n229 | n577 ;
  assign n579 = n228 | n578 ;
  assign n580 = n576 | n579 ;
  assign n581 = n52 & n87 ;
  assign n582 = n450 | n581 ;
  assign n583 = n456 | n582 ;
  assign n584 = n580 | n583 ;
  assign n585 = n572 | n584 ;
  assign n586 = n549 | n585 ;
  assign n587 = n528 | n586 ;
  assign n588 = n113 & n116 ;
  assign n589 = n317 | n588 ;
  assign n590 = n78 & n87 ;
  assign n591 = n87 & n111 ;
  assign n592 = n590 | n591 ;
  assign n593 = n589 | n592 ;
  assign n594 = n86 & n132 ;
  assign n595 = n309 | n594 ;
  assign n596 = n325 | n595 ;
  assign n597 = n593 | n596 ;
  assign n598 = n254 | n305 ;
  assign n599 = n597 | n598 ;
  assign n600 = n35 & n127 ;
  assign n601 = n239 | n600 ;
  assign n602 = n49 & n127 ;
  assign n603 = n461 | n602 ;
  assign n604 = n601 | n603 ;
  assign n605 = n118 | n604 ;
  assign n606 = n170 | n225 ;
  assign n607 = n52 & n98 ;
  assign n608 = ~n38 & n113 ;
  assign n609 = n483 | n608 ;
  assign n610 = n607 | n609 ;
  assign n611 = n606 | n610 ;
  assign n612 = n605 | n611 ;
  assign n613 = n112 | n444 ;
  assign n614 = n363 | n613 ;
  assign n615 = n612 | n614 ;
  assign n616 = n78 & n122 ;
  assign n617 = n416 | n616 ;
  assign n618 = n177 | n617 ;
  assign n619 = n383 | n618 ;
  assign n620 = n209 | n387 ;
  assign n621 = n277 | n447 ;
  assign n622 = n620 | n621 ;
  assign n623 = n102 & n116 ;
  assign n624 = n63 & n109 ;
  assign n625 = n623 | n624 ;
  assign n626 = n332 | n625 ;
  assign n627 = n622 | n626 ;
  assign n628 = n619 | n627 ;
  assign n629 = n615 | n628 ;
  assign n630 = n92 | n192 ;
  assign n631 = n45 & n111 ;
  assign n632 = n280 | n631 ;
  assign n633 = n193 | n283 ;
  assign n634 = n632 | n633 ;
  assign n635 = n443 | n634 ;
  assign n636 = n245 | n312 ;
  assign n637 = n434 | n636 ;
  assign n638 = n65 & n116 ;
  assign n639 = n340 | n638 ;
  assign n640 = n637 | n639 ;
  assign n641 = n635 | n640 ;
  assign n642 = n630 | n641 ;
  assign n643 = n61 & n74 ;
  assign n644 = n66 & n132 ;
  assign n645 = n643 | n644 ;
  assign n646 = n303 | n487 ;
  assign n647 = n645 | n646 ;
  assign n648 = n49 & n63 ;
  assign n649 = n103 | n648 ;
  assign n650 = n457 | n649 ;
  assign n651 = n647 | n650 ;
  assign n652 = n196 | n497 ;
  assign n653 = n126 | n652 ;
  assign n654 = n63 & n84 ;
  assign n655 = n183 | n654 ;
  assign n656 = n131 | n237 ;
  assign n657 = n655 | n656 ;
  assign n658 = n653 | n657 ;
  assign n659 = n651 | n658 ;
  assign n660 = n117 | n418 ;
  assign n661 = n295 | n460 ;
  assign n662 = n660 | n661 ;
  assign n663 = n39 | n424 ;
  assign n664 = n271 | n663 ;
  assign n665 = n662 | n664 ;
  assign n666 = n91 & n132 ;
  assign n667 = n74 & n113 ;
  assign n668 = n666 | n667 ;
  assign n669 = n665 | n668 ;
  assign n670 = n659 | n669 ;
  assign n671 = n642 | n670 ;
  assign n672 = n629 | n671 ;
  assign n673 = n599 | n672 ;
  assign n674 = n587 | n673 ;
  assign n675 = n93 & n150 ;
  assign n676 = n42 & n109 ;
  assign n677 = n675 | n676 ;
  assign n678 = n182 | n677 ;
  assign n679 = n333 | n514 ;
  assign n680 = n184 | n374 ;
  assign n681 = n679 | n680 ;
  assign n682 = n258 | n451 ;
  assign n683 = n274 | n682 ;
  assign n684 = n681 | n683 ;
  assign n685 = n138 | n261 ;
  assign n686 = n124 | n685 ;
  assign n687 = n226 | n686 ;
  assign n688 = n684 | n687 ;
  assign n689 = n78 & n150 ;
  assign n690 = n448 | n689 ;
  assign n691 = n688 | n690 ;
  assign n692 = n678 | n691 ;
  assign n693 = n674 | n692 ;
  assign n694 = ~n38 & n150 ;
  assign n695 = n250 | n694 ;
  assign n696 = n42 & n132 ;
  assign n697 = n193 | n696 ;
  assign n698 = n255 | n406 ;
  assign n699 = n697 | n698 ;
  assign n700 = n104 | n497 ;
  assign n701 = n699 | n700 ;
  assign n702 = n75 | n343 ;
  assign n703 = n114 | n623 ;
  assign n704 = n702 | n703 ;
  assign n705 = n123 | n491 ;
  assign n706 = n483 | n705 ;
  assign n707 = n704 | n706 ;
  assign n708 = n701 | n707 ;
  assign n709 = n695 | n708 ;
  assign n710 = n167 | n568 ;
  assign n711 = n79 | n213 ;
  assign n712 = n710 | n711 ;
  assign n713 = n289 | n364 ;
  assign n714 = n246 | n713 ;
  assign n715 = n712 | n714 ;
  assign n716 = n296 | n715 ;
  assign n717 = n170 | n654 ;
  assign n718 = n154 | n465 ;
  assign n719 = n717 | n718 ;
  assign n720 = n61 & n91 ;
  assign n721 = n443 | n720 ;
  assign n722 = n228 | n588 ;
  assign n723 = n721 | n722 ;
  assign n724 = n719 | n723 ;
  assign n725 = n127 & n132 ;
  assign n726 = n143 & ~n725 ;
  assign n727 = ~n126 & n726 ;
  assign n728 = n142 | n479 ;
  assign n729 = n320 | n444 ;
  assign n730 = n728 | n729 ;
  assign n731 = n727 & ~n730 ;
  assign n732 = ~n724 & n731 ;
  assign n733 = ~n716 & n732 ;
  assign n734 = ~n709 & n733 ;
  assign n735 = n45 & n74 ;
  assign n736 = n233 | n735 ;
  assign n737 = n272 | n447 ;
  assign n738 = n736 | n737 ;
  assign n739 = n240 | n476 ;
  assign n740 = n332 | n739 ;
  assign n741 = n738 | n740 ;
  assign n742 = n734 & ~n741 ;
  assign n743 = n205 | n513 ;
  assign n744 = n517 | n743 ;
  assign n745 = n258 | n399 ;
  assign n746 = n196 | n745 ;
  assign n747 = n744 | n746 ;
  assign n748 = n247 | n270 ;
  assign n749 = n341 | n388 ;
  assign n750 = n660 | n749 ;
  assign n751 = n748 | n750 ;
  assign n752 = n747 | n751 ;
  assign n753 = n192 | n594 ;
  assign n754 = n305 | n624 ;
  assign n755 = n753 | n754 ;
  assign n756 = n752 | n755 ;
  assign n757 = n278 | n511 ;
  assign n758 = n109 & n158 ;
  assign n759 = n124 | n208 ;
  assign n760 = n758 | n759 ;
  assign n761 = n757 | n760 ;
  assign n762 = n52 & n122 ;
  assign n763 = n209 | n762 ;
  assign n764 = n348 | n448 ;
  assign n765 = n763 | n764 ;
  assign n766 = n133 | n249 ;
  assign n767 = n765 | n766 ;
  assign n768 = n761 | n767 ;
  assign n769 = n206 | n262 ;
  assign n770 = n395 | n600 ;
  assign n771 = n769 | n770 ;
  assign n772 = n768 | n771 ;
  assign n773 = n756 | n772 ;
  assign n774 = n176 | n518 ;
  assign n775 = ~n38 & n65 ;
  assign n776 = n92 | n775 ;
  assign n777 = n330 | n487 ;
  assign n778 = n776 | n777 ;
  assign n779 = n141 | n424 ;
  assign n780 = n436 | n779 ;
  assign n781 = n778 | n780 ;
  assign n782 = n774 | n781 ;
  assign n783 = n183 | n461 ;
  assign n784 = n236 | n284 ;
  assign n785 = n783 | n784 ;
  assign n786 = n85 | n574 ;
  assign n787 = n785 | n786 ;
  assign n788 = n592 | n787 ;
  assign n789 = n782 | n788 ;
  assign n790 = n773 | n789 ;
  assign n791 = n742 & ~n790 ;
  assign n792 = n112 | n616 ;
  assign n793 = n514 | n792 ;
  assign n794 = n55 | n793 ;
  assign n795 = n189 | n503 ;
  assign n796 = n226 | n295 ;
  assign n797 = n795 | n796 ;
  assign n798 = n318 | n797 ;
  assign n799 = n794 | n798 ;
  assign n800 = n257 | n355 ;
  assign n801 = n35 & n158 ;
  assign n802 = n675 | n801 ;
  assign n803 = n800 | n802 ;
  assign n804 = n182 | n803 ;
  assign n805 = n799 | n804 ;
  assign n806 = n113 & n127 ;
  assign n807 = n234 | n806 ;
  assign n808 = n64 | n171 ;
  assign n809 = n372 | n416 ;
  assign n810 = n808 | n809 ;
  assign n811 = n288 | n480 ;
  assign n812 = n303 | n811 ;
  assign n813 = n810 | n812 ;
  assign n814 = n118 | n566 ;
  assign n815 = n283 | n405 ;
  assign n816 = n814 | n815 ;
  assign n817 = n813 | n816 ;
  assign n818 = n807 | n817 ;
  assign n819 = n805 | n818 ;
  assign n820 = n52 & n65 ;
  assign n821 = n510 | n820 ;
  assign n822 = n667 | n821 ;
  assign n823 = n819 | n822 ;
  assign n824 = n297 | n457 ;
  assign n825 = ( n163 & n643 ) | ( n163 & ~n824 ) | ( n643 & ~n824 ) ;
  assign n826 = n225 | n824 ;
  assign n827 = n825 | n826 ;
  assign n828 = n823 | n827 ;
  assign n829 = n791 & ~n828 ;
  assign n830 = n693 & ~n829 ;
  assign n831 = ~n693 & n829 ;
  assign n832 = n830 | n831 ;
  assign n833 = n432 | n806 ;
  assign n834 = n348 | n542 ;
  assign n835 = n833 | n834 ;
  assign n836 = n401 | n577 ;
  assign n837 = n204 | n836 ;
  assign n838 = n835 | n837 ;
  assign n839 = n49 & n57 ;
  assign n840 = n284 | n839 ;
  assign n841 = ~n38 & n61 ;
  assign n842 = n456 | n841 ;
  assign n843 = n840 | n842 ;
  assign n844 = n465 | n560 ;
  assign n845 = n413 | n758 ;
  assign n846 = n844 | n845 ;
  assign n847 = n843 | n846 ;
  assign n848 = n838 | n847 ;
  assign n849 = n159 | n179 ;
  assign n850 = n406 | n849 ;
  assign n851 = n90 | n850 ;
  assign n852 = n114 | n190 ;
  assign n853 = n318 | n344 ;
  assign n854 = n263 | n853 ;
  assign n855 = n852 | n854 ;
  assign n856 = n851 | n855 ;
  assign n857 = n104 | n331 ;
  assign n858 = ~n58 & n91 ;
  assign n859 = n801 | n858 ;
  assign n860 = n857 | n859 ;
  assign n861 = n500 | n860 ;
  assign n862 = n626 | n861 ;
  assign n863 = n856 | n862 ;
  assign n864 = n848 | n863 ;
  assign n865 = n671 | n864 ;
  assign n866 = n247 | n775 ;
  assign n867 = n152 | n236 ;
  assign n868 = n866 | n867 ;
  assign n869 = n324 | n395 ;
  assign n870 = n64 | n511 ;
  assign n871 = n869 | n870 ;
  assign n872 = n868 | n871 ;
  assign n873 = n711 | n872 ;
  assign n874 = n865 | n873 ;
  assign n875 = n168 | n590 ;
  assign n876 = n143 & ~n349 ;
  assign n877 = ~n875 & n876 ;
  assign n878 = n355 | n390 ;
  assign n879 = n384 | n878 ;
  assign n880 = n67 | n370 ;
  assign n881 = n449 | n880 ;
  assign n882 = n879 | n881 ;
  assign n883 = n877 & ~n882 ;
  assign n884 = n330 | n762 ;
  assign n885 = n372 | n884 ;
  assign n886 = n42 & n73 ;
  assign n887 = n52 & n73 ;
  assign n888 = n886 | n887 ;
  assign n889 = n240 | n888 ;
  assign n890 = n885 | n889 ;
  assign n891 = n96 | n234 ;
  assign n892 = n890 | n891 ;
  assign n893 = n883 & ~n892 ;
  assign n894 = n575 | n682 ;
  assign n895 = n86 & n102 ;
  assign n896 = n321 | n399 ;
  assign n897 = n895 | n896 ;
  assign n898 = n894 | n897 ;
  assign n899 = n374 | n898 ;
  assign n900 = n296 | n458 ;
  assign n901 = n45 & n57 ;
  assign n902 = n176 | n901 ;
  assign n903 = n900 | n902 ;
  assign n904 = n214 | n725 ;
  assign n905 = n310 | n904 ;
  assign n906 = n903 | n905 ;
  assign n907 = n272 | n381 ;
  assign n908 = n710 | n907 ;
  assign n909 = n906 | n908 ;
  assign n910 = n899 | n909 ;
  assign n911 = n893 & ~n910 ;
  assign n912 = n208 | n441 ;
  assign n913 = n142 | n694 ;
  assign n914 = n912 | n913 ;
  assign n915 = n405 | n914 ;
  assign n916 = n911 & ~n915 ;
  assign n917 = n134 | n257 ;
  assign n918 = n702 | n917 ;
  assign n919 = n250 | n281 ;
  assign n920 = n918 | n919 ;
  assign n921 = n916 & ~n920 ;
  assign n922 = ~n874 & n921 ;
  assign n923 = n92 | n399 ;
  assign n924 = n272 | n689 ;
  assign n925 = n923 | n924 ;
  assign n926 = n143 & ~n347 ;
  assign n927 = ~n639 & n926 ;
  assign n928 = ~n925 & n927 ;
  assign n929 = n278 | n476 ;
  assign n930 = n184 | n501 ;
  assign n931 = n413 | n483 ;
  assign n932 = n930 | n931 ;
  assign n933 = n929 | n932 ;
  assign n934 = n928 & ~n933 ;
  assign n935 = n53 | n372 ;
  assign n936 = n573 | n935 ;
  assign n937 = n460 | n886 ;
  assign n938 = n66 & n113 ;
  assign n939 = n104 | n938 ;
  assign n940 = n937 | n939 ;
  assign n941 = n936 | n940 ;
  assign n942 = n324 | n887 ;
  assign n943 = n332 | n942 ;
  assign n944 = n261 | n574 ;
  assign n945 = n118 | n128 ;
  assign n946 = n944 | n945 ;
  assign n947 = n943 | n946 ;
  assign n948 = n941 | n947 ;
  assign n949 = n934 & ~n948 ;
  assign n950 = n282 | n820 ;
  assign n951 = n112 | n666 ;
  assign n952 = n228 | n341 ;
  assign n953 = n206 | n555 ;
  assign n954 = n952 | n953 ;
  assign n955 = n951 | n954 ;
  assign n956 = n950 | n955 ;
  assign n957 = n344 | n448 ;
  assign n958 = n624 | n957 ;
  assign n959 = n87 & n116 ;
  assign n960 = n405 | n517 ;
  assign n961 = n959 | n960 ;
  assign n962 = n958 | n961 ;
  assign n963 = n131 | n291 ;
  assign n964 = n962 | n963 ;
  assign n965 = n956 | n964 ;
  assign n966 = n432 | n487 ;
  assign n967 = n233 | n667 ;
  assign n968 = n966 | n967 ;
  assign n969 = n607 | n725 ;
  assign n970 = n295 | n969 ;
  assign n971 = n968 | n970 ;
  assign n972 = n254 | n971 ;
  assign n973 = n406 | n839 ;
  assign n974 = n313 | n720 ;
  assign n975 = n973 | n974 ;
  assign n976 = n133 | n196 ;
  assign n977 = n675 | n976 ;
  assign n978 = n975 | n977 ;
  assign n979 = n444 | n801 ;
  assign n980 = n94 | n696 ;
  assign n981 = n979 | n980 ;
  assign n982 = n978 | n981 ;
  assign n983 = n972 | n982 ;
  assign n984 = n965 | n983 ;
  assign n985 = n949 & ~n984 ;
  assign n986 = n381 | n424 ;
  assign n987 = n124 | n212 ;
  assign n988 = n841 | n987 ;
  assign n989 = n986 | n988 ;
  assign n990 = n368 | n989 ;
  assign n991 = n321 | n560 ;
  assign n992 = n317 | n480 ;
  assign n993 = n456 | n992 ;
  assign n994 = n991 | n993 ;
  assign n995 = n269 | n277 ;
  assign n996 = n795 | n995 ;
  assign n997 = n994 | n996 ;
  assign n998 = n990 | n997 ;
  assign n999 = n441 | n577 ;
  assign n1000 = n783 | n999 ;
  assign n1001 = n163 | n477 ;
  assign n1002 = n88 | n458 ;
  assign n1003 = n1001 | n1002 ;
  assign n1004 = n1000 | n1003 ;
  assign n1005 = n374 | n431 ;
  assign n1006 = n247 | n288 ;
  assign n1007 = n1005 | n1006 ;
  assign n1008 = n77 | n644 ;
  assign n1009 = n283 | n343 ;
  assign n1010 = n1008 | n1009 ;
  assign n1011 = n1007 | n1010 ;
  assign n1012 = n1004 | n1011 ;
  assign n1013 = n59 | n245 ;
  assign n1014 = n202 | n602 ;
  assign n1015 = n1013 | n1014 ;
  assign n1016 = n83 | n568 ;
  assign n1017 = n617 | n1016 ;
  assign n1018 = n1015 | n1017 ;
  assign n1019 = n170 | n591 ;
  assign n1020 = n1018 | n1019 ;
  assign n1021 = n1012 | n1020 ;
  assign n1022 = n998 | n1021 ;
  assign n1023 = n123 | n222 ;
  assign n1024 = n192 | n234 ;
  assign n1025 = n1023 | n1024 ;
  assign n1026 = n1022 | n1025 ;
  assign n1027 = n985 & ~n1026 ;
  assign n1028 = n96 | n468 ;
  assign n1029 = n649 | n1028 ;
  assign n1030 = n151 | n518 ;
  assign n1031 = n513 | n775 ;
  assign n1032 = n1030 | n1031 ;
  assign n1033 = n1029 | n1032 ;
  assign n1034 = n401 | n489 ;
  assign n1035 = n79 | n209 ;
  assign n1036 = n1034 | n1035 ;
  assign n1037 = n117 | n1036 ;
  assign n1038 = n1033 | n1037 ;
  assign n1039 = n52 & n61 ;
  assign n1040 = n160 | n1039 ;
  assign n1041 = n1038 | n1040 ;
  assign n1042 = n139 | n1041 ;
  assign n1043 = n1027 & ~n1042 ;
  assign n1044 = n922 | n1043 ;
  assign n1045 = ( ~n693 & n922 ) | ( ~n693 & n1044 ) | ( n922 & n1044 ) ;
  assign n1046 = n832 | n1045 ;
  assign n1047 = n353 & n829 ;
  assign n1048 = n353 | n829 ;
  assign n1049 = ~n1047 & n1048 ;
  assign n1050 = n830 & n1049 ;
  assign n1051 = n1048 & ~n1050 ;
  assign n1052 = ( n1046 & n1047 ) | ( n1046 & n1051 ) | ( n1047 & n1051 ) ;
  assign n1053 = n526 & ~n1052 ;
  assign n1054 = ~n526 & n1052 ;
  assign n1055 = n1053 | n1054 ;
  assign n1822 = n43 & ~n48 ;
  assign n1815 = x28 & ~x29 ;
  assign n1816 = ~x28 & x29 ;
  assign n1817 = n1815 | n1816 ;
  assign n1818 = x26 & ~x27 ;
  assign n1819 = ~x26 & x27 ;
  assign n1820 = n1818 | n1819 ;
  assign n1825 = n1817 & ~n1820 ;
  assign n1826 = ~n1822 & n1825 ;
  assign n1902 = ~n829 & n1826 ;
  assign n1823 = ~n1820 & n1822 ;
  assign n1903 = n352 & n1823 ;
  assign n1904 = ( ~n339 & n1823 ) | ( ~n339 & n1903 ) | ( n1823 & n1903 ) ;
  assign n1905 = n1902 | n1904 ;
  assign n1821 = n1817 & n1820 ;
  assign n1829 = ~n1817 & n1820 ;
  assign n1906 = ~n523 & n1829 ;
  assign n1907 = n1821 | n1906 ;
  assign n1908 = n1905 | n1907 ;
  assign n1909 = ~x29 & n1908 ;
  assign n1910 = n1905 | n1906 ;
  assign n1911 = ~x29 & n1910 ;
  assign n1912 = ( ~n1055 & n1909 ) | ( ~n1055 & n1911 ) | ( n1909 & n1911 ) ;
  assign n1913 = x29 & n1908 ;
  assign n1914 = x29 & ~n1913 ;
  assign n1915 = x29 & n1906 ;
  assign n1916 = ( x29 & n1905 ) | ( x29 & n1915 ) | ( n1905 & n1915 ) ;
  assign n1917 = x29 & ~n1916 ;
  assign n1918 = ( n1055 & n1914 ) | ( n1055 & n1917 ) | ( n1914 & n1917 ) ;
  assign n1919 = n1912 | n1918 ;
  assign n1429 = n461 | n820 ;
  assign n1430 = n291 | n465 ;
  assign n1431 = n1429 | n1430 ;
  assign n1432 = n762 | n1431 ;
  assign n1301 = n347 | n517 ;
  assign n1433 = n257 | n431 ;
  assign n1434 = n1301 | n1433 ;
  assign n1435 = n487 | n1434 ;
  assign n1436 = n134 | n197 ;
  assign n1437 = n478 | n1436 ;
  assign n1438 = n1435 | n1437 ;
  assign n1439 = n189 | n638 ;
  assign n1440 = n306 | n383 ;
  assign n1441 = n1439 | n1440 ;
  assign n1442 = n281 | n895 ;
  assign n1443 = n1441 | n1442 ;
  assign n1444 = n1438 | n1443 ;
  assign n1221 = n77 | n497 ;
  assign n1445 = n83 | n269 ;
  assign n1446 = n1221 | n1445 ;
  assign n1447 = n229 | n608 ;
  assign n1448 = n539 | n1447 ;
  assign n1449 = n1446 | n1448 ;
  assign n1380 = n138 | n375 ;
  assign n1450 = n167 | n228 ;
  assign n1451 = n1380 | n1450 ;
  assign n1452 = n1449 | n1451 ;
  assign n1453 = n418 | n735 ;
  assign n1454 = n143 & ~n272 ;
  assign n1455 = ~n1453 & n1454 ;
  assign n1456 = ~n295 & n1455 ;
  assign n1457 = ~n324 & n1456 ;
  assign n1458 = ~n1452 & n1457 ;
  assign n1459 = ~n1444 & n1458 ;
  assign n1355 = n99 | n214 ;
  assign n1460 = n133 | n332 ;
  assign n1461 = n1355 | n1460 ;
  assign n1462 = n112 | n624 ;
  assign n1463 = n1461 | n1462 ;
  assign n1464 = n177 | n289 ;
  assign n1465 = n480 | n616 ;
  assign n1466 = n720 | n725 ;
  assign n1467 = n1465 | n1466 ;
  assign n1468 = n1464 | n1467 ;
  assign n1469 = n124 | n354 ;
  assign n1470 = n749 | n1469 ;
  assign n1471 = n1468 | n1470 ;
  assign n1472 = n1463 | n1471 ;
  assign n1473 = n46 | n261 ;
  assign n1474 = n226 | n402 ;
  assign n1475 = n1473 | n1474 ;
  assign n1476 = n39 | n435 ;
  assign n1477 = n600 | n1476 ;
  assign n1478 = n1475 | n1477 ;
  assign n1479 = n237 | n254 ;
  assign n1480 = n263 | n1479 ;
  assign n1481 = n1478 | n1480 ;
  assign n1482 = n364 | n696 ;
  assign n1483 = n273 | n310 ;
  assign n1484 = n1482 | n1483 ;
  assign n1303 = n155 | n758 ;
  assign n1485 = n527 | n1303 ;
  assign n1486 = n1484 | n1485 ;
  assign n1487 = n163 | n460 ;
  assign n1488 = n1486 | n1487 ;
  assign n1489 = n1481 | n1488 ;
  assign n1490 = n1472 | n1489 ;
  assign n1491 = n1459 & ~n1490 ;
  assign n1097 = n542 | n858 ;
  assign n1492 = n110 | n1097 ;
  assign n1493 = n88 | n387 ;
  assign n1494 = n331 | n1493 ;
  assign n1495 = n1492 | n1494 ;
  assign n1267 = n198 | n234 ;
  assign n1268 = n390 | n694 ;
  assign n1269 = n1267 | n1268 ;
  assign n1496 = n717 | n757 ;
  assign n1497 = n1269 | n1496 ;
  assign n1498 = n1495 | n1497 ;
  assign n1499 = n206 | n469 ;
  assign n1500 = n190 | n648 ;
  assign n1501 = n1499 | n1500 ;
  assign n1502 = n118 | n1501 ;
  assign n1503 = n551 | n1014 ;
  assign n1504 = n1502 | n1503 ;
  assign n1505 = n1498 | n1504 ;
  assign n1506 = n224 | n836 ;
  assign n1507 = n246 | n806 ;
  assign n1508 = n239 | n1507 ;
  assign n1509 = n1506 | n1508 ;
  assign n1510 = n160 | n344 ;
  assign n1511 = n675 | n1510 ;
  assign n1512 = n1509 | n1511 ;
  assign n1513 = n240 | n374 ;
  assign n1146 = n333 | n886 ;
  assign n1514 = n923 | n1146 ;
  assign n1515 = n297 | n395 ;
  assign n1516 = n560 | n1515 ;
  assign n1517 = n1514 | n1516 ;
  assign n1518 = n1513 | n1517 ;
  assign n1519 = n1512 | n1518 ;
  assign n1520 = n1505 | n1519 ;
  assign n1521 = n288 | n574 ;
  assign n1522 = n417 | n1521 ;
  assign n1523 = n192 | n233 ;
  assign n1524 = n357 | n1523 ;
  assign n1525 = n1522 | n1524 ;
  assign n1526 = n319 | n748 ;
  assign n1527 = n114 | n1526 ;
  assign n1528 = n1525 | n1527 ;
  assign n1172 = n84 & n97 ;
  assign n1529 = n591 | n1172 ;
  assign n1530 = n1528 | n1529 ;
  assign n1531 = n1520 | n1530 ;
  assign n1532 = n1491 & ~n1531 ;
  assign n1533 = ~n1432 & n1532 ;
  assign n1535 = ~n922 & n1043 ;
  assign n1536 = n693 | n1535 ;
  assign n1537 = n693 & n1535 ;
  assign n1538 = n1536 & ~n1537 ;
  assign n1056 = n47 | n72 ;
  assign n1063 = ~x30 & x31 ;
  assign n1064 = ( x30 & ~x31 ) | ( x30 & n1063 ) | ( ~x31 & n1063 ) ;
  assign n1065 = ( ~n1056 & n1063 ) | ( ~n1056 & n1064 ) | ( n1063 & n1064 ) ;
  assign n1539 = ~n922 & n1065 ;
  assign n1059 = x30 & x31 ;
  assign n1060 = ~n1056 & n1059 ;
  assign n1540 = n1042 & n1060 ;
  assign n1541 = ( ~n1027 & n1060 ) | ( ~n1027 & n1540 ) | ( n1060 & n1540 ) ;
  assign n1542 = n1539 | n1541 ;
  assign n1057 = ~x31 & n1056 ;
  assign n1543 = n692 & n1057 ;
  assign n1544 = ( n674 & n1057 ) | ( n674 & n1543 ) | ( n1057 & n1543 ) ;
  assign n1545 = n1542 | n1544 ;
  assign n1062 = x31 & n1056 ;
  assign n1546 = n1062 | n1540 ;
  assign n1547 = n1060 | n1062 ;
  assign n1548 = ( ~n1027 & n1546 ) | ( ~n1027 & n1547 ) | ( n1546 & n1547 ) ;
  assign n1549 = n1539 | n1548 ;
  assign n1550 = n1544 | n1549 ;
  assign n1551 = ( n1538 & n1545 ) | ( n1538 & n1550 ) | ( n1545 & n1550 ) ;
  assign n1920 = n1533 | n1551 ;
  assign n1921 = n1533 & n1551 ;
  assign n1922 = n1920 & ~n1921 ;
  assign n1923 = n1919 & ~n1922 ;
  assign n1924 = ~n1919 & n1922 ;
  assign n1925 = n1923 | n1924 ;
  assign n1206 = ( ~n1046 & n1049 ) | ( ~n1046 & n1050 ) | ( n1049 & n1050 ) ;
  assign n1207 = n830 | n1049 ;
  assign n1208 = n1046 & ~n1207 ;
  assign n1209 = n1206 | n1208 ;
  assign n1926 = ~n829 & n1823 ;
  assign n1927 = n352 & n1829 ;
  assign n1928 = ( ~n339 & n1829 ) | ( ~n339 & n1927 ) | ( n1829 & n1927 ) ;
  assign n1929 = n1926 | n1928 ;
  assign n1930 = n692 & n1826 ;
  assign n1931 = ( n674 & n1826 ) | ( n674 & n1930 ) | ( n1826 & n1930 ) ;
  assign n1932 = n1821 | n1931 ;
  assign n1933 = n1929 | n1932 ;
  assign n1934 = ~x29 & n1933 ;
  assign n1935 = n1929 | n1931 ;
  assign n1936 = ~x29 & n1935 ;
  assign n1937 = ( ~n1209 & n1934 ) | ( ~n1209 & n1936 ) | ( n1934 & n1936 ) ;
  assign n1938 = x29 & n1933 ;
  assign n1939 = x29 & ~n1938 ;
  assign n1940 = x29 & n1931 ;
  assign n1941 = ( x29 & n1929 ) | ( x29 & n1940 ) | ( n1929 & n1940 ) ;
  assign n1942 = x29 & ~n1941 ;
  assign n1943 = ( n1209 & n1939 ) | ( n1209 & n1942 ) | ( n1939 & n1942 ) ;
  assign n1944 = n1937 | n1943 ;
  assign n1945 = n922 & ~n1043 ;
  assign n1946 = n1535 | n1945 ;
  assign n1947 = ~n922 & n1057 ;
  assign n1948 = n1042 & n1065 ;
  assign n1949 = ( ~n1027 & n1065 ) | ( ~n1027 & n1948 ) | ( n1065 & n1948 ) ;
  assign n1950 = n1947 | n1949 ;
  assign n1951 = n1062 | n1949 ;
  assign n1952 = n1947 | n1951 ;
  assign n1953 = ( n1946 & n1950 ) | ( n1946 & n1952 ) | ( n1950 & n1952 ) ;
  assign n1954 = n1944 & n1953 ;
  assign n1955 = n1944 | n1953 ;
  assign n1956 = ~n1954 & n1955 ;
  assign n1553 = n832 & n1045 ;
  assign n1554 = n1046 & ~n1553 ;
  assign n1957 = ~n829 & n1829 ;
  assign n1958 = ~n922 & n1826 ;
  assign n1959 = n1957 | n1958 ;
  assign n1960 = n692 & n1823 ;
  assign n1961 = ( n674 & n1823 ) | ( n674 & n1960 ) | ( n1823 & n1960 ) ;
  assign n1962 = n1959 | n1961 ;
  assign n1963 = n1821 | n1961 ;
  assign n1964 = n1959 | n1963 ;
  assign n1965 = ( n1554 & n1962 ) | ( n1554 & n1964 ) | ( n1962 & n1964 ) ;
  assign n1966 = x29 & n1964 ;
  assign n1967 = x29 & n1962 ;
  assign n1968 = ( n1554 & n1966 ) | ( n1554 & n1967 ) | ( n1966 & n1967 ) ;
  assign n1969 = x29 & ~n1967 ;
  assign n1970 = x29 & ~n1966 ;
  assign n1971 = ( ~n1554 & n1969 ) | ( ~n1554 & n1970 ) | ( n1969 & n1970 ) ;
  assign n1972 = ( n1965 & ~n1968 ) | ( n1965 & n1971 ) | ( ~n1968 & n1971 ) ;
  assign n1973 = ~n922 & n1823 ;
  assign n1974 = n1042 & n1826 ;
  assign n1975 = ( ~n1027 & n1826 ) | ( ~n1027 & n1974 ) | ( n1826 & n1974 ) ;
  assign n1976 = n1973 | n1975 ;
  assign n1977 = n692 & n1829 ;
  assign n1978 = ( n674 & n1829 ) | ( n674 & n1977 ) | ( n1829 & n1977 ) ;
  assign n1979 = n1976 | n1978 ;
  assign n1980 = ( n1538 & n1821 ) | ( n1538 & n1979 ) | ( n1821 & n1979 ) ;
  assign n1981 = ( x29 & ~n1979 ) | ( x29 & n1980 ) | ( ~n1979 & n1980 ) ;
  assign n1982 = ~n1980 & n1981 ;
  assign n1983 = ~n922 & n1829 ;
  assign n1984 = n1042 & n1823 ;
  assign n1985 = ( ~n1027 & n1823 ) | ( ~n1027 & n1984 ) | ( n1823 & n1984 ) ;
  assign n1986 = n1983 | n1985 ;
  assign n1987 = n1821 | n1985 ;
  assign n1988 = n1983 | n1987 ;
  assign n1989 = ( n1946 & n1986 ) | ( n1946 & n1988 ) | ( n1986 & n1988 ) ;
  assign n1990 = ~x29 & n1989 ;
  assign n1991 = n139 & n1820 ;
  assign n1992 = ( n1041 & n1820 ) | ( n1041 & n1991 ) | ( n1820 & n1991 ) ;
  assign n1993 = x29 & ~n1992 ;
  assign n1994 = n1820 | n1991 ;
  assign n1995 = x29 & ~n1994 ;
  assign n1996 = ( n1027 & n1993 ) | ( n1027 & n1995 ) | ( n1993 & n1995 ) ;
  assign n1997 = x29 & n1996 ;
  assign n1998 = ~n1989 & n1997 ;
  assign n1999 = ( n1990 & n1996 ) | ( n1990 & n1998 ) | ( n1996 & n1998 ) ;
  assign n2000 = x29 | n1979 ;
  assign n2001 = n1980 | n2000 ;
  assign n2002 = n1999 & n2001 ;
  assign n2003 = ~x29 & n1999 ;
  assign n2004 = ( n1982 & n2002 ) | ( n1982 & n2003 ) | ( n2002 & n2003 ) ;
  assign n2005 = n1057 | n1062 ;
  assign n2006 = n1041 & n2005 ;
  assign n2007 = ( ~n1027 & n2005 ) | ( ~n1027 & n2006 ) | ( n2005 & n2006 ) ;
  assign n2008 = ( n1972 & n2004 ) | ( n1972 & n2007 ) | ( n2004 & n2007 ) ;
  assign n2009 = n1954 | n2008 ;
  assign n2010 = ( n1954 & n1956 ) | ( n1954 & n2009 ) | ( n1956 & n2009 ) ;
  assign n2011 = ~n1925 & n2010 ;
  assign n2369 = n1925 & ~n2010 ;
  assign n2370 = n2011 | n2369 ;
  assign n1575 = n247 | n654 ;
  assign n1576 = n555 | n735 ;
  assign n1577 = n1575 | n1576 ;
  assign n1578 = n325 | n465 ;
  assign n1579 = n887 | n1578 ;
  assign n1580 = n1577 | n1579 ;
  assign n1581 = n103 | n514 ;
  assign n1582 = n125 | n1581 ;
  assign n1583 = n261 | n456 ;
  assign n1584 = n197 | n375 ;
  assign n1585 = n1583 | n1584 ;
  assign n1586 = n1582 | n1585 ;
  assign n1587 = n1580 | n1586 ;
  assign n1588 = n807 | n1005 ;
  assign n1589 = n153 | n923 ;
  assign n1590 = n1588 | n1589 ;
  assign n1591 = n202 | n483 ;
  assign n1592 = n213 | n590 ;
  assign n1593 = n1591 | n1592 ;
  assign n1594 = n71 | n444 ;
  assign n1595 = n1593 | n1594 ;
  assign n1596 = n1590 | n1595 ;
  assign n1597 = n1587 | n1596 ;
  assign n1598 = n126 | n1597 ;
  assign n1599 = n175 | n648 ;
  assign n1600 = n212 | n270 ;
  assign n1601 = n1599 | n1600 ;
  assign n1602 = n517 | n1601 ;
  assign n1603 = n237 | n623 ;
  assign n1604 = n311 | n1603 ;
  assign n1605 = n694 | n1604 ;
  assign n1606 = n1602 | n1605 ;
  assign n1607 = n395 | n1039 ;
  assign n1118 = n206 | n236 ;
  assign n1608 = n324 | n1118 ;
  assign n1609 = n417 | n1608 ;
  assign n1610 = n1607 | n1609 ;
  assign n1611 = n1606 | n1610 ;
  assign n1612 = n1598 | n1611 ;
  assign n1214 = n79 | n839 ;
  assign n1215 = n154 | n1214 ;
  assign n1331 = n205 | n387 ;
  assign n1332 = n418 | n1331 ;
  assign n1333 = n1215 | n1332 ;
  assign n1334 = n402 | n775 ;
  assign n1335 = n133 | n1334 ;
  assign n1336 = n67 | n1172 ;
  assign n1337 = n1335 | n1336 ;
  assign n1338 = n1333 | n1337 ;
  assign n1339 = n496 | n1338 ;
  assign n1340 = n245 | n257 ;
  assign n1341 = n306 | n354 ;
  assign n1342 = n939 | n1341 ;
  assign n1343 = n1340 | n1342 ;
  assign n1149 = n284 | n435 ;
  assign n1344 = n269 | n344 ;
  assign n1345 = n273 | n801 ;
  assign n1346 = n1344 | n1345 ;
  assign n1347 = n1149 | n1346 ;
  assign n1348 = n1343 | n1347 ;
  assign n1349 = n631 | n725 ;
  assign n1350 = n383 | n666 ;
  assign n1351 = n1349 | n1350 ;
  assign n1352 = n182 | n1351 ;
  assign n1353 = n1348 | n1352 ;
  assign n1354 = n1339 | n1353 ;
  assign n1356 = n256 | n1355 ;
  assign n1357 = n764 | n967 ;
  assign n1358 = n1356 | n1357 ;
  assign n1359 = n341 | n412 ;
  assign n1360 = n1358 | n1359 ;
  assign n1613 = n697 | n728 ;
  assign n1614 = n1303 | n1613 ;
  assign n1362 = n447 | n594 ;
  assign n1363 = n405 | n1362 ;
  assign n1615 = n434 | n858 ;
  assign n1616 = n134 | n1615 ;
  assign n1617 = n1363 | n1616 ;
  assign n1618 = n1614 | n1617 ;
  assign n1619 = n442 | n796 ;
  assign n1620 = n190 | n1619 ;
  assign n1621 = n289 | n355 ;
  assign n1622 = n223 | n280 ;
  assign n1623 = n1621 | n1622 ;
  assign n1624 = n54 | n542 ;
  assign n1625 = n1623 | n1624 ;
  assign n1626 = n1620 | n1625 ;
  assign n1627 = n1618 | n1626 ;
  assign n1628 = n1360 | n1627 ;
  assign n1629 = n1354 | n1628 ;
  assign n1630 = n1612 | n1629 ;
  assign n1631 = n163 | n901 ;
  assign n1632 = n140 | n1631 ;
  assign n1633 = n178 | n192 ;
  assign n1634 = n1632 | n1633 ;
  assign n1635 = n1630 | n1634 ;
  assign n1216 = n269 | n841 ;
  assign n1217 = n577 | n1216 ;
  assign n1218 = ( n503 & ~n1215 ) | ( n503 & n1217 ) | ( ~n1215 & n1217 ) ;
  assign n1219 = n1215 | n1218 ;
  assign n1220 = n356 | n1039 ;
  assign n1222 = n83 | n372 ;
  assign n1223 = n533 | n1222 ;
  assign n1224 = n1221 | n1223 ;
  assign n1225 = n296 | n590 ;
  assign n1226 = n291 | n1225 ;
  assign n1227 = ( ~n1220 & n1224 ) | ( ~n1220 & n1226 ) | ( n1224 & n1226 ) ;
  assign n1228 = n1220 & ~n1226 ;
  assign n1229 = ( n1219 & n1227 ) | ( n1219 & ~n1228 ) | ( n1227 & ~n1228 ) ;
  assign n1230 = n555 | n1220 ;
  assign n1231 = n1229 | n1230 ;
  assign n1232 = n344 | n643 ;
  assign n1233 = n138 | n233 ;
  assign n1234 = n433 | n1233 ;
  assign n1235 = n1232 | n1234 ;
  assign n1086 = n209 | n450 ;
  assign n1087 = n203 | n616 ;
  assign n1088 = n1086 | n1087 ;
  assign n1236 = n771 | n1088 ;
  assign n1237 = n1235 | n1236 ;
  assign n1238 = n364 | n735 ;
  assign n1239 = n239 | n1238 ;
  assign n1240 = n118 | n501 ;
  assign n1241 = n852 | n1240 ;
  assign n1242 = n1239 | n1241 ;
  assign n1243 = n560 | n858 ;
  assign n1244 = n331 | n457 ;
  assign n1245 = n341 | n1244 ;
  assign n1246 = n1243 | n1245 ;
  assign n1247 = n1242 | n1246 ;
  assign n1248 = n1237 | n1247 ;
  assign n1249 = n257 | n483 ;
  assign n1250 = n133 | n1249 ;
  assign n1251 = n246 | n384 ;
  assign n1252 = n980 | n1251 ;
  assign n1253 = n1250 | n1252 ;
  assign n1254 = n289 | n821 ;
  assign n1255 = n178 | n1254 ;
  assign n1256 = n1253 | n1255 ;
  assign n1257 = n1248 | n1256 ;
  assign n1258 = n1231 | n1257 ;
  assign n1274 = n205 | n214 ;
  assign n1275 = n64 | n321 ;
  assign n1276 = n1274 | n1275 ;
  assign n1277 = n320 | n381 ;
  assign n1278 = n1276 | n1277 ;
  assign n1636 = n324 | n468 ;
  assign n1637 = n437 | n675 ;
  assign n1638 = n1636 | n1637 ;
  assign n1639 = n623 | n1638 ;
  assign n1640 = n196 | n198 ;
  assign n1641 = n282 | n1640 ;
  assign n1642 = n155 | n234 ;
  assign n1643 = n1030 | n1642 ;
  assign n1644 = n1641 | n1643 ;
  assign n1645 = n1639 | n1644 ;
  assign n1646 = n363 | n513 ;
  assign n1647 = n695 | n1646 ;
  assign n1648 = n424 | n1647 ;
  assign n1649 = n1645 | n1648 ;
  assign n1650 = n247 | n406 ;
  assign n1651 = n444 | n480 ;
  assign n1652 = n1034 | n1651 ;
  assign n1653 = n333 | n566 ;
  assign n1654 = n230 | n1653 ;
  assign n1655 = n1652 | n1654 ;
  assign n1656 = n1650 | n1655 ;
  assign n1657 = n112 | n192 ;
  assign n1658 = n226 | n469 ;
  assign n1659 = n1657 | n1658 ;
  assign n1114 = n35 & n116 ;
  assign n1660 = n263 | n1114 ;
  assign n1661 = n1659 | n1660 ;
  assign n1662 = n317 | n458 ;
  assign n1663 = n278 | n465 ;
  assign n1664 = n1662 | n1663 ;
  assign n1665 = n330 | n370 ;
  assign n1666 = n354 | n1665 ;
  assign n1667 = n1664 | n1666 ;
  assign n1668 = n1661 | n1667 ;
  assign n1669 = n1656 | n1668 ;
  assign n1670 = n1649 | n1669 ;
  assign n1671 = n1278 | n1670 ;
  assign n1672 = n1258 | n1671 ;
  assign n1165 = n514 | n938 ;
  assign n1673 = n491 | n638 ;
  assign n1674 = n1165 | n1673 ;
  assign n1675 = n369 | n387 ;
  assign n1676 = n1583 | n1675 ;
  assign n1677 = n1674 | n1676 ;
  assign n1678 = n139 | n608 ;
  assign n1679 = n923 | n1678 ;
  assign n1680 = n479 | n1679 ;
  assign n1681 = n1677 | n1680 ;
  assign n1682 = n249 | n654 ;
  assign n1683 = n447 | n901 ;
  assign n1684 = n1682 | n1683 ;
  assign n1685 = n1681 | n1684 ;
  assign n1686 = n274 | n1301 ;
  assign n1687 = n126 | n208 ;
  assign n1688 = n405 | n1687 ;
  assign n1689 = n1686 | n1688 ;
  assign n1690 = n413 | n443 ;
  assign n1691 = n1689 | n1690 ;
  assign n1692 = n303 | n607 ;
  assign n1693 = n128 | n310 ;
  assign n1694 = n1692 | n1693 ;
  assign n1695 = n624 | n959 ;
  assign n1696 = n175 | n1695 ;
  assign n1697 = n1694 | n1696 ;
  assign n1698 = n85 | n775 ;
  assign n1699 = n297 | n594 ;
  assign n1700 = n1698 | n1699 ;
  assign n1701 = n1697 | n1700 ;
  assign n1702 = n1691 | n1701 ;
  assign n1703 = n1685 | n1702 ;
  assign n1704 = n441 | n1521 ;
  assign n1705 = n318 | n1704 ;
  assign n1706 = n1703 | n1705 ;
  assign n1707 = n258 | n1706 ;
  assign n1708 = n1672 | n1707 ;
  assign n1709 = n1635 & n1708 ;
  assign n1710 = n1635 | n1708 ;
  assign n1711 = ~n1709 & n1710 ;
  assign n1134 = n124 | n416 ;
  assign n1135 = n71 | n1134 ;
  assign n1136 = n518 | n696 ;
  assign n1137 = n175 | n1136 ;
  assign n1138 = n1135 | n1137 ;
  assign n1139 = n128 | n349 ;
  assign n1140 = n277 | n443 ;
  assign n1141 = n1139 | n1140 ;
  assign n1142 = n577 | n1141 ;
  assign n1143 = n1138 | n1142 ;
  assign n1712 = n313 | n801 ;
  assign n1713 = n694 | n1712 ;
  assign n1714 = n198 | n555 ;
  assign n1715 = n562 | n1714 ;
  assign n1716 = n1713 | n1715 ;
  assign n1717 = n606 | n1716 ;
  assign n1718 = n1143 | n1717 ;
  assign n1719 = n374 | n643 ;
  assign n1720 = n833 | n1719 ;
  assign n1721 = n304 | n554 ;
  assign n1722 = n1720 | n1721 ;
  assign n1723 = n344 | n527 ;
  assign n1724 = n542 | n1723 ;
  assign n1725 = n142 | n330 ;
  assign n1726 = n94 | n1725 ;
  assign n1727 = n1724 | n1726 ;
  assign n1728 = n1722 | n1727 ;
  assign n1729 = n171 | n189 ;
  assign n1730 = n96 | n270 ;
  assign n1731 = n1729 | n1730 ;
  assign n1732 = n437 | n1731 ;
  assign n1733 = n1728 | n1732 ;
  assign n1734 = n1718 | n1733 ;
  assign n1735 = n160 | n269 ;
  assign n1736 = n283 | n1735 ;
  assign n1737 = n1695 | n1736 ;
  assign n1738 = n401 | n648 ;
  assign n1739 = n154 | n1738 ;
  assign n1740 = n951 | n1739 ;
  assign n1741 = n1737 | n1740 ;
  assign n1742 = n213 | n424 ;
  assign n1743 = n152 | n364 ;
  assign n1744 = n1742 | n1743 ;
  assign n1745 = n197 | n444 ;
  assign n1746 = n676 | n1745 ;
  assign n1747 = n1744 | n1746 ;
  assign n1748 = n703 | n1747 ;
  assign n1749 = n1741 | n1748 ;
  assign n1750 = n256 | n907 ;
  assign n1751 = n906 | n1750 ;
  assign n1752 = n209 | n451 ;
  assign n1753 = n46 | n431 ;
  assign n1754 = n1752 | n1753 ;
  assign n1755 = n1751 | n1754 ;
  assign n1756 = n1749 | n1755 ;
  assign n1757 = n1734 | n1756 ;
  assign n1758 = n851 | n935 ;
  assign n1759 = n1301 | n1380 ;
  assign n1760 = n297 | n1759 ;
  assign n1761 = n746 | n1760 ;
  assign n1762 = n1758 | n1761 ;
  assign n1763 = n192 | n291 ;
  assign n1764 = n469 | n594 ;
  assign n1765 = n1763 | n1764 ;
  assign n1766 = n103 | n1765 ;
  assign n1080 = n190 | n1039 ;
  assign n1767 = n764 | n1080 ;
  assign n1768 = n412 | n418 ;
  assign n1769 = n320 | n1768 ;
  assign n1770 = n1767 | n1769 ;
  assign n1771 = n99 | n193 ;
  assign n1772 = n1447 | n1771 ;
  assign n1773 = n1770 | n1772 ;
  assign n1774 = n1766 | n1773 ;
  assign n1775 = n1762 | n1774 ;
  assign n1776 = n240 | n895 ;
  assign n1777 = n602 | n1675 ;
  assign n1778 = n1608 | n1777 ;
  assign n1779 = n355 | n465 ;
  assign n1780 = n1778 | n1779 ;
  assign n1781 = n1776 | n1780 ;
  assign n1782 = n1775 | n1781 ;
  assign n1783 = n1757 | n1782 ;
  assign n1784 = n502 | n702 ;
  assign n1785 = n208 | n675 ;
  assign n1786 = n292 | n1785 ;
  assign n1787 = n1784 | n1786 ;
  assign n1074 = n233 | n479 ;
  assign n1788 = n644 | n1074 ;
  assign n1789 = n514 | n1788 ;
  assign n1790 = n1787 | n1789 ;
  assign n1791 = n184 | n413 ;
  assign n1792 = n1790 | n1791 ;
  assign n1793 = n182 | n1792 ;
  assign n1794 = n1783 | n1793 ;
  assign n1795 = n1708 & n1794 ;
  assign n1796 = n1708 | n1794 ;
  assign n1797 = ~n1795 & n1796 ;
  assign n1798 = n1795 | n1797 ;
  assign n1799 = n1711 & n1798 ;
  assign n1800 = n1711 & n1795 ;
  assign n1801 = ~n523 & n1794 ;
  assign n1802 = n523 & ~n1794 ;
  assign n1803 = n1801 | n1802 ;
  assign n1804 = n524 & ~n526 ;
  assign n1805 = n1803 | n1804 ;
  assign n1806 = ~n1801 & n1805 ;
  assign n1807 = n524 | n1803 ;
  assign n1808 = ~n1801 & n1807 ;
  assign n1809 = ( n1052 & n1806 ) | ( n1052 & n1808 ) | ( n1806 & n1808 ) ;
  assign n1810 = ( n1799 & n1800 ) | ( n1799 & ~n1809 ) | ( n1800 & ~n1809 ) ;
  assign n1811 = n1711 | n1794 ;
  assign n1812 = n1708 | n1711 ;
  assign n1813 = ( ~n1809 & n1811 ) | ( ~n1809 & n1812 ) | ( n1811 & n1812 ) ;
  assign n1814 = ~n1810 & n1813 ;
  assign n2300 = x23 & ~x24 ;
  assign n2301 = ~x23 & x24 ;
  assign n2302 = n2300 | n2301 ;
  assign n2303 = x25 & ~x26 ;
  assign n2304 = ~x25 & x26 ;
  assign n2305 = n2303 | n2304 ;
  assign n2306 = n2302 & n2305 ;
  assign n2307 = n36 & ~n62 ;
  assign n2308 = ~n2302 & n2307 ;
  assign n2371 = n1708 & n2308 ;
  assign n2311 = ~n2302 & n2305 ;
  assign n2312 = ~n2307 & n2311 ;
  assign n2372 = n1793 & n2312 ;
  assign n2373 = ( n1783 & n2312 ) | ( n1783 & n2372 ) | ( n2312 & n2372 ) ;
  assign n2315 = n2302 & ~n2305 ;
  assign n2374 = n1634 & n2315 ;
  assign n2375 = ( n1630 & n2315 ) | ( n1630 & n2374 ) | ( n2315 & n2374 ) ;
  assign n2376 = n2373 | n2375 ;
  assign n2377 = n2371 | n2376 ;
  assign n2378 = n2306 | n2377 ;
  assign n2379 = n2377 & n2378 ;
  assign n2380 = ( n1814 & n2378 ) | ( n1814 & n2379 ) | ( n2378 & n2379 ) ;
  assign n2381 = x26 & n2379 ;
  assign n2382 = x26 & n2378 ;
  assign n2383 = ( n1814 & n2381 ) | ( n1814 & n2382 ) | ( n2381 & n2382 ) ;
  assign n2384 = x26 & ~n2381 ;
  assign n2385 = x26 & ~n2382 ;
  assign n2386 = ( ~n1814 & n2384 ) | ( ~n1814 & n2385 ) | ( n2384 & n2385 ) ;
  assign n2387 = ( n2380 & ~n2383 ) | ( n2380 & n2386 ) | ( ~n2383 & n2386 ) ;
  assign n2388 = ~n2370 & n2387 ;
  assign n2389 = n2370 | n2388 ;
  assign n2390 = n2370 & n2387 ;
  assign n2391 = n2389 & ~n2390 ;
  assign n2392 = n2004 & ~n2007 ;
  assign n2393 = ~n2004 & n2007 ;
  assign n2394 = n2392 | n2393 ;
  assign n2395 = n1972 & n2394 ;
  assign n2396 = n1972 | n2394 ;
  assign n2397 = ~n2395 & n2396 ;
  assign n1880 = ( n1052 & n1805 ) | ( n1052 & n1807 ) | ( n1805 & n1807 ) ;
  assign n1881 = n1803 & n1804 ;
  assign n1882 = n524 & n1803 ;
  assign n1883 = ( n1052 & n1881 ) | ( n1052 & n1882 ) | ( n1881 & n1882 ) ;
  assign n1884 = n1880 & ~n1883 ;
  assign n2398 = ~n523 & n2308 ;
  assign n2399 = n352 & n2312 ;
  assign n2400 = ( ~n339 & n2312 ) | ( ~n339 & n2399 ) | ( n2312 & n2399 ) ;
  assign n2401 = n1793 & n2315 ;
  assign n2402 = ( n1783 & n2315 ) | ( n1783 & n2401 ) | ( n2315 & n2401 ) ;
  assign n2403 = n2400 | n2402 ;
  assign n2404 = n2398 | n2403 ;
  assign n2405 = n2306 | n2404 ;
  assign n2406 = ( n1884 & n2404 ) | ( n1884 & n2405 ) | ( n2404 & n2405 ) ;
  assign n2407 = x26 & n2405 ;
  assign n2408 = x26 & n2404 ;
  assign n2409 = ( n1884 & n2407 ) | ( n1884 & n2408 ) | ( n2407 & n2408 ) ;
  assign n2410 = x26 & ~n2407 ;
  assign n2411 = x26 & ~n2408 ;
  assign n2412 = ( ~n1884 & n2410 ) | ( ~n1884 & n2411 ) | ( n2410 & n2411 ) ;
  assign n2413 = ( n2406 & ~n2409 ) | ( n2406 & n2412 ) | ( ~n2409 & n2412 ) ;
  assign n2414 = n2397 & n2413 ;
  assign n2415 = ~n2397 & n2413 ;
  assign n2416 = ( n2397 & ~n2414 ) | ( n2397 & n2415 ) | ( ~n2414 & n2415 ) ;
  assign n2417 = ~n829 & n2312 ;
  assign n2418 = n352 & n2308 ;
  assign n2419 = ( ~n339 & n2308 ) | ( ~n339 & n2418 ) | ( n2308 & n2418 ) ;
  assign n2420 = n2417 | n2419 ;
  assign n2421 = ~n523 & n2315 ;
  assign n2422 = n2306 | n2421 ;
  assign n2423 = n2420 | n2422 ;
  assign n2424 = ~x26 & n2423 ;
  assign n2425 = n2420 | n2421 ;
  assign n2426 = ~x26 & n2425 ;
  assign n2427 = ( ~n1055 & n2424 ) | ( ~n1055 & n2426 ) | ( n2424 & n2426 ) ;
  assign n2428 = x26 & n2423 ;
  assign n2429 = x26 & ~n2428 ;
  assign n2430 = x26 & n2421 ;
  assign n2431 = ( x26 & n2420 ) | ( x26 & n2430 ) | ( n2420 & n2430 ) ;
  assign n2432 = x26 & ~n2431 ;
  assign n2433 = ( n1055 & n2429 ) | ( n1055 & n2432 ) | ( n2429 & n2432 ) ;
  assign n2434 = n2427 | n2433 ;
  assign n2435 = n1999 | n2001 ;
  assign n2436 = x29 & ~n1999 ;
  assign n2437 = ( n1982 & n2435 ) | ( n1982 & ~n2436 ) | ( n2435 & ~n2436 ) ;
  assign n2438 = ~n2004 & n2437 ;
  assign n2439 = n2434 & n2438 ;
  assign n2440 = x29 | n1996 ;
  assign n2441 = ( ~n1989 & n1996 ) | ( ~n1989 & n2440 ) | ( n1996 & n2440 ) ;
  assign n2442 = n1990 | n2441 ;
  assign n2443 = ~n1999 & n2442 ;
  assign n2444 = ~n829 & n2308 ;
  assign n2445 = n352 & n2315 ;
  assign n2446 = ( ~n339 & n2315 ) | ( ~n339 & n2445 ) | ( n2315 & n2445 ) ;
  assign n2447 = n2444 | n2446 ;
  assign n2448 = n692 & n2312 ;
  assign n2449 = ( n674 & n2312 ) | ( n674 & n2448 ) | ( n2312 & n2448 ) ;
  assign n2450 = n2447 | n2449 ;
  assign n2451 = n2306 | n2449 ;
  assign n2452 = n2447 | n2451 ;
  assign n2453 = ( ~n1209 & n2450 ) | ( ~n1209 & n2452 ) | ( n2450 & n2452 ) ;
  assign n2454 = ~x26 & n2452 ;
  assign n2455 = ~x26 & n2450 ;
  assign n2456 = ( ~n1209 & n2454 ) | ( ~n1209 & n2455 ) | ( n2454 & n2455 ) ;
  assign n2457 = x26 | n2455 ;
  assign n2458 = x26 | n2454 ;
  assign n2459 = ( ~n1209 & n2457 ) | ( ~n1209 & n2458 ) | ( n2457 & n2458 ) ;
  assign n2460 = ( ~n2453 & n2456 ) | ( ~n2453 & n2459 ) | ( n2456 & n2459 ) ;
  assign n2461 = n2443 & n2460 ;
  assign n2462 = ( ~n1027 & n1992 ) | ( ~n1027 & n1994 ) | ( n1992 & n1994 ) ;
  assign n2463 = ~n922 & n2308 ;
  assign n2464 = n1042 & n2312 ;
  assign n2465 = ( ~n1027 & n2312 ) | ( ~n1027 & n2464 ) | ( n2312 & n2464 ) ;
  assign n2466 = n2463 | n2465 ;
  assign n2467 = n692 & n2315 ;
  assign n2468 = ( n674 & n2315 ) | ( n674 & n2467 ) | ( n2315 & n2467 ) ;
  assign n2469 = n2466 | n2468 ;
  assign n2470 = ( n1538 & n2306 ) | ( n1538 & n2469 ) | ( n2306 & n2469 ) ;
  assign n2471 = ( x26 & ~n2469 ) | ( x26 & n2470 ) | ( ~n2469 & n2470 ) ;
  assign n2472 = ~n2470 & n2471 ;
  assign n2473 = ~n922 & n2315 ;
  assign n2474 = n1042 & n2308 ;
  assign n2475 = ( ~n1027 & n2308 ) | ( ~n1027 & n2474 ) | ( n2308 & n2474 ) ;
  assign n2476 = n2473 | n2475 ;
  assign n2477 = n2306 | n2475 ;
  assign n2478 = n2473 | n2477 ;
  assign n2479 = ( n1946 & n2476 ) | ( n1946 & n2478 ) | ( n2476 & n2478 ) ;
  assign n2480 = ~x26 & n2479 ;
  assign n2481 = n139 & n2302 ;
  assign n2482 = ( n1041 & n2302 ) | ( n1041 & n2481 ) | ( n2302 & n2481 ) ;
  assign n2483 = x26 & ~n2482 ;
  assign n2484 = n2302 | n2481 ;
  assign n2485 = x26 & ~n2484 ;
  assign n2486 = ( n1027 & n2483 ) | ( n1027 & n2485 ) | ( n2483 & n2485 ) ;
  assign n2487 = x26 & n2486 ;
  assign n2488 = ~n2479 & n2487 ;
  assign n2489 = ( n2480 & n2486 ) | ( n2480 & n2488 ) | ( n2486 & n2488 ) ;
  assign n2490 = x26 | n2469 ;
  assign n2491 = n2470 | n2490 ;
  assign n2492 = n2489 & n2491 ;
  assign n2493 = ~x26 & n2489 ;
  assign n2494 = ( n2472 & n2492 ) | ( n2472 & n2493 ) | ( n2492 & n2493 ) ;
  assign n2495 = n2462 & n2494 ;
  assign n2496 = n2494 & ~n2495 ;
  assign n2497 = ~n829 & n2315 ;
  assign n2498 = ~n922 & n2312 ;
  assign n2499 = n2497 | n2498 ;
  assign n2500 = n692 & n2308 ;
  assign n2501 = ( n674 & n2308 ) | ( n674 & n2500 ) | ( n2308 & n2500 ) ;
  assign n2502 = n2499 | n2501 ;
  assign n2503 = n2306 | n2501 ;
  assign n2504 = n2499 | n2503 ;
  assign n2505 = ( n1554 & n2502 ) | ( n1554 & n2504 ) | ( n2502 & n2504 ) ;
  assign n2506 = x26 & n2504 ;
  assign n2507 = x26 & n2502 ;
  assign n2508 = ( n1554 & n2506 ) | ( n1554 & n2507 ) | ( n2506 & n2507 ) ;
  assign n2509 = x26 & ~n2507 ;
  assign n2510 = x26 & ~n2506 ;
  assign n2511 = ( ~n1554 & n2509 ) | ( ~n1554 & n2510 ) | ( n2509 & n2510 ) ;
  assign n2512 = ( n2505 & ~n2508 ) | ( n2505 & n2511 ) | ( ~n2508 & n2511 ) ;
  assign n2513 = n2462 & ~n2494 ;
  assign n2514 = n2512 & n2513 ;
  assign n2515 = ( n2496 & n2512 ) | ( n2496 & n2514 ) | ( n2512 & n2514 ) ;
  assign n2516 = n2495 | n2515 ;
  assign n2517 = n2443 | n2460 ;
  assign n2518 = ~n2461 & n2517 ;
  assign n2519 = n2461 | n2518 ;
  assign n2520 = ( n2461 & n2516 ) | ( n2461 & n2519 ) | ( n2516 & n2519 ) ;
  assign n2521 = n2434 | n2438 ;
  assign n2522 = ~n2439 & n2521 ;
  assign n2523 = n2439 | n2522 ;
  assign n2524 = ( n2439 & n2520 ) | ( n2439 & n2523 ) | ( n2520 & n2523 ) ;
  assign n2525 = n2416 & n2524 ;
  assign n2526 = n2414 | n2525 ;
  assign n2527 = n1956 & n2008 ;
  assign n2528 = n1956 & ~n2527 ;
  assign n1850 = n1797 & ~n1809 ;
  assign n1851 = ~n1797 & n1809 ;
  assign n1852 = n1850 | n1851 ;
  assign n2529 = ~n523 & n2312 ;
  assign n2530 = n1793 & n2308 ;
  assign n2531 = ( n1783 & n2308 ) | ( n1783 & n2530 ) | ( n2308 & n2530 ) ;
  assign n2532 = n2529 | n2531 ;
  assign n2533 = n1708 & n2315 ;
  assign n2535 = n2306 | n2533 ;
  assign n2536 = n2532 | n2535 ;
  assign n2534 = n2532 | n2533 ;
  assign n2537 = n2534 & n2536 ;
  assign n2538 = ( ~n1852 & n2536 ) | ( ~n1852 & n2537 ) | ( n2536 & n2537 ) ;
  assign n2539 = ~x26 & n2537 ;
  assign n2540 = ~x26 & n2536 ;
  assign n2541 = ( ~n1852 & n2539 ) | ( ~n1852 & n2540 ) | ( n2539 & n2540 ) ;
  assign n2542 = x26 | n2539 ;
  assign n2543 = x26 | n2540 ;
  assign n2544 = ( ~n1852 & n2542 ) | ( ~n1852 & n2543 ) | ( n2542 & n2543 ) ;
  assign n2545 = ( ~n2538 & n2541 ) | ( ~n2538 & n2544 ) | ( n2541 & n2544 ) ;
  assign n2546 = ~n1956 & n2008 ;
  assign n2547 = n2545 & n2546 ;
  assign n2548 = ( n2528 & n2545 ) | ( n2528 & n2547 ) | ( n2545 & n2547 ) ;
  assign n2549 = n2545 | n2546 ;
  assign n2550 = n2528 | n2549 ;
  assign n2551 = ~n2548 & n2550 ;
  assign n2552 = n2548 | n2551 ;
  assign n2553 = ( n2526 & n2548 ) | ( n2526 & n2552 ) | ( n2548 & n2552 ) ;
  assign n2554 = ~n2391 & n2553 ;
  assign n2555 = n2388 | n2554 ;
  assign n2012 = n1923 | n2011 ;
  assign n1885 = ~n523 & n1823 ;
  assign n1886 = n352 & n1826 ;
  assign n1887 = ( ~n339 & n1826 ) | ( ~n339 & n1886 ) | ( n1826 & n1886 ) ;
  assign n1888 = n1793 & n1829 ;
  assign n1889 = ( n1783 & n1829 ) | ( n1783 & n1888 ) | ( n1829 & n1888 ) ;
  assign n1890 = n1887 | n1889 ;
  assign n1891 = n1885 | n1890 ;
  assign n1892 = n1821 | n1891 ;
  assign n1893 = ( n1884 & n1891 ) | ( n1884 & n1892 ) | ( n1891 & n1892 ) ;
  assign n1894 = x29 & n1892 ;
  assign n1895 = x29 & n1891 ;
  assign n1896 = ( n1884 & n1894 ) | ( n1884 & n1895 ) | ( n1894 & n1895 ) ;
  assign n1897 = x29 & ~n1894 ;
  assign n1898 = x29 & ~n1895 ;
  assign n1899 = ( ~n1884 & n1897 ) | ( ~n1884 & n1898 ) | ( n1897 & n1898 ) ;
  assign n1900 = ( n1893 & ~n1896 ) | ( n1893 & n1899 ) | ( ~n1896 & n1899 ) ;
  assign n1555 = ~n829 & n1057 ;
  assign n1556 = ~n922 & n1060 ;
  assign n1557 = n1555 | n1556 ;
  assign n1558 = n692 & n1065 ;
  assign n1559 = ( n674 & n1065 ) | ( n674 & n1558 ) | ( n1065 & n1558 ) ;
  assign n1560 = n1557 | n1559 ;
  assign n1561 = n1062 | n1559 ;
  assign n1562 = n1557 | n1561 ;
  assign n1563 = ( n1554 & n1560 ) | ( n1554 & n1562 ) | ( n1560 & n1562 ) ;
  assign n1361 = n1354 | n1360 ;
  assign n1364 = n206 | n250 ;
  assign n1365 = n171 | n202 ;
  assign n1366 = n1364 | n1365 ;
  assign n1367 = n92 | n343 ;
  assign n1368 = n1366 | n1367 ;
  assign n1369 = n395 | n477 ;
  assign n1370 = n390 | n1369 ;
  assign n1371 = n491 | n511 ;
  assign n1372 = n264 | n1371 ;
  assign n1373 = n1370 | n1372 ;
  assign n1374 = n1368 | n1373 ;
  assign n1375 = n1363 | n1374 ;
  assign n1376 = n615 | n1375 ;
  assign n1377 = n1361 | n1376 ;
  assign n1378 = n39 | n437 ;
  assign n1379 = n518 | n1378 ;
  assign n1381 = n85 | n228 ;
  assign n1382 = n1380 | n1381 ;
  assign n1383 = n76 | n1382 ;
  assign n1384 = n155 | n588 ;
  assign n1385 = n441 | n959 ;
  assign n1386 = n280 | n501 ;
  assign n1387 = n1385 | n1386 ;
  assign n1388 = n1384 | n1387 ;
  assign n1389 = n1383 | n1388 ;
  assign n1390 = n382 | n849 ;
  assign n1391 = n1389 | n1390 ;
  assign n1392 = n246 | n401 ;
  assign n1393 = n196 | n1392 ;
  assign n1394 = n321 | n451 ;
  assign n1395 = n661 | n1394 ;
  assign n1396 = n1393 | n1395 ;
  assign n1397 = n305 | n487 ;
  assign n1398 = n689 | n887 ;
  assign n1399 = n143 & ~n644 ;
  assign n1400 = ~n1398 & n1399 ;
  assign n1401 = ~n1397 & n1400 ;
  assign n1402 = ~n1396 & n1401 ;
  assign n1403 = n763 | n1301 ;
  assign n1404 = n340 | n566 ;
  assign n1405 = n124 | n1404 ;
  assign n1406 = n1403 | n1405 ;
  assign n1407 = n310 | n638 ;
  assign n1408 = n1406 | n1407 ;
  assign n1409 = n1402 & ~n1408 ;
  assign n1410 = ~n1391 & n1409 ;
  assign n1411 = ~n1379 & n1410 ;
  assign n1412 = n94 | n364 ;
  assign n1413 = n224 | n1412 ;
  assign n1414 = n183 | n820 ;
  assign n1415 = n355 | n1414 ;
  assign n1416 = n1413 | n1415 ;
  assign n1417 = n131 | n272 ;
  assign n1418 = n476 | n1417 ;
  assign n1419 = n411 | n1418 ;
  assign n1420 = n1416 | n1419 ;
  assign n1421 = n160 | n468 ;
  assign n1422 = n312 | n1421 ;
  assign n1423 = n895 | n1422 ;
  assign n1424 = n624 | n1423 ;
  assign n1425 = n1420 | n1424 ;
  assign n1426 = n1411 & ~n1425 ;
  assign n1427 = ~n1377 & n1426 ;
  assign n1428 = ~n332 & n1427 ;
  assign n1534 = n1428 | n1533 ;
  assign n1552 = ~n1534 & n1551 ;
  assign n1564 = n1428 & n1533 ;
  assign n1565 = ( n1428 & ~n1551 ) | ( n1428 & n1564 ) | ( ~n1551 & n1564 ) ;
  assign n1566 = n1552 | n1565 ;
  assign n1567 = n1563 & ~n1566 ;
  assign n1877 = n1563 & ~n1567 ;
  assign n1878 = n1566 | n1567 ;
  assign n1879 = ~n1877 & n1878 ;
  assign n1901 = ~n1879 & n1900 ;
  assign n2013 = n1900 & ~n1901 ;
  assign n2014 = n1879 | n1900 ;
  assign n2015 = ~n2013 & n2014 ;
  assign n2336 = n2012 & ~n2015 ;
  assign n2337 = ~n2012 & n2015 ;
  assign n2338 = n2336 | n2337 ;
  assign n2023 = n151 | n839 ;
  assign n2204 = n437 | n676 ;
  assign n2205 = n2023 | n2204 ;
  assign n2206 = n880 | n2205 ;
  assign n2207 = n383 | n667 ;
  assign n2208 = n381 | n555 ;
  assign n2209 = n2207 | n2208 ;
  assign n2210 = n155 | n513 ;
  assign n2211 = n2209 | n2210 ;
  assign n2212 = n2206 | n2211 ;
  assign n2213 = n1458 & ~n2212 ;
  assign n2214 = n196 | n841 ;
  assign n2215 = n340 | n574 ;
  assign n2216 = n261 | n1039 ;
  assign n2217 = n1005 | n2216 ;
  assign n2218 = n2215 | n2217 ;
  assign n2219 = n152 | n588 ;
  assign n2220 = n363 | n372 ;
  assign n2221 = n2219 | n2220 ;
  assign n2222 = n436 | n2221 ;
  assign n2223 = n2218 | n2222 ;
  assign n2224 = n2214 | n2223 ;
  assign n2225 = n602 | n648 ;
  assign n2226 = n387 | n959 ;
  assign n2227 = n2225 | n2226 ;
  assign n2228 = n163 | n384 ;
  assign n2229 = n762 | n2228 ;
  assign n2230 = n2227 | n2229 ;
  assign n2231 = n411 | n1114 ;
  assign n2232 = n2230 | n2231 ;
  assign n2233 = n643 | n666 ;
  assign n2234 = n1349 | n2233 ;
  assign n2235 = n178 | n236 ;
  assign n2236 = n820 | n2235 ;
  assign n2237 = n2234 | n2236 ;
  assign n2238 = n189 | n355 ;
  assign n2239 = n2237 | n2238 ;
  assign n2240 = n2232 | n2239 ;
  assign n2241 = n2224 | n2240 ;
  assign n2242 = n2213 & ~n2241 ;
  assign n2243 = n53 | n222 ;
  assign n2244 = n94 | n2243 ;
  assign n2245 = n64 | n895 ;
  assign n2246 = n923 | n2245 ;
  assign n2247 = n2244 | n2246 ;
  assign n2248 = n432 | n590 ;
  assign n2249 = n749 | n2248 ;
  assign n2250 = n1771 | n2249 ;
  assign n2251 = n2247 | n2250 ;
  assign n2117 = n450 | n638 ;
  assign n2252 = n1785 | n2117 ;
  assign n2253 = n318 | n1172 ;
  assign n2254 = n254 | n2253 ;
  assign n2255 = n2252 | n2254 ;
  assign n1163 = n112 | n162 ;
  assign n1164 = n245 | n1163 ;
  assign n2256 = n139 | n234 ;
  assign n2257 = n1164 | n2256 ;
  assign n2258 = n2255 | n2257 ;
  assign n2259 = n2251 | n2258 ;
  assign n2260 = n79 | n85 ;
  assign n2261 = n979 | n2260 ;
  assign n2262 = n321 | n401 ;
  assign n2263 = n2261 | n2262 ;
  assign n2264 = n495 | n2263 ;
  assign n2265 = n2259 | n2264 ;
  assign n2050 = n75 | n456 ;
  assign n2266 = n527 | n2050 ;
  assign n2267 = n1484 | n2266 ;
  assign n2268 = n2265 | n2267 ;
  assign n2269 = n2242 & ~n2268 ;
  assign n2270 = n225 | n332 ;
  assign n2271 = n88 | n124 ;
  assign n2272 = n442 | n2271 ;
  assign n2273 = n46 | n213 ;
  assign n2274 = n510 | n2273 ;
  assign n2275 = n2272 | n2274 ;
  assign n2276 = n59 | n183 ;
  assign n2277 = n118 | n2276 ;
  assign n2278 = n2275 | n2277 ;
  assign n2279 = n2270 | n2278 ;
  assign n2280 = n2269 & ~n2279 ;
  assign n2285 = n1635 & ~n2280 ;
  assign n2286 = ~n1635 & n2280 ;
  assign n2287 = n2285 | n2286 ;
  assign n2288 = n1709 | n1711 ;
  assign n2289 = ( n1709 & n1798 ) | ( n1709 & n2288 ) | ( n1798 & n2288 ) ;
  assign n2290 = ~n2287 & n2289 ;
  assign n2294 = n1709 | n1795 ;
  assign n2295 = ( n1709 & n1711 ) | ( n1709 & n2294 ) | ( n1711 & n2294 ) ;
  assign n2296 = ~n2287 & n2295 ;
  assign n2339 = ( ~n1809 & n2290 ) | ( ~n1809 & n2296 ) | ( n2290 & n2296 ) ;
  assign n2340 = n2287 & ~n2289 ;
  assign n2341 = n2287 & ~n2295 ;
  assign n2342 = ( n1809 & n2340 ) | ( n1809 & n2341 ) | ( n2340 & n2341 ) ;
  assign n2343 = n2339 | n2342 ;
  assign n2344 = n1708 & n2312 ;
  assign n2345 = n1634 & n2308 ;
  assign n2346 = ( n1630 & n2308 ) | ( n1630 & n2345 ) | ( n2308 & n2345 ) ;
  assign n2347 = n2279 & n2315 ;
  assign n2348 = n2306 | n2347 ;
  assign n2349 = n2306 | n2315 ;
  assign n2350 = ( ~n2269 & n2348 ) | ( ~n2269 & n2349 ) | ( n2348 & n2349 ) ;
  assign n2351 = n2346 | n2350 ;
  assign n2352 = n2344 | n2351 ;
  assign n2353 = ( ~n2269 & n2315 ) | ( ~n2269 & n2347 ) | ( n2315 & n2347 ) ;
  assign n2354 = n2346 | n2353 ;
  assign n2355 = n2344 | n2354 ;
  assign n2356 = n2352 & n2355 ;
  assign n2357 = ( ~n2343 & n2352 ) | ( ~n2343 & n2356 ) | ( n2352 & n2356 ) ;
  assign n2358 = ~x26 & n2356 ;
  assign n2359 = ~x26 & n2352 ;
  assign n2360 = ( ~n2343 & n2358 ) | ( ~n2343 & n2359 ) | ( n2358 & n2359 ) ;
  assign n2361 = x26 | n2358 ;
  assign n2362 = x26 | n2359 ;
  assign n2363 = ( ~n2343 & n2361 ) | ( ~n2343 & n2362 ) | ( n2361 & n2362 ) ;
  assign n2364 = ( ~n2357 & n2360 ) | ( ~n2357 & n2363 ) | ( n2360 & n2363 ) ;
  assign n2365 = ~n2338 & n2364 ;
  assign n2366 = n2338 | n2365 ;
  assign n2367 = n2338 & n2364 ;
  assign n2368 = n2366 & ~n2367 ;
  assign n2556 = ~n2368 & n2555 ;
  assign n2980 = n2555 & ~n2556 ;
  assign n2981 = n2368 | n2556 ;
  assign n2982 = ~n2980 & n2981 ;
  assign n2024 = n142 | n435 ;
  assign n2025 = n2023 | n2024 ;
  assign n1286 = n212 | n895 ;
  assign n2026 = n858 | n1286 ;
  assign n2027 = n2025 | n2026 ;
  assign n2028 = n441 | n574 ;
  assign n2029 = n128 | n675 ;
  assign n2030 = n2028 | n2029 ;
  assign n2031 = ( ~n428 & n2027 ) | ( ~n428 & n2030 ) | ( n2027 & n2030 ) ;
  assign n2032 = n164 | n682 ;
  assign n2033 = n143 & ~n2032 ;
  assign n2034 = ~n428 & n2033 ;
  assign n2035 = ~n2031 & n2034 ;
  assign n2036 = n355 | n458 ;
  assign n2037 = n1028 | n1465 ;
  assign n2038 = n637 | n2037 ;
  assign n2039 = n179 | n511 ;
  assign n2040 = n182 | n2039 ;
  assign n2041 = n551 | n2040 ;
  assign n2042 = n2038 | n2041 ;
  assign n2043 = n317 | n901 ;
  assign n2044 = n263 | n2043 ;
  assign n2045 = n2042 | n2044 ;
  assign n1150 = n139 | n208 ;
  assign n1151 = n280 | n1150 ;
  assign n2046 = n1151 | n1342 ;
  assign n2047 = n332 | n500 ;
  assign n2048 = n1436 | n2047 ;
  assign n2049 = n2046 | n2048 ;
  assign n2051 = n71 | n607 ;
  assign n2052 = n2050 | n2051 ;
  assign n2053 = n131 | n775 ;
  assign n2054 = n54 | n2053 ;
  assign n2055 = n2052 | n2054 ;
  assign n2056 = n205 | n591 ;
  assign n2057 = n2055 | n2056 ;
  assign n2058 = n2049 | n2057 ;
  assign n2059 = n2045 | n2058 ;
  assign n2060 = n2036 | n2059 ;
  assign n2061 = n333 | n461 ;
  assign n2062 = n347 | n2061 ;
  assign n2063 = n581 | n667 ;
  assign n2064 = n141 | n2063 ;
  assign n2065 = n2062 | n2064 ;
  assign n2066 = n262 | n348 ;
  assign n2067 = n1714 | n2066 ;
  assign n2068 = n980 | n2067 ;
  assign n2069 = n2065 | n2068 ;
  assign n2070 = n99 | n638 ;
  assign n2071 = n309 | n431 ;
  assign n2072 = n2070 | n2071 ;
  assign n2073 = n254 | n2072 ;
  assign n2074 = n577 | n2073 ;
  assign n2075 = n2069 | n2074 ;
  assign n2076 = n118 | n711 ;
  assign n2077 = n1501 | n2076 ;
  assign n2078 = n274 | n2077 ;
  assign n2079 = n608 | n2078 ;
  assign n2080 = n2075 | n2079 ;
  assign n2081 = n2060 | n2080 ;
  assign n2082 = n2035 & ~n2081 ;
  assign n2083 = n236 | n450 ;
  assign n2084 = n117 | n820 ;
  assign n2085 = n2083 | n2084 ;
  assign n2086 = n320 | n666 ;
  assign n2087 = n432 | n2086 ;
  assign n2088 = n2085 | n2087 ;
  assign n2089 = n103 | n624 ;
  assign n2090 = n2088 | n2089 ;
  assign n2091 = n2082 & ~n2090 ;
  assign n2092 = n950 | n1771 ;
  assign n2093 = n479 | n483 ;
  assign n2094 = n311 | n2093 ;
  assign n2095 = n331 | n676 ;
  assign n2096 = n2094 | n2095 ;
  assign n2097 = n2092 | n2096 ;
  assign n2098 = n679 | n2097 ;
  assign n2099 = n542 | n631 ;
  assign n2100 = n447 | n2099 ;
  assign n1115 = n458 | n1114 ;
  assign n2101 = n399 | n1115 ;
  assign n2102 = n2100 | n2101 ;
  assign n2103 = n198 | n203 ;
  assign n2104 = n269 | n581 ;
  assign n2105 = n272 | n435 ;
  assign n2106 = n2104 | n2105 ;
  assign n2107 = n2103 | n2106 ;
  assign n2108 = n2102 | n2107 ;
  assign n2109 = n88 | n480 ;
  assign n2110 = n54 | n2109 ;
  assign n2111 = n388 | n418 ;
  assign n2112 = n128 | n2111 ;
  assign n2113 = n2110 | n2112 ;
  assign n2114 = n2108 | n2113 ;
  assign n2115 = n2098 | n2114 ;
  assign n2116 = n197 | n434 ;
  assign n2118 = n952 | n2117 ;
  assign n2119 = n405 | n2118 ;
  assign n2120 = n131 | n1039 ;
  assign n2121 = n71 | n491 ;
  assign n2122 = n2120 | n2121 ;
  assign n2123 = n249 | n277 ;
  assign n2124 = n2122 | n2123 ;
  assign n2125 = n2119 | n2124 ;
  assign n2126 = n2116 | n2125 ;
  assign n2127 = n134 | n138 ;
  assign n2128 = n75 | n2127 ;
  assign n2129 = n64 | n461 ;
  assign n2130 = n636 | n2129 ;
  assign n2131 = n2128 | n2130 ;
  assign n2132 = n256 | n711 ;
  assign n2133 = n317 | n2132 ;
  assign n2134 = n2131 | n2133 ;
  assign n2135 = n168 | n644 ;
  assign n2136 = n291 | n402 ;
  assign n2137 = n324 | n443 ;
  assign n2138 = n2136 | n2137 ;
  assign n2139 = n2135 | n2138 ;
  assign n2140 = n2134 | n2139 ;
  assign n2141 = n2126 | n2140 ;
  assign n2142 = n2115 | n2141 ;
  assign n2143 = n510 | n959 ;
  assign n2144 = n1657 | n2143 ;
  assign n2145 = n143 & ~n2144 ;
  assign n2146 = n126 | n292 ;
  assign n2147 = n114 | n468 ;
  assign n2148 = n939 | n2147 ;
  assign n2149 = n205 | n2148 ;
  assign n2150 = ( n2145 & n2146 ) | ( n2145 & n2149 ) | ( n2146 & n2149 ) ;
  assign n2151 = n372 | n689 ;
  assign n2152 = n867 | n2151 ;
  assign n2153 = n184 | n2152 ;
  assign n2154 = n2145 & ~n2153 ;
  assign n2155 = ~n2150 & n2154 ;
  assign n2156 = n59 | n469 ;
  assign n2157 = n561 | n2156 ;
  assign n2158 = n142 | n456 ;
  assign n2159 = n325 | n2158 ;
  assign n2160 = n2157 | n2159 ;
  assign n2161 = n349 | n2160 ;
  assign n2162 = n118 | n222 ;
  assign n2163 = n895 | n2162 ;
  assign n2164 = n779 | n2163 ;
  assign n2165 = n179 | n457 ;
  assign n2166 = n94 | n527 ;
  assign n2167 = n2165 | n2166 ;
  assign n2168 = n1239 | n2167 ;
  assign n2169 = n2164 | n2168 ;
  assign n2170 = n2161 | n2169 ;
  assign n2171 = n2155 & ~n2170 ;
  assign n2172 = n178 | n261 ;
  assign n2173 = n167 | n247 ;
  assign n2174 = n2172 | n2173 ;
  assign n2175 = n297 | n696 ;
  assign n2176 = n501 | n2175 ;
  assign n2177 = n2174 | n2176 ;
  assign n2178 = n283 | n694 ;
  assign n2179 = n2177 | n2178 ;
  assign n2180 = n96 | n250 ;
  assign n2181 = n390 | n568 ;
  assign n2182 = n2180 | n2181 ;
  assign n2183 = n2179 | n2182 ;
  assign n2184 = n2171 & ~n2183 ;
  assign n2185 = ~n2142 & n2184 ;
  assign n2186 = n347 | n432 ;
  assign n2187 = n758 | n2186 ;
  assign n2188 = n330 | n383 ;
  assign n2189 = n1031 | n2188 ;
  assign n2190 = n235 | n979 ;
  assign n2191 = n2189 | n2190 ;
  assign n2192 = n117 | n518 ;
  assign n2193 = n608 | n2192 ;
  assign n2194 = n176 | n2193 ;
  assign n2195 = n2191 | n2194 ;
  assign n2196 = n262 | n725 ;
  assign n2197 = n616 | n2196 ;
  assign n2198 = n2195 | n2197 ;
  assign n2199 = n2187 | n2198 ;
  assign n2200 = n2185 & ~n2199 ;
  assign n2201 = n2091 | n2200 ;
  assign n2281 = n2091 | n2280 ;
  assign n2282 = n2091 & n2280 ;
  assign n2283 = n2281 & ~n2282 ;
  assign n2291 = n2281 & ~n2285 ;
  assign n2292 = ( n2281 & ~n2283 ) | ( n2281 & n2291 ) | ( ~n2283 & n2291 ) ;
  assign n2202 = n2091 & n2200 ;
  assign n2203 = n2201 & ~n2202 ;
  assign n2597 = n2201 & ~n2203 ;
  assign n2598 = ( n2201 & n2292 ) | ( n2201 & n2597 ) | ( n2292 & n2597 ) ;
  assign n2284 = n2281 & ~n2283 ;
  assign n2599 = ( n2201 & n2284 ) | ( n2201 & n2597 ) | ( n2284 & n2597 ) ;
  assign n2600 = ( ~n2290 & n2598 ) | ( ~n2290 & n2599 ) | ( n2598 & n2599 ) ;
  assign n2601 = ( ~n2296 & n2598 ) | ( ~n2296 & n2599 ) | ( n2598 & n2599 ) ;
  assign n2602 = ( n1809 & n2600 ) | ( n1809 & n2601 ) | ( n2600 & n2601 ) ;
  assign n2603 = n151 | n383 ;
  assign n2604 = n577 | n2603 ;
  assign n2605 = n171 | n227 ;
  assign n2606 = n2604 | n2605 ;
  assign n2607 = n96 | n594 ;
  assign n2608 = n184 | n2607 ;
  assign n2609 = n2606 | n2608 ;
  assign n2610 = n162 | n175 ;
  assign n2611 = n330 | n384 ;
  assign n2612 = n2610 | n2611 ;
  assign n2613 = n340 | n2612 ;
  assign n2614 = n176 | n648 ;
  assign n2615 = n1662 | n2614 ;
  assign n2616 = n128 | n2615 ;
  assign n2617 = n46 | n59 ;
  assign n2618 = n229 | n2617 ;
  assign n2619 = n2062 | n2618 ;
  assign n2620 = n2616 | n2619 ;
  assign n2621 = n2613 | n2620 ;
  assign n2622 = n2609 | n2621 ;
  assign n2623 = n414 | n623 ;
  assign n2624 = n222 | n281 ;
  assign n2625 = n198 | n2624 ;
  assign n2626 = n2623 | n2625 ;
  assign n2627 = n389 | n2626 ;
  assign n2628 = n1582 | n1584 ;
  assign n2629 = n2627 | n2628 ;
  assign n2630 = n312 | n991 ;
  assign n2631 = n168 | n1355 ;
  assign n2632 = n2630 | n2631 ;
  assign n2633 = n154 | n694 ;
  assign n2634 = n152 | n1039 ;
  assign n2635 = n206 | n607 ;
  assign n2636 = n2634 | n2635 ;
  assign n2637 = n2633 | n2636 ;
  assign n2638 = n2632 | n2637 ;
  assign n2639 = n306 | n402 ;
  assign n2640 = n806 | n858 ;
  assign n2641 = n2639 | n2640 ;
  assign n2642 = n257 | n320 ;
  assign n2643 = n160 | n2642 ;
  assign n2644 = n2641 | n2643 ;
  assign n2645 = n758 | n2053 ;
  assign n2646 = n406 | n2645 ;
  assign n2647 = n2644 | n2646 ;
  assign n2648 = n2638 | n2647 ;
  assign n2649 = n2629 | n2648 ;
  assign n2650 = n2622 | n2649 ;
  assign n2651 = n114 | n631 ;
  assign n1075 = n237 | n511 ;
  assign n1076 = n1074 | n1075 ;
  assign n1077 = n500 | n1076 ;
  assign n2652 = n369 | n720 ;
  assign n2653 = n600 | n2652 ;
  assign n2654 = n935 | n2653 ;
  assign n2655 = n1077 | n2654 ;
  assign n2656 = n588 | n839 ;
  assign n2657 = n2214 | n2656 ;
  assign n2658 = n39 | n213 ;
  assign n2659 = n118 | n2658 ;
  assign n2660 = n2657 | n2659 ;
  assign n2661 = n250 | n513 ;
  assign n2662 = n448 | n2661 ;
  assign n2663 = n2660 | n2662 ;
  assign n2664 = n2655 | n2663 ;
  assign n2665 = n270 | n491 ;
  assign n2666 = n590 | n2665 ;
  assign n2667 = n419 | n1657 ;
  assign n2668 = n2666 | n2667 ;
  assign n2669 = n697 | n2668 ;
  assign n2670 = n460 | n959 ;
  assign n2671 = n71 | n725 ;
  assign n2672 = n2670 | n2671 ;
  assign n2673 = n273 | n395 ;
  assign n2674 = n2672 | n2673 ;
  assign n2675 = n2669 | n2674 ;
  assign n2676 = n2664 | n2675 ;
  assign n2677 = n2651 | n2676 ;
  assign n2678 = n2650 | n2677 ;
  assign n2679 = n436 | n1336 ;
  assign n2680 = n140 | n503 ;
  assign n2681 = n2679 | n2680 ;
  assign n2682 = n363 | n497 ;
  assign n2683 = n2681 | n2682 ;
  assign n2684 = n849 | n1623 ;
  assign n2685 = n1580 | n2684 ;
  assign n2686 = n2683 | n2685 ;
  assign n2687 = n94 | n189 ;
  assign n2688 = n79 | n2687 ;
  assign n2689 = n644 | n2688 ;
  assign n2690 = n2686 | n2689 ;
  assign n2691 = n104 | n2690 ;
  assign n2692 = n2678 | n2691 ;
  assign n2693 = ~n2200 & n2692 ;
  assign n2694 = n2200 & ~n2692 ;
  assign n2695 = n2693 | n2694 ;
  assign n2983 = n2602 | n2695 ;
  assign n2984 = n2602 & n2695 ;
  assign n2985 = n2983 & ~n2984 ;
  assign n2915 = ~x21 & x22 ;
  assign n2916 = x21 & ~x22 ;
  assign n2917 = n2915 | n2916 ;
  assign n2918 = x20 & ~x21 ;
  assign n2919 = ~x20 & x21 ;
  assign n2920 = n2918 | n2919 ;
  assign n2921 = ~x22 & x23 ;
  assign n2922 = x22 & ~x23 ;
  assign n2923 = n2921 | n2922 ;
  assign n2924 = ~n2920 & n2923 ;
  assign n2925 = ~n2917 & n2924 ;
  assign n2986 = n2090 & n2925 ;
  assign n2987 = ( ~n2082 & n2925 ) | ( ~n2082 & n2986 ) | ( n2925 & n2986 ) ;
  assign n2932 = n2920 & ~n2923 ;
  assign n2988 = n2691 & n2932 ;
  assign n2989 = ( n2678 & n2932 ) | ( n2678 & n2988 ) | ( n2932 & n2988 ) ;
  assign n2928 = n2917 & ~n2920 ;
  assign n2990 = n2199 & n2928 ;
  assign n2991 = ( ~n2185 & n2928 ) | ( ~n2185 & n2990 ) | ( n2928 & n2990 ) ;
  assign n2992 = n2989 | n2991 ;
  assign n2993 = n2987 | n2992 ;
  assign n2936 = n2920 & n2923 ;
  assign n2994 = n2936 | n2993 ;
  assign n2995 = ( n2985 & n2993 ) | ( n2985 & n2994 ) | ( n2993 & n2994 ) ;
  assign n2996 = x23 & n2994 ;
  assign n2997 = x23 & n2993 ;
  assign n2998 = ( n2985 & n2996 ) | ( n2985 & n2997 ) | ( n2996 & n2997 ) ;
  assign n2999 = x23 & ~n2996 ;
  assign n3000 = x23 & ~n2997 ;
  assign n3001 = ( ~n2985 & n2999 ) | ( ~n2985 & n3000 ) | ( n2999 & n3000 ) ;
  assign n3002 = ( n2995 & ~n2998 ) | ( n2995 & n3001 ) | ( ~n2998 & n3001 ) ;
  assign n3003 = ~n2982 & n3002 ;
  assign n3004 = n2982 | n3003 ;
  assign n3005 = n2982 & n3002 ;
  assign n3006 = n3004 & ~n3005 ;
  assign n3007 = n2391 | n2553 ;
  assign n3008 = n2391 & n2553 ;
  assign n3009 = n3007 & ~n3008 ;
  assign n2293 = ( n2284 & ~n2290 ) | ( n2284 & n2292 ) | ( ~n2290 & n2292 ) ;
  assign n2297 = ( n2284 & n2292 ) | ( n2284 & ~n2296 ) | ( n2292 & ~n2296 ) ;
  assign n2298 = ( n1809 & n2293 ) | ( n1809 & n2297 ) | ( n2293 & n2297 ) ;
  assign n2299 = ~n2203 & n2298 ;
  assign n2321 = n2203 & ~n2292 ;
  assign n2322 = n2203 & ~n2284 ;
  assign n2323 = ( n2290 & n2321 ) | ( n2290 & n2322 ) | ( n2321 & n2322 ) ;
  assign n2324 = ( n2296 & n2321 ) | ( n2296 & n2322 ) | ( n2321 & n2322 ) ;
  assign n2325 = ( ~n1809 & n2323 ) | ( ~n1809 & n2324 ) | ( n2323 & n2324 ) ;
  assign n3010 = n2090 & n2928 ;
  assign n3011 = ( ~n2082 & n2928 ) | ( ~n2082 & n3010 ) | ( n2928 & n3010 ) ;
  assign n3012 = n2279 & n2925 ;
  assign n3013 = ( ~n2269 & n2925 ) | ( ~n2269 & n3012 ) | ( n2925 & n3012 ) ;
  assign n3014 = n2199 & n2932 ;
  assign n3015 = ( ~n2185 & n2932 ) | ( ~n2185 & n3014 ) | ( n2932 & n3014 ) ;
  assign n3016 = n3013 | n3015 ;
  assign n3017 = n3011 | n3016 ;
  assign n3018 = n2936 | n3017 ;
  assign n3019 = ( ~n2325 & n3017 ) | ( ~n2325 & n3018 ) | ( n3017 & n3018 ) ;
  assign n3020 = n3017 & n3018 ;
  assign n3021 = ( ~n2299 & n3019 ) | ( ~n2299 & n3020 ) | ( n3019 & n3020 ) ;
  assign n3022 = ~x23 & n3021 ;
  assign n3023 = x23 | n3021 ;
  assign n3024 = ( ~n3021 & n3022 ) | ( ~n3021 & n3023 ) | ( n3022 & n3023 ) ;
  assign n3025 = ~n3009 & n3024 ;
  assign n3026 = n2526 & n2551 ;
  assign n3027 = n2526 & ~n3026 ;
  assign n3028 = ~n2526 & n2551 ;
  assign n3029 = n3027 | n3028 ;
  assign n2560 = n2283 & n2285 ;
  assign n2561 = ( n2283 & n2290 ) | ( n2283 & n2560 ) | ( n2290 & n2560 ) ;
  assign n2562 = ( n2283 & n2296 ) | ( n2283 & n2560 ) | ( n2296 & n2560 ) ;
  assign n2563 = ( ~n1809 & n2561 ) | ( ~n1809 & n2562 ) | ( n2561 & n2562 ) ;
  assign n2564 = n2283 | n2285 ;
  assign n2565 = n2290 | n2564 ;
  assign n2566 = n2296 | n2564 ;
  assign n2567 = ( ~n1809 & n2565 ) | ( ~n1809 & n2566 ) | ( n2565 & n2566 ) ;
  assign n2568 = ~n2563 & n2567 ;
  assign n3030 = n1634 & n2925 ;
  assign n3031 = ( n1630 & n2925 ) | ( n1630 & n3030 ) | ( n2925 & n3030 ) ;
  assign n3032 = n2279 & n2928 ;
  assign n3033 = ( ~n2269 & n2928 ) | ( ~n2269 & n3032 ) | ( n2928 & n3032 ) ;
  assign n3034 = n3031 | n3033 ;
  assign n3035 = n2090 & n2932 ;
  assign n3036 = ( ~n2082 & n2932 ) | ( ~n2082 & n3035 ) | ( n2932 & n3035 ) ;
  assign n3037 = n3034 | n3036 ;
  assign n3038 = n2936 | n3037 ;
  assign n3039 = ( n2568 & n3037 ) | ( n2568 & n3038 ) | ( n3037 & n3038 ) ;
  assign n3040 = x23 & n3038 ;
  assign n3041 = x23 & n3037 ;
  assign n3042 = ( n2568 & n3040 ) | ( n2568 & n3041 ) | ( n3040 & n3041 ) ;
  assign n3043 = x23 & ~n3040 ;
  assign n3044 = x23 & ~n3041 ;
  assign n3045 = ( ~n2568 & n3043 ) | ( ~n2568 & n3044 ) | ( n3043 & n3044 ) ;
  assign n3046 = ( n3039 & ~n3042 ) | ( n3039 & n3045 ) | ( ~n3042 & n3045 ) ;
  assign n3047 = n3028 & n3046 ;
  assign n3048 = ( n3027 & n3046 ) | ( n3027 & n3047 ) | ( n3046 & n3047 ) ;
  assign n3049 = n3029 & ~n3048 ;
  assign n3050 = n2416 | n2524 ;
  assign n3051 = ~n2525 & n3050 ;
  assign n3052 = n1708 & n2925 ;
  assign n3053 = n1634 & n2928 ;
  assign n3054 = ( n1630 & n2928 ) | ( n1630 & n3053 ) | ( n2928 & n3053 ) ;
  assign n3055 = n2279 & n2932 ;
  assign n3056 = ( ~n2269 & n2932 ) | ( ~n2269 & n3055 ) | ( n2932 & n3055 ) ;
  assign n3057 = n3054 | n3056 ;
  assign n3058 = n3052 | n3057 ;
  assign n3059 = n2936 | n3058 ;
  assign n3060 = n3058 & n3059 ;
  assign n3061 = ( ~n2343 & n3059 ) | ( ~n2343 & n3060 ) | ( n3059 & n3060 ) ;
  assign n3062 = ~x23 & n3060 ;
  assign n3063 = ~x23 & n3059 ;
  assign n3064 = ( ~n2343 & n3062 ) | ( ~n2343 & n3063 ) | ( n3062 & n3063 ) ;
  assign n3065 = x23 | n3062 ;
  assign n3066 = x23 | n3063 ;
  assign n3067 = ( ~n2343 & n3065 ) | ( ~n2343 & n3066 ) | ( n3065 & n3066 ) ;
  assign n3068 = ( ~n3061 & n3064 ) | ( ~n3061 & n3067 ) | ( n3064 & n3067 ) ;
  assign n3069 = n3051 & n3068 ;
  assign n3070 = n3051 | n3068 ;
  assign n3071 = ~n3069 & n3070 ;
  assign n3072 = n2516 & n2518 ;
  assign n3073 = n2516 | n2518 ;
  assign n3074 = ~n3072 & n3073 ;
  assign n3075 = ~n523 & n2925 ;
  assign n3076 = n1793 & n2928 ;
  assign n3077 = ( n1783 & n2928 ) | ( n1783 & n3076 ) | ( n2928 & n3076 ) ;
  assign n3078 = n3075 | n3077 ;
  assign n3079 = n1708 & n2932 ;
  assign n3080 = n3078 | n3079 ;
  assign n3081 = n2936 | n3079 ;
  assign n3082 = n3078 | n3081 ;
  assign n3083 = ( ~n1852 & n3080 ) | ( ~n1852 & n3082 ) | ( n3080 & n3082 ) ;
  assign n3084 = ~x23 & n3082 ;
  assign n3085 = ~x23 & n3080 ;
  assign n3086 = ( ~n1852 & n3084 ) | ( ~n1852 & n3085 ) | ( n3084 & n3085 ) ;
  assign n3087 = x23 | n3085 ;
  assign n3088 = x23 | n3084 ;
  assign n3089 = ( ~n1852 & n3087 ) | ( ~n1852 & n3088 ) | ( n3087 & n3088 ) ;
  assign n3090 = ( ~n3083 & n3086 ) | ( ~n3083 & n3089 ) | ( n3086 & n3089 ) ;
  assign n3091 = n3074 & n3090 ;
  assign n3092 = n2512 | n2513 ;
  assign n3093 = n2496 | n3092 ;
  assign n3094 = ~n2515 & n3093 ;
  assign n3095 = ~n523 & n2928 ;
  assign n3096 = n352 & n2925 ;
  assign n3097 = ( ~n339 & n2925 ) | ( ~n339 & n3096 ) | ( n2925 & n3096 ) ;
  assign n3098 = n1793 & n2932 ;
  assign n3099 = ( n1783 & n2932 ) | ( n1783 & n3098 ) | ( n2932 & n3098 ) ;
  assign n3100 = n3097 | n3099 ;
  assign n3101 = n3095 | n3100 ;
  assign n3102 = n2936 | n3101 ;
  assign n3103 = n3101 & n3102 ;
  assign n3104 = ( n1884 & n3102 ) | ( n1884 & n3103 ) | ( n3102 & n3103 ) ;
  assign n3105 = x23 & n3103 ;
  assign n3106 = x23 & n3102 ;
  assign n3107 = ( n1884 & n3105 ) | ( n1884 & n3106 ) | ( n3105 & n3106 ) ;
  assign n3108 = x23 & ~n3105 ;
  assign n3109 = x23 & ~n3106 ;
  assign n3110 = ( ~n1884 & n3108 ) | ( ~n1884 & n3109 ) | ( n3108 & n3109 ) ;
  assign n3111 = ( n3104 & ~n3107 ) | ( n3104 & n3110 ) | ( ~n3107 & n3110 ) ;
  assign n3112 = n3094 & n3111 ;
  assign n3113 = n3094 | n3111 ;
  assign n3114 = ~n3112 & n3113 ;
  assign n3115 = ~n829 & n2925 ;
  assign n3116 = n352 & n2928 ;
  assign n3117 = ( ~n339 & n2928 ) | ( ~n339 & n3116 ) | ( n2928 & n3116 ) ;
  assign n3118 = n3115 | n3117 ;
  assign n3119 = ~n523 & n2932 ;
  assign n3120 = n2936 | n3119 ;
  assign n3121 = n3118 | n3120 ;
  assign n3122 = ~x23 & n3121 ;
  assign n3123 = n3118 | n3119 ;
  assign n3124 = ~x23 & n3123 ;
  assign n3125 = ( ~n1055 & n3122 ) | ( ~n1055 & n3124 ) | ( n3122 & n3124 ) ;
  assign n3126 = x23 & n3121 ;
  assign n3127 = x23 & ~n3126 ;
  assign n3128 = x23 & n3119 ;
  assign n3129 = ( x23 & n3118 ) | ( x23 & n3128 ) | ( n3118 & n3128 ) ;
  assign n3130 = x23 & ~n3129 ;
  assign n3131 = ( n1055 & n3127 ) | ( n1055 & n3130 ) | ( n3127 & n3130 ) ;
  assign n3132 = n3125 | n3131 ;
  assign n3133 = n2489 | n2491 ;
  assign n3134 = x26 & ~n2489 ;
  assign n3135 = ( n2472 & n3133 ) | ( n2472 & ~n3134 ) | ( n3133 & ~n3134 ) ;
  assign n3136 = ~n2494 & n3135 ;
  assign n3137 = n3132 & n3136 ;
  assign n3138 = x26 | n2486 ;
  assign n3139 = ( ~n2479 & n2486 ) | ( ~n2479 & n3138 ) | ( n2486 & n3138 ) ;
  assign n3140 = n2480 | n3139 ;
  assign n3141 = ~n2489 & n3140 ;
  assign n3142 = ~n829 & n2928 ;
  assign n3143 = n352 & n2932 ;
  assign n3144 = ( ~n339 & n2932 ) | ( ~n339 & n3143 ) | ( n2932 & n3143 ) ;
  assign n3145 = n3142 | n3144 ;
  assign n3146 = n692 & n2925 ;
  assign n3147 = ( n674 & n2925 ) | ( n674 & n3146 ) | ( n2925 & n3146 ) ;
  assign n3148 = n3145 | n3147 ;
  assign n3149 = n2936 | n3147 ;
  assign n3150 = n3145 | n3149 ;
  assign n3151 = ( ~n1209 & n3148 ) | ( ~n1209 & n3150 ) | ( n3148 & n3150 ) ;
  assign n3152 = ~x23 & n3150 ;
  assign n3153 = ~x23 & n3148 ;
  assign n3154 = ( ~n1209 & n3152 ) | ( ~n1209 & n3153 ) | ( n3152 & n3153 ) ;
  assign n3155 = x23 | n3153 ;
  assign n3156 = x23 | n3152 ;
  assign n3157 = ( ~n1209 & n3155 ) | ( ~n1209 & n3156 ) | ( n3155 & n3156 ) ;
  assign n3158 = ( ~n3151 & n3154 ) | ( ~n3151 & n3157 ) | ( n3154 & n3157 ) ;
  assign n3159 = n3141 & n3158 ;
  assign n3160 = ( ~n1027 & n2482 ) | ( ~n1027 & n2484 ) | ( n2482 & n2484 ) ;
  assign n3161 = ~n922 & n2928 ;
  assign n3162 = n1042 & n2925 ;
  assign n3163 = ( ~n1027 & n2925 ) | ( ~n1027 & n3162 ) | ( n2925 & n3162 ) ;
  assign n3164 = n3161 | n3163 ;
  assign n3165 = n692 & n2932 ;
  assign n3166 = ( n674 & n2932 ) | ( n674 & n3165 ) | ( n2932 & n3165 ) ;
  assign n3167 = n3164 | n3166 ;
  assign n3168 = ( n1538 & n2936 ) | ( n1538 & n3167 ) | ( n2936 & n3167 ) ;
  assign n3169 = ( x23 & ~n3167 ) | ( x23 & n3168 ) | ( ~n3167 & n3168 ) ;
  assign n3170 = ~n3168 & n3169 ;
  assign n3171 = ~n922 & n2932 ;
  assign n3172 = n1042 & n2928 ;
  assign n3173 = ( ~n1027 & n2928 ) | ( ~n1027 & n3172 ) | ( n2928 & n3172 ) ;
  assign n3174 = n3171 | n3173 ;
  assign n3175 = n2936 | n3173 ;
  assign n3176 = n3171 | n3175 ;
  assign n3177 = ( n1946 & n3174 ) | ( n1946 & n3176 ) | ( n3174 & n3176 ) ;
  assign n3178 = ~x23 & n3177 ;
  assign n3179 = n139 & n2920 ;
  assign n3180 = ( n1041 & n2920 ) | ( n1041 & n3179 ) | ( n2920 & n3179 ) ;
  assign n3181 = x23 & ~n3180 ;
  assign n3182 = n2920 | n3179 ;
  assign n3183 = x23 & ~n3182 ;
  assign n3184 = ( n1027 & n3181 ) | ( n1027 & n3183 ) | ( n3181 & n3183 ) ;
  assign n3185 = x23 & n3184 ;
  assign n3186 = ~n3177 & n3185 ;
  assign n3187 = ( n3178 & n3184 ) | ( n3178 & n3186 ) | ( n3184 & n3186 ) ;
  assign n3188 = x23 | n3167 ;
  assign n3189 = n3168 | n3188 ;
  assign n3190 = n3187 & n3189 ;
  assign n3191 = ~x23 & n3187 ;
  assign n3192 = ( n3170 & n3190 ) | ( n3170 & n3191 ) | ( n3190 & n3191 ) ;
  assign n3193 = n3160 & n3192 ;
  assign n3194 = n3192 & ~n3193 ;
  assign n3195 = ~n829 & n2932 ;
  assign n3196 = ~n922 & n2925 ;
  assign n3197 = n3195 | n3196 ;
  assign n3198 = n692 & n2928 ;
  assign n3199 = ( n674 & n2928 ) | ( n674 & n3198 ) | ( n2928 & n3198 ) ;
  assign n3200 = n3197 | n3199 ;
  assign n3201 = n2936 | n3199 ;
  assign n3202 = n3197 | n3201 ;
  assign n3203 = ( n1554 & n3200 ) | ( n1554 & n3202 ) | ( n3200 & n3202 ) ;
  assign n3204 = x23 & n3202 ;
  assign n3205 = x23 & n3200 ;
  assign n3206 = ( n1554 & n3204 ) | ( n1554 & n3205 ) | ( n3204 & n3205 ) ;
  assign n3207 = x23 & ~n3205 ;
  assign n3208 = x23 & ~n3204 ;
  assign n3209 = ( ~n1554 & n3207 ) | ( ~n1554 & n3208 ) | ( n3207 & n3208 ) ;
  assign n3210 = ( n3203 & ~n3206 ) | ( n3203 & n3209 ) | ( ~n3206 & n3209 ) ;
  assign n3211 = n3160 & ~n3192 ;
  assign n3212 = n3210 & n3211 ;
  assign n3213 = ( n3194 & n3210 ) | ( n3194 & n3212 ) | ( n3210 & n3212 ) ;
  assign n3214 = n3193 | n3213 ;
  assign n3215 = n3141 | n3158 ;
  assign n3216 = ~n3159 & n3215 ;
  assign n3217 = n3159 | n3216 ;
  assign n3218 = ( n3159 & n3214 ) | ( n3159 & n3217 ) | ( n3214 & n3217 ) ;
  assign n3219 = n3132 | n3136 ;
  assign n3220 = ~n3137 & n3219 ;
  assign n3221 = n3137 | n3220 ;
  assign n3222 = ( n3137 & n3218 ) | ( n3137 & n3221 ) | ( n3218 & n3221 ) ;
  assign n3223 = n3114 & n3222 ;
  assign n3224 = n3112 | n3223 ;
  assign n3225 = ~n3074 & n3090 ;
  assign n3226 = ( n3074 & ~n3091 ) | ( n3074 & n3225 ) | ( ~n3091 & n3225 ) ;
  assign n3227 = n3224 & n3226 ;
  assign n3228 = n3091 | n3227 ;
  assign n3229 = n2520 & n2522 ;
  assign n3230 = n2520 | n2522 ;
  assign n3231 = ~n3229 & n3230 ;
  assign n3232 = n1708 & n2928 ;
  assign n3233 = n1793 & n2925 ;
  assign n3234 = ( n1783 & n2925 ) | ( n1783 & n3233 ) | ( n2925 & n3233 ) ;
  assign n3235 = n1634 & n2932 ;
  assign n3236 = ( n1630 & n2932 ) | ( n1630 & n3235 ) | ( n2932 & n3235 ) ;
  assign n3237 = n3234 | n3236 ;
  assign n3238 = n3232 | n3237 ;
  assign n3239 = n2936 | n3238 ;
  assign n3240 = n3238 & n3239 ;
  assign n3241 = ( n1814 & n3239 ) | ( n1814 & n3240 ) | ( n3239 & n3240 ) ;
  assign n3242 = x23 & n3240 ;
  assign n3243 = x23 & n3239 ;
  assign n3244 = ( n1814 & n3242 ) | ( n1814 & n3243 ) | ( n3242 & n3243 ) ;
  assign n3245 = x23 & ~n3242 ;
  assign n3246 = x23 & ~n3243 ;
  assign n3247 = ( ~n1814 & n3245 ) | ( ~n1814 & n3246 ) | ( n3245 & n3246 ) ;
  assign n3248 = ( n3241 & ~n3244 ) | ( n3241 & n3247 ) | ( ~n3244 & n3247 ) ;
  assign n3249 = n3231 & n3248 ;
  assign n3250 = n3231 & ~n3249 ;
  assign n3251 = ~n3231 & n3248 ;
  assign n3252 = n3250 | n3251 ;
  assign n3253 = n3228 & n3252 ;
  assign n3254 = n3071 & n3249 ;
  assign n3255 = ( n3071 & n3253 ) | ( n3071 & n3254 ) | ( n3253 & n3254 ) ;
  assign n3256 = n3069 | n3255 ;
  assign n3257 = ~n3028 & n3046 ;
  assign n3258 = ~n3027 & n3257 ;
  assign n3259 = n3069 & n3258 ;
  assign n3260 = ( n3255 & n3258 ) | ( n3255 & n3259 ) | ( n3258 & n3259 ) ;
  assign n3261 = ( n3049 & n3256 ) | ( n3049 & n3260 ) | ( n3256 & n3260 ) ;
  assign n3262 = n3009 & ~n3024 ;
  assign n3263 = n3025 | n3262 ;
  assign n3264 = n3048 & ~n3263 ;
  assign n3265 = ( n3261 & ~n3263 ) | ( n3261 & n3264 ) | ( ~n3263 & n3264 ) ;
  assign n3266 = n3025 | n3265 ;
  assign n3592 = ~n3006 & n3266 ;
  assign n3593 = n3006 & ~n3266 ;
  assign n3594 = n3592 | n3593 ;
  assign n2696 = n85 | n694 ;
  assign n2697 = n504 | n2696 ;
  assign n2698 = n330 | n480 ;
  assign n2699 = n355 | n2698 ;
  assign n2700 = n2697 | n2699 ;
  assign n2701 = n273 | n2700 ;
  assign n2702 = n138 | n205 ;
  assign n2703 = n313 | n820 ;
  assign n2704 = n2702 | n2703 ;
  assign n2705 = n126 | n577 ;
  assign n2706 = n2704 | n2705 ;
  assign n2707 = n1615 | n1631 ;
  assign n2708 = n344 | n895 ;
  assign n2709 = n405 | n2708 ;
  assign n2710 = n2707 | n2709 ;
  assign n2711 = n717 | n2710 ;
  assign n2712 = n2706 | n2711 ;
  assign n2713 = n77 | n370 ;
  assign n2714 = n2083 | n2713 ;
  assign n2715 = n229 | n2714 ;
  assign n2716 = n645 | n995 ;
  assign n2717 = n530 | n2716 ;
  assign n2718 = n2715 | n2717 ;
  assign n2719 = n2663 | n2718 ;
  assign n2720 = n413 | n676 ;
  assign n2721 = n139 | n262 ;
  assign n2722 = n143 & ~n2721 ;
  assign n2723 = n311 | n979 ;
  assign n2724 = n289 | n458 ;
  assign n2725 = n341 | n2724 ;
  assign n2726 = n2723 | n2725 ;
  assign n2727 = ( n2720 & n2722 ) | ( n2720 & ~n2726 ) | ( n2722 & ~n2726 ) ;
  assign n2728 = ~n2720 & n2727 ;
  assign n2729 = n2720 & n2722 ;
  assign n2730 = ~n2720 & n2729 ;
  assign n2731 = ( ~n2719 & n2728 ) | ( ~n2719 & n2730 ) | ( n2728 & n2730 ) ;
  assign n2732 = ~n2712 & n2731 ;
  assign n2733 = n502 | n639 ;
  assign n2734 = n484 | n1663 ;
  assign n2735 = n2733 | n2734 ;
  assign n2736 = n225 | n675 ;
  assign n2737 = n154 | n2736 ;
  assign n2738 = n67 | n320 ;
  assign n2739 = n234 | n616 ;
  assign n2740 = n2738 | n2739 ;
  assign n2741 = n2737 | n2740 ;
  assign n2742 = n2735 | n2741 ;
  assign n2743 = n303 | n667 ;
  assign n2744 = n562 | n2743 ;
  assign n2745 = n418 | n441 ;
  assign n2746 = n79 | n2745 ;
  assign n2747 = n2744 | n2746 ;
  assign n2748 = n182 | n208 ;
  assign n2749 = n240 | n2748 ;
  assign n2750 = n2747 | n2749 ;
  assign n2751 = n2742 | n2750 ;
  assign n2752 = n291 | n602 ;
  assign n2753 = n437 | n2752 ;
  assign n2754 = n167 | n590 ;
  assign n2755 = n284 | n775 ;
  assign n2756 = n2754 | n2755 ;
  assign n2757 = n134 | n281 ;
  assign n2758 = n206 | n2757 ;
  assign n2759 = n2756 | n2758 ;
  assign n2760 = n2753 | n2759 ;
  assign n2761 = n987 | n2051 ;
  assign n2762 = n763 | n1675 ;
  assign n2763 = n2761 | n2762 ;
  assign n2764 = n412 | n1146 ;
  assign n2765 = n2763 | n2764 ;
  assign n2766 = n2760 | n2765 ;
  assign n2767 = n2751 | n2766 ;
  assign n2768 = n96 | n203 ;
  assign n2769 = n256 | n2768 ;
  assign n2770 = n2244 | n2769 ;
  assign n2771 = n457 | n511 ;
  assign n2772 = n83 | n857 ;
  assign n2773 = n2771 | n2772 ;
  assign n2774 = n2770 | n2773 ;
  assign n2775 = n190 | n383 ;
  assign n2776 = n160 | n306 ;
  assign n2777 = n2775 | n2776 ;
  assign n2778 = n1301 | n2777 ;
  assign n2779 = n1460 | n2778 ;
  assign n2780 = n2774 | n2779 ;
  assign n2781 = n177 | n1030 ;
  assign n2782 = n2780 | n2781 ;
  assign n2783 = n2767 | n2782 ;
  assign n2784 = n2732 & ~n2783 ;
  assign n2785 = ~n2701 & n2784 ;
  assign n2786 = n295 | n404 ;
  assign n2787 = n222 | n289 ;
  assign n2788 = n64 | n437 ;
  assign n2789 = n2787 | n2788 ;
  assign n2790 = n2618 | n2789 ;
  assign n2791 = n718 | n1469 ;
  assign n2792 = n2790 | n2791 ;
  assign n2793 = n2786 | n2792 ;
  assign n2794 = n607 | n895 ;
  assign n2795 = n487 | n2794 ;
  assign n2796 = n371 | n1482 ;
  assign n2797 = n2795 | n2796 ;
  assign n2798 = n189 | n228 ;
  assign n2799 = n213 | n320 ;
  assign n2800 = n2798 | n2799 ;
  assign n2801 = n2797 | n2800 ;
  assign n2802 = n2793 | n2801 ;
  assign n2803 = n412 | n608 ;
  assign n2804 = n77 | n2803 ;
  assign n2805 = n263 | n277 ;
  assign n2806 = n375 | n2805 ;
  assign n2807 = n2804 | n2806 ;
  assign n2808 = n123 | n588 ;
  assign n2809 = n325 | n2808 ;
  assign n2810 = n663 | n2809 ;
  assign n2811 = n2807 | n2810 ;
  assign n2812 = n246 | n297 ;
  assign n2813 = n417 | n2812 ;
  assign n2814 = n255 | n2813 ;
  assign n2815 = n141 | n234 ;
  assign n2816 = n182 | n2815 ;
  assign n2817 = n2814 | n2816 ;
  assign n2818 = n2811 | n2817 ;
  assign n2819 = n355 | n581 ;
  assign n2820 = n502 | n2819 ;
  assign n2821 = n143 & ~n151 ;
  assign n2822 = ~n2820 & n2821 ;
  assign n1307 = n302 | n309 ;
  assign n2823 = n389 | n929 ;
  assign n2824 = n1307 | n2823 ;
  assign n2825 = n2822 & ~n2824 ;
  assign n2826 = ~n2818 & n2825 ;
  assign n2827 = ~n2802 & n2826 ;
  assign n2828 = n480 | n1172 ;
  assign n2829 = n644 | n1039 ;
  assign n2830 = n2828 | n2829 ;
  assign n2831 = n193 | n555 ;
  assign n2832 = n333 | n2831 ;
  assign n2833 = n2830 | n2832 ;
  assign n2834 = n2827 & ~n2833 ;
  assign n2835 = n75 | n284 ;
  assign n2836 = n1719 | n2835 ;
  assign n2837 = n630 | n2836 ;
  assign n2838 = n83 | n313 ;
  assign n2839 = n363 | n762 ;
  assign n2840 = n2838 | n2839 ;
  assign n2841 = n176 | n479 ;
  assign n2842 = n237 | n273 ;
  assign n2843 = n2841 | n2842 ;
  assign n2844 = n2840 | n2843 ;
  assign n2845 = n2837 | n2844 ;
  assign n2846 = n261 | n451 ;
  assign n2847 = n203 | n667 ;
  assign n2848 = n2846 | n2847 ;
  assign n2849 = n110 | n2848 ;
  assign n2850 = n270 | n483 ;
  assign n2851 = n960 | n2850 ;
  assign n2852 = n139 | n254 ;
  assign n2853 = n2851 | n2852 ;
  assign n2854 = n2849 | n2853 ;
  assign n2855 = n2845 | n2854 ;
  assign n2856 = n542 | n594 ;
  assign n2857 = n1404 | n2856 ;
  assign n2858 = n168 | n959 ;
  assign n2859 = n458 | n2858 ;
  assign n2860 = n2857 | n2859 ;
  assign n2861 = n2855 | n2860 ;
  assign n2862 = n134 | n600 ;
  assign n2863 = n372 | n2862 ;
  assign n2864 = n281 | n434 ;
  assign n2865 = n212 | n2864 ;
  assign n2866 = n2863 | n2865 ;
  assign n2867 = n202 | n460 ;
  assign n2868 = n441 | n2867 ;
  assign n2869 = n2866 | n2868 ;
  assign n2870 = n349 | n491 ;
  assign n2871 = n2771 | n2870 ;
  assign n2872 = n196 | n332 ;
  assign n2873 = n2871 | n2872 ;
  assign n2874 = n131 | n591 ;
  assign n2875 = n179 | n654 ;
  assign n2876 = n2874 | n2875 ;
  assign n2877 = n1234 | n2876 ;
  assign n2878 = n2873 | n2877 ;
  assign n2879 = n631 | n638 ;
  assign n2880 = n381 | n2879 ;
  assign n2881 = n721 | n2880 ;
  assign n2882 = n2878 | n2881 ;
  assign n2883 = n2869 | n2882 ;
  assign n2884 = n2861 | n2883 ;
  assign n2885 = n710 | n2884 ;
  assign n2886 = n2834 & ~n2885 ;
  assign n1126 = n390 | n676 ;
  assign n2887 = n288 | n841 ;
  assign n2888 = n1126 | n2887 ;
  assign n2889 = n208 | n344 ;
  assign n2890 = n272 | n2889 ;
  assign n2891 = n2888 | n2890 ;
  assign n2892 = n184 | n577 ;
  assign n2893 = n2891 | n2892 ;
  assign n2894 = n2886 & ~n2893 ;
  assign n2895 = n2785 | n2894 ;
  assign n2896 = n2785 & n2894 ;
  assign n2897 = n2895 & ~n2896 ;
  assign n2898 = n2692 & ~n2785 ;
  assign n2899 = ~n2692 & n2785 ;
  assign n2900 = n2898 | n2899 ;
  assign n2901 = n2693 | n2898 ;
  assign n2902 = ( n2898 & ~n2900 ) | ( n2898 & n2901 ) | ( ~n2900 & n2901 ) ;
  assign n2903 = n2897 & n2902 ;
  assign n3444 = n465 | n594 ;
  assign n3445 = n318 | n624 ;
  assign n3446 = n77 | n160 ;
  assign n3447 = n3445 | n3446 ;
  assign n3448 = n3444 | n3447 ;
  assign n3449 = n2221 | n3448 ;
  assign n3450 = n257 | n654 ;
  assign n3451 = n833 | n3450 ;
  assign n3452 = n239 | n273 ;
  assign n3453 = n3451 | n3452 ;
  assign n3454 = n513 | n689 ;
  assign n3455 = n254 | n3454 ;
  assign n3456 = n3453 | n3455 ;
  assign n3457 = n3449 | n3456 ;
  assign n3458 = n2651 | n3457 ;
  assign n3459 = n167 | n258 ;
  assign n3460 = n154 | n226 ;
  assign n3461 = n3459 | n3460 ;
  assign n3462 = n110 | n3461 ;
  assign n3463 = n1393 | n3462 ;
  assign n3464 = n1368 | n3463 ;
  assign n3465 = n240 | n839 ;
  assign n3466 = n2841 | n3465 ;
  assign n3467 = n214 | n347 ;
  assign n3468 = n841 | n3467 ;
  assign n3469 = n3466 | n3468 ;
  assign n3470 = n489 | n666 ;
  assign n3471 = n762 | n3470 ;
  assign n3472 = n573 | n3471 ;
  assign n3473 = n3469 | n3472 ;
  assign n3474 = n364 | n608 ;
  assign n3475 = n416 | n510 ;
  assign n3476 = n3474 | n3475 ;
  assign n3477 = n59 | n725 ;
  assign n3478 = n302 | n3477 ;
  assign n3479 = n3476 | n3478 ;
  assign n3480 = n3473 | n3479 ;
  assign n3481 = n3464 | n3480 ;
  assign n3482 = n3458 | n3481 ;
  assign n3483 = n2060 | n3482 ;
  assign n3484 = n212 | n447 ;
  assign n3485 = n333 | n3484 ;
  assign n3486 = n478 | n1637 ;
  assign n3487 = n3485 | n3486 ;
  assign n3488 = n112 | n1172 ;
  assign n3489 = n64 | n313 ;
  assign n3490 = n3488 | n3489 ;
  assign n3491 = n229 | n405 ;
  assign n3492 = n1243 | n3491 ;
  assign n3493 = n3490 | n3492 ;
  assign n3494 = n3487 | n3493 ;
  assign n3495 = n170 | n1114 ;
  assign n3496 = n1607 | n3495 ;
  assign n3497 = n2117 | n3496 ;
  assign n3498 = n2192 | n3497 ;
  assign n3499 = n3494 | n3498 ;
  assign n3500 = n445 | n3499 ;
  assign n3501 = n123 | n183 ;
  assign n3502 = n88 | n356 ;
  assign n3503 = n3501 | n3502 ;
  assign n3504 = n381 | n895 ;
  assign n3505 = n126 | n3504 ;
  assign n3506 = n3503 | n3505 ;
  assign n3507 = n3500 | n3506 ;
  assign n3508 = n3483 | n3507 ;
  assign n3515 = ~n2894 & n3508 ;
  assign n3516 = n2894 & ~n3508 ;
  assign n3517 = n3515 | n3516 ;
  assign n3518 = n2895 | n3517 ;
  assign n3519 = ( ~n2903 & n3517 ) | ( ~n2903 & n3518 ) | ( n3517 & n3518 ) ;
  assign n2904 = ~n2898 & n2900 ;
  assign n2905 = n2897 & ~n2904 ;
  assign n3520 = ( ~n2905 & n3517 ) | ( ~n2905 & n3518 ) | ( n3517 & n3518 ) ;
  assign n3521 = n3519 | n3520 ;
  assign n3523 = ( n2695 & n3519 ) | ( n2695 & n3520 ) | ( n3519 & n3520 ) ;
  assign n3595 = ( n2602 & n3521 ) | ( n2602 & n3523 ) | ( n3521 & n3523 ) ;
  assign n3596 = n2895 & ~n2903 ;
  assign n3597 = n2895 & ~n2905 ;
  assign n3598 = n3596 | n3597 ;
  assign n3599 = n3517 & n3598 ;
  assign n3600 = ( n2695 & n3596 ) | ( n2695 & n3597 ) | ( n3596 & n3597 ) ;
  assign n3601 = n3517 & n3600 ;
  assign n3602 = ( n2602 & n3599 ) | ( n2602 & n3601 ) | ( n3599 & n3601 ) ;
  assign n3603 = n3595 & ~n3602 ;
  assign n3531 = x19 & ~x20 ;
  assign n3532 = ~x19 & x20 ;
  assign n3533 = n3531 | n3532 ;
  assign n3534 = x17 & ~x18 ;
  assign n3535 = ~x17 & x18 ;
  assign n3536 = n3534 | n3535 ;
  assign n3537 = n3533 & n3536 ;
  assign n3538 = ~x18 & x19 ;
  assign n3539 = x18 & ~x19 ;
  assign n3540 = n3538 | n3539 ;
  assign n3541 = ~n3536 & n3540 ;
  assign n3604 = n2893 & n3541 ;
  assign n3605 = ( ~n2886 & n3541 ) | ( ~n2886 & n3604 ) | ( n3541 & n3604 ) ;
  assign n3543 = n3533 & ~n3536 ;
  assign n3544 = ~n3540 & n3543 ;
  assign n3606 = n2701 & n3544 ;
  assign n3607 = ( ~n2784 & n3544 ) | ( ~n2784 & n3606 ) | ( n3544 & n3606 ) ;
  assign n3547 = ~n3533 & n3536 ;
  assign n3608 = n3507 & n3547 ;
  assign n3609 = ( n3483 & n3547 ) | ( n3483 & n3608 ) | ( n3547 & n3608 ) ;
  assign n3610 = n3607 | n3609 ;
  assign n3611 = n3605 | n3610 ;
  assign n3612 = n3537 | n3611 ;
  assign n3613 = n3611 & n3612 ;
  assign n3614 = ( n3603 & n3612 ) | ( n3603 & n3613 ) | ( n3612 & n3613 ) ;
  assign n3615 = x20 & n3613 ;
  assign n3616 = x20 & n3612 ;
  assign n3617 = ( n3603 & n3615 ) | ( n3603 & n3616 ) | ( n3615 & n3616 ) ;
  assign n3618 = x20 & ~n3615 ;
  assign n3619 = x20 & ~n3616 ;
  assign n3620 = ( ~n3603 & n3618 ) | ( ~n3603 & n3619 ) | ( n3618 & n3619 ) ;
  assign n3621 = ( n3614 & ~n3617 ) | ( n3614 & n3620 ) | ( ~n3617 & n3620 ) ;
  assign n3622 = ~n3594 & n3621 ;
  assign n3623 = n3594 | n3622 ;
  assign n3624 = n3594 & n3621 ;
  assign n3625 = n3623 & ~n3624 ;
  assign n3626 = ~n3048 & n3263 ;
  assign n3627 = ~n3261 & n3626 ;
  assign n3628 = n3265 | n3627 ;
  assign n2906 = ( ~n2695 & n2903 ) | ( ~n2695 & n2905 ) | ( n2903 & n2905 ) ;
  assign n2907 = n2903 & n2905 ;
  assign n2908 = ( ~n2602 & n2906 ) | ( ~n2602 & n2907 ) | ( n2906 & n2907 ) ;
  assign n2909 = n2902 & ~n2904 ;
  assign n2910 = n2897 | n2909 ;
  assign n2911 = ( n2695 & ~n2902 ) | ( n2695 & n2904 ) | ( ~n2902 & n2904 ) ;
  assign n2912 = ~n2897 & n2911 ;
  assign n2913 = ( n2602 & ~n2910 ) | ( n2602 & n2912 ) | ( ~n2910 & n2912 ) ;
  assign n2914 = n2908 | n2913 ;
  assign n3629 = n2691 & n3544 ;
  assign n3630 = ( n2678 & n3544 ) | ( n2678 & n3629 ) | ( n3544 & n3629 ) ;
  assign n3631 = n2701 & n3541 ;
  assign n3632 = ( ~n2784 & n3541 ) | ( ~n2784 & n3631 ) | ( n3541 & n3631 ) ;
  assign n3633 = n3630 | n3632 ;
  assign n3634 = n2893 & n3547 ;
  assign n3635 = ( ~n2886 & n3547 ) | ( ~n2886 & n3634 ) | ( n3547 & n3634 ) ;
  assign n3636 = n3633 | n3635 ;
  assign n3637 = n3537 | n3636 ;
  assign n3638 = n3636 & n3637 ;
  assign n3639 = ( ~n2914 & n3637 ) | ( ~n2914 & n3638 ) | ( n3637 & n3638 ) ;
  assign n3640 = ~x20 & n3638 ;
  assign n3641 = ~x20 & n3637 ;
  assign n3642 = ( ~n2914 & n3640 ) | ( ~n2914 & n3641 ) | ( n3640 & n3641 ) ;
  assign n3643 = x20 | n3640 ;
  assign n3644 = x20 | n3641 ;
  assign n3645 = ( ~n2914 & n3643 ) | ( ~n2914 & n3644 ) | ( n3643 & n3644 ) ;
  assign n3646 = ( ~n3639 & n3642 ) | ( ~n3639 & n3645 ) | ( n3642 & n3645 ) ;
  assign n3647 = ~n3628 & n3646 ;
  assign n3648 = n3628 | n3647 ;
  assign n3649 = n3628 & n3646 ;
  assign n3650 = n3648 & ~n3649 ;
  assign n3651 = n3069 | n3258 ;
  assign n3652 = n3255 | n3651 ;
  assign n3653 = n3049 | n3652 ;
  assign n3654 = ~n3261 & n3653 ;
  assign n2953 = n2693 & ~n2900 ;
  assign n2954 = ( n2695 & n2900 ) | ( n2695 & ~n2953 ) | ( n2900 & ~n2953 ) ;
  assign n2955 = ~n2900 & n2953 ;
  assign n2956 = ( n2602 & n2954 ) | ( n2602 & ~n2955 ) | ( n2954 & ~n2955 ) ;
  assign n2957 = ~n2693 & n2900 ;
  assign n2958 = n2695 & n2957 ;
  assign n2959 = ( n2602 & n2957 ) | ( n2602 & n2958 ) | ( n2957 & n2958 ) ;
  assign n2960 = n2956 & ~n2959 ;
  assign n3655 = n2701 & n3547 ;
  assign n3656 = ( ~n2784 & n3547 ) | ( ~n2784 & n3655 ) | ( n3547 & n3655 ) ;
  assign n3657 = n2691 & n3541 ;
  assign n3658 = ( n2678 & n3541 ) | ( n2678 & n3657 ) | ( n3541 & n3657 ) ;
  assign n3659 = n3656 | n3658 ;
  assign n3660 = n2199 & n3544 ;
  assign n3661 = ( ~n2185 & n3544 ) | ( ~n2185 & n3660 ) | ( n3544 & n3660 ) ;
  assign n3662 = n3659 | n3661 ;
  assign n3663 = n3537 | n3661 ;
  assign n3664 = n3659 | n3663 ;
  assign n3665 = ( n2960 & n3662 ) | ( n2960 & n3664 ) | ( n3662 & n3664 ) ;
  assign n3666 = x20 & n3664 ;
  assign n3667 = x20 & n3662 ;
  assign n3668 = ( n2960 & n3666 ) | ( n2960 & n3667 ) | ( n3666 & n3667 ) ;
  assign n3669 = x20 & ~n3667 ;
  assign n3670 = x20 & ~n3666 ;
  assign n3671 = ( ~n2960 & n3669 ) | ( ~n2960 & n3670 ) | ( n3669 & n3670 ) ;
  assign n3672 = ( n3665 & ~n3668 ) | ( n3665 & n3671 ) | ( ~n3668 & n3671 ) ;
  assign n3673 = n3654 & n3672 ;
  assign n3674 = n3654 & ~n3673 ;
  assign n3675 = ~n3654 & n3672 ;
  assign n3676 = n3674 | n3675 ;
  assign n3677 = n3071 | n3249 ;
  assign n3678 = n3253 | n3677 ;
  assign n3679 = ~n3255 & n3678 ;
  assign n3680 = n2090 & n3544 ;
  assign n3681 = ( ~n2082 & n3544 ) | ( ~n2082 & n3680 ) | ( n3544 & n3680 ) ;
  assign n3682 = n2691 & n3547 ;
  assign n3683 = ( n2678 & n3547 ) | ( n2678 & n3682 ) | ( n3547 & n3682 ) ;
  assign n3684 = n2199 & n3541 ;
  assign n3685 = ( ~n2185 & n3541 ) | ( ~n2185 & n3684 ) | ( n3541 & n3684 ) ;
  assign n3686 = n3683 | n3685 ;
  assign n3687 = n3681 | n3686 ;
  assign n3688 = n3537 | n3687 ;
  assign n3689 = ( n2985 & n3687 ) | ( n2985 & n3688 ) | ( n3687 & n3688 ) ;
  assign n3690 = x20 & n3688 ;
  assign n3691 = x20 & n3687 ;
  assign n3692 = ( n2985 & n3690 ) | ( n2985 & n3691 ) | ( n3690 & n3691 ) ;
  assign n3693 = x20 & ~n3690 ;
  assign n3694 = x20 & ~n3691 ;
  assign n3695 = ( ~n2985 & n3693 ) | ( ~n2985 & n3694 ) | ( n3693 & n3694 ) ;
  assign n3696 = ( n3689 & ~n3692 ) | ( n3689 & n3695 ) | ( ~n3692 & n3695 ) ;
  assign n3697 = n3679 & n3696 ;
  assign n3698 = ~n3228 & n3252 ;
  assign n3699 = n3228 & ~n3252 ;
  assign n3700 = n3698 | n3699 ;
  assign n3701 = n2090 & n3541 ;
  assign n3702 = ( ~n2082 & n3541 ) | ( ~n2082 & n3701 ) | ( n3541 & n3701 ) ;
  assign n3703 = n2279 & n3544 ;
  assign n3704 = ( ~n2269 & n3544 ) | ( ~n2269 & n3703 ) | ( n3544 & n3703 ) ;
  assign n3705 = n2199 & n3547 ;
  assign n3706 = ( ~n2185 & n3547 ) | ( ~n2185 & n3705 ) | ( n3547 & n3705 ) ;
  assign n3707 = n3704 | n3706 ;
  assign n3708 = n3702 | n3707 ;
  assign n3709 = n3537 | n3708 ;
  assign n3710 = ( ~n2325 & n3708 ) | ( ~n2325 & n3709 ) | ( n3708 & n3709 ) ;
  assign n3711 = n3708 & n3709 ;
  assign n3712 = ( ~n2299 & n3710 ) | ( ~n2299 & n3711 ) | ( n3710 & n3711 ) ;
  assign n3713 = ~x20 & n3712 ;
  assign n3714 = x20 | n3712 ;
  assign n3715 = ( ~n3712 & n3713 ) | ( ~n3712 & n3714 ) | ( n3713 & n3714 ) ;
  assign n3716 = n3700 & n3715 ;
  assign n3717 = n3700 | n3715 ;
  assign n3718 = ~n3716 & n3717 ;
  assign n3719 = n3224 | n3226 ;
  assign n3720 = ~n3227 & n3719 ;
  assign n3721 = n1634 & n3544 ;
  assign n3722 = ( n1630 & n3544 ) | ( n1630 & n3721 ) | ( n3544 & n3721 ) ;
  assign n3723 = n2279 & n3541 ;
  assign n3724 = ( ~n2269 & n3541 ) | ( ~n2269 & n3723 ) | ( n3541 & n3723 ) ;
  assign n3725 = n3722 | n3724 ;
  assign n3726 = n2090 & n3547 ;
  assign n3727 = ( ~n2082 & n3547 ) | ( ~n2082 & n3726 ) | ( n3547 & n3726 ) ;
  assign n3728 = n3725 | n3727 ;
  assign n3729 = n3537 | n3728 ;
  assign n3730 = n3728 & n3729 ;
  assign n3731 = ( n2568 & n3729 ) | ( n2568 & n3730 ) | ( n3729 & n3730 ) ;
  assign n3732 = x20 & n3730 ;
  assign n3733 = x20 & n3729 ;
  assign n3734 = ( n2568 & n3732 ) | ( n2568 & n3733 ) | ( n3732 & n3733 ) ;
  assign n3735 = x20 & ~n3732 ;
  assign n3736 = x20 & ~n3733 ;
  assign n3737 = ( ~n2568 & n3735 ) | ( ~n2568 & n3736 ) | ( n3735 & n3736 ) ;
  assign n3738 = ( n3731 & ~n3734 ) | ( n3731 & n3737 ) | ( ~n3734 & n3737 ) ;
  assign n3739 = n3720 & n3738 ;
  assign n3740 = n3114 | n3222 ;
  assign n3741 = ~n3223 & n3740 ;
  assign n3742 = n1708 & n3544 ;
  assign n3743 = n1634 & n3541 ;
  assign n3744 = ( n1630 & n3541 ) | ( n1630 & n3743 ) | ( n3541 & n3743 ) ;
  assign n3745 = n2279 & n3547 ;
  assign n3746 = ( ~n2269 & n3547 ) | ( ~n2269 & n3745 ) | ( n3547 & n3745 ) ;
  assign n3747 = n3744 | n3746 ;
  assign n3748 = n3742 | n3747 ;
  assign n3749 = n3537 | n3748 ;
  assign n3750 = n3748 & n3749 ;
  assign n3751 = ( ~n2343 & n3749 ) | ( ~n2343 & n3750 ) | ( n3749 & n3750 ) ;
  assign n3752 = ~x20 & n3750 ;
  assign n3753 = ~x20 & n3749 ;
  assign n3754 = ( ~n2343 & n3752 ) | ( ~n2343 & n3753 ) | ( n3752 & n3753 ) ;
  assign n3755 = x20 | n3752 ;
  assign n3756 = x20 | n3753 ;
  assign n3757 = ( ~n2343 & n3755 ) | ( ~n2343 & n3756 ) | ( n3755 & n3756 ) ;
  assign n3758 = ( ~n3751 & n3754 ) | ( ~n3751 & n3757 ) | ( n3754 & n3757 ) ;
  assign n3759 = n3741 & n3758 ;
  assign n3760 = n3218 & n3220 ;
  assign n3761 = n3218 | n3220 ;
  assign n3762 = ~n3760 & n3761 ;
  assign n3763 = n1708 & n3541 ;
  assign n3764 = n1793 & n3544 ;
  assign n3765 = ( n1783 & n3544 ) | ( n1783 & n3764 ) | ( n3544 & n3764 ) ;
  assign n3766 = n1634 & n3547 ;
  assign n3767 = ( n1630 & n3547 ) | ( n1630 & n3766 ) | ( n3547 & n3766 ) ;
  assign n3768 = n3765 | n3767 ;
  assign n3769 = n3763 | n3768 ;
  assign n3770 = n3537 | n3769 ;
  assign n3771 = n3769 & n3770 ;
  assign n3772 = ( n1814 & n3770 ) | ( n1814 & n3771 ) | ( n3770 & n3771 ) ;
  assign n3773 = x20 & n3771 ;
  assign n3774 = x20 & n3770 ;
  assign n3775 = ( n1814 & n3773 ) | ( n1814 & n3774 ) | ( n3773 & n3774 ) ;
  assign n3776 = x20 & ~n3773 ;
  assign n3777 = x20 & ~n3774 ;
  assign n3778 = ( ~n1814 & n3776 ) | ( ~n1814 & n3777 ) | ( n3776 & n3777 ) ;
  assign n3779 = ( n3772 & ~n3775 ) | ( n3772 & n3778 ) | ( ~n3775 & n3778 ) ;
  assign n3780 = n3762 & n3779 ;
  assign n3781 = n3214 & n3216 ;
  assign n3782 = n3214 | n3216 ;
  assign n3783 = ~n3781 & n3782 ;
  assign n3784 = ~n523 & n3544 ;
  assign n3785 = n1793 & n3541 ;
  assign n3786 = ( n1783 & n3541 ) | ( n1783 & n3785 ) | ( n3541 & n3785 ) ;
  assign n3787 = n3784 | n3786 ;
  assign n3788 = n1708 & n3547 ;
  assign n3789 = n3787 | n3788 ;
  assign n3790 = n3537 | n3788 ;
  assign n3791 = n3787 | n3790 ;
  assign n3792 = ( ~n1852 & n3789 ) | ( ~n1852 & n3791 ) | ( n3789 & n3791 ) ;
  assign n3793 = ~x20 & n3791 ;
  assign n3794 = ~x20 & n3789 ;
  assign n3795 = ( ~n1852 & n3793 ) | ( ~n1852 & n3794 ) | ( n3793 & n3794 ) ;
  assign n3796 = x20 | n3794 ;
  assign n3797 = x20 | n3793 ;
  assign n3798 = ( ~n1852 & n3796 ) | ( ~n1852 & n3797 ) | ( n3796 & n3797 ) ;
  assign n3799 = ( ~n3792 & n3795 ) | ( ~n3792 & n3798 ) | ( n3795 & n3798 ) ;
  assign n3800 = n3783 & n3799 ;
  assign n3801 = n3210 | n3211 ;
  assign n3802 = n3194 | n3801 ;
  assign n3803 = ~n3213 & n3802 ;
  assign n3804 = ~n523 & n3541 ;
  assign n3805 = n352 & n3544 ;
  assign n3806 = ( ~n339 & n3544 ) | ( ~n339 & n3805 ) | ( n3544 & n3805 ) ;
  assign n3807 = n1793 & n3547 ;
  assign n3808 = ( n1783 & n3547 ) | ( n1783 & n3807 ) | ( n3547 & n3807 ) ;
  assign n3809 = n3806 | n3808 ;
  assign n3810 = n3804 | n3809 ;
  assign n3811 = n3537 | n3810 ;
  assign n3812 = n3810 & n3811 ;
  assign n3813 = ( n1884 & n3811 ) | ( n1884 & n3812 ) | ( n3811 & n3812 ) ;
  assign n3814 = x20 & n3812 ;
  assign n3815 = x20 & n3811 ;
  assign n3816 = ( n1884 & n3814 ) | ( n1884 & n3815 ) | ( n3814 & n3815 ) ;
  assign n3817 = x20 & ~n3814 ;
  assign n3818 = x20 & ~n3815 ;
  assign n3819 = ( ~n1884 & n3817 ) | ( ~n1884 & n3818 ) | ( n3817 & n3818 ) ;
  assign n3820 = ( n3813 & ~n3816 ) | ( n3813 & n3819 ) | ( ~n3816 & n3819 ) ;
  assign n3821 = n3803 & n3820 ;
  assign n3822 = n3803 | n3820 ;
  assign n3823 = ~n3821 & n3822 ;
  assign n3824 = ~n829 & n3544 ;
  assign n3825 = n352 & n3541 ;
  assign n3826 = ( ~n339 & n3541 ) | ( ~n339 & n3825 ) | ( n3541 & n3825 ) ;
  assign n3827 = n3824 | n3826 ;
  assign n3828 = ~n523 & n3547 ;
  assign n3829 = n3537 | n3828 ;
  assign n3830 = n3827 | n3829 ;
  assign n3831 = ~x20 & n3830 ;
  assign n3832 = n3827 | n3828 ;
  assign n3833 = ~x20 & n3832 ;
  assign n3834 = ( ~n1055 & n3831 ) | ( ~n1055 & n3833 ) | ( n3831 & n3833 ) ;
  assign n3835 = x20 & n3830 ;
  assign n3836 = x20 & ~n3835 ;
  assign n3837 = x20 & n3828 ;
  assign n3838 = ( x20 & n3827 ) | ( x20 & n3837 ) | ( n3827 & n3837 ) ;
  assign n3839 = x20 & ~n3838 ;
  assign n3840 = ( n1055 & n3836 ) | ( n1055 & n3839 ) | ( n3836 & n3839 ) ;
  assign n3841 = n3834 | n3840 ;
  assign n3842 = n3187 | n3189 ;
  assign n3843 = x23 & ~n3187 ;
  assign n3844 = ( n3170 & n3842 ) | ( n3170 & ~n3843 ) | ( n3842 & ~n3843 ) ;
  assign n3845 = ~n3192 & n3844 ;
  assign n3846 = n3841 & n3845 ;
  assign n3847 = x23 | n3184 ;
  assign n3848 = ( ~n3177 & n3184 ) | ( ~n3177 & n3847 ) | ( n3184 & n3847 ) ;
  assign n3849 = n3178 | n3848 ;
  assign n3850 = ~n3187 & n3849 ;
  assign n3851 = ~n829 & n3541 ;
  assign n3852 = n352 & n3547 ;
  assign n3853 = ( ~n339 & n3547 ) | ( ~n339 & n3852 ) | ( n3547 & n3852 ) ;
  assign n3854 = n3851 | n3853 ;
  assign n3855 = n692 & n3544 ;
  assign n3856 = ( n674 & n3544 ) | ( n674 & n3855 ) | ( n3544 & n3855 ) ;
  assign n3857 = n3854 | n3856 ;
  assign n3858 = n3537 | n3856 ;
  assign n3859 = n3854 | n3858 ;
  assign n3860 = ( ~n1209 & n3857 ) | ( ~n1209 & n3859 ) | ( n3857 & n3859 ) ;
  assign n3861 = ~x20 & n3859 ;
  assign n3862 = ~x20 & n3857 ;
  assign n3863 = ( ~n1209 & n3861 ) | ( ~n1209 & n3862 ) | ( n3861 & n3862 ) ;
  assign n3864 = x20 | n3862 ;
  assign n3865 = x20 | n3861 ;
  assign n3866 = ( ~n1209 & n3864 ) | ( ~n1209 & n3865 ) | ( n3864 & n3865 ) ;
  assign n3867 = ( ~n3860 & n3863 ) | ( ~n3860 & n3866 ) | ( n3863 & n3866 ) ;
  assign n3868 = n3850 & n3867 ;
  assign n3869 = ( ~n1027 & n3180 ) | ( ~n1027 & n3182 ) | ( n3180 & n3182 ) ;
  assign n3870 = ~n922 & n3541 ;
  assign n3871 = n1042 & n3544 ;
  assign n3872 = ( ~n1027 & n3544 ) | ( ~n1027 & n3871 ) | ( n3544 & n3871 ) ;
  assign n3873 = n3870 | n3872 ;
  assign n3874 = n692 & n3547 ;
  assign n3875 = ( n674 & n3547 ) | ( n674 & n3874 ) | ( n3547 & n3874 ) ;
  assign n3876 = n3873 | n3875 ;
  assign n3877 = ( n1538 & n3537 ) | ( n1538 & n3876 ) | ( n3537 & n3876 ) ;
  assign n3878 = ( x20 & ~n3876 ) | ( x20 & n3877 ) | ( ~n3876 & n3877 ) ;
  assign n3879 = ~n3877 & n3878 ;
  assign n3880 = ~n922 & n3547 ;
  assign n3881 = n1042 & n3541 ;
  assign n3882 = ( ~n1027 & n3541 ) | ( ~n1027 & n3881 ) | ( n3541 & n3881 ) ;
  assign n3883 = n3880 | n3882 ;
  assign n3884 = n3537 | n3882 ;
  assign n3885 = n3880 | n3884 ;
  assign n3886 = ( n1946 & n3883 ) | ( n1946 & n3885 ) | ( n3883 & n3885 ) ;
  assign n3887 = ~x20 & n3886 ;
  assign n3888 = n139 & n3536 ;
  assign n3889 = ( n1041 & n3536 ) | ( n1041 & n3888 ) | ( n3536 & n3888 ) ;
  assign n3890 = x20 & ~n3889 ;
  assign n3891 = n3536 | n3888 ;
  assign n3892 = x20 & ~n3891 ;
  assign n3893 = ( n1027 & n3890 ) | ( n1027 & n3892 ) | ( n3890 & n3892 ) ;
  assign n3894 = x20 & n3893 ;
  assign n3895 = ~n3886 & n3894 ;
  assign n3896 = ( n3887 & n3893 ) | ( n3887 & n3895 ) | ( n3893 & n3895 ) ;
  assign n3897 = x20 | n3876 ;
  assign n3898 = n3877 | n3897 ;
  assign n3899 = n3896 & n3898 ;
  assign n3900 = ~x20 & n3896 ;
  assign n3901 = ( n3879 & n3899 ) | ( n3879 & n3900 ) | ( n3899 & n3900 ) ;
  assign n3902 = n3869 & n3901 ;
  assign n3903 = n3901 & ~n3902 ;
  assign n3904 = ~n829 & n3547 ;
  assign n3905 = ~n922 & n3544 ;
  assign n3906 = n3904 | n3905 ;
  assign n3907 = n692 & n3541 ;
  assign n3908 = ( n674 & n3541 ) | ( n674 & n3907 ) | ( n3541 & n3907 ) ;
  assign n3909 = n3906 | n3908 ;
  assign n3910 = n3537 | n3908 ;
  assign n3911 = n3906 | n3910 ;
  assign n3912 = ( n1554 & n3909 ) | ( n1554 & n3911 ) | ( n3909 & n3911 ) ;
  assign n3913 = x20 & n3911 ;
  assign n3914 = x20 & n3909 ;
  assign n3915 = ( n1554 & n3913 ) | ( n1554 & n3914 ) | ( n3913 & n3914 ) ;
  assign n3916 = x20 & ~n3914 ;
  assign n3917 = x20 & ~n3913 ;
  assign n3918 = ( ~n1554 & n3916 ) | ( ~n1554 & n3917 ) | ( n3916 & n3917 ) ;
  assign n3919 = ( n3912 & ~n3915 ) | ( n3912 & n3918 ) | ( ~n3915 & n3918 ) ;
  assign n3920 = n3869 & ~n3901 ;
  assign n3921 = n3919 & n3920 ;
  assign n3922 = ( n3903 & n3919 ) | ( n3903 & n3921 ) | ( n3919 & n3921 ) ;
  assign n3923 = n3902 | n3922 ;
  assign n3924 = n3850 | n3867 ;
  assign n3925 = ~n3868 & n3924 ;
  assign n3926 = n3868 | n3925 ;
  assign n3927 = ( n3868 & n3923 ) | ( n3868 & n3926 ) | ( n3923 & n3926 ) ;
  assign n3928 = n3841 | n3845 ;
  assign n3929 = ~n3846 & n3928 ;
  assign n3930 = n3846 | n3929 ;
  assign n3931 = ( n3846 & n3927 ) | ( n3846 & n3930 ) | ( n3927 & n3930 ) ;
  assign n3932 = n3823 & n3931 ;
  assign n3933 = n3821 | n3932 ;
  assign n3934 = ~n3783 & n3799 ;
  assign n3935 = ( n3783 & ~n3800 ) | ( n3783 & n3934 ) | ( ~n3800 & n3934 ) ;
  assign n3936 = n3933 & n3935 ;
  assign n3937 = n3800 | n3936 ;
  assign n3938 = n3762 & ~n3780 ;
  assign n3939 = ~n3762 & n3779 ;
  assign n3940 = n3938 | n3939 ;
  assign n3941 = n3937 & n3940 ;
  assign n3942 = n3780 | n3941 ;
  assign n3943 = n3741 & ~n3759 ;
  assign n3944 = ~n3741 & n3758 ;
  assign n3945 = n3943 | n3944 ;
  assign n3946 = n3759 | n3945 ;
  assign n3947 = ( n3759 & n3942 ) | ( n3759 & n3946 ) | ( n3942 & n3946 ) ;
  assign n3948 = n3720 | n3738 ;
  assign n3949 = ~n3739 & n3948 ;
  assign n3950 = n3739 | n3949 ;
  assign n3951 = ( n3739 & n3947 ) | ( n3739 & n3950 ) | ( n3947 & n3950 ) ;
  assign n3952 = n3718 & n3951 ;
  assign n3953 = n3716 | n3952 ;
  assign n3954 = ~n3679 & n3696 ;
  assign n3955 = ( n3679 & ~n3697 ) | ( n3679 & n3954 ) | ( ~n3697 & n3954 ) ;
  assign n3956 = n3697 | n3955 ;
  assign n3957 = ( n3697 & n3953 ) | ( n3697 & n3956 ) | ( n3953 & n3956 ) ;
  assign n3958 = n3673 | n3957 ;
  assign n3959 = ( n3673 & n3676 ) | ( n3673 & n3958 ) | ( n3676 & n3958 ) ;
  assign n3960 = ~n3650 & n3959 ;
  assign n3961 = n3647 | n3960 ;
  assign n3962 = n3622 | n3961 ;
  assign n3963 = ( n3622 & ~n3625 ) | ( n3622 & n3962 ) | ( ~n3625 & n3962 ) ;
  assign n3267 = n3003 | n3266 ;
  assign n3268 = ( n3003 & ~n3006 ) | ( n3003 & n3267 ) | ( ~n3006 & n3267 ) ;
  assign n2557 = n2365 | n2556 ;
  assign n1568 = n1552 | n1567 ;
  assign n1210 = ~n829 & n1065 ;
  assign n1211 = n692 & n1060 ;
  assign n1212 = ( n674 & n1060 ) | ( n674 & n1211 ) | ( n1060 & n1211 ) ;
  assign n1213 = n1210 | n1212 ;
  assign n1259 = n124 | n443 ;
  assign n1260 = n375 | n1259 ;
  assign n1261 = n764 | n801 ;
  assign n1262 = n1260 | n1261 ;
  assign n1263 = n333 | n1262 ;
  assign n1264 = n159 | n176 ;
  assign n1265 = n496 | n1264 ;
  assign n1266 = n637 | n1265 ;
  assign n1270 = n46 | n418 ;
  assign n1271 = n1269 | n1270 ;
  assign n1272 = n1266 | n1271 ;
  assign n1273 = n1263 | n1272 ;
  assign n1279 = n1273 | n1278 ;
  assign n1280 = n213 | n667 ;
  assign n1281 = n343 | n1280 ;
  assign n1282 = n162 | n591 ;
  assign n1283 = n340 | n431 ;
  assign n1284 = n1282 | n1283 ;
  assign n1285 = n1281 | n1284 ;
  assign n1287 = n223 | n388 ;
  assign n1288 = n1286 | n1287 ;
  assign n1289 = n460 | n1288 ;
  assign n1290 = n1285 | n1289 ;
  assign n1291 = n167 | n588 ;
  assign n1292 = n170 | n720 ;
  assign n1293 = n1291 | n1292 ;
  assign n1294 = n270 | n1293 ;
  assign n1295 = n151 | n1294 ;
  assign n1296 = n1290 | n1295 ;
  assign n1297 = n784 | n1296 ;
  assign n1298 = n1279 | n1297 ;
  assign n1299 = n1258 | n1298 ;
  assign n1300 = n272 | n513 ;
  assign n1302 = n680 | n1301 ;
  assign n1304 = n134 | n183 ;
  assign n1305 = n1303 | n1304 ;
  assign n1306 = n1302 | n1305 ;
  assign n1308 = n451 | n1307 ;
  assign n1309 = n222 | n1308 ;
  assign n1310 = n1306 | n1309 ;
  assign n1311 = n123 | n237 ;
  assign n1312 = n1310 | n1311 ;
  assign n1313 = n1300 | n1312 ;
  assign n1314 = n1299 | n1313 ;
  assign n1315 = n352 & n1057 ;
  assign n1316 = ( ~n339 & n1057 ) | ( ~n339 & n1315 ) | ( n1057 & n1315 ) ;
  assign n1317 = n1062 | n1316 ;
  assign n1318 = n1314 & n1317 ;
  assign n1319 = ( n1213 & n1314 ) | ( n1213 & n1318 ) | ( n1314 & n1318 ) ;
  assign n1320 = n1314 & n1316 ;
  assign n1321 = ( n1213 & n1314 ) | ( n1213 & n1320 ) | ( n1314 & n1320 ) ;
  assign n1322 = ( ~n1209 & n1319 ) | ( ~n1209 & n1321 ) | ( n1319 & n1321 ) ;
  assign n1323 = n1213 | n1316 ;
  assign n1324 = n1213 | n1317 ;
  assign n1325 = ( ~n1209 & n1323 ) | ( ~n1209 & n1324 ) | ( n1323 & n1324 ) ;
  assign n1326 = ~n1322 & n1325 ;
  assign n1327 = n1314 & ~n1324 ;
  assign n1328 = n1314 & ~n1323 ;
  assign n1329 = ( n1209 & n1327 ) | ( n1209 & n1328 ) | ( n1327 & n1328 ) ;
  assign n1330 = n1326 | n1329 ;
  assign n1847 = n1330 | n1568 ;
  assign n1848 = ~n1330 & n1847 ;
  assign n1849 = ( ~n1568 & n1847 ) | ( ~n1568 & n1848 ) | ( n1847 & n1848 ) ;
  assign n1853 = ~n523 & n1826 ;
  assign n1854 = n1793 & n1823 ;
  assign n1855 = ( n1783 & n1823 ) | ( n1783 & n1854 ) | ( n1823 & n1854 ) ;
  assign n1856 = n1853 | n1855 ;
  assign n1857 = n1708 & n1829 ;
  assign n1858 = n1856 | n1857 ;
  assign n1859 = n1821 | n1857 ;
  assign n1860 = n1856 | n1859 ;
  assign n1861 = ( ~n1852 & n1858 ) | ( ~n1852 & n1860 ) | ( n1858 & n1860 ) ;
  assign n1862 = ~x29 & n1860 ;
  assign n1863 = ~x29 & n1858 ;
  assign n1864 = ( ~n1852 & n1862 ) | ( ~n1852 & n1863 ) | ( n1862 & n1863 ) ;
  assign n1865 = x29 | n1863 ;
  assign n1866 = x29 | n1862 ;
  assign n1867 = ( ~n1852 & n1865 ) | ( ~n1852 & n1866 ) | ( n1865 & n1866 ) ;
  assign n1868 = ( ~n1861 & n1864 ) | ( ~n1861 & n1867 ) | ( n1864 & n1867 ) ;
  assign n1869 = n1847 & n1868 ;
  assign n1870 = ~n1568 & n1868 ;
  assign n1871 = ( n1848 & n1869 ) | ( n1848 & n1870 ) | ( n1869 & n1870 ) ;
  assign n1872 = n1849 & ~n1871 ;
  assign n1873 = ~n1847 & n1868 ;
  assign n1874 = n1568 & n1868 ;
  assign n1875 = ( ~n1848 & n1873 ) | ( ~n1848 & n1874 ) | ( n1873 & n1874 ) ;
  assign n1876 = n1872 | n1875 ;
  assign n2016 = ~n1901 & n2015 ;
  assign n2017 = ( n1901 & n2012 ) | ( n1901 & ~n2016 ) | ( n2012 & ~n2016 ) ;
  assign n2018 = n1876 & n2017 ;
  assign n2558 = n1876 | n2017 ;
  assign n2559 = ~n2018 & n2558 ;
  assign n2569 = n1634 & n2312 ;
  assign n2570 = ( n1630 & n2312 ) | ( n1630 & n2569 ) | ( n2312 & n2569 ) ;
  assign n2571 = n2279 & n2308 ;
  assign n2572 = ( ~n2269 & n2308 ) | ( ~n2269 & n2571 ) | ( n2308 & n2571 ) ;
  assign n2573 = n2570 | n2572 ;
  assign n2574 = n2090 & n2315 ;
  assign n2575 = ( ~n2082 & n2315 ) | ( ~n2082 & n2574 ) | ( n2315 & n2574 ) ;
  assign n2576 = n2573 | n2575 ;
  assign n2577 = n2306 | n2576 ;
  assign n2578 = n2576 & n2577 ;
  assign n2579 = ( n2568 & n2577 ) | ( n2568 & n2578 ) | ( n2577 & n2578 ) ;
  assign n2580 = x26 & n2578 ;
  assign n2581 = x26 & n2577 ;
  assign n2582 = ( n2568 & n2580 ) | ( n2568 & n2581 ) | ( n2580 & n2581 ) ;
  assign n2583 = x26 & ~n2580 ;
  assign n2584 = x26 & ~n2581 ;
  assign n2585 = ( ~n2568 & n2583 ) | ( ~n2568 & n2584 ) | ( n2583 & n2584 ) ;
  assign n2586 = ( n2579 & ~n2582 ) | ( n2579 & n2585 ) | ( ~n2582 & n2585 ) ;
  assign n2587 = n2559 & n2586 ;
  assign n2588 = n2559 & ~n2587 ;
  assign n2589 = ~n2559 & n2586 ;
  assign n2590 = n2588 | n2589 ;
  assign n2950 = ~n2557 & n2590 ;
  assign n2951 = n2557 & ~n2590 ;
  assign n2952 = n2950 | n2951 ;
  assign n2961 = n2701 & n2932 ;
  assign n2962 = ( ~n2784 & n2932 ) | ( ~n2784 & n2961 ) | ( n2932 & n2961 ) ;
  assign n2963 = n2691 & n2928 ;
  assign n2964 = ( n2678 & n2928 ) | ( n2678 & n2963 ) | ( n2928 & n2963 ) ;
  assign n2965 = n2962 | n2964 ;
  assign n2966 = n2199 & n2925 ;
  assign n2967 = ( ~n2185 & n2925 ) | ( ~n2185 & n2966 ) | ( n2925 & n2966 ) ;
  assign n2968 = n2965 | n2967 ;
  assign n2969 = n2936 | n2967 ;
  assign n2970 = n2965 | n2969 ;
  assign n2971 = ( n2960 & n2968 ) | ( n2960 & n2970 ) | ( n2968 & n2970 ) ;
  assign n2972 = x23 & n2970 ;
  assign n2973 = x23 & n2968 ;
  assign n2974 = ( n2960 & n2972 ) | ( n2960 & n2973 ) | ( n2972 & n2973 ) ;
  assign n2975 = x23 & ~n2973 ;
  assign n2976 = x23 & ~n2972 ;
  assign n2977 = ( ~n2960 & n2975 ) | ( ~n2960 & n2976 ) | ( n2975 & n2976 ) ;
  assign n2978 = ( n2971 & ~n2974 ) | ( n2971 & n2977 ) | ( ~n2974 & n2977 ) ;
  assign n2979 = n2952 & n2978 ;
  assign n3269 = n2952 | n2978 ;
  assign n3270 = ~n2979 & n3269 ;
  assign n3563 = n3268 & n3270 ;
  assign n3564 = n3268 | n3270 ;
  assign n3565 = ~n3563 & n3564 ;
  assign n3276 = n263 | n518 ;
  assign n3277 = n162 | n418 ;
  assign n3278 = n811 | n3277 ;
  assign n3279 = n64 | n1300 ;
  assign n3280 = n3278 | n3279 ;
  assign n3281 = n3276 | n3280 ;
  assign n3282 = n246 | n591 ;
  assign n3283 = n228 | n460 ;
  assign n3284 = n3282 | n3283 ;
  assign n3285 = n171 | n178 ;
  assign n3286 = n631 | n3285 ;
  assign n3287 = n3284 | n3286 ;
  assign n3288 = n142 | n901 ;
  assign n3289 = ( n133 & n468 ) | ( n133 & ~n3288 ) | ( n468 & ~n3288 ) ;
  assign n3290 = n3288 | n3289 ;
  assign n3291 = n3287 | n3290 ;
  assign n3292 = n245 | n3291 ;
  assign n3293 = n177 | n282 ;
  assign n3294 = n226 | n1678 ;
  assign n3295 = n3293 | n3294 ;
  assign n3296 = n118 | n305 ;
  assign n3297 = n2146 | n3296 ;
  assign n3298 = n689 | n858 ;
  assign n3299 = n3297 | n3298 ;
  assign n3300 = n3295 | n3299 ;
  assign n3301 = n324 | n3300 ;
  assign n3302 = n3292 | n3301 ;
  assign n3303 = n3281 | n3302 ;
  assign n3304 = n110 | n183 ;
  assign n3305 = n1394 | n3304 ;
  assign n3306 = n2623 | n3305 ;
  assign n3307 = n1760 | n3306 ;
  assign n3308 = n284 | n1039 ;
  assign n3309 = n240 | n269 ;
  assign n3310 = n3308 | n3309 ;
  assign n3311 = n254 | n3310 ;
  assign n3312 = n343 | n675 ;
  assign n3313 = n128 | n190 ;
  assign n3314 = n3312 | n3313 ;
  assign n3315 = n3311 | n3314 ;
  assign n3316 = n3307 | n3315 ;
  assign n3317 = n1286 | n3316 ;
  assign n3318 = n445 | n478 ;
  assign n3319 = n2863 | n3318 ;
  assign n3320 = n479 | n574 ;
  assign n3321 = n401 | n510 ;
  assign n3322 = n3320 | n3321 ;
  assign n3323 = n3319 | n3322 ;
  assign n1193 = n309 | n424 ;
  assign n3324 = n568 | n886 ;
  assign n3325 = n1193 | n3324 ;
  assign n3326 = n487 | n3325 ;
  assign n3327 = n1287 | n3326 ;
  assign n3328 = n3323 | n3327 ;
  assign n3329 = n939 | n1126 ;
  assign n3330 = n77 | n624 ;
  assign n3331 = n152 | n3330 ;
  assign n3332 = n3329 | n3331 ;
  assign n3333 = n616 | n801 ;
  assign n3334 = n694 | n3333 ;
  assign n3335 = n3332 | n3334 ;
  assign n3336 = n3328 | n3335 ;
  assign n3337 = n3317 | n3336 ;
  assign n3338 = n3303 | n3337 ;
  assign n3339 = n357 | n807 ;
  assign n3340 = n2809 | n3339 ;
  assign n3341 = n99 | n432 ;
  assign n3342 = n469 | n3341 ;
  assign n3343 = n198 | n3342 ;
  assign n3344 = n3340 | n3343 ;
  assign n3345 = n354 | n3344 ;
  assign n1116 = n46 | n247 ;
  assign n3346 = n370 | n457 ;
  assign n3347 = n255 | n3346 ;
  assign n3348 = n1116 | n3347 ;
  assign n3349 = n160 | n735 ;
  assign n3350 = n514 | n3349 ;
  assign n3351 = n643 | n839 ;
  assign n3352 = n213 | n1114 ;
  assign n3353 = n3351 | n3352 ;
  assign n3354 = n3350 | n3353 ;
  assign n3355 = n348 | n887 ;
  assign n3356 = n3354 | n3355 ;
  assign n3357 = n3348 | n3356 ;
  assign n3358 = n296 | n602 ;
  assign n3359 = n438 | n3358 ;
  assign n3360 = n141 | n262 ;
  assign n3361 = n3359 | n3360 ;
  assign n3362 = n273 | n283 ;
  assign n3363 = n117 | n644 ;
  assign n3364 = n501 | n560 ;
  assign n3365 = n3363 | n3364 ;
  assign n3366 = ( ~n3361 & n3362 ) | ( ~n3361 & n3365 ) | ( n3362 & n3365 ) ;
  assign n3367 = n103 | n250 ;
  assign n3368 = n333 | n3367 ;
  assign n3369 = n3361 | n3368 ;
  assign n3370 = n3366 | n3369 ;
  assign n3371 = n3357 | n3370 ;
  assign n3372 = n197 | n225 ;
  assign n3373 = n758 | n3372 ;
  assign n3374 = n402 | n725 ;
  assign n3375 = n239 | n3374 ;
  assign n3376 = n406 | n489 ;
  assign n3377 = n2047 | n3376 ;
  assign n3378 = n3375 | n3377 ;
  assign n3379 = n163 | n387 ;
  assign n3380 = n447 | n3379 ;
  assign n3381 = n3378 | n3380 ;
  assign n3382 = n3373 | n3381 ;
  assign n3383 = n849 | n3382 ;
  assign n3384 = n3371 | n3383 ;
  assign n3385 = n3345 | n3384 ;
  assign n3386 = n3338 | n3385 ;
  assign n3509 = n3386 & n3508 ;
  assign n3510 = n3386 | n3508 ;
  assign n3511 = ~n3509 & n3510 ;
  assign n3522 = ~n3515 & n3521 ;
  assign n3524 = ~n3515 & n3523 ;
  assign n3525 = ( n2602 & n3522 ) | ( n2602 & n3524 ) | ( n3522 & n3524 ) ;
  assign n3566 = n3511 & ~n3525 ;
  assign n3567 = ~n3511 & n3525 ;
  assign n3568 = n3566 | n3567 ;
  assign n3569 = n2893 & n3544 ;
  assign n3570 = ( ~n2886 & n3544 ) | ( ~n2886 & n3569 ) | ( n3544 & n3569 ) ;
  assign n3571 = n3507 & n3541 ;
  assign n3572 = ( n3483 & n3541 ) | ( n3483 & n3571 ) | ( n3541 & n3571 ) ;
  assign n3573 = n3570 | n3572 ;
  assign n3574 = n3537 | n3547 ;
  assign n3575 = ( n3386 & n3537 ) | ( n3386 & n3574 ) | ( n3537 & n3574 ) ;
  assign n3576 = n3573 | n3575 ;
  assign n3577 = n3386 & n3547 ;
  assign n3578 = n3573 | n3577 ;
  assign n3579 = n3576 & n3578 ;
  assign n3580 = ( ~n3568 & n3576 ) | ( ~n3568 & n3579 ) | ( n3576 & n3579 ) ;
  assign n3581 = ~x20 & n3579 ;
  assign n3582 = ~x20 & n3576 ;
  assign n3583 = ( ~n3568 & n3581 ) | ( ~n3568 & n3582 ) | ( n3581 & n3582 ) ;
  assign n3584 = x20 | n3581 ;
  assign n3585 = x20 | n3582 ;
  assign n3586 = ( ~n3568 & n3584 ) | ( ~n3568 & n3585 ) | ( n3584 & n3585 ) ;
  assign n3587 = ( ~n3580 & n3583 ) | ( ~n3580 & n3586 ) | ( n3583 & n3586 ) ;
  assign n3588 = n3565 & n3587 ;
  assign n3589 = n3565 & ~n3588 ;
  assign n3590 = ~n3565 & n3587 ;
  assign n3591 = n3589 | n3590 ;
  assign n3964 = n3591 & n3963 ;
  assign n4519 = n3963 & ~n3964 ;
  assign n4520 = n3591 & ~n3964 ;
  assign n4521 = n4519 | n4520 ;
  assign n4142 = n590 | n608 ;
  assign n4143 = n3323 | n3326 ;
  assign n4144 = n296 | n456 ;
  assign n4145 = n291 | n841 ;
  assign n4146 = n4144 | n4145 ;
  assign n4147 = n767 | n4146 ;
  assign n4148 = n2613 | n4147 ;
  assign n4149 = n4143 | n4148 ;
  assign n4150 = n4142 | n4149 ;
  assign n4151 = n341 | n418 ;
  assign n4152 = n239 | n313 ;
  assign n4153 = n4151 | n4152 ;
  assign n4154 = n720 | n1126 ;
  assign n4155 = n4153 | n4154 ;
  assign n4156 = n432 | n489 ;
  assign n4157 = n689 | n4156 ;
  assign n4158 = n4155 | n4157 ;
  assign n4159 = n2649 | n4158 ;
  assign n4160 = n4150 | n4159 ;
  assign n4161 = n702 | n967 ;
  assign n4162 = n170 | n483 ;
  assign n4163 = n542 | n4162 ;
  assign n4164 = n4161 | n4163 ;
  assign n4165 = n92 | n395 ;
  assign n4166 = n302 | n4165 ;
  assign n4167 = n234 | n4166 ;
  assign n4168 = n4164 | n4167 ;
  assign n4169 = n305 | n4168 ;
  assign n4170 = n497 | n500 ;
  assign n4171 = n744 | n4170 ;
  assign n4172 = n3445 | n3485 ;
  assign n4173 = n4171 | n4172 ;
  assign n4174 = n262 | n284 ;
  assign n4175 = ( n1013 & n1785 ) | ( n1013 & ~n4174 ) | ( n1785 & ~n4174 ) ;
  assign n4176 = n4174 | n4175 ;
  assign n4177 = n303 | n381 ;
  assign n4178 = n4176 | n4177 ;
  assign n4179 = n4173 | n4178 ;
  assign n4180 = n53 | n236 ;
  assign n4181 = n317 | n503 ;
  assign n4182 = n1030 | n4181 ;
  assign n4183 = n4180 | n4182 ;
  assign n4184 = n94 | n278 ;
  assign n3430 = n110 | n588 ;
  assign n4185 = n167 | n735 ;
  assign n4186 = n3430 | n4185 ;
  assign n4187 = n4184 | n4186 ;
  assign n4188 = n4183 | n4187 ;
  assign n4189 = n527 | n1484 ;
  assign n4190 = n1661 | n4189 ;
  assign n4191 = n4188 | n4190 ;
  assign n4192 = n4179 | n4191 ;
  assign n4193 = n190 | n331 ;
  assign n4194 = n39 | n355 ;
  assign n4195 = n4193 | n4194 ;
  assign n4196 = n225 | n4195 ;
  assign n4197 = n117 | n325 ;
  assign n4198 = n2117 | n4197 ;
  assign n4199 = n2040 | n4198 ;
  assign n4200 = n140 | n202 ;
  assign n4201 = n959 | n4200 ;
  assign n4202 = n4199 | n4201 ;
  assign n4203 = n4196 | n4202 ;
  assign n4204 = n4192 | n4203 ;
  assign n4205 = n4169 | n4204 ;
  assign n4206 = n4160 | n4205 ;
  assign n4305 = n448 | n1355 ;
  assign n4306 = n203 | n901 ;
  assign n4307 = n1303 | n4306 ;
  assign n4308 = n4305 | n4307 ;
  assign n4309 = n249 | n938 ;
  assign n4310 = n237 | n517 ;
  assign n4311 = n4309 | n4310 ;
  assign n4312 = n222 | n959 ;
  assign n4313 = n527 | n560 ;
  assign n4314 = n4312 | n4313 ;
  assign n4315 = n4311 | n4314 ;
  assign n4316 = n4308 | n4315 ;
  assign n4317 = n2248 | n4316 ;
  assign n4318 = n663 | n1615 ;
  assign n4319 = n2040 | n4318 ;
  assign n4320 = n71 | n90 ;
  assign n4321 = n4319 | n4320 ;
  assign n4322 = n4317 | n4321 ;
  assign n4323 = n937 | n1380 ;
  assign n4324 = n92 | n1005 ;
  assign n4325 = n4323 | n4324 ;
  assign n4326 = n291 | n4325 ;
  assign n4257 = n356 | n820 ;
  assign n4258 = n305 | n4257 ;
  assign n4400 = n1370 | n4258 ;
  assign n4401 = n1346 | n4400 ;
  assign n4402 = n53 | n591 ;
  assign n4403 = n666 | n841 ;
  assign n4404 = n4402 | n4403 ;
  assign n4405 = n141 | n160 ;
  assign n4406 = n4404 | n4405 ;
  assign n4407 = n4401 | n4406 ;
  assign n4408 = n4326 | n4407 ;
  assign n4409 = n4322 | n4408 ;
  assign n4410 = n349 | n581 ;
  assign n4411 = n1714 | n4410 ;
  assign n4412 = n371 | n649 ;
  assign n4413 = n4411 | n4412 ;
  assign n4293 = n324 | n542 ;
  assign n4414 = n321 | n631 ;
  assign n4415 = n4293 | n4414 ;
  assign n4416 = n110 | n689 ;
  assign n4417 = n2805 | n4416 ;
  assign n4418 = n4415 | n4417 ;
  assign n4419 = n4413 | n4418 ;
  assign n4420 = n2609 | n4419 ;
  assign n4421 = n4409 | n4420 ;
  assign n4422 = n550 | n1465 ;
  assign n4423 = n124 | n239 ;
  assign n4424 = n401 | n4423 ;
  assign n4425 = n4422 | n4424 ;
  assign n4426 = n281 | n348 ;
  assign n4427 = n4425 | n4426 ;
  assign n4428 = n742 & ~n4427 ;
  assign n4429 = ~n4421 & n4428 ;
  assign n4436 = n4206 & ~n4429 ;
  assign n4437 = ~n4206 & n4429 ;
  assign n4438 = n4436 | n4437 ;
  assign n3387 = n937 | n2050 ;
  assign n3388 = n331 | n3387 ;
  assign n1127 = n600 | n901 ;
  assign n3389 = n94 | n369 ;
  assign n3390 = n281 | n3389 ;
  assign n3391 = n1127 | n3390 ;
  assign n3392 = n3388 | n3391 ;
  assign n3393 = n39 | n160 ;
  assign n3394 = n212 | n258 ;
  assign n3395 = n821 | n3394 ;
  assign n3396 = n3393 | n3395 ;
  assign n3397 = n877 & ~n3396 ;
  assign n3398 = ~n3392 & n3397 ;
  assign n3399 = n807 | n3360 ;
  assign n3400 = n3359 | n3399 ;
  assign n3401 = n550 | n3400 ;
  assign n3402 = n179 | n292 ;
  assign n3403 = n1005 | n3402 ;
  assign n3404 = n77 | n513 ;
  assign n3405 = n3403 | n3404 ;
  assign n3406 = n3401 | n3405 ;
  assign n3407 = n3398 & ~n3406 ;
  assign n3408 = ~n659 & n3407 ;
  assign n3409 = n291 | n489 ;
  assign n3410 = n263 | n527 ;
  assign n3411 = n3409 | n3410 ;
  assign n3412 = n272 | n416 ;
  assign n3413 = n381 | n480 ;
  assign n3414 = n198 | n3413 ;
  assign n3415 = n3412 | n3414 ;
  assign n3416 = n1617 | n3415 ;
  assign n3417 = n3411 | n3416 ;
  assign n3418 = n1360 | n3417 ;
  assign n3419 = n1354 | n3418 ;
  assign n3420 = n3408 & ~n3419 ;
  assign n3421 = n309 | n450 ;
  assign n3422 = n468 | n3421 ;
  assign n3423 = n2840 | n3422 ;
  assign n3424 = n696 | n735 ;
  assign n3425 = n372 | n1114 ;
  assign n3426 = n128 | n246 ;
  assign n3427 = n3425 | n3426 ;
  assign n3428 = n3424 | n3427 ;
  assign n3429 = n3423 | n3428 ;
  assign n3431 = n401 | n566 ;
  assign n3432 = n3430 | n3431 ;
  assign n3433 = n608 | n3432 ;
  assign n3434 = n574 | n3433 ;
  assign n3435 = n3429 | n3434 ;
  assign n3436 = n388 | n720 ;
  assign n3437 = n465 | n501 ;
  assign n3438 = n3436 | n3437 ;
  assign n3439 = n3435 | n3438 ;
  assign n3440 = n3420 & ~n3439 ;
  assign n4207 = ~n3440 & n4206 ;
  assign n3441 = n3386 & ~n3440 ;
  assign n3442 = ~n3386 & n3440 ;
  assign n3443 = n3441 | n3442 ;
  assign n4213 = n3441 | n3509 ;
  assign n4214 = ( n3441 & ~n3443 ) | ( n3441 & n4213 ) | ( ~n3443 & n4213 ) ;
  assign n4208 = n3440 & ~n4206 ;
  assign n4209 = n4207 | n4208 ;
  assign n4439 = ~n4207 & n4209 ;
  assign n4440 = ( n4207 & n4214 ) | ( n4207 & ~n4439 ) | ( n4214 & ~n4439 ) ;
  assign n4441 = ~n4438 & n4440 ;
  assign n3512 = n3509 | n3511 ;
  assign n4210 = ~n3441 & n3443 ;
  assign n4211 = ( n3441 & n3512 ) | ( n3441 & ~n4210 ) | ( n3512 & ~n4210 ) ;
  assign n4444 = n4438 | n4439 ;
  assign n4445 = n4207 & ~n4438 ;
  assign n4446 = ( n4211 & ~n4444 ) | ( n4211 & n4445 ) | ( ~n4444 & n4445 ) ;
  assign n4522 = ( ~n3525 & n4441 ) | ( ~n3525 & n4446 ) | ( n4441 & n4446 ) ;
  assign n4523 = ( n4207 & n4211 ) | ( n4207 & ~n4439 ) | ( n4211 & ~n4439 ) ;
  assign n4524 = n4438 & ~n4523 ;
  assign n4525 = n4438 & ~n4440 ;
  assign n4526 = ( n3525 & n4524 ) | ( n3525 & n4525 ) | ( n4524 & n4525 ) ;
  assign n4527 = n4522 | n4526 ;
  assign n4456 = ~x15 & x16 ;
  assign n4457 = x15 & ~x16 ;
  assign n4458 = n4456 | n4457 ;
  assign n4459 = x14 & ~x15 ;
  assign n4460 = ~x14 & x15 ;
  assign n4461 = n4459 | n4460 ;
  assign n4468 = n4458 & ~n4461 ;
  assign n4528 = n4206 & n4468 ;
  assign n4462 = x16 & ~x17 ;
  assign n4463 = ~x16 & x17 ;
  assign n4464 = n4462 | n4463 ;
  assign n4471 = n4461 & ~n4464 ;
  assign n4529 = ~n4429 & n4471 ;
  assign n4465 = ~n4461 & n4464 ;
  assign n4466 = ~n4458 & n4465 ;
  assign n4530 = n3439 & n4466 ;
  assign n4531 = ( ~n3420 & n4466 ) | ( ~n3420 & n4530 ) | ( n4466 & n4530 ) ;
  assign n4532 = n4529 | n4531 ;
  assign n4533 = n4528 | n4532 ;
  assign n4475 = n4461 & n4464 ;
  assign n4534 = n4475 | n4528 ;
  assign n4535 = n4532 | n4534 ;
  assign n4536 = ( ~n4527 & n4533 ) | ( ~n4527 & n4535 ) | ( n4533 & n4535 ) ;
  assign n4537 = ~x17 & n4535 ;
  assign n4538 = ~x17 & n4533 ;
  assign n4539 = ( ~n4527 & n4537 ) | ( ~n4527 & n4538 ) | ( n4537 & n4538 ) ;
  assign n4540 = x17 | n4538 ;
  assign n4541 = x17 | n4537 ;
  assign n4542 = ( ~n4527 & n4540 ) | ( ~n4527 & n4541 ) | ( n4540 & n4541 ) ;
  assign n4543 = ( ~n4536 & n4539 ) | ( ~n4536 & n4542 ) | ( n4539 & n4542 ) ;
  assign n4544 = n4521 & n4543 ;
  assign n4545 = n4521 & ~n4544 ;
  assign n4546 = ~n4521 & n4543 ;
  assign n4547 = n4545 | n4546 ;
  assign n4548 = ~n3625 & n3961 ;
  assign n4549 = n3625 | n4548 ;
  assign n4212 = ~n4209 & n4211 ;
  assign n4215 = ~n4209 & n4214 ;
  assign n4216 = ( ~n3525 & n4212 ) | ( ~n3525 & n4215 ) | ( n4212 & n4215 ) ;
  assign n4217 = n4209 & ~n4211 ;
  assign n4218 = n4209 & ~n4214 ;
  assign n4219 = ( n3525 & n4217 ) | ( n3525 & n4218 ) | ( n4217 & n4218 ) ;
  assign n4220 = n4216 | n4219 ;
  assign n4552 = n4206 & n4471 ;
  assign n4553 = n3386 & n4466 ;
  assign n4554 = n3439 & n4468 ;
  assign n4555 = ( ~n3420 & n4468 ) | ( ~n3420 & n4554 ) | ( n4468 & n4554 ) ;
  assign n4556 = n4553 | n4555 ;
  assign n4557 = n4552 | n4556 ;
  assign n4558 = n4475 | n4552 ;
  assign n4559 = n4556 | n4558 ;
  assign n4560 = ( ~n4220 & n4557 ) | ( ~n4220 & n4559 ) | ( n4557 & n4559 ) ;
  assign n4561 = ~x17 & n4559 ;
  assign n4562 = ~x17 & n4557 ;
  assign n4563 = ( ~n4220 & n4561 ) | ( ~n4220 & n4562 ) | ( n4561 & n4562 ) ;
  assign n4564 = x17 | n4562 ;
  assign n4565 = x17 | n4561 ;
  assign n4566 = ( ~n4220 & n4564 ) | ( ~n4220 & n4565 ) | ( n4564 & n4565 ) ;
  assign n4567 = ( ~n4560 & n4563 ) | ( ~n4560 & n4566 ) | ( n4563 & n4566 ) ;
  assign n4550 = n3625 & n3961 ;
  assign n4568 = n4550 & n4567 ;
  assign n4569 = ( ~n4549 & n4567 ) | ( ~n4549 & n4568 ) | ( n4567 & n4568 ) ;
  assign n4551 = n4549 & ~n4550 ;
  assign n4570 = n4551 | n4569 ;
  assign n4571 = ~n4550 & n4567 ;
  assign n4572 = n4549 & n4571 ;
  assign n4573 = n4570 & ~n4572 ;
  assign n4574 = n3959 & ~n3960 ;
  assign n4575 = n3650 | n3960 ;
  assign n4576 = ~n4574 & n4575 ;
  assign n3513 = ~n3443 & n3512 ;
  assign n3514 = ~n3443 & n3509 ;
  assign n3526 = ( n3513 & n3514 ) | ( n3513 & ~n3525 ) | ( n3514 & ~n3525 ) ;
  assign n3527 = ~n3386 & n3443 ;
  assign n3528 = n3443 & ~n3508 ;
  assign n3529 = ( n3525 & n3527 ) | ( n3525 & n3528 ) | ( n3527 & n3528 ) ;
  assign n3530 = n3526 | n3529 ;
  assign n4577 = n3386 & n4468 ;
  assign n4578 = n3507 & n4466 ;
  assign n4579 = ( n3483 & n4466 ) | ( n3483 & n4578 ) | ( n4466 & n4578 ) ;
  assign n4580 = n3439 & n4471 ;
  assign n4581 = ( ~n3420 & n4471 ) | ( ~n3420 & n4580 ) | ( n4471 & n4580 ) ;
  assign n4582 = n4579 | n4581 ;
  assign n4583 = n4577 | n4582 ;
  assign n4584 = n4475 | n4583 ;
  assign n4585 = ( ~n3530 & n4583 ) | ( ~n3530 & n4584 ) | ( n4583 & n4584 ) ;
  assign n4586 = ~x17 & n4584 ;
  assign n4587 = ~x17 & n4583 ;
  assign n4588 = ( ~n3530 & n4586 ) | ( ~n3530 & n4587 ) | ( n4586 & n4587 ) ;
  assign n4589 = x17 | n4586 ;
  assign n4590 = x17 | n4587 ;
  assign n4591 = ( ~n3530 & n4589 ) | ( ~n3530 & n4590 ) | ( n4589 & n4590 ) ;
  assign n4592 = ( ~n4585 & n4588 ) | ( ~n4585 & n4591 ) | ( n4588 & n4591 ) ;
  assign n4593 = ~n4576 & n4592 ;
  assign n4594 = n4576 | n4593 ;
  assign n4595 = n4576 & n4592 ;
  assign n4596 = n4594 & ~n4595 ;
  assign n4597 = n3676 & n3957 ;
  assign n4598 = n3676 & ~n4597 ;
  assign n4601 = n2893 & n4466 ;
  assign n4602 = ( ~n2886 & n4466 ) | ( ~n2886 & n4601 ) | ( n4466 & n4601 ) ;
  assign n4603 = n3507 & n4468 ;
  assign n4604 = ( n3483 & n4468 ) | ( n3483 & n4603 ) | ( n4468 & n4603 ) ;
  assign n4605 = n4602 | n4604 ;
  assign n4606 = n3386 & n4471 ;
  assign n4607 = n4605 | n4606 ;
  assign n4608 = n4475 | n4606 ;
  assign n4609 = n4605 | n4608 ;
  assign n4610 = ( ~n3568 & n4607 ) | ( ~n3568 & n4609 ) | ( n4607 & n4609 ) ;
  assign n4611 = ~x17 & n4609 ;
  assign n4612 = ~x17 & n4607 ;
  assign n4613 = ( ~n3568 & n4611 ) | ( ~n3568 & n4612 ) | ( n4611 & n4612 ) ;
  assign n4614 = x17 | n4612 ;
  assign n4615 = x17 | n4611 ;
  assign n4616 = ( ~n3568 & n4614 ) | ( ~n3568 & n4615 ) | ( n4614 & n4615 ) ;
  assign n4617 = ( ~n4610 & n4613 ) | ( ~n4610 & n4616 ) | ( n4613 & n4616 ) ;
  assign n4599 = ~n3676 & n3957 ;
  assign n4618 = n4599 & n4617 ;
  assign n4619 = ( n4598 & n4617 ) | ( n4598 & n4618 ) | ( n4617 & n4618 ) ;
  assign n4600 = n4598 | n4599 ;
  assign n4620 = n4600 & ~n4619 ;
  assign n4621 = ~n4599 & n4617 ;
  assign n4622 = ~n4598 & n4621 ;
  assign n4623 = n4620 | n4622 ;
  assign n4624 = n3718 | n3951 ;
  assign n4625 = ~n3952 & n4624 ;
  assign n4626 = n2691 & n4466 ;
  assign n4627 = ( n2678 & n4466 ) | ( n2678 & n4626 ) | ( n4466 & n4626 ) ;
  assign n4628 = n2701 & n4468 ;
  assign n4629 = ( ~n2784 & n4468 ) | ( ~n2784 & n4628 ) | ( n4468 & n4628 ) ;
  assign n4630 = n4627 | n4629 ;
  assign n4631 = n2893 & n4471 ;
  assign n4632 = ( ~n2886 & n4471 ) | ( ~n2886 & n4631 ) | ( n4471 & n4631 ) ;
  assign n4633 = n4630 | n4632 ;
  assign n4634 = n4475 | n4633 ;
  assign n4635 = n4633 & n4634 ;
  assign n4636 = ( ~n2914 & n4634 ) | ( ~n2914 & n4635 ) | ( n4634 & n4635 ) ;
  assign n4637 = ~x17 & n4635 ;
  assign n4638 = ~x17 & n4634 ;
  assign n4639 = ( ~n2914 & n4637 ) | ( ~n2914 & n4638 ) | ( n4637 & n4638 ) ;
  assign n4640 = x17 | n4637 ;
  assign n4641 = x17 | n4638 ;
  assign n4642 = ( ~n2914 & n4640 ) | ( ~n2914 & n4641 ) | ( n4640 & n4641 ) ;
  assign n4643 = ( ~n4636 & n4639 ) | ( ~n4636 & n4642 ) | ( n4639 & n4642 ) ;
  assign n4644 = n4625 & n4643 ;
  assign n4645 = n3953 & n3955 ;
  assign n4646 = n3953 | n3955 ;
  assign n4647 = ~n4645 & n4646 ;
  assign n4648 = n2893 & n4468 ;
  assign n4649 = ( ~n2886 & n4468 ) | ( ~n2886 & n4648 ) | ( n4468 & n4648 ) ;
  assign n4650 = n2701 & n4466 ;
  assign n4651 = ( ~n2784 & n4466 ) | ( ~n2784 & n4650 ) | ( n4466 & n4650 ) ;
  assign n4652 = n3507 & n4471 ;
  assign n4653 = ( n3483 & n4471 ) | ( n3483 & n4652 ) | ( n4471 & n4652 ) ;
  assign n4654 = n4651 | n4653 ;
  assign n4655 = n4649 | n4654 ;
  assign n4656 = n4475 | n4655 ;
  assign n4657 = n4655 & n4656 ;
  assign n4658 = ( n3603 & n4656 ) | ( n3603 & n4657 ) | ( n4656 & n4657 ) ;
  assign n4659 = x17 & n4657 ;
  assign n4660 = x17 & n4656 ;
  assign n4661 = ( n3603 & n4659 ) | ( n3603 & n4660 ) | ( n4659 & n4660 ) ;
  assign n4662 = x17 & ~n4659 ;
  assign n4663 = x17 & ~n4660 ;
  assign n4664 = ( ~n3603 & n4662 ) | ( ~n3603 & n4663 ) | ( n4662 & n4663 ) ;
  assign n4665 = ( n4658 & ~n4661 ) | ( n4658 & n4664 ) | ( ~n4661 & n4664 ) ;
  assign n4666 = n4647 & n4665 ;
  assign n4667 = n4647 | n4665 ;
  assign n4668 = ~n4666 & n4667 ;
  assign n4669 = n4644 & n4668 ;
  assign n4670 = n4666 | n4668 ;
  assign n4671 = n4625 & ~n4644 ;
  assign n4672 = ~n4625 & n4643 ;
  assign n4673 = n4671 | n4672 ;
  assign n4674 = n3947 & n3949 ;
  assign n4675 = n3947 | n3949 ;
  assign n4676 = ~n4674 & n4675 ;
  assign n4677 = n2701 & n4471 ;
  assign n4678 = ( ~n2784 & n4471 ) | ( ~n2784 & n4677 ) | ( n4471 & n4677 ) ;
  assign n4679 = n2691 & n4468 ;
  assign n4680 = ( n2678 & n4468 ) | ( n2678 & n4679 ) | ( n4468 & n4679 ) ;
  assign n4681 = n4678 | n4680 ;
  assign n4682 = n2199 & n4466 ;
  assign n4683 = ( ~n2185 & n4466 ) | ( ~n2185 & n4682 ) | ( n4466 & n4682 ) ;
  assign n4684 = n4681 | n4683 ;
  assign n4685 = n4475 | n4683 ;
  assign n4686 = n4681 | n4685 ;
  assign n4687 = ( n2960 & n4684 ) | ( n2960 & n4686 ) | ( n4684 & n4686 ) ;
  assign n4688 = x17 & n4686 ;
  assign n4689 = x17 & n4684 ;
  assign n4690 = ( n2960 & n4688 ) | ( n2960 & n4689 ) | ( n4688 & n4689 ) ;
  assign n4691 = x17 & ~n4689 ;
  assign n4692 = x17 & ~n4688 ;
  assign n4693 = ( ~n2960 & n4691 ) | ( ~n2960 & n4692 ) | ( n4691 & n4692 ) ;
  assign n4694 = ( n4687 & ~n4690 ) | ( n4687 & n4693 ) | ( ~n4690 & n4693 ) ;
  assign n4695 = n4676 & n4694 ;
  assign n4696 = n3942 & n3945 ;
  assign n4697 = n3942 & ~n4696 ;
  assign n4700 = n2090 & n4466 ;
  assign n4701 = ( ~n2082 & n4466 ) | ( ~n2082 & n4700 ) | ( n4466 & n4700 ) ;
  assign n4702 = n2691 & n4471 ;
  assign n4703 = ( n2678 & n4471 ) | ( n2678 & n4702 ) | ( n4471 & n4702 ) ;
  assign n4704 = n2199 & n4468 ;
  assign n4705 = ( ~n2185 & n4468 ) | ( ~n2185 & n4704 ) | ( n4468 & n4704 ) ;
  assign n4706 = n4703 | n4705 ;
  assign n4707 = n4701 | n4706 ;
  assign n4708 = n4475 | n4707 ;
  assign n4709 = ( n2985 & n4707 ) | ( n2985 & n4708 ) | ( n4707 & n4708 ) ;
  assign n4710 = x17 & n4708 ;
  assign n4711 = x17 & n4707 ;
  assign n4712 = ( n2985 & n4710 ) | ( n2985 & n4711 ) | ( n4710 & n4711 ) ;
  assign n4713 = x17 & ~n4710 ;
  assign n4714 = x17 & ~n4711 ;
  assign n4715 = ( ~n2985 & n4713 ) | ( ~n2985 & n4714 ) | ( n4713 & n4714 ) ;
  assign n4716 = ( n4709 & ~n4712 ) | ( n4709 & n4715 ) | ( ~n4712 & n4715 ) ;
  assign n4698 = ~n3942 & n3945 ;
  assign n4717 = n4698 & n4716 ;
  assign n4718 = ( n4697 & n4716 ) | ( n4697 & n4717 ) | ( n4716 & n4717 ) ;
  assign n4699 = n4697 | n4698 ;
  assign n4719 = n4699 & ~n4718 ;
  assign n4720 = ~n4698 & n4716 ;
  assign n4721 = ~n4697 & n4720 ;
  assign n4722 = n4719 | n4721 ;
  assign n4723 = ~n3937 & n3940 ;
  assign n4724 = n3937 & ~n3940 ;
  assign n4725 = n4723 | n4724 ;
  assign n4726 = n2090 & n4468 ;
  assign n4727 = ( ~n2082 & n4468 ) | ( ~n2082 & n4726 ) | ( n4468 & n4726 ) ;
  assign n4728 = n2279 & n4466 ;
  assign n4729 = ( ~n2269 & n4466 ) | ( ~n2269 & n4728 ) | ( n4466 & n4728 ) ;
  assign n4730 = n2199 & n4471 ;
  assign n4731 = ( ~n2185 & n4471 ) | ( ~n2185 & n4730 ) | ( n4471 & n4730 ) ;
  assign n4732 = n4729 | n4731 ;
  assign n4733 = n4727 | n4732 ;
  assign n4734 = n4475 | n4733 ;
  assign n4735 = ( ~n2325 & n4733 ) | ( ~n2325 & n4734 ) | ( n4733 & n4734 ) ;
  assign n4736 = n4733 & n4734 ;
  assign n4737 = ( ~n2299 & n4735 ) | ( ~n2299 & n4736 ) | ( n4735 & n4736 ) ;
  assign n4738 = ~x17 & n4737 ;
  assign n4739 = x17 | n4737 ;
  assign n4740 = ( ~n4737 & n4738 ) | ( ~n4737 & n4739 ) | ( n4738 & n4739 ) ;
  assign n4741 = n4725 & n4740 ;
  assign n4742 = n4725 | n4740 ;
  assign n4743 = ~n4741 & n4742 ;
  assign n4744 = n3933 | n3935 ;
  assign n4745 = ~n3936 & n4744 ;
  assign n4746 = n1634 & n4466 ;
  assign n4747 = ( n1630 & n4466 ) | ( n1630 & n4746 ) | ( n4466 & n4746 ) ;
  assign n4748 = n2279 & n4468 ;
  assign n4749 = ( ~n2269 & n4468 ) | ( ~n2269 & n4748 ) | ( n4468 & n4748 ) ;
  assign n4750 = n4747 | n4749 ;
  assign n4751 = n2090 & n4471 ;
  assign n4752 = ( ~n2082 & n4471 ) | ( ~n2082 & n4751 ) | ( n4471 & n4751 ) ;
  assign n4753 = n4750 | n4752 ;
  assign n4754 = n4475 | n4753 ;
  assign n4755 = n4753 & n4754 ;
  assign n4756 = ( n2568 & n4754 ) | ( n2568 & n4755 ) | ( n4754 & n4755 ) ;
  assign n4757 = x17 & n4755 ;
  assign n4758 = x17 & n4754 ;
  assign n4759 = ( n2568 & n4757 ) | ( n2568 & n4758 ) | ( n4757 & n4758 ) ;
  assign n4760 = x17 & ~n4757 ;
  assign n4761 = x17 & ~n4758 ;
  assign n4762 = ( ~n2568 & n4760 ) | ( ~n2568 & n4761 ) | ( n4760 & n4761 ) ;
  assign n4763 = ( n4756 & ~n4759 ) | ( n4756 & n4762 ) | ( ~n4759 & n4762 ) ;
  assign n4764 = n4745 & n4763 ;
  assign n4765 = n3823 | n3931 ;
  assign n4766 = ~n3932 & n4765 ;
  assign n4767 = n1708 & n4466 ;
  assign n4768 = n1634 & n4468 ;
  assign n4769 = ( n1630 & n4468 ) | ( n1630 & n4768 ) | ( n4468 & n4768 ) ;
  assign n4770 = n2279 & n4471 ;
  assign n4771 = ( ~n2269 & n4471 ) | ( ~n2269 & n4770 ) | ( n4471 & n4770 ) ;
  assign n4772 = n4769 | n4771 ;
  assign n4773 = n4767 | n4772 ;
  assign n4774 = n4475 | n4773 ;
  assign n4775 = n4773 & n4774 ;
  assign n4776 = ( ~n2343 & n4774 ) | ( ~n2343 & n4775 ) | ( n4774 & n4775 ) ;
  assign n4777 = ~x17 & n4775 ;
  assign n4778 = ~x17 & n4774 ;
  assign n4779 = ( ~n2343 & n4777 ) | ( ~n2343 & n4778 ) | ( n4777 & n4778 ) ;
  assign n4780 = x17 | n4777 ;
  assign n4781 = x17 | n4778 ;
  assign n4782 = ( ~n2343 & n4780 ) | ( ~n2343 & n4781 ) | ( n4780 & n4781 ) ;
  assign n4783 = ( ~n4776 & n4779 ) | ( ~n4776 & n4782 ) | ( n4779 & n4782 ) ;
  assign n4784 = n4766 & n4783 ;
  assign n4785 = n3927 & n3929 ;
  assign n4786 = n3927 | n3929 ;
  assign n4787 = ~n4785 & n4786 ;
  assign n4788 = n1708 & n4468 ;
  assign n4789 = n1793 & n4466 ;
  assign n4790 = ( n1783 & n4466 ) | ( n1783 & n4789 ) | ( n4466 & n4789 ) ;
  assign n4791 = n1634 & n4471 ;
  assign n4792 = ( n1630 & n4471 ) | ( n1630 & n4791 ) | ( n4471 & n4791 ) ;
  assign n4793 = n4790 | n4792 ;
  assign n4794 = n4788 | n4793 ;
  assign n4795 = n4475 | n4794 ;
  assign n4796 = n4794 & n4795 ;
  assign n4797 = ( n1814 & n4795 ) | ( n1814 & n4796 ) | ( n4795 & n4796 ) ;
  assign n4798 = x17 & n4796 ;
  assign n4799 = x17 & n4795 ;
  assign n4800 = ( n1814 & n4798 ) | ( n1814 & n4799 ) | ( n4798 & n4799 ) ;
  assign n4801 = x17 & ~n4798 ;
  assign n4802 = x17 & ~n4799 ;
  assign n4803 = ( ~n1814 & n4801 ) | ( ~n1814 & n4802 ) | ( n4801 & n4802 ) ;
  assign n4804 = ( n4797 & ~n4800 ) | ( n4797 & n4803 ) | ( ~n4800 & n4803 ) ;
  assign n4805 = n4787 & n4804 ;
  assign n4806 = n3923 & n3925 ;
  assign n4807 = n3923 | n3925 ;
  assign n4808 = ~n4806 & n4807 ;
  assign n4809 = ~n523 & n4466 ;
  assign n4810 = n1793 & n4468 ;
  assign n4811 = ( n1783 & n4468 ) | ( n1783 & n4810 ) | ( n4468 & n4810 ) ;
  assign n4812 = n4809 | n4811 ;
  assign n4813 = n1708 & n4471 ;
  assign n4814 = n4812 | n4813 ;
  assign n4815 = n4475 | n4813 ;
  assign n4816 = n4812 | n4815 ;
  assign n4817 = ( ~n1852 & n4814 ) | ( ~n1852 & n4816 ) | ( n4814 & n4816 ) ;
  assign n4818 = ~x17 & n4816 ;
  assign n4819 = ~x17 & n4814 ;
  assign n4820 = ( ~n1852 & n4818 ) | ( ~n1852 & n4819 ) | ( n4818 & n4819 ) ;
  assign n4821 = x17 | n4819 ;
  assign n4822 = x17 | n4818 ;
  assign n4823 = ( ~n1852 & n4821 ) | ( ~n1852 & n4822 ) | ( n4821 & n4822 ) ;
  assign n4824 = ( ~n4817 & n4820 ) | ( ~n4817 & n4823 ) | ( n4820 & n4823 ) ;
  assign n4825 = n4808 & n4824 ;
  assign n4826 = n3919 | n3920 ;
  assign n4827 = n3903 | n4826 ;
  assign n4828 = ~n3922 & n4827 ;
  assign n4829 = ~n523 & n4468 ;
  assign n4830 = n352 & n4466 ;
  assign n4831 = ( ~n339 & n4466 ) | ( ~n339 & n4830 ) | ( n4466 & n4830 ) ;
  assign n4832 = n1793 & n4471 ;
  assign n4833 = ( n1783 & n4471 ) | ( n1783 & n4832 ) | ( n4471 & n4832 ) ;
  assign n4834 = n4831 | n4833 ;
  assign n4835 = n4829 | n4834 ;
  assign n4836 = n4475 | n4835 ;
  assign n4837 = n4835 & n4836 ;
  assign n4838 = ( n1884 & n4836 ) | ( n1884 & n4837 ) | ( n4836 & n4837 ) ;
  assign n4839 = x17 & n4837 ;
  assign n4840 = x17 & n4836 ;
  assign n4841 = ( n1884 & n4839 ) | ( n1884 & n4840 ) | ( n4839 & n4840 ) ;
  assign n4842 = x17 & ~n4839 ;
  assign n4843 = x17 & ~n4840 ;
  assign n4844 = ( ~n1884 & n4842 ) | ( ~n1884 & n4843 ) | ( n4842 & n4843 ) ;
  assign n4845 = ( n4838 & ~n4841 ) | ( n4838 & n4844 ) | ( ~n4841 & n4844 ) ;
  assign n4846 = n4828 & n4845 ;
  assign n4847 = n4828 | n4845 ;
  assign n4848 = ~n4846 & n4847 ;
  assign n4849 = ~n829 & n4466 ;
  assign n4850 = n352 & n4468 ;
  assign n4851 = ( ~n339 & n4468 ) | ( ~n339 & n4850 ) | ( n4468 & n4850 ) ;
  assign n4852 = n4849 | n4851 ;
  assign n4853 = ~n523 & n4471 ;
  assign n4854 = n4475 | n4853 ;
  assign n4855 = n4852 | n4854 ;
  assign n4856 = ~x17 & n4855 ;
  assign n4857 = n4852 | n4853 ;
  assign n4858 = ~x17 & n4857 ;
  assign n4859 = ( ~n1055 & n4856 ) | ( ~n1055 & n4858 ) | ( n4856 & n4858 ) ;
  assign n4860 = x17 & n4855 ;
  assign n4861 = x17 & ~n4860 ;
  assign n4862 = x17 & n4853 ;
  assign n4863 = ( x17 & n4852 ) | ( x17 & n4862 ) | ( n4852 & n4862 ) ;
  assign n4864 = x17 & ~n4863 ;
  assign n4865 = ( n1055 & n4861 ) | ( n1055 & n4864 ) | ( n4861 & n4864 ) ;
  assign n4866 = n4859 | n4865 ;
  assign n4867 = n3896 | n3898 ;
  assign n4868 = x20 & ~n3896 ;
  assign n4869 = ( n3879 & n4867 ) | ( n3879 & ~n4868 ) | ( n4867 & ~n4868 ) ;
  assign n4870 = ~n3901 & n4869 ;
  assign n4871 = n4866 & n4870 ;
  assign n4872 = x20 | n3893 ;
  assign n4873 = ( ~n3886 & n3893 ) | ( ~n3886 & n4872 ) | ( n3893 & n4872 ) ;
  assign n4874 = n3887 | n4873 ;
  assign n4875 = ~n3896 & n4874 ;
  assign n4876 = ~n829 & n4468 ;
  assign n4877 = n352 & n4471 ;
  assign n4878 = ( ~n339 & n4471 ) | ( ~n339 & n4877 ) | ( n4471 & n4877 ) ;
  assign n4879 = n4876 | n4878 ;
  assign n4880 = n692 & n4466 ;
  assign n4881 = ( n674 & n4466 ) | ( n674 & n4880 ) | ( n4466 & n4880 ) ;
  assign n4882 = n4879 | n4881 ;
  assign n4883 = n4475 | n4881 ;
  assign n4884 = n4879 | n4883 ;
  assign n4885 = ( ~n1209 & n4882 ) | ( ~n1209 & n4884 ) | ( n4882 & n4884 ) ;
  assign n4886 = ~x17 & n4884 ;
  assign n4887 = ~x17 & n4882 ;
  assign n4888 = ( ~n1209 & n4886 ) | ( ~n1209 & n4887 ) | ( n4886 & n4887 ) ;
  assign n4889 = x17 | n4887 ;
  assign n4890 = x17 | n4886 ;
  assign n4891 = ( ~n1209 & n4889 ) | ( ~n1209 & n4890 ) | ( n4889 & n4890 ) ;
  assign n4892 = ( ~n4885 & n4888 ) | ( ~n4885 & n4891 ) | ( n4888 & n4891 ) ;
  assign n4893 = n4875 & n4892 ;
  assign n4894 = ( ~n1027 & n3889 ) | ( ~n1027 & n3891 ) | ( n3889 & n3891 ) ;
  assign n4895 = ~n922 & n4468 ;
  assign n4896 = n1042 & n4466 ;
  assign n4897 = ( ~n1027 & n4466 ) | ( ~n1027 & n4896 ) | ( n4466 & n4896 ) ;
  assign n4898 = n4895 | n4897 ;
  assign n4899 = n692 & n4471 ;
  assign n4900 = ( n674 & n4471 ) | ( n674 & n4899 ) | ( n4471 & n4899 ) ;
  assign n4901 = n4898 | n4900 ;
  assign n4902 = ( n1538 & n4475 ) | ( n1538 & n4901 ) | ( n4475 & n4901 ) ;
  assign n4903 = ( x17 & ~n4901 ) | ( x17 & n4902 ) | ( ~n4901 & n4902 ) ;
  assign n4904 = ~n4902 & n4903 ;
  assign n4905 = ~n922 & n4471 ;
  assign n4906 = n1042 & n4468 ;
  assign n4907 = ( ~n1027 & n4468 ) | ( ~n1027 & n4906 ) | ( n4468 & n4906 ) ;
  assign n4908 = n4905 | n4907 ;
  assign n4909 = n4475 | n4907 ;
  assign n4910 = n4905 | n4909 ;
  assign n4911 = ( n1946 & n4908 ) | ( n1946 & n4910 ) | ( n4908 & n4910 ) ;
  assign n4912 = ~x17 & n4911 ;
  assign n4913 = n139 & n4461 ;
  assign n4914 = ( n1041 & n4461 ) | ( n1041 & n4913 ) | ( n4461 & n4913 ) ;
  assign n4915 = x17 & ~n4914 ;
  assign n4916 = n4461 | n4913 ;
  assign n4917 = x17 & ~n4916 ;
  assign n4918 = ( n1027 & n4915 ) | ( n1027 & n4917 ) | ( n4915 & n4917 ) ;
  assign n4919 = x17 & n4918 ;
  assign n4920 = ~n4911 & n4919 ;
  assign n4921 = ( n4912 & n4918 ) | ( n4912 & n4920 ) | ( n4918 & n4920 ) ;
  assign n4922 = x17 | n4901 ;
  assign n4923 = n4902 | n4922 ;
  assign n4924 = n4921 & n4923 ;
  assign n4925 = ~x17 & n4921 ;
  assign n4926 = ( n4904 & n4924 ) | ( n4904 & n4925 ) | ( n4924 & n4925 ) ;
  assign n4927 = n4894 & n4926 ;
  assign n4928 = n4926 & ~n4927 ;
  assign n4929 = ~n829 & n4471 ;
  assign n4930 = ~n922 & n4466 ;
  assign n4931 = n4929 | n4930 ;
  assign n4932 = n692 & n4468 ;
  assign n4933 = ( n674 & n4468 ) | ( n674 & n4932 ) | ( n4468 & n4932 ) ;
  assign n4934 = n4931 | n4933 ;
  assign n4935 = n4475 | n4933 ;
  assign n4936 = n4931 | n4935 ;
  assign n4937 = ( n1554 & n4934 ) | ( n1554 & n4936 ) | ( n4934 & n4936 ) ;
  assign n4938 = x17 & n4936 ;
  assign n4939 = x17 & n4934 ;
  assign n4940 = ( n1554 & n4938 ) | ( n1554 & n4939 ) | ( n4938 & n4939 ) ;
  assign n4941 = x17 & ~n4939 ;
  assign n4942 = x17 & ~n4938 ;
  assign n4943 = ( ~n1554 & n4941 ) | ( ~n1554 & n4942 ) | ( n4941 & n4942 ) ;
  assign n4944 = ( n4937 & ~n4940 ) | ( n4937 & n4943 ) | ( ~n4940 & n4943 ) ;
  assign n4945 = n4894 & ~n4926 ;
  assign n4946 = n4944 & n4945 ;
  assign n4947 = ( n4928 & n4944 ) | ( n4928 & n4946 ) | ( n4944 & n4946 ) ;
  assign n4948 = n4927 | n4947 ;
  assign n4949 = n4875 | n4892 ;
  assign n4950 = ~n4893 & n4949 ;
  assign n4951 = n4893 | n4950 ;
  assign n4952 = ( n4893 & n4948 ) | ( n4893 & n4951 ) | ( n4948 & n4951 ) ;
  assign n4953 = n4866 | n4870 ;
  assign n4954 = ~n4871 & n4953 ;
  assign n4955 = n4871 | n4954 ;
  assign n4956 = ( n4871 & n4952 ) | ( n4871 & n4955 ) | ( n4952 & n4955 ) ;
  assign n4957 = n4848 & n4956 ;
  assign n4958 = n4846 | n4957 ;
  assign n4959 = ~n4808 & n4824 ;
  assign n4960 = ( n4808 & ~n4825 ) | ( n4808 & n4959 ) | ( ~n4825 & n4959 ) ;
  assign n4961 = n4958 & n4960 ;
  assign n4962 = n4825 | n4961 ;
  assign n4963 = n4787 & ~n4805 ;
  assign n4964 = ~n4787 & n4804 ;
  assign n4965 = n4963 | n4964 ;
  assign n4966 = n4962 & n4965 ;
  assign n4967 = n4805 | n4966 ;
  assign n4968 = n4766 & ~n4784 ;
  assign n4969 = ~n4766 & n4783 ;
  assign n4970 = n4968 | n4969 ;
  assign n4971 = n4784 | n4970 ;
  assign n4972 = ( n4784 & n4967 ) | ( n4784 & n4971 ) | ( n4967 & n4971 ) ;
  assign n4973 = n4745 | n4763 ;
  assign n4974 = ~n4764 & n4973 ;
  assign n4975 = n4764 | n4974 ;
  assign n4976 = ( n4764 & n4972 ) | ( n4764 & n4975 ) | ( n4972 & n4975 ) ;
  assign n4977 = n4743 & n4976 ;
  assign n4978 = n4741 | n4977 ;
  assign n4979 = n4718 | n4978 ;
  assign n4980 = ( n4718 & n4722 ) | ( n4718 & n4979 ) | ( n4722 & n4979 ) ;
  assign n4981 = ~n4676 & n4694 ;
  assign n4982 = ( n4676 & ~n4695 ) | ( n4676 & n4981 ) | ( ~n4695 & n4981 ) ;
  assign n4983 = n4695 | n4982 ;
  assign n4984 = ( n4695 & n4980 ) | ( n4695 & n4983 ) | ( n4980 & n4983 ) ;
  assign n4985 = n4673 & n4984 ;
  assign n4986 = n4666 | n4985 ;
  assign n4987 = ( n4669 & n4670 ) | ( n4669 & n4986 ) | ( n4670 & n4986 ) ;
  assign n4988 = n4619 | n4987 ;
  assign n4989 = ( n4619 & n4623 ) | ( n4619 & n4988 ) | ( n4623 & n4988 ) ;
  assign n4990 = n4593 | n4989 ;
  assign n4991 = ( n4593 & ~n4596 ) | ( n4593 & n4990 ) | ( ~n4596 & n4990 ) ;
  assign n4992 = n4569 | n4991 ;
  assign n4993 = ( n4569 & ~n4573 ) | ( n4569 & n4992 ) | ( ~n4573 & n4992 ) ;
  assign n4994 = n4544 | n4993 ;
  assign n4995 = ( n4544 & n4547 ) | ( n4544 & n4994 ) | ( n4547 & n4994 ) ;
  assign n3965 = n3588 | n3964 ;
  assign n2591 = n2587 | n2590 ;
  assign n2592 = ( n2557 & n2587 ) | ( n2557 & n2591 ) | ( n2587 & n2591 ) ;
  assign n1569 = n1322 | n1568 ;
  assign n1570 = ( n1322 & n1330 ) | ( n1322 & n1569 ) | ( n1330 & n1569 ) ;
  assign n1058 = ~n523 & n1057 ;
  assign n1061 = ~n829 & n1060 ;
  assign n1066 = n352 & n1065 ;
  assign n1067 = ( ~n339 & n1065 ) | ( ~n339 & n1066 ) | ( n1065 & n1066 ) ;
  assign n1068 = n1062 | n1067 ;
  assign n1069 = n1061 | n1068 ;
  assign n1070 = n1058 | n1069 ;
  assign n1071 = n1061 | n1067 ;
  assign n1072 = n1058 | n1071 ;
  assign n1073 = ( ~n1055 & n1070 ) | ( ~n1055 & n1072 ) | ( n1070 & n1072 ) ;
  assign n1078 = n288 | n434 ;
  assign n1079 = n325 | n1078 ;
  assign n1081 = n104 | n594 ;
  assign n1082 = n1080 | n1081 ;
  assign n1083 = n1079 | n1082 ;
  assign n1084 = n1077 | n1083 ;
  assign n1085 = n90 | n1084 ;
  assign n1089 = n183 | n527 ;
  assign n1090 = n303 | n1089 ;
  assign n1091 = n1088 | n1090 ;
  assign n1092 = n240 | n305 ;
  assign n1093 = n413 | n1092 ;
  assign n1094 = n1091 | n1093 ;
  assign n1095 = n406 | n602 ;
  assign n1096 = n418 | n1095 ;
  assign n1098 = n110 | n114 ;
  assign n1099 = n1097 | n1098 ;
  assign n1100 = n1096 | n1099 ;
  assign n1101 = n192 | n343 ;
  assign n1102 = n143 & ~n332 ;
  assign n1103 = ~n1101 & n1102 ;
  assign n1104 = ~n1100 & n1103 ;
  assign n1105 = ~n1094 & n1104 ;
  assign n1106 = ~n1085 & n1105 ;
  assign n1107 = n246 | n258 ;
  assign n1108 = n269 | n341 ;
  assign n1109 = n1107 | n1108 ;
  assign n1110 = n447 | n513 ;
  assign n1111 = n895 | n1110 ;
  assign n1112 = n1109 | n1111 ;
  assign n1113 = n1106 & ~n1112 ;
  assign n1117 = n1115 | n1116 ;
  assign n1119 = n324 | n608 ;
  assign n1120 = n1118 | n1119 ;
  assign n1121 = n152 | n171 ;
  assign n1122 = n1120 | n1121 ;
  assign n1123 = n1117 | n1122 ;
  assign n1124 = n154 | n568 ;
  assign n1125 = n581 | n1124 ;
  assign n1128 = n1126 | n1127 ;
  assign n1129 = n1125 | n1128 ;
  assign n1130 = n383 | n456 ;
  assign n1131 = n1129 | n1130 ;
  assign n1132 = n1123 | n1131 ;
  assign n1133 = n225 | n437 ;
  assign n1144 = n1133 | n1143 ;
  assign n1145 = n1132 | n1144 ;
  assign n1147 = n824 | n1146 ;
  assign n1148 = n254 | n1147 ;
  assign n1152 = n1149 | n1151 ;
  assign n1153 = n1148 | n1152 ;
  assign n1154 = n170 | n321 ;
  assign n1155 = n979 | n1154 ;
  assign n1156 = n302 | n1155 ;
  assign n1157 = n384 | n643 ;
  assign n1158 = n711 | n1157 ;
  assign n1159 = n99 | n448 ;
  assign n1160 = n1158 | n1159 ;
  assign n1161 = n1156 | n1160 ;
  assign n1162 = n1153 | n1161 ;
  assign n1166 = n654 | n689 ;
  assign n1167 = n1165 | n1166 ;
  assign n1168 = n1164 | n1167 ;
  assign n1169 = n278 | n762 ;
  assign n1170 = n196 | n1169 ;
  assign n1171 = n405 | n497 ;
  assign n1173 = n590 | n1172 ;
  assign n1174 = n1171 | n1173 ;
  assign n1175 = n1170 | n1174 ;
  assign n1176 = n1168 | n1175 ;
  assign n1177 = n274 | n966 ;
  assign n1178 = n480 | n503 ;
  assign n1179 = n296 | n1178 ;
  assign n1180 = n1177 | n1179 ;
  assign n1181 = n465 | n725 ;
  assign n1182 = n39 | n59 ;
  assign n1183 = n1181 | n1182 ;
  assign n1184 = n363 | n468 ;
  assign n1185 = n1183 | n1184 ;
  assign n1186 = n1180 | n1185 ;
  assign n1187 = n1176 | n1186 ;
  assign n1188 = n1162 | n1187 ;
  assign n1189 = n1145 | n1188 ;
  assign n1190 = n1113 & ~n1189 ;
  assign n1191 = n291 | n451 ;
  assign n1192 = n133 | n1191 ;
  assign n1194 = n566 | n1193 ;
  assign n1195 = n1192 | n1194 ;
  assign n1196 = n1190 & ~n1195 ;
  assign n1197 = n1058 & ~n1196 ;
  assign n1198 = ( n1069 & ~n1196 ) | ( n1069 & n1197 ) | ( ~n1196 & n1197 ) ;
  assign n1199 = ( n1071 & ~n1196 ) | ( n1071 & n1197 ) | ( ~n1196 & n1197 ) ;
  assign n1200 = ( ~n1055 & n1198 ) | ( ~n1055 & n1199 ) | ( n1198 & n1199 ) ;
  assign n1201 = n1073 & ~n1200 ;
  assign n1202 = n1072 | n1196 ;
  assign n1203 = n1070 | n1196 ;
  assign n1204 = ( ~n1055 & n1202 ) | ( ~n1055 & n1203 ) | ( n1202 & n1203 ) ;
  assign n1205 = ~n1201 & n1204 ;
  assign n1571 = ~n1205 & n1570 ;
  assign n1572 = n1570 & ~n1571 ;
  assign n1573 = n1205 | n1571 ;
  assign n1574 = ~n1572 & n1573 ;
  assign n1824 = n1708 & n1823 ;
  assign n1827 = n1793 & n1826 ;
  assign n1828 = ( n1783 & n1826 ) | ( n1783 & n1827 ) | ( n1826 & n1827 ) ;
  assign n1830 = n1634 & n1829 ;
  assign n1831 = ( n1630 & n1829 ) | ( n1630 & n1830 ) | ( n1829 & n1830 ) ;
  assign n1832 = n1828 | n1831 ;
  assign n1833 = n1824 | n1832 ;
  assign n1834 = n1821 | n1833 ;
  assign n1835 = ( n1814 & n1833 ) | ( n1814 & n1834 ) | ( n1833 & n1834 ) ;
  assign n1836 = x29 & n1834 ;
  assign n1837 = x29 & n1833 ;
  assign n1838 = ( n1814 & n1836 ) | ( n1814 & n1837 ) | ( n1836 & n1837 ) ;
  assign n1839 = x29 & ~n1836 ;
  assign n1840 = x29 & ~n1837 ;
  assign n1841 = ( ~n1814 & n1839 ) | ( ~n1814 & n1840 ) | ( n1839 & n1840 ) ;
  assign n1842 = ( n1835 & ~n1838 ) | ( n1835 & n1841 ) | ( ~n1838 & n1841 ) ;
  assign n1843 = ~n1574 & n1842 ;
  assign n1844 = n1574 | n1843 ;
  assign n1845 = n1574 & n1842 ;
  assign n1846 = n1844 & ~n1845 ;
  assign n2019 = n1871 | n2018 ;
  assign n2020 = ~n1846 & n2019 ;
  assign n2021 = n1846 & ~n2019 ;
  assign n2022 = n2020 | n2021 ;
  assign n2309 = n2090 & n2308 ;
  assign n2310 = ( ~n2082 & n2308 ) | ( ~n2082 & n2309 ) | ( n2308 & n2309 ) ;
  assign n2313 = n2279 & n2312 ;
  assign n2314 = ( ~n2269 & n2312 ) | ( ~n2269 & n2313 ) | ( n2312 & n2313 ) ;
  assign n2316 = n2199 & n2315 ;
  assign n2317 = ( ~n2185 & n2315 ) | ( ~n2185 & n2316 ) | ( n2315 & n2316 ) ;
  assign n2318 = n2314 | n2317 ;
  assign n2319 = n2310 | n2318 ;
  assign n2320 = n2306 | n2319 ;
  assign n2326 = ( n2319 & n2320 ) | ( n2319 & ~n2325 ) | ( n2320 & ~n2325 ) ;
  assign n2327 = n2319 & n2320 ;
  assign n2328 = ( ~n2299 & n2326 ) | ( ~n2299 & n2327 ) | ( n2326 & n2327 ) ;
  assign n2329 = ~x26 & n2328 ;
  assign n2330 = x26 | n2328 ;
  assign n2331 = ( ~n2328 & n2329 ) | ( ~n2328 & n2330 ) | ( n2329 & n2330 ) ;
  assign n2332 = ~n2022 & n2331 ;
  assign n2333 = n2022 | n2332 ;
  assign n2334 = n2022 & n2331 ;
  assign n2335 = n2333 & ~n2334 ;
  assign n2593 = ~n2335 & n2592 ;
  assign n2594 = n2592 & ~n2593 ;
  assign n2595 = n2335 | n2593 ;
  assign n2596 = ~n2594 & n2595 ;
  assign n2926 = n2691 & n2925 ;
  assign n2927 = ( n2678 & n2925 ) | ( n2678 & n2926 ) | ( n2925 & n2926 ) ;
  assign n2929 = n2701 & n2928 ;
  assign n2930 = ( ~n2784 & n2928 ) | ( ~n2784 & n2929 ) | ( n2928 & n2929 ) ;
  assign n2931 = n2927 | n2930 ;
  assign n2933 = n2893 & n2932 ;
  assign n2934 = ( ~n2886 & n2932 ) | ( ~n2886 & n2933 ) | ( n2932 & n2933 ) ;
  assign n2935 = n2931 | n2934 ;
  assign n2937 = n2935 | n2936 ;
  assign n2938 = ( ~n2914 & n2935 ) | ( ~n2914 & n2937 ) | ( n2935 & n2937 ) ;
  assign n2939 = ~x23 & n2937 ;
  assign n2940 = ~x23 & n2935 ;
  assign n2941 = ( ~n2914 & n2939 ) | ( ~n2914 & n2940 ) | ( n2939 & n2940 ) ;
  assign n2942 = x23 | n2939 ;
  assign n2943 = x23 | n2940 ;
  assign n2944 = ( ~n2914 & n2942 ) | ( ~n2914 & n2943 ) | ( n2942 & n2943 ) ;
  assign n2945 = ( ~n2938 & n2941 ) | ( ~n2938 & n2944 ) | ( n2941 & n2944 ) ;
  assign n2946 = ~n2596 & n2945 ;
  assign n2947 = n2596 | n2946 ;
  assign n2948 = n2596 & n2945 ;
  assign n2949 = n2947 & ~n2948 ;
  assign n3271 = n2979 | n3270 ;
  assign n3272 = ( n2979 & n3268 ) | ( n2979 & n3271 ) | ( n3268 & n3271 ) ;
  assign n3273 = ~n2949 & n3272 ;
  assign n3274 = n2949 & ~n3272 ;
  assign n3275 = n3273 | n3274 ;
  assign n3542 = n3386 & n3541 ;
  assign n3545 = n3507 & n3544 ;
  assign n3546 = ( n3483 & n3544 ) | ( n3483 & n3545 ) | ( n3544 & n3545 ) ;
  assign n3548 = n3439 & n3547 ;
  assign n3549 = ( ~n3420 & n3547 ) | ( ~n3420 & n3548 ) | ( n3547 & n3548 ) ;
  assign n3550 = n3546 | n3549 ;
  assign n3551 = n3542 | n3550 ;
  assign n3552 = n3537 | n3551 ;
  assign n3553 = n3551 & n3552 ;
  assign n3554 = ( ~n3530 & n3552 ) | ( ~n3530 & n3553 ) | ( n3552 & n3553 ) ;
  assign n3555 = ~x20 & n3553 ;
  assign n3556 = ~x20 & n3552 ;
  assign n3557 = ( ~n3530 & n3555 ) | ( ~n3530 & n3556 ) | ( n3555 & n3556 ) ;
  assign n3558 = x20 | n3555 ;
  assign n3559 = x20 | n3556 ;
  assign n3560 = ( ~n3530 & n3558 ) | ( ~n3530 & n3559 ) | ( n3558 & n3559 ) ;
  assign n3561 = ( ~n3554 & n3557 ) | ( ~n3554 & n3560 ) | ( n3557 & n3560 ) ;
  assign n3562 = ~n3275 & n3561 ;
  assign n3966 = n3275 | n3562 ;
  assign n3967 = n3275 & n3561 ;
  assign n3968 = n3966 & ~n3967 ;
  assign n4492 = n3965 | n3968 ;
  assign n4493 = n3965 & n3968 ;
  assign n4494 = n4492 & ~n4493 ;
  assign n4327 = n313 | n497 ;
  assign n4328 = n347 | n4327 ;
  assign n4329 = n175 | n607 ;
  assign n4330 = n1307 | n4329 ;
  assign n4331 = n4328 | n4330 ;
  assign n4332 = n717 | n4331 ;
  assign n4333 = n682 | n728 ;
  assign n4334 = n332 | n501 ;
  assign n4335 = n695 | n4334 ;
  assign n4336 = n4333 | n4335 ;
  assign n4337 = n4332 | n4336 ;
  assign n4338 = n4326 | n4337 ;
  assign n4339 = n4322 | n4338 ;
  assign n4340 = n363 | n459 ;
  assign n4341 = n240 | n245 ;
  assign n4342 = n1286 | n4341 ;
  assign n4343 = n4340 | n4342 ;
  assign n4344 = n289 | n667 ;
  assign n4345 = n4184 | n4344 ;
  assign n4346 = n4343 | n4345 ;
  assign n4347 = n292 | n412 ;
  assign n4348 = n213 | n638 ;
  assign n4349 = n4347 | n4348 ;
  assign n4350 = n402 | n4349 ;
  assign n4351 = n887 | n4350 ;
  assign n4352 = n4346 | n4351 ;
  assign n4353 = n297 | n491 ;
  assign n4354 = n280 | n4353 ;
  assign n4355 = ( n720 & ~n885 ) | ( n720 & n4354 ) | ( ~n885 & n4354 ) ;
  assign n4356 = n159 | n885 ;
  assign n4357 = n4355 | n4356 ;
  assign n4358 = n4352 | n4357 ;
  assign n4359 = n382 | n4358 ;
  assign n4360 = n4339 | n4359 ;
  assign n4361 = n262 | n331 ;
  assign n4362 = n395 | n469 ;
  assign n4363 = n4361 | n4362 ;
  assign n4364 = n312 | n4363 ;
  assign n3984 = n318 | n591 ;
  assign n4365 = n2256 | n3984 ;
  assign n4366 = n4364 | n4365 ;
  assign n4367 = n435 | n623 ;
  assign n4368 = n1473 | n4367 ;
  assign n4369 = n283 | n574 ;
  assign n4370 = n364 | n4369 ;
  assign n4371 = n4368 | n4370 ;
  assign n4372 = n205 | n388 ;
  assign n4373 = n447 | n643 ;
  assign n4374 = n4372 | n4373 ;
  assign n4375 = n4371 | n4374 ;
  assign n4376 = n4366 | n4375 ;
  assign n4377 = n1215 | n1349 ;
  assign n4378 = n1218 | n4377 ;
  assign n4379 = n679 | n4378 ;
  assign n4380 = n4376 | n4379 ;
  assign n4381 = n151 | n675 ;
  assign n4382 = n126 | n4381 ;
  assign n4249 = n123 | n225 ;
  assign n4383 = n67 | n384 ;
  assign n4384 = n4249 | n4383 ;
  assign n4385 = n141 | n223 ;
  assign n4386 = n305 | n4385 ;
  assign n4387 = n4384 | n4386 ;
  assign n4388 = n4382 | n4387 ;
  assign n4389 = n256 | n4388 ;
  assign n4390 = n4380 | n4389 ;
  assign n4391 = n284 | n317 ;
  assign n4392 = n702 | n4391 ;
  assign n4393 = n190 | n624 ;
  assign n4394 = n4392 | n4393 ;
  assign n4395 = n4390 | n4394 ;
  assign n4396 = n4360 | n4395 ;
  assign n4430 = n4396 & ~n4429 ;
  assign n4431 = ~n4396 & n4429 ;
  assign n4432 = n4430 | n4431 ;
  assign n4442 = n4436 | n4441 ;
  assign n4495 = ~n4432 & n4442 ;
  assign n4447 = n4436 | n4446 ;
  assign n4496 = ~n4432 & n4447 ;
  assign n4497 = ( ~n3525 & n4495 ) | ( ~n3525 & n4496 ) | ( n4495 & n4496 ) ;
  assign n4498 = n4432 & ~n4442 ;
  assign n4499 = n4432 & ~n4447 ;
  assign n4500 = ( n3525 & n4498 ) | ( n3525 & n4499 ) | ( n4498 & n4499 ) ;
  assign n4501 = n4497 | n4500 ;
  assign n4502 = ~n4429 & n4468 ;
  assign n4503 = n4466 | n4468 ;
  assign n4504 = ( ~n4429 & n4466 ) | ( ~n4429 & n4503 ) | ( n4466 & n4503 ) ;
  assign n4505 = ( n4206 & n4502 ) | ( n4206 & n4504 ) | ( n4502 & n4504 ) ;
  assign n4506 = n4396 & n4471 ;
  assign n4507 = n4505 | n4506 ;
  assign n4508 = n4475 | n4506 ;
  assign n4509 = n4505 | n4508 ;
  assign n4510 = ( ~n4501 & n4507 ) | ( ~n4501 & n4509 ) | ( n4507 & n4509 ) ;
  assign n4511 = ~x17 & n4509 ;
  assign n4512 = ~x17 & n4507 ;
  assign n4513 = ( ~n4501 & n4511 ) | ( ~n4501 & n4512 ) | ( n4511 & n4512 ) ;
  assign n4514 = x17 | n4512 ;
  assign n4515 = x17 | n4511 ;
  assign n4516 = ( ~n4501 & n4514 ) | ( ~n4501 & n4515 ) | ( n4514 & n4515 ) ;
  assign n4517 = ( ~n4510 & n4513 ) | ( ~n4510 & n4516 ) | ( n4513 & n4516 ) ;
  assign n4518 = ~n4494 & n4517 ;
  assign n4996 = n4494 & ~n4517 ;
  assign n4997 = n4518 | n4996 ;
  assign n5256 = n4995 & ~n4997 ;
  assign n5257 = ~n4995 & n4997 ;
  assign n5258 = n5256 | n5257 ;
  assign n5123 = n364 | n370 ;
  assign n5124 = n2135 | n5123 ;
  assign n5125 = n99 | n387 ;
  assign n5126 = n184 | n5125 ;
  assign n5127 = n5124 | n5126 ;
  assign n5128 = n577 | n5127 ;
  assign n5129 = n71 | n4319 ;
  assign n5130 = n175 | n450 ;
  assign n5131 = n702 | n5130 ;
  assign n5132 = n513 | n5131 ;
  assign n5133 = n128 | n348 ;
  assign n5134 = n2204 | n5133 ;
  assign n5135 = n5132 | n5134 ;
  assign n5136 = n5129 | n5135 ;
  assign n5137 = n141 | n483 ;
  assign n5138 = n118 | n487 ;
  assign n5139 = n5137 | n5138 ;
  assign n5140 = n2100 | n5139 ;
  assign n5141 = n245 | n318 ;
  assign n5142 = n1163 | n5141 ;
  assign n5143 = n5140 | n5142 ;
  assign n5144 = n170 | n331 ;
  assign n5145 = n247 | n510 ;
  assign n5146 = n5144 | n5145 ;
  assign n5147 = n402 | n5146 ;
  assign n5148 = n131 | n273 ;
  assign n5149 = n5147 | n5148 ;
  assign n5150 = n5143 | n5149 ;
  assign n5151 = n5136 | n5150 ;
  assign n5152 = n5128 | n5151 ;
  assign n5153 = n300 | n1384 ;
  assign n5028 = n77 | n317 ;
  assign n5029 = n2803 | n5028 ;
  assign n5030 = n451 | n5029 ;
  assign n5154 = n476 | n2156 ;
  assign n5155 = n5030 | n5154 ;
  assign n5156 = n5153 | n5155 ;
  assign n5157 = n92 | n183 ;
  assign n5158 = n489 | n5157 ;
  assign n5159 = n189 | n1695 ;
  assign n5160 = n5158 | n5159 ;
  assign n5161 = n79 | n341 ;
  assign n5162 = n354 | n413 ;
  assign n5163 = n5161 | n5162 ;
  assign n5164 = n5160 | n5163 ;
  assign n5165 = n256 | n888 ;
  assign n5166 = n504 | n5165 ;
  assign n5167 = n5164 | n5166 ;
  assign n5168 = n5156 | n5167 ;
  assign n5169 = n264 | n1016 ;
  assign n5170 = n602 | n5169 ;
  assign n5171 = n775 | n4249 ;
  assign n5172 = n257 | n5171 ;
  assign n5173 = n5170 | n5172 ;
  assign n5174 = n735 | n5173 ;
  assign n5175 = ( n133 & n160 ) | ( n133 & ~n376 ) | ( n160 & ~n376 ) ;
  assign n5176 = n376 | n5175 ;
  assign n5177 = n5174 | n5176 ;
  assign n5178 = n5168 | n5177 ;
  assign n5179 = n5152 | n5178 ;
  assign n5180 = n206 | n333 ;
  assign n5181 = n46 | n591 ;
  assign n5182 = n465 | n694 ;
  assign n5183 = n5181 | n5182 ;
  assign n5184 = n551 | n2147 ;
  assign n5185 = n5183 | n5184 ;
  assign n5186 = n1523 | n1607 ;
  assign n5187 = n406 | n5186 ;
  assign n5188 = n5185 | n5187 ;
  assign n5189 = n441 | n841 ;
  assign n5190 = n239 | n5189 ;
  assign n5191 = n5188 | n5190 ;
  assign n5192 = n5180 | n5191 ;
  assign n5193 = n5179 | n5192 ;
  assign n5003 = n435 | n607 ;
  assign n5004 = n354 | n5003 ;
  assign n5005 = n53 | n457 ;
  assign n5006 = n344 | n5005 ;
  assign n5007 = n1605 | n5006 ;
  assign n5008 = n701 | n5007 ;
  assign n5009 = n3494 | n5008 ;
  assign n5010 = n46 | n138 ;
  assign n5011 = n239 | n5010 ;
  assign n5012 = n441 | n3313 ;
  assign n5013 = n5011 | n5012 ;
  assign n5014 = n295 | n381 ;
  assign n5015 = n1220 | n5014 ;
  assign n5016 = n155 | n5015 ;
  assign n5017 = n5013 | n5016 ;
  assign n5018 = n2053 | n5017 ;
  assign n5019 = n274 | n297 ;
  assign n5020 = n294 | n5019 ;
  assign n5021 = n820 | n1404 ;
  assign n5022 = n644 | n5021 ;
  assign n5023 = n5020 | n5022 ;
  assign n5024 = n5018 | n5023 ;
  assign n5025 = n5009 | n5024 ;
  assign n5026 = n5004 | n5025 ;
  assign n5027 = n773 | n788 ;
  assign n5031 = n3388 | n5030 ;
  assign n5032 = n774 | n5031 ;
  assign n5033 = n732 & ~n4419 ;
  assign n5034 = ~n5032 & n5033 ;
  assign n5035 = ~n636 & n5034 ;
  assign n5036 = ~n5027 & n5035 ;
  assign n5037 = ~n5026 & n5036 ;
  assign n5109 = n88 | n178 ;
  assign n5110 = n134 | n222 ;
  assign n5111 = n5109 | n5110 ;
  assign n5112 = n71 | n489 ;
  assign n5113 = n302 | n5112 ;
  assign n5114 = n5111 | n5113 ;
  assign n5115 = n254 | n363 ;
  assign n5116 = n676 | n5115 ;
  assign n5117 = n5114 | n5116 ;
  assign n5199 = n5037 & ~n5117 ;
  assign n5200 = n5193 & ~n5199 ;
  assign n5201 = ~n5193 & n5199 ;
  assign n5202 = n5200 | n5201 ;
  assign n4245 = n255 | n514 ;
  assign n4246 = n269 | n762 ;
  assign n4247 = n203 | n4246 ;
  assign n4248 = n1464 | n4247 ;
  assign n4250 = n2696 | n4249 ;
  assign n4251 = n412 | n480 ;
  assign n4252 = n458 | n4251 ;
  assign n4253 = n4250 | n4252 ;
  assign n4254 = ( ~n2676 & n4248 ) | ( ~n2676 & n4253 ) | ( n4248 & n4253 ) ;
  assign n4255 = n561 | n2676 ;
  assign n4256 = n4254 | n4255 ;
  assign n4259 = n152 | n979 ;
  assign n4260 = n4258 | n4259 ;
  assign n4261 = n226 | n456 ;
  assign n4262 = n310 | n447 ;
  assign n4263 = n4261 | n4262 ;
  assign n4264 = n4260 | n4263 ;
  assign n4265 = n317 | n388 ;
  assign n4266 = n133 | n4265 ;
  assign n4267 = n279 | n779 ;
  assign n4268 = n4266 | n4267 ;
  assign n4269 = n1521 | n4268 ;
  assign n4270 = n4264 | n4269 ;
  assign n4271 = n406 | n631 ;
  assign n4272 = n952 | n4271 ;
  assign n4273 = n272 | n306 ;
  assign n4274 = n155 | n4273 ;
  assign n4275 = n4272 | n4274 ;
  assign n4276 = n1304 | n1404 ;
  assign n4277 = n703 | n3467 ;
  assign n4278 = n682 | n4277 ;
  assign n4279 = n4276 | n4278 ;
  assign n4280 = n4275 | n4279 ;
  assign n4281 = n4270 | n4280 ;
  assign n4282 = n886 | n4281 ;
  assign n4283 = n2743 | n3282 ;
  assign n4284 = n450 | n735 ;
  assign n4285 = n666 | n4284 ;
  assign n4286 = n4283 | n4285 ;
  assign n4287 = n142 | n4286 ;
  assign n4288 = n222 | n938 ;
  assign n4289 = n1124 | n4288 ;
  assign n4290 = n370 | n435 ;
  assign n4291 = n349 | n4290 ;
  assign n4292 = n4289 | n4291 ;
  assign n4294 = n234 | n254 ;
  assign n4295 = n374 | n4294 ;
  assign n4296 = n4293 | n4295 ;
  assign n4297 = n4292 | n4296 ;
  assign n4298 = n4287 | n4297 ;
  assign n4299 = n264 | n387 ;
  assign n4300 = n83 | n4299 ;
  assign n4301 = n4298 | n4300 ;
  assign n4302 = n4282 | n4301 ;
  assign n4303 = n4256 | n4302 ;
  assign n4304 = n4245 | n4303 ;
  assign n5194 = n4304 & n5193 ;
  assign n4397 = n4304 & n4396 ;
  assign n4398 = n4304 | n4396 ;
  assign n4399 = ~n4397 & n4398 ;
  assign n5207 = n4397 | n4430 ;
  assign n5208 = ( n4397 & n4399 ) | ( n4397 & n5207 ) | ( n4399 & n5207 ) ;
  assign n5195 = n4304 | n5193 ;
  assign n5196 = ~n5194 & n5195 ;
  assign n5209 = n5194 | n5196 ;
  assign n5210 = ( n5194 & n5208 ) | ( n5194 & n5209 ) | ( n5208 & n5209 ) ;
  assign n5259 = ~n5202 & n5210 ;
  assign n4433 = ~n4430 & n4432 ;
  assign n4434 = n4399 & ~n4433 ;
  assign n5197 = n4397 & n5196 ;
  assign n5198 = ( n4434 & n5196 ) | ( n4434 & n5197 ) | ( n5196 & n5197 ) ;
  assign n5203 = n5194 & ~n5202 ;
  assign n5260 = ( n5198 & ~n5202 ) | ( n5198 & n5203 ) | ( ~n5202 & n5203 ) ;
  assign n5261 = ( n4442 & n5259 ) | ( n4442 & n5260 ) | ( n5259 & n5260 ) ;
  assign n5262 = ( n4447 & n5259 ) | ( n4447 & n5260 ) | ( n5259 & n5260 ) ;
  assign n5263 = ( ~n3525 & n5261 ) | ( ~n3525 & n5262 ) | ( n5261 & n5262 ) ;
  assign n5264 = n5194 | n5198 ;
  assign n5265 = ( n4447 & n5210 ) | ( n4447 & n5264 ) | ( n5210 & n5264 ) ;
  assign n5266 = n5202 & ~n5265 ;
  assign n5267 = ( n4442 & n5210 ) | ( n4442 & n5264 ) | ( n5210 & n5264 ) ;
  assign n5268 = n5202 & ~n5267 ;
  assign n5269 = ( n3525 & n5266 ) | ( n3525 & n5268 ) | ( n5266 & n5268 ) ;
  assign n5270 = n5263 | n5269 ;
  assign n5228 = ~x12 & x13 ;
  assign n5229 = x12 & ~x13 ;
  assign n5230 = n5228 | n5229 ;
  assign n5221 = x11 & ~x12 ;
  assign n5222 = ~x11 & x12 ;
  assign n5223 = n5221 | n5222 ;
  assign n5224 = x13 & ~x14 ;
  assign n5225 = ~x13 & x14 ;
  assign n5226 = n5224 | n5225 ;
  assign n5236 = ~n5223 & n5226 ;
  assign n5237 = ~n5230 & n5236 ;
  assign n5271 = n4245 & n5237 ;
  assign n5272 = ( n4303 & n5237 ) | ( n4303 & n5271 ) | ( n5237 & n5271 ) ;
  assign n5231 = ~n5223 & n5230 ;
  assign n5273 = n5192 & n5231 ;
  assign n5274 = ( n5179 & n5231 ) | ( n5179 & n5273 ) | ( n5231 & n5273 ) ;
  assign n5275 = n5272 | n5274 ;
  assign n5227 = n5223 & n5226 ;
  assign n5234 = n5223 & ~n5226 ;
  assign n5276 = n5117 & n5234 ;
  assign n5277 = n5227 | n5276 ;
  assign n5278 = n5227 | n5234 ;
  assign n5279 = ( ~n5037 & n5277 ) | ( ~n5037 & n5278 ) | ( n5277 & n5278 ) ;
  assign n5280 = n5275 | n5279 ;
  assign n5281 = ( ~n5037 & n5234 ) | ( ~n5037 & n5276 ) | ( n5234 & n5276 ) ;
  assign n5282 = n5275 | n5281 ;
  assign n5283 = n5280 & n5282 ;
  assign n5284 = ( ~n5270 & n5280 ) | ( ~n5270 & n5283 ) | ( n5280 & n5283 ) ;
  assign n5285 = ~x14 & n5283 ;
  assign n5286 = ~x14 & n5280 ;
  assign n5287 = ( ~n5270 & n5285 ) | ( ~n5270 & n5286 ) | ( n5285 & n5286 ) ;
  assign n5288 = x14 | n5285 ;
  assign n5289 = x14 | n5286 ;
  assign n5290 = ( ~n5270 & n5288 ) | ( ~n5270 & n5289 ) | ( n5288 & n5289 ) ;
  assign n5291 = ( ~n5284 & n5287 ) | ( ~n5284 & n5290 ) | ( n5287 & n5290 ) ;
  assign n5292 = ~n5258 & n5291 ;
  assign n5293 = n4547 & n4993 ;
  assign n5294 = n4547 | n4993 ;
  assign n5295 = ~n5293 & n5294 ;
  assign n5296 = n5196 & n5208 ;
  assign n5297 = ( n4442 & n5198 ) | ( n4442 & n5296 ) | ( n5198 & n5296 ) ;
  assign n5298 = ( n4447 & n5198 ) | ( n4447 & n5296 ) | ( n5198 & n5296 ) ;
  assign n5299 = ( ~n3525 & n5297 ) | ( ~n3525 & n5298 ) | ( n5297 & n5298 ) ;
  assign n5300 = n4397 | n4434 ;
  assign n5301 = ( n4447 & n5208 ) | ( n4447 & n5300 ) | ( n5208 & n5300 ) ;
  assign n5302 = n5196 | n5301 ;
  assign n5303 = ( n4442 & n5208 ) | ( n4442 & n5300 ) | ( n5208 & n5300 ) ;
  assign n5304 = n5196 | n5303 ;
  assign n5305 = ( ~n3525 & n5302 ) | ( ~n3525 & n5304 ) | ( n5302 & n5304 ) ;
  assign n5306 = ~n5299 & n5305 ;
  assign n5307 = n4396 & n5237 ;
  assign n5308 = n4245 & n5231 ;
  assign n5309 = ( n4303 & n5231 ) | ( n4303 & n5308 ) | ( n5231 & n5308 ) ;
  assign n5310 = n5307 | n5309 ;
  assign n5311 = n5192 & n5234 ;
  assign n5312 = ( n5179 & n5234 ) | ( n5179 & n5311 ) | ( n5234 & n5311 ) ;
  assign n5314 = n5227 | n5312 ;
  assign n5315 = n5310 | n5314 ;
  assign n5313 = n5310 | n5312 ;
  assign n5316 = n5313 & n5315 ;
  assign n5317 = ( n5306 & n5315 ) | ( n5306 & n5316 ) | ( n5315 & n5316 ) ;
  assign n5318 = x14 & n5316 ;
  assign n5319 = x14 & n5315 ;
  assign n5320 = ( n5306 & n5318 ) | ( n5306 & n5319 ) | ( n5318 & n5319 ) ;
  assign n5321 = x14 & ~n5318 ;
  assign n5322 = x14 & ~n5319 ;
  assign n5323 = ( ~n5306 & n5321 ) | ( ~n5306 & n5322 ) | ( n5321 & n5322 ) ;
  assign n5324 = ( n5317 & ~n5320 ) | ( n5317 & n5323 ) | ( ~n5320 & n5323 ) ;
  assign n5325 = n5295 & n5324 ;
  assign n5326 = n5295 & ~n5325 ;
  assign n5327 = ~n5295 & n5324 ;
  assign n5328 = n5326 | n5327 ;
  assign n5329 = ~n4573 & n4991 ;
  assign n5330 = n4573 & ~n4991 ;
  assign n5331 = n5329 | n5330 ;
  assign n4435 = n4399 & n4430 ;
  assign n4443 = ( n4434 & n4435 ) | ( n4434 & n4442 ) | ( n4435 & n4442 ) ;
  assign n4448 = ( n4434 & n4435 ) | ( n4434 & n4447 ) | ( n4435 & n4447 ) ;
  assign n4449 = ( ~n3525 & n4443 ) | ( ~n3525 & n4448 ) | ( n4443 & n4448 ) ;
  assign n4450 = ( n4396 & ~n4429 ) | ( n4396 & n4447 ) | ( ~n4429 & n4447 ) ;
  assign n4451 = n4399 | n4450 ;
  assign n4452 = ( n4396 & ~n4429 ) | ( n4396 & n4442 ) | ( ~n4429 & n4442 ) ;
  assign n4453 = n4399 | n4452 ;
  assign n4454 = ( ~n3525 & n4451 ) | ( ~n3525 & n4453 ) | ( n4451 & n4453 ) ;
  assign n4455 = ~n4449 & n4454 ;
  assign n5332 = ~n4429 & n5237 ;
  assign n5333 = n4396 & n5231 ;
  assign n5334 = n5332 | n5333 ;
  assign n5335 = n4245 & n5234 ;
  assign n5336 = ( n4303 & n5234 ) | ( n4303 & n5335 ) | ( n5234 & n5335 ) ;
  assign n5338 = n5227 | n5336 ;
  assign n5339 = n5334 | n5338 ;
  assign n5337 = n5334 | n5336 ;
  assign n5340 = n5337 & n5339 ;
  assign n5341 = ( n4455 & n5339 ) | ( n4455 & n5340 ) | ( n5339 & n5340 ) ;
  assign n5342 = x14 & n5340 ;
  assign n5343 = x14 & n5339 ;
  assign n5344 = ( n4455 & n5342 ) | ( n4455 & n5343 ) | ( n5342 & n5343 ) ;
  assign n5345 = x14 & ~n5342 ;
  assign n5346 = x14 & ~n5343 ;
  assign n5347 = ( ~n4455 & n5345 ) | ( ~n4455 & n5346 ) | ( n5345 & n5346 ) ;
  assign n5348 = ( n5341 & ~n5344 ) | ( n5341 & n5347 ) | ( ~n5344 & n5347 ) ;
  assign n5349 = ~n5331 & n5348 ;
  assign n5350 = n5331 | n5349 ;
  assign n5351 = n5331 & n5348 ;
  assign n5352 = n5350 & ~n5351 ;
  assign n5353 = ~n4596 & n4989 ;
  assign n5354 = n4596 & ~n4989 ;
  assign n5355 = n5353 | n5354 ;
  assign n5356 = ~n4429 & n5231 ;
  assign n5357 = n5231 | n5237 ;
  assign n5358 = ( ~n4429 & n5237 ) | ( ~n4429 & n5357 ) | ( n5237 & n5357 ) ;
  assign n5359 = ( n4206 & n5356 ) | ( n4206 & n5358 ) | ( n5356 & n5358 ) ;
  assign n5360 = n4396 & n5234 ;
  assign n5362 = n5227 | n5360 ;
  assign n5363 = n5359 | n5362 ;
  assign n5361 = n5359 | n5360 ;
  assign n5364 = n5361 & n5363 ;
  assign n5365 = ( ~n4501 & n5363 ) | ( ~n4501 & n5364 ) | ( n5363 & n5364 ) ;
  assign n5366 = ~x14 & n5364 ;
  assign n5367 = ~x14 & n5363 ;
  assign n5368 = ( ~n4501 & n5366 ) | ( ~n4501 & n5367 ) | ( n5366 & n5367 ) ;
  assign n5369 = x14 | n5366 ;
  assign n5370 = x14 | n5367 ;
  assign n5371 = ( ~n4501 & n5369 ) | ( ~n4501 & n5370 ) | ( n5369 & n5370 ) ;
  assign n5372 = ( ~n5365 & n5368 ) | ( ~n5365 & n5371 ) | ( n5368 & n5371 ) ;
  assign n5373 = ~n5355 & n5372 ;
  assign n5374 = n5355 | n5373 ;
  assign n5375 = n5355 & n5372 ;
  assign n5376 = n5374 & ~n5375 ;
  assign n5377 = n4623 & n4987 ;
  assign n5378 = n4623 | n4987 ;
  assign n5379 = ~n5377 & n5378 ;
  assign n5380 = n4206 & n5231 ;
  assign n5381 = ~n4429 & n5234 ;
  assign n5382 = n3439 & n5237 ;
  assign n5383 = ( ~n3420 & n5237 ) | ( ~n3420 & n5382 ) | ( n5237 & n5382 ) ;
  assign n5384 = n5381 | n5383 ;
  assign n5385 = n5380 | n5384 ;
  assign n5386 = n5227 | n5380 ;
  assign n5387 = n5384 | n5386 ;
  assign n5388 = ( ~n4527 & n5385 ) | ( ~n4527 & n5387 ) | ( n5385 & n5387 ) ;
  assign n5389 = ~x14 & n5387 ;
  assign n5390 = ~x14 & n5385 ;
  assign n5391 = ( ~n4527 & n5389 ) | ( ~n4527 & n5390 ) | ( n5389 & n5390 ) ;
  assign n5392 = x14 | n5390 ;
  assign n5393 = x14 | n5389 ;
  assign n5394 = ( ~n4527 & n5392 ) | ( ~n4527 & n5393 ) | ( n5392 & n5393 ) ;
  assign n5395 = ( ~n5388 & n5391 ) | ( ~n5388 & n5394 ) | ( n5391 & n5394 ) ;
  assign n5396 = n5379 & n5395 ;
  assign n5397 = n5379 & ~n5396 ;
  assign n5398 = ~n5379 & n5395 ;
  assign n5399 = n5397 | n5398 ;
  assign n5400 = ( n4668 & n4669 ) | ( n4668 & n4985 ) | ( n4669 & n4985 ) ;
  assign n5401 = n4644 | n4668 ;
  assign n5402 = n4985 | n5401 ;
  assign n5403 = ~n5400 & n5402 ;
  assign n5404 = n4206 & n5234 ;
  assign n5405 = n3386 & n5237 ;
  assign n5406 = n3439 & n5231 ;
  assign n5407 = ( ~n3420 & n5231 ) | ( ~n3420 & n5406 ) | ( n5231 & n5406 ) ;
  assign n5408 = n5405 | n5407 ;
  assign n5409 = n5404 | n5408 ;
  assign n5410 = n5227 | n5404 ;
  assign n5411 = n5408 | n5410 ;
  assign n5412 = ( ~n4220 & n5409 ) | ( ~n4220 & n5411 ) | ( n5409 & n5411 ) ;
  assign n5413 = ~x14 & n5411 ;
  assign n5414 = ~x14 & n5409 ;
  assign n5415 = ( ~n4220 & n5413 ) | ( ~n4220 & n5414 ) | ( n5413 & n5414 ) ;
  assign n5416 = x14 | n5414 ;
  assign n5417 = x14 | n5413 ;
  assign n5418 = ( ~n4220 & n5416 ) | ( ~n4220 & n5417 ) | ( n5416 & n5417 ) ;
  assign n5419 = ( ~n5412 & n5415 ) | ( ~n5412 & n5418 ) | ( n5415 & n5418 ) ;
  assign n5420 = n5403 & n5419 ;
  assign n5421 = n4984 & ~n4985 ;
  assign n5422 = n4673 & ~n4985 ;
  assign n5423 = n5421 | n5422 ;
  assign n5424 = n3386 & n5231 ;
  assign n5425 = n3507 & n5237 ;
  assign n5426 = ( n3483 & n5237 ) | ( n3483 & n5425 ) | ( n5237 & n5425 ) ;
  assign n5427 = n3439 & n5234 ;
  assign n5428 = ( ~n3420 & n5234 ) | ( ~n3420 & n5427 ) | ( n5234 & n5427 ) ;
  assign n5429 = n5426 | n5428 ;
  assign n5430 = n5424 | n5429 ;
  assign n5431 = n5227 | n5430 ;
  assign n5432 = ( ~n3530 & n5430 ) | ( ~n3530 & n5431 ) | ( n5430 & n5431 ) ;
  assign n5433 = ~x14 & n5431 ;
  assign n5434 = ~x14 & n5430 ;
  assign n5435 = ( ~n3530 & n5433 ) | ( ~n3530 & n5434 ) | ( n5433 & n5434 ) ;
  assign n5436 = x14 | n5433 ;
  assign n5437 = x14 | n5434 ;
  assign n5438 = ( ~n3530 & n5436 ) | ( ~n3530 & n5437 ) | ( n5436 & n5437 ) ;
  assign n5439 = ( ~n5432 & n5435 ) | ( ~n5432 & n5438 ) | ( n5435 & n5438 ) ;
  assign n5440 = n5423 & n5439 ;
  assign n5441 = n5423 & ~n5440 ;
  assign n5442 = ~n5423 & n5439 ;
  assign n5443 = n5441 | n5442 ;
  assign n5444 = n4980 & n4982 ;
  assign n5445 = n4980 | n4982 ;
  assign n5446 = ~n5444 & n5445 ;
  assign n5447 = n2893 & n5237 ;
  assign n5448 = ( ~n2886 & n5237 ) | ( ~n2886 & n5447 ) | ( n5237 & n5447 ) ;
  assign n5449 = n3507 & n5231 ;
  assign n5450 = ( n3483 & n5231 ) | ( n3483 & n5449 ) | ( n5231 & n5449 ) ;
  assign n5451 = n5448 | n5450 ;
  assign n5452 = n3386 & n5234 ;
  assign n5454 = n5227 | n5452 ;
  assign n5455 = n5451 | n5454 ;
  assign n5453 = n5451 | n5452 ;
  assign n5456 = n5453 & n5455 ;
  assign n5457 = ( ~n3568 & n5455 ) | ( ~n3568 & n5456 ) | ( n5455 & n5456 ) ;
  assign n5458 = ~x14 & n5456 ;
  assign n5459 = ~x14 & n5455 ;
  assign n5460 = ( ~n3568 & n5458 ) | ( ~n3568 & n5459 ) | ( n5458 & n5459 ) ;
  assign n5461 = x14 | n5458 ;
  assign n5462 = x14 | n5459 ;
  assign n5463 = ( ~n3568 & n5461 ) | ( ~n3568 & n5462 ) | ( n5461 & n5462 ) ;
  assign n5464 = ( ~n5457 & n5460 ) | ( ~n5457 & n5463 ) | ( n5460 & n5463 ) ;
  assign n5465 = n5446 & n5464 ;
  assign n5466 = n4743 | n4976 ;
  assign n5467 = ~n4977 & n5466 ;
  assign n5468 = n2691 & n5237 ;
  assign n5469 = ( n2678 & n5237 ) | ( n2678 & n5468 ) | ( n5237 & n5468 ) ;
  assign n5470 = n2701 & n5231 ;
  assign n5471 = ( ~n2784 & n5231 ) | ( ~n2784 & n5470 ) | ( n5231 & n5470 ) ;
  assign n5472 = n5469 | n5471 ;
  assign n5473 = n2893 & n5234 ;
  assign n5474 = ( ~n2886 & n5234 ) | ( ~n2886 & n5473 ) | ( n5234 & n5473 ) ;
  assign n5475 = n5472 | n5474 ;
  assign n5476 = n5227 | n5475 ;
  assign n5477 = n5475 & n5476 ;
  assign n5478 = ( ~n2914 & n5476 ) | ( ~n2914 & n5477 ) | ( n5476 & n5477 ) ;
  assign n5479 = ~x14 & n5477 ;
  assign n5480 = ~x14 & n5476 ;
  assign n5481 = ( ~n2914 & n5479 ) | ( ~n2914 & n5480 ) | ( n5479 & n5480 ) ;
  assign n5482 = x14 | n5479 ;
  assign n5483 = x14 | n5480 ;
  assign n5484 = ( ~n2914 & n5482 ) | ( ~n2914 & n5483 ) | ( n5482 & n5483 ) ;
  assign n5485 = ( ~n5478 & n5481 ) | ( ~n5478 & n5484 ) | ( n5481 & n5484 ) ;
  assign n5486 = n5467 & n5485 ;
  assign n5487 = n5467 & ~n5486 ;
  assign n5488 = ~n5467 & n5485 ;
  assign n5489 = n5487 | n5488 ;
  assign n5490 = n4972 & n4974 ;
  assign n5491 = n4972 | n4974 ;
  assign n5492 = ~n5490 & n5491 ;
  assign n5493 = n2701 & n5234 ;
  assign n5494 = ( ~n2784 & n5234 ) | ( ~n2784 & n5493 ) | ( n5234 & n5493 ) ;
  assign n5495 = n2691 & n5231 ;
  assign n5496 = ( n2678 & n5231 ) | ( n2678 & n5495 ) | ( n5231 & n5495 ) ;
  assign n5497 = n5494 | n5496 ;
  assign n5498 = n2199 & n5237 ;
  assign n5499 = ( ~n2185 & n5237 ) | ( ~n2185 & n5498 ) | ( n5237 & n5498 ) ;
  assign n5500 = n5497 | n5499 ;
  assign n5501 = n5227 | n5499 ;
  assign n5502 = n5497 | n5501 ;
  assign n5503 = ( n2960 & n5500 ) | ( n2960 & n5502 ) | ( n5500 & n5502 ) ;
  assign n5504 = x14 & n5502 ;
  assign n5505 = x14 & n5500 ;
  assign n5506 = ( n2960 & n5504 ) | ( n2960 & n5505 ) | ( n5504 & n5505 ) ;
  assign n5507 = x14 & ~n5505 ;
  assign n5508 = x14 & ~n5504 ;
  assign n5509 = ( ~n2960 & n5507 ) | ( ~n2960 & n5508 ) | ( n5507 & n5508 ) ;
  assign n5510 = ( n5503 & ~n5506 ) | ( n5503 & n5509 ) | ( ~n5506 & n5509 ) ;
  assign n5511 = n5492 & n5510 ;
  assign n5512 = n4967 & n4970 ;
  assign n5513 = n4967 & ~n5512 ;
  assign n5516 = n2090 & n5237 ;
  assign n5517 = ( ~n2082 & n5237 ) | ( ~n2082 & n5516 ) | ( n5237 & n5516 ) ;
  assign n5518 = n2691 & n5234 ;
  assign n5519 = ( n2678 & n5234 ) | ( n2678 & n5518 ) | ( n5234 & n5518 ) ;
  assign n5520 = n2199 & n5231 ;
  assign n5521 = ( ~n2185 & n5231 ) | ( ~n2185 & n5520 ) | ( n5231 & n5520 ) ;
  assign n5522 = n5519 | n5521 ;
  assign n5523 = n5517 | n5522 ;
  assign n5524 = n5227 | n5523 ;
  assign n5525 = ( n2985 & n5523 ) | ( n2985 & n5524 ) | ( n5523 & n5524 ) ;
  assign n5526 = x14 & n5524 ;
  assign n5527 = x14 & n5523 ;
  assign n5528 = ( n2985 & n5526 ) | ( n2985 & n5527 ) | ( n5526 & n5527 ) ;
  assign n5529 = x14 & ~n5526 ;
  assign n5530 = x14 & ~n5527 ;
  assign n5531 = ( ~n2985 & n5529 ) | ( ~n2985 & n5530 ) | ( n5529 & n5530 ) ;
  assign n5532 = ( n5525 & ~n5528 ) | ( n5525 & n5531 ) | ( ~n5528 & n5531 ) ;
  assign n5514 = ~n4967 & n4970 ;
  assign n5533 = n5514 & n5532 ;
  assign n5534 = ( n5513 & n5532 ) | ( n5513 & n5533 ) | ( n5532 & n5533 ) ;
  assign n5515 = n5513 | n5514 ;
  assign n5535 = n5515 & ~n5534 ;
  assign n5536 = ~n5514 & n5532 ;
  assign n5537 = ~n5513 & n5536 ;
  assign n5538 = n5535 | n5537 ;
  assign n5539 = ~n4962 & n4965 ;
  assign n5540 = n4962 & ~n4965 ;
  assign n5541 = n5539 | n5540 ;
  assign n5542 = n2090 & n5231 ;
  assign n5543 = ( ~n2082 & n5231 ) | ( ~n2082 & n5542 ) | ( n5231 & n5542 ) ;
  assign n5544 = n2279 & n5237 ;
  assign n5545 = ( ~n2269 & n5237 ) | ( ~n2269 & n5544 ) | ( n5237 & n5544 ) ;
  assign n5546 = n2199 & n5234 ;
  assign n5547 = ( ~n2185 & n5234 ) | ( ~n2185 & n5546 ) | ( n5234 & n5546 ) ;
  assign n5548 = n5545 | n5547 ;
  assign n5549 = n5543 | n5548 ;
  assign n5550 = n5227 | n5549 ;
  assign n5551 = ( ~n2325 & n5549 ) | ( ~n2325 & n5550 ) | ( n5549 & n5550 ) ;
  assign n5552 = n5549 & n5550 ;
  assign n5553 = ( ~n2299 & n5551 ) | ( ~n2299 & n5552 ) | ( n5551 & n5552 ) ;
  assign n5554 = ~x14 & n5553 ;
  assign n5555 = x14 | n5553 ;
  assign n5556 = ( ~n5553 & n5554 ) | ( ~n5553 & n5555 ) | ( n5554 & n5555 ) ;
  assign n5557 = n5541 & n5556 ;
  assign n5558 = n5541 | n5556 ;
  assign n5559 = ~n5557 & n5558 ;
  assign n5560 = n4958 | n4960 ;
  assign n5561 = ~n4961 & n5560 ;
  assign n5562 = n1634 & n5237 ;
  assign n5563 = ( n1630 & n5237 ) | ( n1630 & n5562 ) | ( n5237 & n5562 ) ;
  assign n5564 = n2279 & n5231 ;
  assign n5565 = ( ~n2269 & n5231 ) | ( ~n2269 & n5564 ) | ( n5231 & n5564 ) ;
  assign n5566 = n5563 | n5565 ;
  assign n5567 = n2090 & n5234 ;
  assign n5568 = ( ~n2082 & n5234 ) | ( ~n2082 & n5567 ) | ( n5234 & n5567 ) ;
  assign n5569 = n5566 | n5568 ;
  assign n5570 = n5227 | n5569 ;
  assign n5571 = n5569 & n5570 ;
  assign n5572 = ( n2568 & n5570 ) | ( n2568 & n5571 ) | ( n5570 & n5571 ) ;
  assign n5573 = x14 & n5571 ;
  assign n5574 = x14 & n5570 ;
  assign n5575 = ( n2568 & n5573 ) | ( n2568 & n5574 ) | ( n5573 & n5574 ) ;
  assign n5576 = x14 & ~n5573 ;
  assign n5577 = x14 & ~n5574 ;
  assign n5578 = ( ~n2568 & n5576 ) | ( ~n2568 & n5577 ) | ( n5576 & n5577 ) ;
  assign n5579 = ( n5572 & ~n5575 ) | ( n5572 & n5578 ) | ( ~n5575 & n5578 ) ;
  assign n5580 = n5561 & n5579 ;
  assign n5581 = n4848 | n4956 ;
  assign n5582 = ~n4957 & n5581 ;
  assign n5583 = n1708 & n5237 ;
  assign n5584 = n1634 & n5231 ;
  assign n5585 = ( n1630 & n5231 ) | ( n1630 & n5584 ) | ( n5231 & n5584 ) ;
  assign n5586 = n2279 & n5234 ;
  assign n5587 = ( ~n2269 & n5234 ) | ( ~n2269 & n5586 ) | ( n5234 & n5586 ) ;
  assign n5588 = n5585 | n5587 ;
  assign n5589 = n5583 | n5588 ;
  assign n5590 = n5227 | n5589 ;
  assign n5591 = n5589 & n5590 ;
  assign n5592 = ( ~n2343 & n5590 ) | ( ~n2343 & n5591 ) | ( n5590 & n5591 ) ;
  assign n5593 = ~x14 & n5591 ;
  assign n5594 = ~x14 & n5590 ;
  assign n5595 = ( ~n2343 & n5593 ) | ( ~n2343 & n5594 ) | ( n5593 & n5594 ) ;
  assign n5596 = x14 | n5593 ;
  assign n5597 = x14 | n5594 ;
  assign n5598 = ( ~n2343 & n5596 ) | ( ~n2343 & n5597 ) | ( n5596 & n5597 ) ;
  assign n5599 = ( ~n5592 & n5595 ) | ( ~n5592 & n5598 ) | ( n5595 & n5598 ) ;
  assign n5600 = n5582 & n5599 ;
  assign n5601 = n4952 & n4954 ;
  assign n5602 = n4952 | n4954 ;
  assign n5603 = ~n5601 & n5602 ;
  assign n5604 = n1708 & n5231 ;
  assign n5605 = n1793 & n5237 ;
  assign n5606 = ( n1783 & n5237 ) | ( n1783 & n5605 ) | ( n5237 & n5605 ) ;
  assign n5607 = n1634 & n5234 ;
  assign n5608 = ( n1630 & n5234 ) | ( n1630 & n5607 ) | ( n5234 & n5607 ) ;
  assign n5609 = n5606 | n5608 ;
  assign n5610 = n5604 | n5609 ;
  assign n5611 = n5227 | n5610 ;
  assign n5612 = n5610 & n5611 ;
  assign n5613 = ( n1814 & n5611 ) | ( n1814 & n5612 ) | ( n5611 & n5612 ) ;
  assign n5614 = x14 & n5612 ;
  assign n5615 = x14 & n5611 ;
  assign n5616 = ( n1814 & n5614 ) | ( n1814 & n5615 ) | ( n5614 & n5615 ) ;
  assign n5617 = x14 & ~n5614 ;
  assign n5618 = x14 & ~n5615 ;
  assign n5619 = ( ~n1814 & n5617 ) | ( ~n1814 & n5618 ) | ( n5617 & n5618 ) ;
  assign n5620 = ( n5613 & ~n5616 ) | ( n5613 & n5619 ) | ( ~n5616 & n5619 ) ;
  assign n5621 = n5603 & n5620 ;
  assign n5622 = n4948 & n4950 ;
  assign n5623 = n4948 | n4950 ;
  assign n5624 = ~n5622 & n5623 ;
  assign n5625 = ~n523 & n5237 ;
  assign n5626 = n1793 & n5231 ;
  assign n5627 = ( n1783 & n5231 ) | ( n1783 & n5626 ) | ( n5231 & n5626 ) ;
  assign n5628 = n5625 | n5627 ;
  assign n5629 = n1708 & n5234 ;
  assign n5630 = n5628 | n5629 ;
  assign n5631 = n5227 | n5629 ;
  assign n5632 = n5628 | n5631 ;
  assign n5633 = ( ~n1852 & n5630 ) | ( ~n1852 & n5632 ) | ( n5630 & n5632 ) ;
  assign n5634 = ~x14 & n5632 ;
  assign n5635 = ~x14 & n5630 ;
  assign n5636 = ( ~n1852 & n5634 ) | ( ~n1852 & n5635 ) | ( n5634 & n5635 ) ;
  assign n5637 = x14 | n5635 ;
  assign n5638 = x14 | n5634 ;
  assign n5639 = ( ~n1852 & n5637 ) | ( ~n1852 & n5638 ) | ( n5637 & n5638 ) ;
  assign n5640 = ( ~n5633 & n5636 ) | ( ~n5633 & n5639 ) | ( n5636 & n5639 ) ;
  assign n5641 = n5624 & n5640 ;
  assign n5642 = n4944 | n4945 ;
  assign n5643 = n4928 | n5642 ;
  assign n5644 = ~n4947 & n5643 ;
  assign n5645 = ~n523 & n5231 ;
  assign n5646 = n352 & n5237 ;
  assign n5647 = ( ~n339 & n5237 ) | ( ~n339 & n5646 ) | ( n5237 & n5646 ) ;
  assign n5648 = n1793 & n5234 ;
  assign n5649 = ( n1783 & n5234 ) | ( n1783 & n5648 ) | ( n5234 & n5648 ) ;
  assign n5650 = n5647 | n5649 ;
  assign n5651 = n5645 | n5650 ;
  assign n5652 = n5227 | n5651 ;
  assign n5653 = n5651 & n5652 ;
  assign n5654 = ( n1884 & n5652 ) | ( n1884 & n5653 ) | ( n5652 & n5653 ) ;
  assign n5655 = x14 & n5653 ;
  assign n5656 = x14 & n5652 ;
  assign n5657 = ( n1884 & n5655 ) | ( n1884 & n5656 ) | ( n5655 & n5656 ) ;
  assign n5658 = x14 & ~n5655 ;
  assign n5659 = x14 & ~n5656 ;
  assign n5660 = ( ~n1884 & n5658 ) | ( ~n1884 & n5659 ) | ( n5658 & n5659 ) ;
  assign n5661 = ( n5654 & ~n5657 ) | ( n5654 & n5660 ) | ( ~n5657 & n5660 ) ;
  assign n5662 = n5644 & n5661 ;
  assign n5663 = n5644 | n5661 ;
  assign n5664 = ~n5662 & n5663 ;
  assign n5665 = ~n829 & n5237 ;
  assign n5666 = n352 & n5231 ;
  assign n5667 = ( ~n339 & n5231 ) | ( ~n339 & n5666 ) | ( n5231 & n5666 ) ;
  assign n5668 = n5665 | n5667 ;
  assign n5669 = ~n523 & n5234 ;
  assign n5670 = n5227 | n5669 ;
  assign n5671 = n5668 | n5670 ;
  assign n5672 = ~x14 & n5671 ;
  assign n5673 = n5668 | n5669 ;
  assign n5674 = ~x14 & n5673 ;
  assign n5675 = ( ~n1055 & n5672 ) | ( ~n1055 & n5674 ) | ( n5672 & n5674 ) ;
  assign n5676 = x14 & n5671 ;
  assign n5677 = x14 & ~n5676 ;
  assign n5678 = x14 & n5669 ;
  assign n5679 = ( x14 & n5668 ) | ( x14 & n5678 ) | ( n5668 & n5678 ) ;
  assign n5680 = x14 & ~n5679 ;
  assign n5681 = ( n1055 & n5677 ) | ( n1055 & n5680 ) | ( n5677 & n5680 ) ;
  assign n5682 = n5675 | n5681 ;
  assign n5683 = n4921 | n4923 ;
  assign n5684 = x17 & ~n4921 ;
  assign n5685 = ( n4904 & n5683 ) | ( n4904 & ~n5684 ) | ( n5683 & ~n5684 ) ;
  assign n5686 = ~n4926 & n5685 ;
  assign n5687 = n5682 & n5686 ;
  assign n5688 = x17 | n4918 ;
  assign n5689 = ( ~n4911 & n4918 ) | ( ~n4911 & n5688 ) | ( n4918 & n5688 ) ;
  assign n5690 = n4912 | n5689 ;
  assign n5691 = ~n4921 & n5690 ;
  assign n5692 = ~n829 & n5231 ;
  assign n5693 = n352 & n5234 ;
  assign n5694 = ( ~n339 & n5234 ) | ( ~n339 & n5693 ) | ( n5234 & n5693 ) ;
  assign n5695 = n5692 | n5694 ;
  assign n5696 = n692 & n5237 ;
  assign n5697 = ( n674 & n5237 ) | ( n674 & n5696 ) | ( n5237 & n5696 ) ;
  assign n5698 = n5695 | n5697 ;
  assign n5699 = n5227 | n5697 ;
  assign n5700 = n5695 | n5699 ;
  assign n5701 = ( ~n1209 & n5698 ) | ( ~n1209 & n5700 ) | ( n5698 & n5700 ) ;
  assign n5702 = ~x14 & n5700 ;
  assign n5703 = ~x14 & n5698 ;
  assign n5704 = ( ~n1209 & n5702 ) | ( ~n1209 & n5703 ) | ( n5702 & n5703 ) ;
  assign n5705 = x14 | n5703 ;
  assign n5706 = x14 | n5702 ;
  assign n5707 = ( ~n1209 & n5705 ) | ( ~n1209 & n5706 ) | ( n5705 & n5706 ) ;
  assign n5708 = ( ~n5701 & n5704 ) | ( ~n5701 & n5707 ) | ( n5704 & n5707 ) ;
  assign n5709 = n5691 & n5708 ;
  assign n5710 = ( ~n1027 & n4914 ) | ( ~n1027 & n4916 ) | ( n4914 & n4916 ) ;
  assign n5711 = ~n922 & n5231 ;
  assign n5712 = n1042 & n5237 ;
  assign n5713 = ( ~n1027 & n5237 ) | ( ~n1027 & n5712 ) | ( n5237 & n5712 ) ;
  assign n5714 = n5711 | n5713 ;
  assign n5715 = n692 & n5234 ;
  assign n5716 = ( n674 & n5234 ) | ( n674 & n5715 ) | ( n5234 & n5715 ) ;
  assign n5717 = n5714 | n5716 ;
  assign n5718 = ( n1538 & n5227 ) | ( n1538 & n5717 ) | ( n5227 & n5717 ) ;
  assign n5719 = ( x14 & ~n5717 ) | ( x14 & n5718 ) | ( ~n5717 & n5718 ) ;
  assign n5720 = ~n5718 & n5719 ;
  assign n5721 = ~n922 & n5234 ;
  assign n5722 = n1042 & n5231 ;
  assign n5723 = ( ~n1027 & n5231 ) | ( ~n1027 & n5722 ) | ( n5231 & n5722 ) ;
  assign n5724 = n5721 | n5723 ;
  assign n5725 = n5227 | n5723 ;
  assign n5726 = n5721 | n5725 ;
  assign n5727 = ( n1946 & n5724 ) | ( n1946 & n5726 ) | ( n5724 & n5726 ) ;
  assign n5728 = ~x14 & n5727 ;
  assign n5729 = n139 & n5223 ;
  assign n5730 = ( n1041 & n5223 ) | ( n1041 & n5729 ) | ( n5223 & n5729 ) ;
  assign n5731 = x14 & ~n5730 ;
  assign n5732 = n5223 | n5729 ;
  assign n5733 = x14 & ~n5732 ;
  assign n5734 = ( n1027 & n5731 ) | ( n1027 & n5733 ) | ( n5731 & n5733 ) ;
  assign n5735 = x14 & n5734 ;
  assign n5736 = ~n5727 & n5735 ;
  assign n5737 = ( n5728 & n5734 ) | ( n5728 & n5736 ) | ( n5734 & n5736 ) ;
  assign n5738 = x14 | n5717 ;
  assign n5739 = n5718 | n5738 ;
  assign n5740 = n5737 & n5739 ;
  assign n5741 = ~x14 & n5737 ;
  assign n5742 = ( n5720 & n5740 ) | ( n5720 & n5741 ) | ( n5740 & n5741 ) ;
  assign n5743 = n5710 & n5742 ;
  assign n5744 = n5742 & ~n5743 ;
  assign n5745 = ~n829 & n5234 ;
  assign n5746 = ~n922 & n5237 ;
  assign n5747 = n5745 | n5746 ;
  assign n5748 = n692 & n5231 ;
  assign n5749 = ( n674 & n5231 ) | ( n674 & n5748 ) | ( n5231 & n5748 ) ;
  assign n5750 = n5747 | n5749 ;
  assign n5751 = n5227 | n5749 ;
  assign n5752 = n5747 | n5751 ;
  assign n5753 = ( n1554 & n5750 ) | ( n1554 & n5752 ) | ( n5750 & n5752 ) ;
  assign n5754 = x14 & n5752 ;
  assign n5755 = x14 & n5750 ;
  assign n5756 = ( n1554 & n5754 ) | ( n1554 & n5755 ) | ( n5754 & n5755 ) ;
  assign n5757 = x14 & ~n5755 ;
  assign n5758 = x14 & ~n5754 ;
  assign n5759 = ( ~n1554 & n5757 ) | ( ~n1554 & n5758 ) | ( n5757 & n5758 ) ;
  assign n5760 = ( n5753 & ~n5756 ) | ( n5753 & n5759 ) | ( ~n5756 & n5759 ) ;
  assign n5761 = n5710 & ~n5742 ;
  assign n5762 = n5760 & n5761 ;
  assign n5763 = ( n5744 & n5760 ) | ( n5744 & n5762 ) | ( n5760 & n5762 ) ;
  assign n5764 = n5743 | n5763 ;
  assign n5765 = n5691 | n5708 ;
  assign n5766 = ~n5709 & n5765 ;
  assign n5767 = n5709 | n5766 ;
  assign n5768 = ( n5709 & n5764 ) | ( n5709 & n5767 ) | ( n5764 & n5767 ) ;
  assign n5769 = n5682 | n5686 ;
  assign n5770 = ~n5687 & n5769 ;
  assign n5771 = n5687 | n5770 ;
  assign n5772 = ( n5687 & n5768 ) | ( n5687 & n5771 ) | ( n5768 & n5771 ) ;
  assign n5773 = n5664 & n5772 ;
  assign n5774 = n5662 | n5773 ;
  assign n5775 = ~n5624 & n5640 ;
  assign n5776 = ( n5624 & ~n5641 ) | ( n5624 & n5775 ) | ( ~n5641 & n5775 ) ;
  assign n5777 = n5774 & n5776 ;
  assign n5778 = n5641 | n5777 ;
  assign n5779 = n5603 & ~n5621 ;
  assign n5780 = ~n5603 & n5620 ;
  assign n5781 = n5779 | n5780 ;
  assign n5782 = n5778 & n5781 ;
  assign n5783 = n5621 | n5782 ;
  assign n5784 = n5582 & ~n5600 ;
  assign n5785 = ~n5582 & n5599 ;
  assign n5786 = n5784 | n5785 ;
  assign n5787 = n5600 | n5786 ;
  assign n5788 = ( n5600 & n5783 ) | ( n5600 & n5787 ) | ( n5783 & n5787 ) ;
  assign n5789 = n5561 | n5579 ;
  assign n5790 = ~n5580 & n5789 ;
  assign n5791 = n5580 | n5790 ;
  assign n5792 = ( n5580 & n5788 ) | ( n5580 & n5791 ) | ( n5788 & n5791 ) ;
  assign n5793 = n5559 & n5792 ;
  assign n5794 = n5557 | n5793 ;
  assign n5795 = n5534 | n5794 ;
  assign n5796 = ( n5534 & n5538 ) | ( n5534 & n5795 ) | ( n5538 & n5795 ) ;
  assign n5797 = ~n5492 & n5510 ;
  assign n5798 = ( n5492 & ~n5511 ) | ( n5492 & n5797 ) | ( ~n5511 & n5797 ) ;
  assign n5799 = n5511 | n5798 ;
  assign n5800 = ( n5511 & n5796 ) | ( n5511 & n5799 ) | ( n5796 & n5799 ) ;
  assign n5801 = n5489 & n5800 ;
  assign n5802 = n5486 | n5801 ;
  assign n5803 = n4722 & n4978 ;
  assign n5804 = n4722 | n4978 ;
  assign n5805 = ~n5803 & n5804 ;
  assign n5806 = n2893 & n5231 ;
  assign n5807 = ( ~n2886 & n5231 ) | ( ~n2886 & n5806 ) | ( n5231 & n5806 ) ;
  assign n5808 = n2701 & n5237 ;
  assign n5809 = ( ~n2784 & n5237 ) | ( ~n2784 & n5808 ) | ( n5237 & n5808 ) ;
  assign n5810 = n3507 & n5234 ;
  assign n5811 = ( n3483 & n5234 ) | ( n3483 & n5810 ) | ( n5234 & n5810 ) ;
  assign n5812 = n5809 | n5811 ;
  assign n5813 = n5807 | n5812 ;
  assign n5814 = n5227 | n5813 ;
  assign n5815 = n5813 & n5814 ;
  assign n5816 = ( n3603 & n5814 ) | ( n3603 & n5815 ) | ( n5814 & n5815 ) ;
  assign n5817 = x14 & n5815 ;
  assign n5818 = x14 & n5814 ;
  assign n5819 = ( n3603 & n5817 ) | ( n3603 & n5818 ) | ( n5817 & n5818 ) ;
  assign n5820 = x14 & ~n5817 ;
  assign n5821 = x14 & ~n5818 ;
  assign n5822 = ( ~n3603 & n5820 ) | ( ~n3603 & n5821 ) | ( n5820 & n5821 ) ;
  assign n5823 = ( n5816 & ~n5819 ) | ( n5816 & n5822 ) | ( ~n5819 & n5822 ) ;
  assign n5824 = n5805 & n5823 ;
  assign n5825 = n5805 & ~n5824 ;
  assign n5826 = ~n5805 & n5823 ;
  assign n5827 = n5825 | n5826 ;
  assign n5828 = n5802 & n5827 ;
  assign n5829 = n5446 | n5464 ;
  assign n5830 = ~n5465 & n5829 ;
  assign n5831 = n5824 & n5830 ;
  assign n5832 = ( n5828 & n5830 ) | ( n5828 & n5831 ) | ( n5830 & n5831 ) ;
  assign n5833 = n5465 | n5832 ;
  assign n5834 = n5443 & n5833 ;
  assign n5835 = ~n5403 & n5419 ;
  assign n5836 = ( n5403 & ~n5420 ) | ( n5403 & n5835 ) | ( ~n5420 & n5835 ) ;
  assign n5837 = n5440 & n5836 ;
  assign n5838 = ( n5834 & n5836 ) | ( n5834 & n5837 ) | ( n5836 & n5837 ) ;
  assign n5839 = n5420 | n5838 ;
  assign n5840 = n5399 & n5839 ;
  assign n5841 = n5396 | n5840 ;
  assign n5842 = ~n5376 & n5841 ;
  assign n5843 = n5373 | n5842 ;
  assign n5844 = ~n5352 & n5843 ;
  assign n5845 = n5349 | n5844 ;
  assign n5846 = n5328 & n5845 ;
  assign n5847 = n5325 | n5846 ;
  assign n5848 = n5258 | n5292 ;
  assign n5849 = n5258 & n5291 ;
  assign n5850 = n5848 & ~n5849 ;
  assign n5851 = ~n5292 & n5850 ;
  assign n5852 = ( n5292 & n5847 ) | ( n5292 & ~n5851 ) | ( n5847 & ~n5851 ) ;
  assign n3969 = n3965 & ~n3968 ;
  assign n3970 = n3562 | n3969 ;
  assign n3971 = n2332 | n2593 ;
  assign n3972 = n1057 & n1793 ;
  assign n3973 = ( n1057 & n1783 ) | ( n1057 & n3972 ) | ( n1783 & n3972 ) ;
  assign n3974 = ~n523 & n1065 ;
  assign n3975 = n352 & n1060 ;
  assign n3976 = ( ~n339 & n1060 ) | ( ~n339 & n3975 ) | ( n1060 & n3975 ) ;
  assign n3977 = n1062 | n3976 ;
  assign n3978 = n3974 | n3977 ;
  assign n3979 = n3973 | n3978 ;
  assign n3980 = n3973 | n3976 ;
  assign n3981 = n3974 | n3980 ;
  assign n3982 = ( n1884 & n3979 ) | ( n1884 & n3981 ) | ( n3979 & n3981 ) ;
  assign n3983 = n347 | n666 ;
  assign n3985 = n3362 | n3984 ;
  assign n3986 = n555 | n762 ;
  assign n3987 = n64 | n500 ;
  assign n3988 = n3986 | n3987 ;
  assign n3989 = n3985 | n3988 ;
  assign n3990 = n1657 | n1725 ;
  assign n3991 = n703 | n3990 ;
  assign n3992 = n3989 | n3991 ;
  assign n3993 = n77 | n233 ;
  assign n3994 = n390 | n3993 ;
  assign n3995 = n594 | n602 ;
  assign n3996 = n1404 | n3995 ;
  assign n3997 = n2040 | n3996 ;
  assign n3998 = n3994 | n3997 ;
  assign n3999 = n3992 | n3998 ;
  assign n4000 = n979 | n1251 ;
  assign n4001 = n1222 | n2835 ;
  assign n4002 = n4000 | n4001 ;
  assign n4003 = n117 | n190 ;
  assign n4004 = n1005 | n4003 ;
  assign n4005 = n1469 | n4004 ;
  assign n4006 = n4002 | n4005 ;
  assign n4007 = n67 | n735 ;
  assign n4008 = n1607 | n4007 ;
  assign n4009 = n223 | n324 ;
  assign n4010 = n2135 | n4009 ;
  assign n4011 = n4008 | n4010 ;
  assign n4012 = n929 | n4011 ;
  assign n4013 = n4006 | n4012 ;
  assign n4014 = n3999 | n4013 ;
  assign n4015 = n3983 | n4014 ;
  assign n4016 = n383 | n479 ;
  assign n4017 = n531 | n4016 ;
  assign n4018 = n406 | n461 ;
  assign n4019 = n325 | n624 ;
  assign n4020 = n4018 | n4019 ;
  assign n4021 = n4017 | n4020 ;
  assign n4022 = n260 | n369 ;
  assign n4023 = n4021 | n4022 ;
  assign n4024 = n491 | n725 ;
  assign n4025 = n4023 | n4024 ;
  assign n4026 = n263 | n1478 ;
  assign n4027 = n133 | n1114 ;
  assign n4028 = n212 | n4027 ;
  assign n4029 = n321 | n654 ;
  assign n4030 = n518 | n4029 ;
  assign n4031 = n4028 | n4030 ;
  assign n4032 = n1436 | n2768 ;
  assign n4033 = n4031 | n4032 ;
  assign n4034 = n4026 | n4033 ;
  assign n4035 = n575 | n1171 ;
  assign n4036 = n205 | n648 ;
  assign n4037 = n331 | n4036 ;
  assign n4038 = n4035 | n4037 ;
  assign n4039 = n465 | n643 ;
  assign n4040 = n448 | n568 ;
  assign n4041 = n4039 | n4040 ;
  assign n4042 = n4038 | n4041 ;
  assign n4043 = n4034 | n4042 ;
  assign n4044 = n4025 | n4043 ;
  assign n4045 = n4015 | n4044 ;
  assign n4046 = n110 | n126 ;
  assign n4047 = n433 | n4046 ;
  assign n4048 = n88 | n901 ;
  assign n4049 = n483 | n4048 ;
  assign n4050 = n4047 | n4049 ;
  assign n4051 = n281 | n621 ;
  assign n4052 = n4050 | n4051 ;
  assign n4053 = n4045 | n4052 ;
  assign n4054 = n3981 & n4053 ;
  assign n4055 = n3973 & n4053 ;
  assign n4056 = ( n3978 & n4053 ) | ( n3978 & n4055 ) | ( n4053 & n4055 ) ;
  assign n4057 = ( n1884 & n4054 ) | ( n1884 & n4056 ) | ( n4054 & n4056 ) ;
  assign n4058 = n3982 & ~n4057 ;
  assign n4059 = ~n3979 & n4053 ;
  assign n4060 = ~n3981 & n4053 ;
  assign n4061 = ( ~n1884 & n4059 ) | ( ~n1884 & n4060 ) | ( n4059 & n4060 ) ;
  assign n4062 = n4058 | n4061 ;
  assign n4063 = n1200 & n4062 ;
  assign n4064 = ( n1571 & n4062 ) | ( n1571 & n4063 ) | ( n4062 & n4063 ) ;
  assign n4065 = n1200 | n4062 ;
  assign n4066 = n1571 | n4065 ;
  assign n4067 = ~n4064 & n4066 ;
  assign n4068 = n1708 & n1826 ;
  assign n4069 = n1634 & n1823 ;
  assign n4070 = ( n1630 & n1823 ) | ( n1630 & n4069 ) | ( n1823 & n4069 ) ;
  assign n4071 = n1829 & n2279 ;
  assign n4072 = ( n1829 & ~n2269 ) | ( n1829 & n4071 ) | ( ~n2269 & n4071 ) ;
  assign n4073 = n4070 | n4072 ;
  assign n4074 = n4068 | n4073 ;
  assign n4075 = n1821 | n4074 ;
  assign n4076 = n4074 & n4075 ;
  assign n4077 = ( ~n2343 & n4075 ) | ( ~n2343 & n4076 ) | ( n4075 & n4076 ) ;
  assign n4078 = ~x29 & n4076 ;
  assign n4079 = ~x29 & n4075 ;
  assign n4080 = ( ~n2343 & n4078 ) | ( ~n2343 & n4079 ) | ( n4078 & n4079 ) ;
  assign n4081 = x29 | n4078 ;
  assign n4082 = x29 | n4079 ;
  assign n4083 = ( ~n2343 & n4081 ) | ( ~n2343 & n4082 ) | ( n4081 & n4082 ) ;
  assign n4084 = ( ~n4077 & n4080 ) | ( ~n4077 & n4083 ) | ( n4080 & n4083 ) ;
  assign n4085 = n4067 & n4084 ;
  assign n4086 = n4067 | n4084 ;
  assign n4087 = ~n4085 & n4086 ;
  assign n4088 = n1843 & n4087 ;
  assign n4089 = ( n2020 & n4087 ) | ( n2020 & n4088 ) | ( n4087 & n4088 ) ;
  assign n4090 = n1843 | n4087 ;
  assign n4091 = n2020 | n4090 ;
  assign n4092 = ~n4089 & n4091 ;
  assign n4093 = n2090 & n2312 ;
  assign n4094 = ( ~n2082 & n2312 ) | ( ~n2082 & n4093 ) | ( n2312 & n4093 ) ;
  assign n4095 = n2315 & n2691 ;
  assign n4096 = ( n2315 & n2678 ) | ( n2315 & n4095 ) | ( n2678 & n4095 ) ;
  assign n4097 = n2199 & n2308 ;
  assign n4098 = ( ~n2185 & n2308 ) | ( ~n2185 & n4097 ) | ( n2308 & n4097 ) ;
  assign n4099 = n4096 | n4098 ;
  assign n4100 = n4094 | n4099 ;
  assign n4101 = n2306 | n4100 ;
  assign n4102 = ( n2985 & n4100 ) | ( n2985 & n4101 ) | ( n4100 & n4101 ) ;
  assign n4103 = x26 & n4101 ;
  assign n4104 = x26 & n4100 ;
  assign n4105 = ( n2985 & n4103 ) | ( n2985 & n4104 ) | ( n4103 & n4104 ) ;
  assign n4106 = x26 & ~n4103 ;
  assign n4107 = x26 & ~n4104 ;
  assign n4108 = ( ~n2985 & n4106 ) | ( ~n2985 & n4107 ) | ( n4106 & n4107 ) ;
  assign n4109 = ( n4102 & ~n4105 ) | ( n4102 & n4108 ) | ( ~n4105 & n4108 ) ;
  assign n4110 = n4092 & n4109 ;
  assign n4111 = n4092 & ~n4110 ;
  assign n4112 = ~n4092 & n4109 ;
  assign n4113 = n4111 | n4112 ;
  assign n4114 = ~n3971 & n4113 ;
  assign n4115 = n3971 & ~n4113 ;
  assign n4116 = n4114 | n4115 ;
  assign n4117 = n2893 & n2928 ;
  assign n4118 = ( ~n2886 & n2928 ) | ( ~n2886 & n4117 ) | ( n2928 & n4117 ) ;
  assign n4119 = n2701 & n2925 ;
  assign n4120 = ( ~n2784 & n2925 ) | ( ~n2784 & n4119 ) | ( n2925 & n4119 ) ;
  assign n4121 = n2932 & n3507 ;
  assign n4122 = ( n2932 & n3483 ) | ( n2932 & n4121 ) | ( n3483 & n4121 ) ;
  assign n4123 = n4120 | n4122 ;
  assign n4124 = n4118 | n4123 ;
  assign n4125 = n2936 | n4124 ;
  assign n4126 = ( n3603 & n4124 ) | ( n3603 & n4125 ) | ( n4124 & n4125 ) ;
  assign n4127 = x23 & n4125 ;
  assign n4128 = x23 & n4124 ;
  assign n4129 = ( n3603 & n4127 ) | ( n3603 & n4128 ) | ( n4127 & n4128 ) ;
  assign n4130 = x23 & ~n4127 ;
  assign n4131 = x23 & ~n4128 ;
  assign n4132 = ( ~n3603 & n4130 ) | ( ~n3603 & n4131 ) | ( n4130 & n4131 ) ;
  assign n4133 = ( n4126 & ~n4129 ) | ( n4126 & n4132 ) | ( ~n4129 & n4132 ) ;
  assign n4134 = n4116 & n4133 ;
  assign n4135 = n4116 | n4133 ;
  assign n4136 = ~n4134 & n4135 ;
  assign n4137 = n2946 | n3272 ;
  assign n4138 = ( n2946 & ~n2949 ) | ( n2946 & n4137 ) | ( ~n2949 & n4137 ) ;
  assign n4139 = n4136 & n4138 ;
  assign n4140 = n4136 | n4138 ;
  assign n4141 = ~n4139 & n4140 ;
  assign n4221 = n3547 & n4206 ;
  assign n4222 = n3386 & n3544 ;
  assign n4223 = n3439 & n3541 ;
  assign n4224 = ( ~n3420 & n3541 ) | ( ~n3420 & n4223 ) | ( n3541 & n4223 ) ;
  assign n4225 = n4222 | n4224 ;
  assign n4226 = n4221 | n4225 ;
  assign n4227 = n3537 | n4221 ;
  assign n4228 = n4225 | n4227 ;
  assign n4229 = ( ~n4220 & n4226 ) | ( ~n4220 & n4228 ) | ( n4226 & n4228 ) ;
  assign n4230 = ~x20 & n4228 ;
  assign n4231 = ~x20 & n4226 ;
  assign n4232 = ( ~n4220 & n4230 ) | ( ~n4220 & n4231 ) | ( n4230 & n4231 ) ;
  assign n4233 = x20 | n4231 ;
  assign n4234 = x20 | n4230 ;
  assign n4235 = ( ~n4220 & n4233 ) | ( ~n4220 & n4234 ) | ( n4233 & n4234 ) ;
  assign n4236 = ( ~n4229 & n4232 ) | ( ~n4229 & n4235 ) | ( n4232 & n4235 ) ;
  assign n4237 = n4141 & n4236 ;
  assign n4238 = n4141 & ~n4237 ;
  assign n4239 = ~n4141 & n4236 ;
  assign n4240 = n4238 | n4239 ;
  assign n4241 = n3970 & n4240 ;
  assign n4242 = n3970 & ~n4241 ;
  assign n4243 = ~n3970 & n4240 ;
  assign n4244 = n4242 | n4243 ;
  assign n4467 = ~n4429 & n4466 ;
  assign n4469 = n4396 & n4468 ;
  assign n4470 = n4467 | n4469 ;
  assign n4472 = n4245 & n4471 ;
  assign n4473 = ( n4303 & n4471 ) | ( n4303 & n4472 ) | ( n4471 & n4472 ) ;
  assign n4474 = n4470 | n4473 ;
  assign n4476 = n4473 | n4475 ;
  assign n4477 = n4470 | n4476 ;
  assign n4478 = ( n4455 & n4474 ) | ( n4455 & n4477 ) | ( n4474 & n4477 ) ;
  assign n4479 = x17 & n4477 ;
  assign n4480 = x17 & n4474 ;
  assign n4481 = ( n4455 & n4479 ) | ( n4455 & n4480 ) | ( n4479 & n4480 ) ;
  assign n4482 = x17 & ~n4480 ;
  assign n4483 = x17 & ~n4479 ;
  assign n4484 = ( ~n4455 & n4482 ) | ( ~n4455 & n4483 ) | ( n4482 & n4483 ) ;
  assign n4485 = ( n4478 & ~n4481 ) | ( n4478 & n4484 ) | ( ~n4481 & n4484 ) ;
  assign n4486 = n4243 & n4485 ;
  assign n4487 = ( n4242 & n4485 ) | ( n4242 & n4486 ) | ( n4485 & n4486 ) ;
  assign n4488 = n4244 & ~n4487 ;
  assign n4489 = ~n4243 & n4485 ;
  assign n4490 = ~n4242 & n4489 ;
  assign n4491 = n4488 | n4490 ;
  assign n4998 = ~n4518 & n4997 ;
  assign n4999 = ( n4518 & n4995 ) | ( n4518 & ~n4998 ) | ( n4995 & ~n4998 ) ;
  assign n5000 = n4491 & n4999 ;
  assign n5001 = n4491 | n4999 ;
  assign n5002 = ~n5000 & n5001 ;
  assign n5038 = n134 | n616 ;
  assign n5039 = n207 | n5038 ;
  assign n5040 = n776 | n5039 ;
  assign n5041 = n53 | n841 ;
  assign n5042 = n966 | n5041 ;
  assign n5043 = n951 | n5042 ;
  assign n5044 = n5040 | n5043 ;
  assign n5045 = n3281 | n5044 ;
  assign n5046 = n259 | n4293 ;
  assign n5047 = n503 | n1662 ;
  assign n5048 = n5046 | n5047 ;
  assign n5049 = n388 | n5048 ;
  assign n5050 = n77 | n5049 ;
  assign n5051 = n5045 | n5050 ;
  assign n5052 = n451 | n588 ;
  assign n5053 = n2116 | n5052 ;
  assign n5054 = n477 | n959 ;
  assign n5055 = n214 | n5054 ;
  assign n5056 = n5053 | n5055 ;
  assign n5057 = n332 | n5056 ;
  assign n5058 = n196 | n527 ;
  assign n5059 = n705 | n5058 ;
  assign n5060 = n382 | n5059 ;
  assign n5061 = n1602 | n5060 ;
  assign n5062 = n5057 | n5061 ;
  assign n5063 = n937 | n4046 ;
  assign n5064 = n79 | n168 ;
  assign n5065 = n510 | n5064 ;
  assign n5066 = n5063 | n5065 ;
  assign n5067 = n209 | n476 ;
  assign n5068 = n302 | n5067 ;
  assign n5069 = n152 | n167 ;
  assign n5070 = n2874 | n5069 ;
  assign n5071 = n5068 | n5070 ;
  assign n5072 = n306 | n479 ;
  assign n5073 = n383 | n395 ;
  assign n5074 = n624 | n1114 ;
  assign n5075 = n5073 | n5074 ;
  assign n5076 = n5072 | n5075 ;
  assign n5077 = n5071 | n5076 ;
  assign n5078 = n5066 | n5077 ;
  assign n5079 = n5062 | n5078 ;
  assign n5080 = n5051 | n5079 ;
  assign n5081 = n445 | n496 ;
  assign n5082 = n387 | n643 ;
  assign n5083 = n222 | n5082 ;
  assign n5084 = n5081 | n5083 ;
  assign n5085 = n151 | n468 ;
  assign n5086 = n192 | n401 ;
  assign n5087 = n103 | n295 ;
  assign n5088 = n5086 | n5087 ;
  assign n5089 = n5085 | n5088 ;
  assign n5090 = n5084 | n5089 ;
  assign n5091 = n601 | n602 ;
  assign n5092 = n88 | n171 ;
  assign n5093 = n161 | n5092 ;
  assign n5094 = n5091 | n5093 ;
  assign n5095 = n5090 | n5094 ;
  assign n5096 = n533 | n1081 ;
  assign n5097 = n289 | n631 ;
  assign n5098 = n560 | n5097 ;
  assign n5099 = n5096 | n5098 ;
  assign n5100 = n75 | n5099 ;
  assign n5101 = n484 | n5100 ;
  assign n5102 = n5095 | n5101 ;
  assign n5103 = n282 | n1126 ;
  assign n5104 = n183 | n236 ;
  assign n5105 = n141 | n5104 ;
  assign n5106 = n5103 | n5105 ;
  assign n5107 = n5102 | n5106 ;
  assign n5108 = n5080 | n5107 ;
  assign n5118 = n5108 & n5117 ;
  assign n5119 = ( ~n5037 & n5108 ) | ( ~n5037 & n5118 ) | ( n5108 & n5118 ) ;
  assign n5120 = n5108 | n5117 ;
  assign n5121 = n5037 & ~n5120 ;
  assign n5122 = n5119 | n5121 ;
  assign n5204 = n5200 | n5203 ;
  assign n5205 = ~n5200 & n5202 ;
  assign n5206 = ( n5198 & n5204 ) | ( n5198 & ~n5205 ) | ( n5204 & ~n5205 ) ;
  assign n5211 = ( n5200 & ~n5205 ) | ( n5200 & n5210 ) | ( ~n5205 & n5210 ) ;
  assign n5212 = ( n4447 & n5206 ) | ( n4447 & n5211 ) | ( n5206 & n5211 ) ;
  assign n5213 = ~n5122 & n5212 ;
  assign n5214 = ( n4442 & n5206 ) | ( n4442 & n5211 ) | ( n5206 & n5211 ) ;
  assign n5215 = ~n5122 & n5214 ;
  assign n5216 = ( ~n3525 & n5213 ) | ( ~n3525 & n5215 ) | ( n5213 & n5215 ) ;
  assign n5217 = n5122 & ~n5212 ;
  assign n5218 = n5122 & ~n5214 ;
  assign n5219 = ( n3525 & n5217 ) | ( n3525 & n5218 ) | ( n5217 & n5218 ) ;
  assign n5220 = n5216 | n5219 ;
  assign n5232 = n5117 & n5231 ;
  assign n5233 = ( ~n5037 & n5231 ) | ( ~n5037 & n5232 ) | ( n5231 & n5232 ) ;
  assign n5235 = n5108 & n5234 ;
  assign n5238 = n5192 & n5237 ;
  assign n5239 = ( n5179 & n5237 ) | ( n5179 & n5238 ) | ( n5237 & n5238 ) ;
  assign n5240 = n5235 | n5239 ;
  assign n5241 = n5233 | n5240 ;
  assign n5242 = n5227 | n5241 ;
  assign n5243 = n5241 & n5242 ;
  assign n5244 = ( ~n5220 & n5242 ) | ( ~n5220 & n5243 ) | ( n5242 & n5243 ) ;
  assign n5245 = ~x14 & n5243 ;
  assign n5246 = ~x14 & n5242 ;
  assign n5247 = ( ~n5220 & n5245 ) | ( ~n5220 & n5246 ) | ( n5245 & n5246 ) ;
  assign n5248 = x14 | n5245 ;
  assign n5249 = x14 | n5246 ;
  assign n5250 = ( ~n5220 & n5248 ) | ( ~n5220 & n5249 ) | ( n5248 & n5249 ) ;
  assign n5251 = ( ~n5244 & n5247 ) | ( ~n5244 & n5250 ) | ( n5247 & n5250 ) ;
  assign n5252 = n5002 & n5251 ;
  assign n5253 = n5002 & ~n5252 ;
  assign n5254 = ~n5002 & n5251 ;
  assign n5255 = n5253 | n5254 ;
  assign n5853 = n5255 & n5852 ;
  assign n5854 = n5852 & ~n5853 ;
  assign n5855 = n5255 & ~n5853 ;
  assign n5856 = n5854 | n5855 ;
  assign n5857 = n263 | n568 ;
  assign n5858 = n224 | n1482 ;
  assign n5859 = n1713 | n5858 ;
  assign n5860 = n320 | n1172 ;
  assign n5861 = n2066 | n3467 ;
  assign n5862 = n5860 | n5861 ;
  assign n5863 = n5859 | n5862 ;
  assign n5864 = n357 | n4197 ;
  assign n5865 = n177 | n1166 ;
  assign n5866 = n5864 | n5865 ;
  assign n5867 = n901 | n938 ;
  assign n5868 = n139 | n372 ;
  assign n5869 = n5867 | n5868 ;
  assign n5870 = n126 | n468 ;
  assign n5871 = n5869 | n5870 ;
  assign n5872 = n5866 | n5871 ;
  assign n5873 = n5863 | n5872 ;
  assign n5874 = n758 | n5873 ;
  assign n5875 = n446 | n452 ;
  assign n5876 = n59 | n291 ;
  assign n5877 = n305 | n5876 ;
  assign n5878 = n143 & ~n675 ;
  assign n5879 = ~n601 & n5878 ;
  assign n5880 = ~n5877 & n5879 ;
  assign n5881 = ~n230 & n5880 ;
  assign n5882 = ~n5875 & n5881 ;
  assign n5883 = n173 | n185 ;
  assign n5884 = n166 | n5883 ;
  assign n5885 = n5882 & ~n5884 ;
  assign n5886 = ~n3999 & n5885 ;
  assign n5887 = ~n5874 & n5886 ;
  assign n5888 = n2115 | n2122 ;
  assign n5889 = n290 | n1240 ;
  assign n5890 = n460 | n888 ;
  assign n5891 = n5889 | n5890 ;
  assign n5892 = n249 | n2050 ;
  assign n5893 = n1251 | n5892 ;
  assign n5894 = n5891 | n5893 ;
  assign n5895 = n1171 | n2233 ;
  assign n5896 = n416 | n5895 ;
  assign n5897 = n5894 | n5896 ;
  assign n5898 = n5888 | n5897 ;
  assign n5899 = n5887 & ~n5898 ;
  assign n5900 = ~n5857 & n5899 ;
  assign n5901 = n284 | n489 ;
  assign n5902 = n995 | n5901 ;
  assign n5903 = n112 | n331 ;
  assign n5904 = n320 | n5903 ;
  assign n5905 = n5902 | n5904 ;
  assign n5906 = n182 | n206 ;
  assign n5907 = n5905 | n5906 ;
  assign n5908 = n381 | n775 ;
  assign n5909 = n4249 | n5908 ;
  assign n5910 = n958 | n5909 ;
  assign n5911 = n85 | n608 ;
  assign n5912 = n340 | n689 ;
  assign n5913 = n5911 | n5912 ;
  assign n5914 = n208 | n616 ;
  assign n5915 = n555 | n5914 ;
  assign n5916 = n5913 | n5915 ;
  assign n5917 = n5910 | n5916 ;
  assign n5918 = n5907 | n5917 ;
  assign n5919 = n1479 | n5918 ;
  assign n5920 = n223 | n476 ;
  assign n5921 = n2156 | n5920 ;
  assign n5922 = n443 | n5921 ;
  assign n5923 = n77 | n887 ;
  assign n5924 = n1643 | n5923 ;
  assign n5925 = n5922 | n5924 ;
  assign n5926 = n386 | n1636 ;
  assign n5927 = n5925 | n5926 ;
  assign n5928 = n159 | n198 ;
  assign n5929 = n979 | n5928 ;
  assign n5930 = n236 | n987 ;
  assign n5931 = n5929 | n5930 ;
  assign n5932 = n139 | n370 ;
  assign n5933 = n2129 | n5932 ;
  assign n5934 = n5931 | n5933 ;
  assign n5935 = n1521 | n1631 ;
  assign n5936 = n1016 | n2233 ;
  assign n5937 = n5935 | n5936 ;
  assign n5938 = n128 | n399 ;
  assign n5939 = n5937 | n5938 ;
  assign n5940 = n5934 | n5939 ;
  assign n5941 = n5927 | n5940 ;
  assign n5942 = n5919 | n5941 ;
  assign n5943 = n292 | n510 ;
  assign n5944 = n190 | n325 ;
  assign n5945 = n5943 | n5944 ;
  assign n5946 = n103 | n305 ;
  assign n5947 = n138 | n302 ;
  assign n5948 = n5946 | n5947 ;
  assign n5949 = n757 | n2204 ;
  assign n5950 = n5948 | n5949 ;
  assign n5951 = n5945 | n5950 ;
  assign n5952 = n214 | n1172 ;
  assign n5953 = n1615 | n5952 ;
  assign n5954 = n356 | n566 ;
  assign n5955 = n312 | n5954 ;
  assign n5956 = n5953 | n5955 ;
  assign n5957 = n4046 | n5956 ;
  assign n5958 = n5951 | n5957 ;
  assign n5959 = n679 | n5958 ;
  assign n5960 = n280 | n354 ;
  assign n5961 = n2665 | n5960 ;
  assign n5962 = n375 | n5961 ;
  assign n5963 = n1742 | n3312 ;
  assign n5964 = n588 | n5963 ;
  assign n5965 = n5962 | n5964 ;
  assign n5966 = n483 | n959 ;
  assign n5967 = n176 | n291 ;
  assign n5968 = n5966 | n5967 ;
  assign n5969 = n255 | n5968 ;
  assign n5970 = n432 | n5969 ;
  assign n5971 = n5965 | n5970 ;
  assign n5972 = n1035 | n1607 ;
  assign n5973 = n591 | n952 ;
  assign n5974 = n5972 | n5973 ;
  assign n5975 = n154 | n725 ;
  assign n5976 = n5974 | n5975 ;
  assign n5977 = n5971 | n5976 ;
  assign n5978 = n5959 | n5977 ;
  assign n5979 = n5942 | n5978 ;
  assign n5980 = n295 | n560 ;
  assign n5981 = n500 | n5980 ;
  assign n5982 = n192 | n696 ;
  assign n5983 = n162 | n841 ;
  assign n5984 = n504 | n5983 ;
  assign n5985 = n2653 | n5984 ;
  assign n5986 = n246 | n667 ;
  assign n5987 = n222 | n631 ;
  assign n5988 = n5986 | n5987 ;
  assign n5989 = n321 | n402 ;
  assign n5990 = n184 | n347 ;
  assign n5991 = n5989 | n5990 ;
  assign n5992 = n5988 | n5991 ;
  assign n5993 = n5985 | n5992 ;
  assign n5994 = n311 | n480 ;
  assign n5995 = n5993 | n5994 ;
  assign n5996 = n5982 | n5995 ;
  assign n5997 = n5981 | n5996 ;
  assign n5998 = n5979 | n5997 ;
  assign n5999 = ~n5900 & n5998 ;
  assign n6000 = n5900 & ~n5998 ;
  assign n6001 = n5999 | n6000 ;
  assign n6002 = n5108 & n5998 ;
  assign n6003 = n5108 | n5998 ;
  assign n6004 = ~n6002 & n6003 ;
  assign n6005 = n5119 | n6002 ;
  assign n6006 = ( n6002 & n6004 ) | ( n6002 & n6005 ) | ( n6004 & n6005 ) ;
  assign n6007 = ~n6001 & n6006 ;
  assign n6008 = n175 | n178 ;
  assign n6009 = n2875 | n6008 ;
  assign n6010 = n852 | n3412 ;
  assign n6011 = n760 | n6010 ;
  assign n6012 = n6009 | n6011 ;
  assign n6013 = n986 | n1650 ;
  assign n6014 = n226 | n292 ;
  assign n6015 = n2188 | n6014 ;
  assign n6016 = n6013 | n6015 ;
  assign n6017 = n6012 | n6016 ;
  assign n6018 = n357 | n411 ;
  assign n6019 = n1030 | n1675 ;
  assign n6020 = n6018 | n6019 ;
  assign n6021 = n319 | n6020 ;
  assign n6022 = n103 | n189 ;
  assign n6023 = n104 | n517 ;
  assign n6024 = n6022 | n6023 ;
  assign n6025 = n254 | n500 ;
  assign n6026 = n6024 | n6025 ;
  assign n6027 = n6021 | n6026 ;
  assign n6028 = n6017 | n6027 ;
  assign n6029 = n249 | n631 ;
  assign n6030 = n384 | n503 ;
  assign n6031 = n6029 | n6030 ;
  assign n6032 = n2215 | n6031 ;
  assign n6033 = n155 | n450 ;
  assign n6034 = n1035 | n6033 ;
  assign n6035 = n6032 | n6034 ;
  assign n6036 = n419 | n966 ;
  assign n6037 = n234 | n1172 ;
  assign n6038 = n6036 | n6037 ;
  assign n6039 = n2710 | n6038 ;
  assign n6040 = n6035 | n6039 ;
  assign n6041 = n313 | n458 ;
  assign n6042 = n666 | n6041 ;
  assign n6043 = n377 | n6042 ;
  assign n6044 = n160 | n325 ;
  assign n6045 = n143 & ~n250 ;
  assign n6046 = ~n6044 & n6045 ;
  assign n6047 = ~n212 & n6046 ;
  assign n6048 = ~n6043 & n6047 ;
  assign n6049 = ~n1657 & n6048 ;
  assign n6050 = ~n6040 & n6049 ;
  assign n6051 = ~n6028 & n6050 ;
  assign n6052 = n171 | n193 ;
  assign n6053 = n302 | n332 ;
  assign n6054 = n6052 | n6053 ;
  assign n6055 = n261 | n539 ;
  assign n6056 = n6054 | n6055 ;
  assign n6057 = n154 | n196 ;
  assign n6058 = n245 | n6057 ;
  assign n6059 = n85 | n959 ;
  assign n6060 = n92 | n801 ;
  assign n6061 = n6059 | n6060 ;
  assign n6062 = n6058 | n6061 ;
  assign n6063 = n6056 | n6062 ;
  assign n6064 = n123 | n388 ;
  assign n6065 = n3296 | n6064 ;
  assign n6066 = n497 | n6065 ;
  assign n6067 = n279 | n645 ;
  assign n6068 = n1250 | n6067 ;
  assign n6069 = n6066 | n6068 ;
  assign n6070 = n6063 | n6069 ;
  assign n6071 = n139 | n607 ;
  assign n6072 = n142 | n689 ;
  assign n6073 = n6071 | n6072 ;
  assign n6074 = n184 | n6073 ;
  assign n6075 = n364 | n938 ;
  assign n6076 = n550 | n6075 ;
  assign n6077 = n162 | n441 ;
  assign n6078 = n134 | n6077 ;
  assign n6079 = n6076 | n6078 ;
  assign n6080 = n6074 | n6079 ;
  assign n6081 = n6070 | n6080 ;
  assign n6082 = n821 | n1126 ;
  assign n6083 = n83 | n289 ;
  assign n6084 = n444 | n6083 ;
  assign n6085 = n6082 | n6084 ;
  assign n6086 = n96 | n183 ;
  assign n6087 = n281 | n6086 ;
  assign n6088 = n675 | n6087 ;
  assign n6089 = n6085 | n6088 ;
  assign n6090 = n6081 | n6089 ;
  assign n6091 = n6051 & ~n6090 ;
  assign n6092 = n5857 & ~n6091 ;
  assign n6093 = ( n5899 & n6091 ) | ( n5899 & ~n6092 ) | ( n6091 & ~n6092 ) ;
  assign n6094 = ~n5857 & n6091 ;
  assign n6095 = n5899 & n6094 ;
  assign n6096 = n6093 & ~n6095 ;
  assign n6097 = n5999 & n6096 ;
  assign n6098 = ( n6007 & n6096 ) | ( n6007 & n6097 ) | ( n6096 & n6097 ) ;
  assign n6099 = n6002 | n6004 ;
  assign n6100 = ~n6001 & n6099 ;
  assign n6101 = ( n6096 & n6097 ) | ( n6096 & n6100 ) | ( n6097 & n6100 ) ;
  assign n6102 = ( n5216 & n6098 ) | ( n5216 & n6101 ) | ( n6098 & n6101 ) ;
  assign n6103 = n5999 | n6100 ;
  assign n6104 = n6096 | n6103 ;
  assign n6105 = n5999 | n6007 ;
  assign n6106 = n6096 | n6105 ;
  assign n6107 = ( n5216 & n6104 ) | ( n5216 & n6106 ) | ( n6104 & n6106 ) ;
  assign n6108 = ~n6102 & n6107 ;
  assign n6112 = x8 & ~x9 ;
  assign n6113 = ~x8 & x9 ;
  assign n6114 = n6112 | n6113 ;
  assign n6116 = ~x9 & x10 ;
  assign n6117 = x9 & ~x10 ;
  assign n6118 = n6116 | n6117 ;
  assign n6119 = ~n6114 & n6118 ;
  assign n6120 = n5857 & n6119 ;
  assign n6121 = ( ~n5899 & n6119 ) | ( ~n5899 & n6120 ) | ( n6119 & n6120 ) ;
  assign n6109 = x10 & ~x11 ;
  assign n6110 = ~x10 & x11 ;
  assign n6111 = n6109 | n6110 ;
  assign n6122 = ~n6111 & n6114 ;
  assign n6123 = ~n6091 & n6122 ;
  assign n6124 = n6111 & ~n6114 ;
  assign n6125 = ~n6118 & n6124 ;
  assign n6126 = n5997 & n6125 ;
  assign n6127 = ( n5979 & n6125 ) | ( n5979 & n6126 ) | ( n6125 & n6126 ) ;
  assign n6128 = n6123 | n6127 ;
  assign n6129 = n6121 | n6128 ;
  assign n6115 = n6111 & n6114 ;
  assign n6130 = n6115 | n6129 ;
  assign n6131 = ( n6108 & n6129 ) | ( n6108 & n6130 ) | ( n6129 & n6130 ) ;
  assign n6132 = x11 & n6130 ;
  assign n6133 = x11 & n6129 ;
  assign n6134 = ( n6108 & n6132 ) | ( n6108 & n6133 ) | ( n6132 & n6133 ) ;
  assign n6135 = x11 & ~n6132 ;
  assign n6136 = x11 & ~n6133 ;
  assign n6137 = ( ~n6108 & n6135 ) | ( ~n6108 & n6136 ) | ( n6135 & n6136 ) ;
  assign n6138 = ( n6131 & ~n6134 ) | ( n6131 & n6137 ) | ( ~n6134 & n6137 ) ;
  assign n6139 = n5856 & n6138 ;
  assign n6140 = n5856 & ~n6139 ;
  assign n6141 = ~n5856 & n6138 ;
  assign n6142 = n6140 | n6141 ;
  assign n6143 = n5847 & ~n5850 ;
  assign n6144 = n5847 & ~n6143 ;
  assign n6147 = ( n5216 & n6007 ) | ( n5216 & n6100 ) | ( n6007 & n6100 ) ;
  assign n6148 = n6001 & ~n6006 ;
  assign n6149 = n6001 & ~n6099 ;
  assign n6150 = ( ~n5216 & n6148 ) | ( ~n5216 & n6149 ) | ( n6148 & n6149 ) ;
  assign n6151 = n6147 | n6150 ;
  assign n6152 = n5108 & n6125 ;
  assign n6153 = n5997 & n6119 ;
  assign n6154 = ( n5979 & n6119 ) | ( n5979 & n6153 ) | ( n6119 & n6153 ) ;
  assign n6155 = n6152 | n6154 ;
  assign n6156 = n5857 & n6122 ;
  assign n6157 = ( ~n5899 & n6122 ) | ( ~n5899 & n6156 ) | ( n6122 & n6156 ) ;
  assign n6158 = n6155 | n6157 ;
  assign n6159 = n6115 | n6158 ;
  assign n6160 = ( ~n6151 & n6158 ) | ( ~n6151 & n6159 ) | ( n6158 & n6159 ) ;
  assign n6161 = ~x11 & n6159 ;
  assign n6162 = ~x11 & n6158 ;
  assign n6163 = ( ~n6151 & n6161 ) | ( ~n6151 & n6162 ) | ( n6161 & n6162 ) ;
  assign n6164 = x11 | n6161 ;
  assign n6165 = x11 | n6162 ;
  assign n6166 = ( ~n6151 & n6164 ) | ( ~n6151 & n6165 ) | ( n6164 & n6165 ) ;
  assign n6167 = ( ~n6160 & n6163 ) | ( ~n6160 & n6166 ) | ( n6163 & n6166 ) ;
  assign n6145 = n5847 | n5850 ;
  assign n6168 = ~n6145 & n6167 ;
  assign n6169 = ( n6144 & n6167 ) | ( n6144 & n6168 ) | ( n6167 & n6168 ) ;
  assign n6146 = ~n6144 & n6145 ;
  assign n6170 = n6146 | n6169 ;
  assign n6171 = n6145 & n6167 ;
  assign n6172 = ~n6144 & n6171 ;
  assign n6173 = n6170 & ~n6172 ;
  assign n6174 = ~n5328 & n5845 ;
  assign n6175 = n5328 & ~n5845 ;
  assign n6176 = n6174 | n6175 ;
  assign n6177 = n5119 & n6004 ;
  assign n6178 = ( n5216 & n6004 ) | ( n5216 & n6177 ) | ( n6004 & n6177 ) ;
  assign n6179 = n5119 | n6004 ;
  assign n6180 = n5216 | n6179 ;
  assign n6181 = ~n6178 & n6180 ;
  assign n6182 = n5117 & n6125 ;
  assign n6183 = ( ~n5037 & n6125 ) | ( ~n5037 & n6182 ) | ( n6125 & n6182 ) ;
  assign n6184 = n5108 & n6119 ;
  assign n6185 = n5997 & n6122 ;
  assign n6186 = ( n5979 & n6122 ) | ( n5979 & n6185 ) | ( n6122 & n6185 ) ;
  assign n6187 = n6184 | n6186 ;
  assign n6188 = n6183 | n6187 ;
  assign n6189 = n6115 | n6188 ;
  assign n6190 = ( n6181 & n6188 ) | ( n6181 & n6189 ) | ( n6188 & n6189 ) ;
  assign n6191 = x11 & n6189 ;
  assign n6192 = x11 & n6188 ;
  assign n6193 = ( n6181 & n6191 ) | ( n6181 & n6192 ) | ( n6191 & n6192 ) ;
  assign n6194 = x11 & ~n6191 ;
  assign n6195 = x11 & ~n6192 ;
  assign n6196 = ( ~n6181 & n6194 ) | ( ~n6181 & n6195 ) | ( n6194 & n6195 ) ;
  assign n6197 = ( n6190 & ~n6193 ) | ( n6190 & n6196 ) | ( ~n6193 & n6196 ) ;
  assign n6198 = n6176 & n6197 ;
  assign n6199 = n6176 | n6197 ;
  assign n6200 = ~n6198 & n6199 ;
  assign n6201 = n5352 & n5843 ;
  assign n6202 = n5352 | n5843 ;
  assign n6203 = ~n6201 & n6202 ;
  assign n6204 = n5117 & n6119 ;
  assign n6205 = ( ~n5037 & n6119 ) | ( ~n5037 & n6204 ) | ( n6119 & n6204 ) ;
  assign n6206 = n5108 & n6122 ;
  assign n6207 = n5192 & n6125 ;
  assign n6208 = ( n5179 & n6125 ) | ( n5179 & n6207 ) | ( n6125 & n6207 ) ;
  assign n6209 = n6206 | n6208 ;
  assign n6210 = n6205 | n6209 ;
  assign n6211 = n6115 | n6210 ;
  assign n6212 = ( ~n5220 & n6210 ) | ( ~n5220 & n6211 ) | ( n6210 & n6211 ) ;
  assign n6213 = ~x11 & n6211 ;
  assign n6214 = ~x11 & n6210 ;
  assign n6215 = ( ~n5220 & n6213 ) | ( ~n5220 & n6214 ) | ( n6213 & n6214 ) ;
  assign n6216 = x11 | n6213 ;
  assign n6217 = x11 | n6214 ;
  assign n6218 = ( ~n5220 & n6216 ) | ( ~n5220 & n6217 ) | ( n6216 & n6217 ) ;
  assign n6219 = ( ~n6212 & n6215 ) | ( ~n6212 & n6218 ) | ( n6215 & n6218 ) ;
  assign n6220 = ~n6203 & n6219 ;
  assign n6221 = n6203 & ~n6219 ;
  assign n6222 = n6220 | n6221 ;
  assign n6223 = n5376 & n5841 ;
  assign n6224 = n5376 | n5841 ;
  assign n6225 = ~n6223 & n6224 ;
  assign n6226 = n4245 & n6125 ;
  assign n6227 = ( n4303 & n6125 ) | ( n4303 & n6226 ) | ( n6125 & n6226 ) ;
  assign n6228 = n5192 & n6119 ;
  assign n6229 = ( n5179 & n6119 ) | ( n5179 & n6228 ) | ( n6119 & n6228 ) ;
  assign n6230 = n6227 | n6229 ;
  assign n6231 = n5117 & n6122 ;
  assign n6232 = ( ~n5037 & n6122 ) | ( ~n5037 & n6231 ) | ( n6122 & n6231 ) ;
  assign n6233 = n6230 | n6232 ;
  assign n6234 = n6115 | n6232 ;
  assign n6235 = n6230 | n6234 ;
  assign n6236 = ( ~n5270 & n6233 ) | ( ~n5270 & n6235 ) | ( n6233 & n6235 ) ;
  assign n6237 = ~x11 & n6235 ;
  assign n6238 = ~x11 & n6233 ;
  assign n6239 = ( ~n5270 & n6237 ) | ( ~n5270 & n6238 ) | ( n6237 & n6238 ) ;
  assign n6240 = x11 | n6238 ;
  assign n6241 = x11 | n6237 ;
  assign n6242 = ( ~n5270 & n6240 ) | ( ~n5270 & n6241 ) | ( n6240 & n6241 ) ;
  assign n6243 = ( ~n6236 & n6239 ) | ( ~n6236 & n6242 ) | ( n6239 & n6242 ) ;
  assign n6244 = ~n6225 & n6243 ;
  assign n6245 = n6225 & ~n6243 ;
  assign n6246 = n6244 | n6245 ;
  assign n6247 = ~n5399 & n5839 ;
  assign n6248 = n5399 & ~n5839 ;
  assign n6249 = n6247 | n6248 ;
  assign n6250 = n4396 & n6125 ;
  assign n6251 = n4245 & n6119 ;
  assign n6252 = ( n4303 & n6119 ) | ( n4303 & n6251 ) | ( n6119 & n6251 ) ;
  assign n6253 = n6250 | n6252 ;
  assign n6254 = n5192 & n6122 ;
  assign n6255 = ( n5179 & n6122 ) | ( n5179 & n6254 ) | ( n6122 & n6254 ) ;
  assign n6256 = n6253 | n6255 ;
  assign n6257 = n6115 | n6255 ;
  assign n6258 = n6253 | n6257 ;
  assign n6259 = ( n5306 & n6256 ) | ( n5306 & n6258 ) | ( n6256 & n6258 ) ;
  assign n6260 = x11 & n6258 ;
  assign n6261 = x11 & n6256 ;
  assign n6262 = ( n5306 & n6260 ) | ( n5306 & n6261 ) | ( n6260 & n6261 ) ;
  assign n6263 = x11 & ~n6261 ;
  assign n6264 = x11 & ~n6260 ;
  assign n6265 = ( ~n5306 & n6263 ) | ( ~n5306 & n6264 ) | ( n6263 & n6264 ) ;
  assign n6266 = ( n6259 & ~n6262 ) | ( n6259 & n6265 ) | ( ~n6262 & n6265 ) ;
  assign n6267 = n6249 & n6266 ;
  assign n6268 = n5440 | n5836 ;
  assign n6269 = n5834 | n6268 ;
  assign n6270 = ~n5838 & n6269 ;
  assign n6271 = ~n4429 & n6125 ;
  assign n6272 = n4396 & n6119 ;
  assign n6273 = n6271 | n6272 ;
  assign n6274 = n4245 & n6122 ;
  assign n6275 = ( n4303 & n6122 ) | ( n4303 & n6274 ) | ( n6122 & n6274 ) ;
  assign n6277 = n6115 | n6275 ;
  assign n6278 = n6273 | n6277 ;
  assign n6276 = n6273 | n6275 ;
  assign n6279 = n6276 & n6278 ;
  assign n6280 = ( n4455 & n6278 ) | ( n4455 & n6279 ) | ( n6278 & n6279 ) ;
  assign n6281 = x11 & n6279 ;
  assign n6282 = x11 & n6278 ;
  assign n6283 = ( n4455 & n6281 ) | ( n4455 & n6282 ) | ( n6281 & n6282 ) ;
  assign n6284 = x11 & ~n6281 ;
  assign n6285 = x11 & ~n6282 ;
  assign n6286 = ( ~n4455 & n6284 ) | ( ~n4455 & n6285 ) | ( n6284 & n6285 ) ;
  assign n6287 = ( n6280 & ~n6283 ) | ( n6280 & n6286 ) | ( ~n6283 & n6286 ) ;
  assign n6288 = n6270 & n6287 ;
  assign n6289 = n6270 | n6287 ;
  assign n6290 = ~n6288 & n6289 ;
  assign n6291 = n5443 | n5833 ;
  assign n6292 = ~n5834 & n6291 ;
  assign n6293 = ~n4429 & n6119 ;
  assign n6294 = n6119 | n6125 ;
  assign n6295 = ( ~n4429 & n6125 ) | ( ~n4429 & n6294 ) | ( n6125 & n6294 ) ;
  assign n6296 = ( n4206 & n6293 ) | ( n4206 & n6295 ) | ( n6293 & n6295 ) ;
  assign n6297 = n4396 & n6122 ;
  assign n6299 = n6115 | n6297 ;
  assign n6300 = n6296 | n6299 ;
  assign n6298 = n6296 | n6297 ;
  assign n6301 = n6298 & n6300 ;
  assign n6302 = ( ~n4501 & n6300 ) | ( ~n4501 & n6301 ) | ( n6300 & n6301 ) ;
  assign n6303 = ~x11 & n6301 ;
  assign n6304 = ~x11 & n6300 ;
  assign n6305 = ( ~n4501 & n6303 ) | ( ~n4501 & n6304 ) | ( n6303 & n6304 ) ;
  assign n6306 = x11 | n6303 ;
  assign n6307 = x11 | n6304 ;
  assign n6308 = ( ~n4501 & n6306 ) | ( ~n4501 & n6307 ) | ( n6306 & n6307 ) ;
  assign n6309 = ( ~n6302 & n6305 ) | ( ~n6302 & n6308 ) | ( n6305 & n6308 ) ;
  assign n6310 = n6292 & n6309 ;
  assign n6311 = n6292 & ~n6310 ;
  assign n6312 = ~n6292 & n6309 ;
  assign n6313 = n6311 | n6312 ;
  assign n6314 = n5824 | n5830 ;
  assign n6315 = n5828 | n6314 ;
  assign n6316 = ~n5832 & n6315 ;
  assign n6317 = n4206 & n6119 ;
  assign n6318 = ~n4429 & n6122 ;
  assign n6319 = n3439 & n6125 ;
  assign n6320 = ( ~n3420 & n6125 ) | ( ~n3420 & n6319 ) | ( n6125 & n6319 ) ;
  assign n6321 = n6318 | n6320 ;
  assign n6322 = n6317 | n6321 ;
  assign n6323 = n6115 | n6317 ;
  assign n6324 = n6321 | n6323 ;
  assign n6325 = ( ~n4527 & n6322 ) | ( ~n4527 & n6324 ) | ( n6322 & n6324 ) ;
  assign n6326 = ~x11 & n6324 ;
  assign n6327 = ~x11 & n6322 ;
  assign n6328 = ( ~n4527 & n6326 ) | ( ~n4527 & n6327 ) | ( n6326 & n6327 ) ;
  assign n6329 = x11 | n6327 ;
  assign n6330 = x11 | n6326 ;
  assign n6331 = ( ~n4527 & n6329 ) | ( ~n4527 & n6330 ) | ( n6329 & n6330 ) ;
  assign n6332 = ( ~n6325 & n6328 ) | ( ~n6325 & n6331 ) | ( n6328 & n6331 ) ;
  assign n6333 = n6316 & n6332 ;
  assign n6334 = n5827 & ~n5828 ;
  assign n6335 = n5802 & ~n5827 ;
  assign n6336 = n6334 | n6335 ;
  assign n6337 = n4206 & n6122 ;
  assign n6338 = n3386 & n6125 ;
  assign n6339 = n3439 & n6119 ;
  assign n6340 = ( ~n3420 & n6119 ) | ( ~n3420 & n6339 ) | ( n6119 & n6339 ) ;
  assign n6341 = n6338 | n6340 ;
  assign n6342 = n6337 | n6341 ;
  assign n6343 = n6115 | n6337 ;
  assign n6344 = n6341 | n6343 ;
  assign n6345 = ( ~n4220 & n6342 ) | ( ~n4220 & n6344 ) | ( n6342 & n6344 ) ;
  assign n6346 = ~x11 & n6344 ;
  assign n6347 = ~x11 & n6342 ;
  assign n6348 = ( ~n4220 & n6346 ) | ( ~n4220 & n6347 ) | ( n6346 & n6347 ) ;
  assign n6349 = x11 | n6347 ;
  assign n6350 = x11 | n6346 ;
  assign n6351 = ( ~n4220 & n6349 ) | ( ~n4220 & n6350 ) | ( n6349 & n6350 ) ;
  assign n6352 = ( ~n6345 & n6348 ) | ( ~n6345 & n6351 ) | ( n6348 & n6351 ) ;
  assign n6353 = n6335 & n6352 ;
  assign n6354 = ( n6334 & n6352 ) | ( n6334 & n6353 ) | ( n6352 & n6353 ) ;
  assign n6355 = n6336 & ~n6354 ;
  assign n6356 = ~n6335 & n6352 ;
  assign n6357 = ~n6334 & n6356 ;
  assign n6358 = n6355 | n6357 ;
  assign n6359 = n5800 & ~n5801 ;
  assign n6360 = n5489 & ~n5801 ;
  assign n6361 = n6359 | n6360 ;
  assign n6362 = n3386 & n6119 ;
  assign n6363 = n3507 & n6125 ;
  assign n6364 = ( n3483 & n6125 ) | ( n3483 & n6363 ) | ( n6125 & n6363 ) ;
  assign n6365 = n3439 & n6122 ;
  assign n6366 = ( ~n3420 & n6122 ) | ( ~n3420 & n6365 ) | ( n6122 & n6365 ) ;
  assign n6367 = n6364 | n6366 ;
  assign n6368 = n6362 | n6367 ;
  assign n6369 = n6115 | n6368 ;
  assign n6370 = ( ~n3530 & n6368 ) | ( ~n3530 & n6369 ) | ( n6368 & n6369 ) ;
  assign n6371 = ~x11 & n6369 ;
  assign n6372 = ~x11 & n6368 ;
  assign n6373 = ( ~n3530 & n6371 ) | ( ~n3530 & n6372 ) | ( n6371 & n6372 ) ;
  assign n6374 = x11 | n6371 ;
  assign n6375 = x11 | n6372 ;
  assign n6376 = ( ~n3530 & n6374 ) | ( ~n3530 & n6375 ) | ( n6374 & n6375 ) ;
  assign n6377 = ( ~n6370 & n6373 ) | ( ~n6370 & n6376 ) | ( n6373 & n6376 ) ;
  assign n6378 = n6361 & n6377 ;
  assign n6379 = n6361 & ~n6378 ;
  assign n6380 = ~n6361 & n6377 ;
  assign n6381 = n6379 | n6380 ;
  assign n6382 = n5796 & n5798 ;
  assign n6383 = n5796 | n5798 ;
  assign n6384 = ~n6382 & n6383 ;
  assign n6385 = n2893 & n6125 ;
  assign n6386 = ( ~n2886 & n6125 ) | ( ~n2886 & n6385 ) | ( n6125 & n6385 ) ;
  assign n6387 = n3507 & n6119 ;
  assign n6388 = ( n3483 & n6119 ) | ( n3483 & n6387 ) | ( n6119 & n6387 ) ;
  assign n6389 = n6386 | n6388 ;
  assign n6390 = n3386 & n6122 ;
  assign n6392 = n6115 | n6390 ;
  assign n6393 = n6389 | n6392 ;
  assign n6391 = n6389 | n6390 ;
  assign n6394 = n6391 & n6393 ;
  assign n6395 = ( ~n3568 & n6393 ) | ( ~n3568 & n6394 ) | ( n6393 & n6394 ) ;
  assign n6396 = ~x11 & n6394 ;
  assign n6397 = ~x11 & n6393 ;
  assign n6398 = ( ~n3568 & n6396 ) | ( ~n3568 & n6397 ) | ( n6396 & n6397 ) ;
  assign n6399 = x11 | n6396 ;
  assign n6400 = x11 | n6397 ;
  assign n6401 = ( ~n3568 & n6399 ) | ( ~n3568 & n6400 ) | ( n6399 & n6400 ) ;
  assign n6402 = ( ~n6395 & n6398 ) | ( ~n6395 & n6401 ) | ( n6398 & n6401 ) ;
  assign n6403 = n6384 & n6402 ;
  assign n6404 = n5559 | n5792 ;
  assign n6405 = ~n5793 & n6404 ;
  assign n6406 = n2691 & n6125 ;
  assign n6407 = ( n2678 & n6125 ) | ( n2678 & n6406 ) | ( n6125 & n6406 ) ;
  assign n6408 = n2701 & n6119 ;
  assign n6409 = ( ~n2784 & n6119 ) | ( ~n2784 & n6408 ) | ( n6119 & n6408 ) ;
  assign n6410 = n6407 | n6409 ;
  assign n6411 = n2893 & n6122 ;
  assign n6412 = ( ~n2886 & n6122 ) | ( ~n2886 & n6411 ) | ( n6122 & n6411 ) ;
  assign n6413 = n6410 | n6412 ;
  assign n6414 = n6115 | n6413 ;
  assign n6415 = n6413 & n6414 ;
  assign n6416 = ( ~n2914 & n6414 ) | ( ~n2914 & n6415 ) | ( n6414 & n6415 ) ;
  assign n6417 = ~x11 & n6415 ;
  assign n6418 = ~x11 & n6414 ;
  assign n6419 = ( ~n2914 & n6417 ) | ( ~n2914 & n6418 ) | ( n6417 & n6418 ) ;
  assign n6420 = x11 | n6417 ;
  assign n6421 = x11 | n6418 ;
  assign n6422 = ( ~n2914 & n6420 ) | ( ~n2914 & n6421 ) | ( n6420 & n6421 ) ;
  assign n6423 = ( ~n6416 & n6419 ) | ( ~n6416 & n6422 ) | ( n6419 & n6422 ) ;
  assign n6424 = n6405 & n6423 ;
  assign n6425 = n6405 & ~n6424 ;
  assign n6426 = ~n6405 & n6423 ;
  assign n6427 = n6425 | n6426 ;
  assign n6428 = n5788 & n5790 ;
  assign n6429 = n5788 | n5790 ;
  assign n6430 = ~n6428 & n6429 ;
  assign n6431 = n2701 & n6122 ;
  assign n6432 = ( ~n2784 & n6122 ) | ( ~n2784 & n6431 ) | ( n6122 & n6431 ) ;
  assign n6433 = n2691 & n6119 ;
  assign n6434 = ( n2678 & n6119 ) | ( n2678 & n6433 ) | ( n6119 & n6433 ) ;
  assign n6435 = n6432 | n6434 ;
  assign n6436 = n2199 & n6125 ;
  assign n6437 = ( ~n2185 & n6125 ) | ( ~n2185 & n6436 ) | ( n6125 & n6436 ) ;
  assign n6438 = n6435 | n6437 ;
  assign n6439 = n6115 | n6437 ;
  assign n6440 = n6435 | n6439 ;
  assign n6441 = ( n2960 & n6438 ) | ( n2960 & n6440 ) | ( n6438 & n6440 ) ;
  assign n6442 = x11 & n6440 ;
  assign n6443 = x11 & n6438 ;
  assign n6444 = ( n2960 & n6442 ) | ( n2960 & n6443 ) | ( n6442 & n6443 ) ;
  assign n6445 = x11 & ~n6443 ;
  assign n6446 = x11 & ~n6442 ;
  assign n6447 = ( ~n2960 & n6445 ) | ( ~n2960 & n6446 ) | ( n6445 & n6446 ) ;
  assign n6448 = ( n6441 & ~n6444 ) | ( n6441 & n6447 ) | ( ~n6444 & n6447 ) ;
  assign n6449 = n6430 & n6448 ;
  assign n6450 = n5783 & n5786 ;
  assign n6451 = n5783 & ~n6450 ;
  assign n6454 = n2090 & n6125 ;
  assign n6455 = ( ~n2082 & n6125 ) | ( ~n2082 & n6454 ) | ( n6125 & n6454 ) ;
  assign n6456 = n2691 & n6122 ;
  assign n6457 = ( n2678 & n6122 ) | ( n2678 & n6456 ) | ( n6122 & n6456 ) ;
  assign n6458 = n2199 & n6119 ;
  assign n6459 = ( ~n2185 & n6119 ) | ( ~n2185 & n6458 ) | ( n6119 & n6458 ) ;
  assign n6460 = n6457 | n6459 ;
  assign n6461 = n6455 | n6460 ;
  assign n6462 = n6115 | n6461 ;
  assign n6463 = ( n2985 & n6461 ) | ( n2985 & n6462 ) | ( n6461 & n6462 ) ;
  assign n6464 = x11 & n6462 ;
  assign n6465 = x11 & n6461 ;
  assign n6466 = ( n2985 & n6464 ) | ( n2985 & n6465 ) | ( n6464 & n6465 ) ;
  assign n6467 = x11 & ~n6464 ;
  assign n6468 = x11 & ~n6465 ;
  assign n6469 = ( ~n2985 & n6467 ) | ( ~n2985 & n6468 ) | ( n6467 & n6468 ) ;
  assign n6470 = ( n6463 & ~n6466 ) | ( n6463 & n6469 ) | ( ~n6466 & n6469 ) ;
  assign n6452 = ~n5783 & n5786 ;
  assign n6471 = n6452 & n6470 ;
  assign n6472 = ( n6451 & n6470 ) | ( n6451 & n6471 ) | ( n6470 & n6471 ) ;
  assign n6453 = n6451 | n6452 ;
  assign n6473 = n6453 & ~n6472 ;
  assign n6474 = ~n6452 & n6470 ;
  assign n6475 = ~n6451 & n6474 ;
  assign n6476 = n6473 | n6475 ;
  assign n6477 = ~n5778 & n5781 ;
  assign n6478 = n5778 & ~n5781 ;
  assign n6479 = n6477 | n6478 ;
  assign n6480 = n2090 & n6119 ;
  assign n6481 = ( ~n2082 & n6119 ) | ( ~n2082 & n6480 ) | ( n6119 & n6480 ) ;
  assign n6482 = n2279 & n6125 ;
  assign n6483 = ( ~n2269 & n6125 ) | ( ~n2269 & n6482 ) | ( n6125 & n6482 ) ;
  assign n6484 = n2199 & n6122 ;
  assign n6485 = ( ~n2185 & n6122 ) | ( ~n2185 & n6484 ) | ( n6122 & n6484 ) ;
  assign n6486 = n6483 | n6485 ;
  assign n6487 = n6481 | n6486 ;
  assign n6488 = n6115 | n6487 ;
  assign n6489 = ( ~n2325 & n6487 ) | ( ~n2325 & n6488 ) | ( n6487 & n6488 ) ;
  assign n6490 = n6487 & n6488 ;
  assign n6491 = ( ~n2299 & n6489 ) | ( ~n2299 & n6490 ) | ( n6489 & n6490 ) ;
  assign n6492 = ~x11 & n6491 ;
  assign n6493 = x11 | n6491 ;
  assign n6494 = ( ~n6491 & n6492 ) | ( ~n6491 & n6493 ) | ( n6492 & n6493 ) ;
  assign n6495 = n6479 & n6494 ;
  assign n6496 = n6479 | n6494 ;
  assign n6497 = ~n6495 & n6496 ;
  assign n6498 = n5774 | n5776 ;
  assign n6499 = ~n5777 & n6498 ;
  assign n6500 = n1634 & n6125 ;
  assign n6501 = ( n1630 & n6125 ) | ( n1630 & n6500 ) | ( n6125 & n6500 ) ;
  assign n6502 = n2279 & n6119 ;
  assign n6503 = ( ~n2269 & n6119 ) | ( ~n2269 & n6502 ) | ( n6119 & n6502 ) ;
  assign n6504 = n6501 | n6503 ;
  assign n6505 = n2090 & n6122 ;
  assign n6506 = ( ~n2082 & n6122 ) | ( ~n2082 & n6505 ) | ( n6122 & n6505 ) ;
  assign n6507 = n6504 | n6506 ;
  assign n6508 = n6115 | n6507 ;
  assign n6509 = n6507 & n6508 ;
  assign n6510 = ( n2568 & n6508 ) | ( n2568 & n6509 ) | ( n6508 & n6509 ) ;
  assign n6511 = x11 & n6509 ;
  assign n6512 = x11 & n6508 ;
  assign n6513 = ( n2568 & n6511 ) | ( n2568 & n6512 ) | ( n6511 & n6512 ) ;
  assign n6514 = x11 & ~n6511 ;
  assign n6515 = x11 & ~n6512 ;
  assign n6516 = ( ~n2568 & n6514 ) | ( ~n2568 & n6515 ) | ( n6514 & n6515 ) ;
  assign n6517 = ( n6510 & ~n6513 ) | ( n6510 & n6516 ) | ( ~n6513 & n6516 ) ;
  assign n6518 = n6499 & n6517 ;
  assign n6519 = n5664 | n5772 ;
  assign n6520 = ~n5773 & n6519 ;
  assign n6521 = n1708 & n6125 ;
  assign n6522 = n1634 & n6119 ;
  assign n6523 = ( n1630 & n6119 ) | ( n1630 & n6522 ) | ( n6119 & n6522 ) ;
  assign n6524 = n2279 & n6122 ;
  assign n6525 = ( ~n2269 & n6122 ) | ( ~n2269 & n6524 ) | ( n6122 & n6524 ) ;
  assign n6526 = n6523 | n6525 ;
  assign n6527 = n6521 | n6526 ;
  assign n6528 = n6115 | n6527 ;
  assign n6529 = n6527 & n6528 ;
  assign n6530 = ( ~n2343 & n6528 ) | ( ~n2343 & n6529 ) | ( n6528 & n6529 ) ;
  assign n6531 = ~x11 & n6529 ;
  assign n6532 = ~x11 & n6528 ;
  assign n6533 = ( ~n2343 & n6531 ) | ( ~n2343 & n6532 ) | ( n6531 & n6532 ) ;
  assign n6534 = x11 | n6531 ;
  assign n6535 = x11 | n6532 ;
  assign n6536 = ( ~n2343 & n6534 ) | ( ~n2343 & n6535 ) | ( n6534 & n6535 ) ;
  assign n6537 = ( ~n6530 & n6533 ) | ( ~n6530 & n6536 ) | ( n6533 & n6536 ) ;
  assign n6538 = n6520 & n6537 ;
  assign n6539 = n5768 & n5770 ;
  assign n6540 = n5768 | n5770 ;
  assign n6541 = ~n6539 & n6540 ;
  assign n6542 = n1708 & n6119 ;
  assign n6543 = n1793 & n6125 ;
  assign n6544 = ( n1783 & n6125 ) | ( n1783 & n6543 ) | ( n6125 & n6543 ) ;
  assign n6545 = n1634 & n6122 ;
  assign n6546 = ( n1630 & n6122 ) | ( n1630 & n6545 ) | ( n6122 & n6545 ) ;
  assign n6547 = n6544 | n6546 ;
  assign n6548 = n6542 | n6547 ;
  assign n6549 = n6115 | n6548 ;
  assign n6550 = n6548 & n6549 ;
  assign n6551 = ( n1814 & n6549 ) | ( n1814 & n6550 ) | ( n6549 & n6550 ) ;
  assign n6552 = x11 & n6550 ;
  assign n6553 = x11 & n6549 ;
  assign n6554 = ( n1814 & n6552 ) | ( n1814 & n6553 ) | ( n6552 & n6553 ) ;
  assign n6555 = x11 & ~n6552 ;
  assign n6556 = x11 & ~n6553 ;
  assign n6557 = ( ~n1814 & n6555 ) | ( ~n1814 & n6556 ) | ( n6555 & n6556 ) ;
  assign n6558 = ( n6551 & ~n6554 ) | ( n6551 & n6557 ) | ( ~n6554 & n6557 ) ;
  assign n6559 = n6541 & n6558 ;
  assign n6560 = n5764 & n5766 ;
  assign n6561 = n5764 | n5766 ;
  assign n6562 = ~n6560 & n6561 ;
  assign n6563 = ~n523 & n6125 ;
  assign n6564 = n1793 & n6119 ;
  assign n6565 = ( n1783 & n6119 ) | ( n1783 & n6564 ) | ( n6119 & n6564 ) ;
  assign n6566 = n6563 | n6565 ;
  assign n6567 = n1708 & n6122 ;
  assign n6568 = n6566 | n6567 ;
  assign n6569 = n6115 | n6567 ;
  assign n6570 = n6566 | n6569 ;
  assign n6571 = ( ~n1852 & n6568 ) | ( ~n1852 & n6570 ) | ( n6568 & n6570 ) ;
  assign n6572 = ~x11 & n6570 ;
  assign n6573 = ~x11 & n6568 ;
  assign n6574 = ( ~n1852 & n6572 ) | ( ~n1852 & n6573 ) | ( n6572 & n6573 ) ;
  assign n6575 = x11 | n6573 ;
  assign n6576 = x11 | n6572 ;
  assign n6577 = ( ~n1852 & n6575 ) | ( ~n1852 & n6576 ) | ( n6575 & n6576 ) ;
  assign n6578 = ( ~n6571 & n6574 ) | ( ~n6571 & n6577 ) | ( n6574 & n6577 ) ;
  assign n6579 = n6562 & n6578 ;
  assign n6580 = n5760 | n5761 ;
  assign n6581 = n5744 | n6580 ;
  assign n6582 = ~n5763 & n6581 ;
  assign n6583 = ~n523 & n6119 ;
  assign n6584 = n352 & n6125 ;
  assign n6585 = ( ~n339 & n6125 ) | ( ~n339 & n6584 ) | ( n6125 & n6584 ) ;
  assign n6586 = n1793 & n6122 ;
  assign n6587 = ( n1783 & n6122 ) | ( n1783 & n6586 ) | ( n6122 & n6586 ) ;
  assign n6588 = n6585 | n6587 ;
  assign n6589 = n6583 | n6588 ;
  assign n6590 = n6115 | n6589 ;
  assign n6591 = n6589 & n6590 ;
  assign n6592 = ( n1884 & n6590 ) | ( n1884 & n6591 ) | ( n6590 & n6591 ) ;
  assign n6593 = x11 & n6591 ;
  assign n6594 = x11 & n6590 ;
  assign n6595 = ( n1884 & n6593 ) | ( n1884 & n6594 ) | ( n6593 & n6594 ) ;
  assign n6596 = x11 & ~n6593 ;
  assign n6597 = x11 & ~n6594 ;
  assign n6598 = ( ~n1884 & n6596 ) | ( ~n1884 & n6597 ) | ( n6596 & n6597 ) ;
  assign n6599 = ( n6592 & ~n6595 ) | ( n6592 & n6598 ) | ( ~n6595 & n6598 ) ;
  assign n6600 = n6582 & n6599 ;
  assign n6601 = n6582 | n6599 ;
  assign n6602 = ~n6600 & n6601 ;
  assign n6603 = ~n829 & n6125 ;
  assign n6604 = n352 & n6119 ;
  assign n6605 = ( ~n339 & n6119 ) | ( ~n339 & n6604 ) | ( n6119 & n6604 ) ;
  assign n6606 = n6603 | n6605 ;
  assign n6607 = ~n523 & n6122 ;
  assign n6608 = n6115 | n6607 ;
  assign n6609 = n6606 | n6608 ;
  assign n6610 = ~x11 & n6609 ;
  assign n6611 = n6606 | n6607 ;
  assign n6612 = ~x11 & n6611 ;
  assign n6613 = ( ~n1055 & n6610 ) | ( ~n1055 & n6612 ) | ( n6610 & n6612 ) ;
  assign n6614 = x11 & n6609 ;
  assign n6615 = x11 & ~n6614 ;
  assign n6616 = x11 & n6607 ;
  assign n6617 = ( x11 & n6606 ) | ( x11 & n6616 ) | ( n6606 & n6616 ) ;
  assign n6618 = x11 & ~n6617 ;
  assign n6619 = ( n1055 & n6615 ) | ( n1055 & n6618 ) | ( n6615 & n6618 ) ;
  assign n6620 = n6613 | n6619 ;
  assign n6621 = n5737 | n5739 ;
  assign n6622 = x14 & ~n5737 ;
  assign n6623 = ( n5720 & n6621 ) | ( n5720 & ~n6622 ) | ( n6621 & ~n6622 ) ;
  assign n6624 = ~n5742 & n6623 ;
  assign n6625 = n6620 & n6624 ;
  assign n6626 = x14 | n5734 ;
  assign n6627 = ( ~n5727 & n5734 ) | ( ~n5727 & n6626 ) | ( n5734 & n6626 ) ;
  assign n6628 = n5728 | n6627 ;
  assign n6629 = ~n5737 & n6628 ;
  assign n6630 = ~n829 & n6119 ;
  assign n6631 = n352 & n6122 ;
  assign n6632 = ( ~n339 & n6122 ) | ( ~n339 & n6631 ) | ( n6122 & n6631 ) ;
  assign n6633 = n6630 | n6632 ;
  assign n6634 = n692 & n6125 ;
  assign n6635 = ( n674 & n6125 ) | ( n674 & n6634 ) | ( n6125 & n6634 ) ;
  assign n6636 = n6633 | n6635 ;
  assign n6637 = n6115 | n6635 ;
  assign n6638 = n6633 | n6637 ;
  assign n6639 = ( ~n1209 & n6636 ) | ( ~n1209 & n6638 ) | ( n6636 & n6638 ) ;
  assign n6640 = ~x11 & n6638 ;
  assign n6641 = ~x11 & n6636 ;
  assign n6642 = ( ~n1209 & n6640 ) | ( ~n1209 & n6641 ) | ( n6640 & n6641 ) ;
  assign n6643 = x11 | n6641 ;
  assign n6644 = x11 | n6640 ;
  assign n6645 = ( ~n1209 & n6643 ) | ( ~n1209 & n6644 ) | ( n6643 & n6644 ) ;
  assign n6646 = ( ~n6639 & n6642 ) | ( ~n6639 & n6645 ) | ( n6642 & n6645 ) ;
  assign n6647 = n6629 & n6646 ;
  assign n6648 = ( ~n1027 & n5730 ) | ( ~n1027 & n5732 ) | ( n5730 & n5732 ) ;
  assign n6649 = ~n922 & n6119 ;
  assign n6650 = n1042 & n6125 ;
  assign n6651 = ( ~n1027 & n6125 ) | ( ~n1027 & n6650 ) | ( n6125 & n6650 ) ;
  assign n6652 = n6649 | n6651 ;
  assign n6653 = n692 & n6122 ;
  assign n6654 = ( n674 & n6122 ) | ( n674 & n6653 ) | ( n6122 & n6653 ) ;
  assign n6655 = n6652 | n6654 ;
  assign n6656 = ( n1538 & n6115 ) | ( n1538 & n6655 ) | ( n6115 & n6655 ) ;
  assign n6657 = ( x11 & ~n6655 ) | ( x11 & n6656 ) | ( ~n6655 & n6656 ) ;
  assign n6658 = ~n6656 & n6657 ;
  assign n6659 = ~n922 & n6122 ;
  assign n6660 = n1042 & n6119 ;
  assign n6661 = ( ~n1027 & n6119 ) | ( ~n1027 & n6660 ) | ( n6119 & n6660 ) ;
  assign n6662 = n6659 | n6661 ;
  assign n6663 = n6115 | n6661 ;
  assign n6664 = n6659 | n6663 ;
  assign n6665 = ( n1946 & n6662 ) | ( n1946 & n6664 ) | ( n6662 & n6664 ) ;
  assign n6666 = ~x11 & n6665 ;
  assign n6667 = n139 & n6114 ;
  assign n6668 = ( n1041 & n6114 ) | ( n1041 & n6667 ) | ( n6114 & n6667 ) ;
  assign n6669 = x11 & ~n6668 ;
  assign n6670 = n6114 | n6667 ;
  assign n6671 = x11 & ~n6670 ;
  assign n6672 = ( n1027 & n6669 ) | ( n1027 & n6671 ) | ( n6669 & n6671 ) ;
  assign n6673 = x11 & n6672 ;
  assign n6674 = ~n6665 & n6673 ;
  assign n6675 = ( n6666 & n6672 ) | ( n6666 & n6674 ) | ( n6672 & n6674 ) ;
  assign n6676 = x11 | n6655 ;
  assign n6677 = n6656 | n6676 ;
  assign n6678 = n6675 & n6677 ;
  assign n6679 = ~x11 & n6675 ;
  assign n6680 = ( n6658 & n6678 ) | ( n6658 & n6679 ) | ( n6678 & n6679 ) ;
  assign n6681 = n6648 & n6680 ;
  assign n6682 = n6680 & ~n6681 ;
  assign n6683 = ~n829 & n6122 ;
  assign n6684 = ~n922 & n6125 ;
  assign n6685 = n6683 | n6684 ;
  assign n6686 = n692 & n6119 ;
  assign n6687 = ( n674 & n6119 ) | ( n674 & n6686 ) | ( n6119 & n6686 ) ;
  assign n6688 = n6685 | n6687 ;
  assign n6689 = n6115 | n6687 ;
  assign n6690 = n6685 | n6689 ;
  assign n6691 = ( n1554 & n6688 ) | ( n1554 & n6690 ) | ( n6688 & n6690 ) ;
  assign n6692 = x11 & n6690 ;
  assign n6693 = x11 & n6688 ;
  assign n6694 = ( n1554 & n6692 ) | ( n1554 & n6693 ) | ( n6692 & n6693 ) ;
  assign n6695 = x11 & ~n6693 ;
  assign n6696 = x11 & ~n6692 ;
  assign n6697 = ( ~n1554 & n6695 ) | ( ~n1554 & n6696 ) | ( n6695 & n6696 ) ;
  assign n6698 = ( n6691 & ~n6694 ) | ( n6691 & n6697 ) | ( ~n6694 & n6697 ) ;
  assign n6699 = n6648 & ~n6680 ;
  assign n6700 = n6698 & n6699 ;
  assign n6701 = ( n6682 & n6698 ) | ( n6682 & n6700 ) | ( n6698 & n6700 ) ;
  assign n6702 = n6681 | n6701 ;
  assign n6703 = n6629 | n6646 ;
  assign n6704 = ~n6647 & n6703 ;
  assign n6705 = n6647 | n6704 ;
  assign n6706 = ( n6647 & n6702 ) | ( n6647 & n6705 ) | ( n6702 & n6705 ) ;
  assign n6707 = n6620 | n6624 ;
  assign n6708 = ~n6625 & n6707 ;
  assign n6709 = n6625 | n6708 ;
  assign n6710 = ( n6625 & n6706 ) | ( n6625 & n6709 ) | ( n6706 & n6709 ) ;
  assign n6711 = n6602 & n6710 ;
  assign n6712 = n6600 | n6711 ;
  assign n6713 = ~n6562 & n6578 ;
  assign n6714 = ( n6562 & ~n6579 ) | ( n6562 & n6713 ) | ( ~n6579 & n6713 ) ;
  assign n6715 = n6712 & n6714 ;
  assign n6716 = n6579 | n6715 ;
  assign n6717 = n6541 & ~n6559 ;
  assign n6718 = ~n6541 & n6558 ;
  assign n6719 = n6717 | n6718 ;
  assign n6720 = n6716 & n6719 ;
  assign n6721 = n6559 | n6720 ;
  assign n6722 = n6520 & ~n6538 ;
  assign n6723 = ~n6520 & n6537 ;
  assign n6724 = n6722 | n6723 ;
  assign n6725 = n6538 | n6724 ;
  assign n6726 = ( n6538 & n6721 ) | ( n6538 & n6725 ) | ( n6721 & n6725 ) ;
  assign n6727 = n6499 | n6517 ;
  assign n6728 = ~n6518 & n6727 ;
  assign n6729 = n6518 | n6728 ;
  assign n6730 = ( n6518 & n6726 ) | ( n6518 & n6729 ) | ( n6726 & n6729 ) ;
  assign n6731 = n6497 & n6730 ;
  assign n6732 = n6495 | n6731 ;
  assign n6733 = n6472 | n6732 ;
  assign n6734 = ( n6472 & n6476 ) | ( n6472 & n6733 ) | ( n6476 & n6733 ) ;
  assign n6735 = ~n6430 & n6448 ;
  assign n6736 = ( n6430 & ~n6449 ) | ( n6430 & n6735 ) | ( ~n6449 & n6735 ) ;
  assign n6737 = n6449 | n6736 ;
  assign n6738 = ( n6449 & n6734 ) | ( n6449 & n6737 ) | ( n6734 & n6737 ) ;
  assign n6739 = n6427 & n6738 ;
  assign n6740 = n6424 | n6739 ;
  assign n6741 = n5538 & n5794 ;
  assign n6742 = n5538 | n5794 ;
  assign n6743 = ~n6741 & n6742 ;
  assign n6744 = n2893 & n6119 ;
  assign n6745 = ( ~n2886 & n6119 ) | ( ~n2886 & n6744 ) | ( n6119 & n6744 ) ;
  assign n6746 = n2701 & n6125 ;
  assign n6747 = ( ~n2784 & n6125 ) | ( ~n2784 & n6746 ) | ( n6125 & n6746 ) ;
  assign n6748 = n3507 & n6122 ;
  assign n6749 = ( n3483 & n6122 ) | ( n3483 & n6748 ) | ( n6122 & n6748 ) ;
  assign n6750 = n6747 | n6749 ;
  assign n6751 = n6745 | n6750 ;
  assign n6752 = n6115 | n6751 ;
  assign n6753 = n6751 & n6752 ;
  assign n6754 = ( n3603 & n6752 ) | ( n3603 & n6753 ) | ( n6752 & n6753 ) ;
  assign n6755 = x11 & n6753 ;
  assign n6756 = x11 & n6752 ;
  assign n6757 = ( n3603 & n6755 ) | ( n3603 & n6756 ) | ( n6755 & n6756 ) ;
  assign n6758 = x11 & ~n6755 ;
  assign n6759 = x11 & ~n6756 ;
  assign n6760 = ( ~n3603 & n6758 ) | ( ~n3603 & n6759 ) | ( n6758 & n6759 ) ;
  assign n6761 = ( n6754 & ~n6757 ) | ( n6754 & n6760 ) | ( ~n6757 & n6760 ) ;
  assign n6762 = n6743 & n6761 ;
  assign n6763 = n6743 & ~n6762 ;
  assign n6764 = ~n6743 & n6761 ;
  assign n6765 = n6763 | n6764 ;
  assign n6766 = n6740 & n6765 ;
  assign n6767 = n6384 | n6402 ;
  assign n6768 = ~n6403 & n6767 ;
  assign n6769 = n6762 & n6768 ;
  assign n6770 = ( n6766 & n6768 ) | ( n6766 & n6769 ) | ( n6768 & n6769 ) ;
  assign n6771 = n6403 | n6770 ;
  assign n6772 = n6381 & n6771 ;
  assign n6773 = n6378 | n6772 ;
  assign n6774 = n6358 & n6773 ;
  assign n6775 = ~n6316 & n6332 ;
  assign n6776 = ( n6316 & ~n6333 ) | ( n6316 & n6775 ) | ( ~n6333 & n6775 ) ;
  assign n6777 = n6354 & n6776 ;
  assign n6778 = ( n6774 & n6776 ) | ( n6774 & n6777 ) | ( n6776 & n6777 ) ;
  assign n6779 = n6333 | n6778 ;
  assign n6780 = n6313 & n6779 ;
  assign n6781 = n6290 & n6310 ;
  assign n6782 = ( n6290 & n6780 ) | ( n6290 & n6781 ) | ( n6780 & n6781 ) ;
  assign n6783 = n6288 | n6782 ;
  assign n6784 = n6249 | n6266 ;
  assign n6785 = ~n6267 & n6784 ;
  assign n6786 = n6267 | n6785 ;
  assign n6787 = ( n6267 & n6783 ) | ( n6267 & n6786 ) | ( n6783 & n6786 ) ;
  assign n6788 = ~n6246 & n6787 ;
  assign n6789 = n6244 | n6788 ;
  assign n6790 = ~n6222 & n6789 ;
  assign n6791 = n6220 | n6790 ;
  assign n6792 = n6200 & n6791 ;
  assign n6793 = n6198 | n6792 ;
  assign n6794 = n6169 | n6793 ;
  assign n6795 = ( n6169 & ~n6173 ) | ( n6169 & n6794 ) | ( ~n6173 & n6794 ) ;
  assign n6796 = n6142 & n6795 ;
  assign n6797 = n6142 | n6795 ;
  assign n6798 = ~n6796 & n6797 ;
  assign n6799 = n1464 | n4000 ;
  assign n6800 = n126 | n229 ;
  assign n6801 = n5946 | n6800 ;
  assign n6802 = n3393 | n6801 ;
  assign n6803 = n6799 | n6802 ;
  assign n6804 = n2248 | n6803 ;
  assign n6805 = n457 | n648 ;
  assign n6806 = n923 | n6805 ;
  assign n6807 = n456 | n6806 ;
  assign n6808 = n224 | n2743 ;
  assign n6809 = n261 | n1282 ;
  assign n6810 = n6808 | n6809 ;
  assign n6811 = n309 | n370 ;
  assign n6812 = n363 | n6811 ;
  assign n6813 = n6810 | n6812 ;
  assign n6814 = n6807 | n6813 ;
  assign n6815 = n6804 | n6814 ;
  assign n6816 = n551 | n1394 ;
  assign n6817 = n274 | n710 ;
  assign n6818 = n6816 | n6817 ;
  assign n6819 = n249 | n313 ;
  assign n6820 = n6818 | n6819 ;
  assign n6821 = n6815 | n6820 ;
  assign n6822 = n450 | n469 ;
  assign n6823 = n1303 | n6822 ;
  assign n6824 = n240 | n6823 ;
  assign n6825 = n123 | n297 ;
  assign n6826 = n71 | n6825 ;
  assign n6827 = n142 | n263 ;
  assign n6828 = n6826 | n6827 ;
  assign n6829 = n6824 | n6828 ;
  assign n6830 = n1301 | n5058 ;
  assign n6831 = n118 | n302 ;
  assign n6832 = n431 | n6831 ;
  assign n6833 = n6830 | n6832 ;
  assign n6834 = n354 | n405 ;
  assign n6835 = n6833 | n6834 ;
  assign n6836 = n6829 | n6835 ;
  assign n6837 = n340 | n369 ;
  assign n6838 = n193 | n206 ;
  assign n6839 = n6837 | n6838 ;
  assign n6840 = n6836 | n6839 ;
  assign n6841 = n6821 | n6840 ;
  assign n6842 = n53 | n806 ;
  assign n6843 = n210 | n6842 ;
  assign n6844 = n341 | n6843 ;
  assign n6845 = n702 | n1465 ;
  assign n6846 = n205 | n6845 ;
  assign n6847 = n143 & ~n588 ;
  assign n6848 = ~n159 & n6847 ;
  assign n6849 = n1127 | n1719 ;
  assign n6850 = n6848 & ~n6849 ;
  assign n6851 = ~n6846 & n6850 ;
  assign n6852 = ~n6844 & n6851 ;
  assign n6853 = n476 | n1039 ;
  assign n6854 = n364 | n375 ;
  assign n6855 = n6853 | n6854 ;
  assign n6856 = n461 | n510 ;
  assign n6857 = n344 | n6856 ;
  assign n6858 = n6855 | n6857 ;
  assign n6859 = n281 | n306 ;
  assign n6860 = n5860 | n6859 ;
  assign n6861 = n6858 | n6860 ;
  assign n6862 = n288 | n317 ;
  assign n6863 = n190 | n312 ;
  assign n6864 = n6862 | n6863 ;
  assign n6865 = n154 | n577 ;
  assign n6866 = n6864 | n6865 ;
  assign n6867 = n6861 | n6866 ;
  assign n6868 = n6852 & ~n6867 ;
  assign n6869 = ~n1002 & n6868 ;
  assign n6870 = n138 | n477 ;
  assign n6871 = n250 | n6870 ;
  assign n6872 = n69 | n6871 ;
  assign n6873 = n406 | n483 ;
  assign n6874 = n1136 | n6873 ;
  assign n6875 = n131 | n152 ;
  assign n6876 = n5014 | n6875 ;
  assign n6877 = n6874 | n6876 ;
  assign n6878 = n6872 | n6877 ;
  assign n6879 = n1031 | n3986 ;
  assign n6880 = n1479 | n6879 ;
  assign n6881 = n1304 | n6880 ;
  assign n6882 = n6878 | n6881 ;
  assign n6883 = n6869 & ~n6882 ;
  assign n6884 = ~n6841 & n6883 ;
  assign n6885 = n292 | n748 ;
  assign n6886 = n566 | n5182 ;
  assign n6887 = n6885 | n6886 ;
  assign n6888 = n212 | n348 ;
  assign n6889 = n6887 | n6888 ;
  assign n6890 = n6884 & ~n6889 ;
  assign n6891 = n375 | n578 ;
  assign n6892 = n2023 | n6891 ;
  assign n6893 = n1639 | n6892 ;
  assign n6894 = n257 | n284 ;
  assign n6895 = n444 | n465 ;
  assign n6896 = n6894 | n6895 ;
  assign n6897 = n237 | n304 ;
  assign n6898 = n6896 | n6897 ;
  assign n6899 = n292 | n344 ;
  assign n6900 = n476 | n501 ;
  assign n6901 = n6899 | n6900 ;
  assign n6902 = ( ~n156 & n6898 ) | ( ~n156 & n6901 ) | ( n6898 & n6901 ) ;
  assign n6903 = n156 & ~n6901 ;
  assign n6904 = ( n6893 & n6902 ) | ( n6893 & ~n6903 ) | ( n6902 & ~n6903 ) ;
  assign n6905 = n156 | n6904 ;
  assign n6906 = n83 | n806 ;
  assign n6907 = n1251 | n6906 ;
  assign n6908 = n270 | n3501 ;
  assign n6909 = n6907 | n6908 ;
  assign n6910 = n395 | n6909 ;
  assign n6911 = n414 | n2748 ;
  assign n6912 = n405 | n503 ;
  assign n6913 = n443 | n6912 ;
  assign n6914 = n6911 | n6913 ;
  assign n6915 = n103 | n321 ;
  assign n6916 = n1385 | n6915 ;
  assign n6917 = n2167 | n6916 ;
  assign n6918 = n6914 | n6917 ;
  assign n6919 = n6910 | n6918 ;
  assign n6920 = n2801 | n6919 ;
  assign n6921 = n6905 | n6920 ;
  assign n6922 = n5888 | n6921 ;
  assign n6923 = n178 | n349 ;
  assign n6924 = n159 | n600 ;
  assign n6925 = n6923 | n6924 ;
  assign n6926 = n225 | n6925 ;
  assign n6927 = n1283 | n2128 ;
  assign n6928 = n6926 | n6927 ;
  assign n6929 = n118 | n3376 ;
  assign n6930 = n1501 | n6929 ;
  assign n6931 = n6928 | n6930 ;
  assign n6932 = n511 | n735 ;
  assign n6933 = n2192 | n6932 ;
  assign n6934 = n296 | n1035 ;
  assign n6935 = n6933 | n6934 ;
  assign n6936 = n163 | n6935 ;
  assign n6937 = n513 | n6936 ;
  assign n6938 = n6931 | n6937 ;
  assign n6939 = n114 | n288 ;
  assign n6940 = n6938 | n6939 ;
  assign n6941 = n176 | n638 ;
  assign n6942 = n236 | n313 ;
  assign n6943 = n6941 | n6942 ;
  assign n6944 = n306 | n694 ;
  assign n6945 = n263 | n6944 ;
  assign n6946 = n6943 | n6945 ;
  assign n6947 = n245 | n254 ;
  assign n6948 = n6946 | n6947 ;
  assign n6949 = n6940 | n6948 ;
  assign n6950 = n6922 | n6949 ;
  assign n6951 = ~n6890 & n6950 ;
  assign n6952 = n6890 & ~n6950 ;
  assign n6953 = n6951 | n6952 ;
  assign n6954 = n2215 | n5983 ;
  assign n6955 = n441 | n1301 ;
  assign n6956 = n6954 | n6955 ;
  assign n6957 = n117 | n465 ;
  assign n6958 = n193 | n623 ;
  assign n6959 = n6957 | n6958 ;
  assign n6960 = n6956 | n6959 ;
  assign n6961 = n4170 | n5133 ;
  assign n6962 = n1222 | n1499 ;
  assign n6963 = n6961 | n6962 ;
  assign n6964 = n6960 | n6963 ;
  assign n6965 = n411 | n5860 ;
  assign n6966 = n317 | n3430 ;
  assign n6967 = n6965 | n6966 ;
  assign n6968 = n79 | n233 ;
  assign n6969 = n6967 | n6968 ;
  assign n6970 = n5090 | n6969 ;
  assign n6971 = n6964 | n6970 ;
  assign n6972 = n67 | n255 ;
  assign n6973 = n1124 | n6972 ;
  assign n6974 = n1115 | n6973 ;
  assign n6975 = n64 | n959 ;
  assign n6976 = n644 | n6975 ;
  assign n6977 = n407 | n6976 ;
  assign n6978 = n6974 | n6977 ;
  assign n6979 = n514 | n775 ;
  assign n6980 = n305 | n6979 ;
  assign n6981 = n412 | n6980 ;
  assign n6982 = n303 | n6981 ;
  assign n6983 = n6978 | n6982 ;
  assign n6984 = n6971 | n6983 ;
  assign n6985 = n402 | n511 ;
  assign n6986 = n5006 | n6985 ;
  assign n6987 = n138 | n437 ;
  assign n6988 = n952 | n6987 ;
  assign n6989 = n777 | n6988 ;
  assign n6990 = n6986 | n6989 ;
  assign n6991 = n160 | n858 ;
  assign n6992 = n2235 | n6991 ;
  assign n6993 = n1081 | n1742 ;
  assign n6994 = n2651 | n6993 ;
  assign n6995 = n6992 | n6994 ;
  assign n6996 = n6990 | n6995 ;
  assign n6997 = n1447 | n4410 ;
  assign n6998 = n262 | n638 ;
  assign n6999 = n226 | n6998 ;
  assign n7000 = n6997 | n6999 ;
  assign n7001 = n324 | n513 ;
  assign n7002 = n4246 | n5092 ;
  assign n7003 = n7001 | n7002 ;
  assign n7004 = n7000 | n7003 ;
  assign n7005 = n2051 | n4249 ;
  assign n7006 = n168 | n696 ;
  assign n7007 = n272 | n7006 ;
  assign n7008 = n7005 | n7007 ;
  assign n7009 = n7004 | n7008 ;
  assign n7010 = n6996 | n7009 ;
  assign n7011 = n159 | n356 ;
  assign n7012 = n99 | n390 ;
  assign n7013 = n617 | n7012 ;
  assign n7014 = n7011 | n7013 ;
  assign n7015 = n131 | n249 ;
  assign n7016 = n155 | n7015 ;
  assign n7017 = n5923 | n7016 ;
  assign n7018 = n7014 | n7017 ;
  assign n7019 = n1436 | n5945 ;
  assign n7020 = n555 | n7019 ;
  assign n7021 = n7018 | n7020 ;
  assign n7022 = n7010 | n7021 ;
  assign n7023 = n6984 | n7022 ;
  assign n7024 = n75 | n126 ;
  assign n7025 = n489 | n591 ;
  assign n7026 = n7024 | n7025 ;
  assign n7027 = n250 | n363 ;
  assign n7028 = n476 | n7027 ;
  assign n7029 = n7026 | n7028 ;
  assign n7030 = n1394 | n2666 ;
  assign n7031 = n7029 | n7030 ;
  assign n7032 = n484 | n3445 ;
  assign n7033 = n163 | n7032 ;
  assign n7034 = n310 | n7033 ;
  assign n7035 = n7031 | n7034 ;
  assign n7036 = n675 | n7035 ;
  assign n7037 = n7023 | n7036 ;
  assign n7038 = n6950 & n7037 ;
  assign n7039 = ~n6953 & n7038 ;
  assign n7040 = n6950 | n7037 ;
  assign n7041 = ~n7038 & n7040 ;
  assign n7042 = ~n6091 & n7037 ;
  assign n7043 = n6093 & ~n6097 ;
  assign n7044 = n6093 & ~n6096 ;
  assign n7045 = ( ~n6007 & n7043 ) | ( ~n6007 & n7044 ) | ( n7043 & n7044 ) ;
  assign n7046 = n6091 & ~n7037 ;
  assign n7047 = n7042 | n7046 ;
  assign n7048 = ~n7042 & n7047 ;
  assign n7049 = ( ~n7042 & n7045 ) | ( ~n7042 & n7048 ) | ( n7045 & n7048 ) ;
  assign n7050 = n7041 & ~n7049 ;
  assign n7051 = ( ~n6953 & n7039 ) | ( ~n6953 & n7050 ) | ( n7039 & n7050 ) ;
  assign n7052 = ( ~n6100 & n7043 ) | ( ~n6100 & n7044 ) | ( n7043 & n7044 ) ;
  assign n7053 = ( ~n7042 & n7048 ) | ( ~n7042 & n7052 ) | ( n7048 & n7052 ) ;
  assign n7054 = n7041 & ~n7053 ;
  assign n7055 = ( ~n6953 & n7039 ) | ( ~n6953 & n7054 ) | ( n7039 & n7054 ) ;
  assign n7056 = ( n5216 & n7051 ) | ( n5216 & n7055 ) | ( n7051 & n7055 ) ;
  assign n7057 = n6953 & ~n7038 ;
  assign n7058 = ~n7050 & n7057 ;
  assign n7059 = ~n7054 & n7057 ;
  assign n7060 = ( ~n5216 & n7058 ) | ( ~n5216 & n7059 ) | ( n7058 & n7059 ) ;
  assign n7061 = n7056 | n7060 ;
  assign n7062 = ~x6 & x7 ;
  assign n7063 = x6 & ~x7 ;
  assign n7064 = n7062 | n7063 ;
  assign n7065 = x5 & ~x6 ;
  assign n7066 = ~x5 & x6 ;
  assign n7067 = n7065 | n7066 ;
  assign n7068 = n7064 & ~n7067 ;
  assign n7069 = n6950 & n7068 ;
  assign n7070 = x7 & ~x8 ;
  assign n7071 = ~x7 & x8 ;
  assign n7072 = n7070 | n7071 ;
  assign n7073 = ~n7067 & n7072 ;
  assign n7074 = ~n7064 & n7073 ;
  assign n7075 = n7036 & n7074 ;
  assign n7076 = ( n7023 & n7074 ) | ( n7023 & n7075 ) | ( n7074 & n7075 ) ;
  assign n7077 = n7069 | n7076 ;
  assign n7078 = n7067 & n7072 ;
  assign n7079 = n7067 & ~n7072 ;
  assign n7080 = n6889 & n7079 ;
  assign n7081 = n7078 | n7080 ;
  assign n7082 = n7078 | n7079 ;
  assign n7083 = ( ~n6884 & n7081 ) | ( ~n6884 & n7082 ) | ( n7081 & n7082 ) ;
  assign n7084 = n7077 | n7083 ;
  assign n7085 = ( ~n6884 & n7079 ) | ( ~n6884 & n7080 ) | ( n7079 & n7080 ) ;
  assign n7086 = n7077 | n7085 ;
  assign n7087 = n7084 & n7086 ;
  assign n7088 = ( ~n7061 & n7084 ) | ( ~n7061 & n7087 ) | ( n7084 & n7087 ) ;
  assign n7089 = ~x8 & n7087 ;
  assign n7090 = ~x8 & n7084 ;
  assign n7091 = ( ~n7061 & n7089 ) | ( ~n7061 & n7090 ) | ( n7089 & n7090 ) ;
  assign n7092 = x8 | n7089 ;
  assign n7093 = x8 | n7090 ;
  assign n7094 = ( ~n7061 & n7092 ) | ( ~n7061 & n7093 ) | ( n7092 & n7093 ) ;
  assign n7095 = ( ~n7088 & n7091 ) | ( ~n7088 & n7094 ) | ( n7091 & n7094 ) ;
  assign n7096 = n6798 & n7095 ;
  assign n7097 = n6798 & ~n7096 ;
  assign n7098 = ~n6798 & n7095 ;
  assign n7099 = n7097 | n7098 ;
  assign n7100 = ~n6173 & n6793 ;
  assign n7101 = n6173 & ~n6793 ;
  assign n7102 = n7100 | n7101 ;
  assign n7103 = ( n5216 & n7050 ) | ( n5216 & n7054 ) | ( n7050 & n7054 ) ;
  assign n7104 = ~n7041 & n7053 ;
  assign n7105 = ~n7041 & n7049 ;
  assign n7106 = ( ~n5216 & n7104 ) | ( ~n5216 & n7105 ) | ( n7104 & n7105 ) ;
  assign n7107 = n7103 | n7106 ;
  assign n7108 = ~n6091 & n7074 ;
  assign n7109 = n7036 & n7068 ;
  assign n7110 = ( n7023 & n7068 ) | ( n7023 & n7109 ) | ( n7068 & n7109 ) ;
  assign n7111 = n7108 | n7110 ;
  assign n7112 = n6950 & n7079 ;
  assign n7113 = n7111 | n7112 ;
  assign n7114 = n7078 | n7113 ;
  assign n7115 = n7113 & n7114 ;
  assign n7116 = ( ~n7107 & n7114 ) | ( ~n7107 & n7115 ) | ( n7114 & n7115 ) ;
  assign n7117 = ~x8 & n7115 ;
  assign n7118 = ~x8 & n7114 ;
  assign n7119 = ( ~n7107 & n7117 ) | ( ~n7107 & n7118 ) | ( n7117 & n7118 ) ;
  assign n7120 = x8 | n7117 ;
  assign n7121 = x8 | n7118 ;
  assign n7122 = ( ~n7107 & n7120 ) | ( ~n7107 & n7121 ) | ( n7120 & n7121 ) ;
  assign n7123 = ( ~n7116 & n7119 ) | ( ~n7116 & n7122 ) | ( n7119 & n7122 ) ;
  assign n7124 = ~n7102 & n7123 ;
  assign n7125 = n7102 | n7124 ;
  assign n7126 = n7102 & n7123 ;
  assign n7127 = n7125 & ~n7126 ;
  assign n7128 = n6200 | n6791 ;
  assign n7129 = ~n6792 & n7128 ;
  assign n7130 = n7045 | n7047 ;
  assign n7131 = n7047 | n7052 ;
  assign n7132 = ( ~n5216 & n7130 ) | ( ~n5216 & n7131 ) | ( n7130 & n7131 ) ;
  assign n7133 = n7047 & n7052 ;
  assign n7134 = n7045 & n7047 ;
  assign n7135 = ( ~n5216 & n7133 ) | ( ~n5216 & n7134 ) | ( n7133 & n7134 ) ;
  assign n7136 = n7132 & ~n7135 ;
  assign n7137 = n5857 & n7074 ;
  assign n7138 = ( ~n5899 & n7074 ) | ( ~n5899 & n7137 ) | ( n7074 & n7137 ) ;
  assign n7139 = ~n6091 & n7068 ;
  assign n7140 = n7036 & n7079 ;
  assign n7141 = ( n7023 & n7079 ) | ( n7023 & n7140 ) | ( n7079 & n7140 ) ;
  assign n7142 = n7139 | n7141 ;
  assign n7143 = n7138 | n7142 ;
  assign n7144 = n7078 | n7143 ;
  assign n7145 = n7143 & n7144 ;
  assign n7146 = ( n7136 & n7144 ) | ( n7136 & n7145 ) | ( n7144 & n7145 ) ;
  assign n7147 = x8 & n7145 ;
  assign n7148 = x8 & n7144 ;
  assign n7149 = ( n7136 & n7147 ) | ( n7136 & n7148 ) | ( n7147 & n7148 ) ;
  assign n7150 = x8 & ~n7147 ;
  assign n7151 = x8 & ~n7148 ;
  assign n7152 = ( ~n7136 & n7150 ) | ( ~n7136 & n7151 ) | ( n7150 & n7151 ) ;
  assign n7153 = ( n7146 & ~n7149 ) | ( n7146 & n7152 ) | ( ~n7149 & n7152 ) ;
  assign n7154 = n7129 & n7153 ;
  assign n7155 = n6222 & ~n6789 ;
  assign n7156 = n6790 | n7155 ;
  assign n7157 = n5857 & n7068 ;
  assign n7158 = ( ~n5899 & n7068 ) | ( ~n5899 & n7157 ) | ( n7068 & n7157 ) ;
  assign n7159 = ~n6091 & n7079 ;
  assign n7160 = n5997 & n7074 ;
  assign n7161 = ( n5979 & n7074 ) | ( n5979 & n7160 ) | ( n7074 & n7160 ) ;
  assign n7162 = n7159 | n7161 ;
  assign n7163 = n7158 | n7162 ;
  assign n7164 = n7078 | n7163 ;
  assign n7165 = n7163 & n7164 ;
  assign n7166 = ( n6108 & n7164 ) | ( n6108 & n7165 ) | ( n7164 & n7165 ) ;
  assign n7167 = x8 & n7165 ;
  assign n7168 = x8 & n7164 ;
  assign n7169 = ( n6108 & n7167 ) | ( n6108 & n7168 ) | ( n7167 & n7168 ) ;
  assign n7170 = x8 & ~n7167 ;
  assign n7171 = x8 & ~n7168 ;
  assign n7172 = ( ~n6108 & n7170 ) | ( ~n6108 & n7171 ) | ( n7170 & n7171 ) ;
  assign n7173 = ( n7166 & ~n7169 ) | ( n7166 & n7172 ) | ( ~n7169 & n7172 ) ;
  assign n7174 = ~n7156 & n7173 ;
  assign n7175 = n6246 & ~n6787 ;
  assign n7176 = n6788 | n7175 ;
  assign n7177 = n5108 & n7074 ;
  assign n7178 = n5997 & n7068 ;
  assign n7179 = ( n5979 & n7068 ) | ( n5979 & n7178 ) | ( n7068 & n7178 ) ;
  assign n7180 = n7177 | n7179 ;
  assign n7181 = n5857 & n7079 ;
  assign n7182 = ( ~n5899 & n7079 ) | ( ~n5899 & n7181 ) | ( n7079 & n7181 ) ;
  assign n7183 = n7180 | n7182 ;
  assign n7184 = n7078 | n7183 ;
  assign n7185 = n7183 & n7184 ;
  assign n7186 = ( ~n6151 & n7184 ) | ( ~n6151 & n7185 ) | ( n7184 & n7185 ) ;
  assign n7187 = ~x8 & n7185 ;
  assign n7188 = ~x8 & n7184 ;
  assign n7189 = ( ~n6151 & n7187 ) | ( ~n6151 & n7188 ) | ( n7187 & n7188 ) ;
  assign n7190 = x8 | n7187 ;
  assign n7191 = x8 | n7188 ;
  assign n7192 = ( ~n6151 & n7190 ) | ( ~n6151 & n7191 ) | ( n7190 & n7191 ) ;
  assign n7193 = ( ~n7186 & n7189 ) | ( ~n7186 & n7192 ) | ( n7189 & n7192 ) ;
  assign n7194 = ~n7176 & n7193 ;
  assign n7195 = n7176 | n7194 ;
  assign n7196 = n7176 & n7193 ;
  assign n7197 = n7195 & ~n7196 ;
  assign n7198 = n6783 & n6785 ;
  assign n7199 = n6783 | n6785 ;
  assign n7200 = ~n7198 & n7199 ;
  assign n7201 = n5117 & n7074 ;
  assign n7202 = ( ~n5037 & n7074 ) | ( ~n5037 & n7201 ) | ( n7074 & n7201 ) ;
  assign n7203 = n5108 & n7068 ;
  assign n7204 = n5997 & n7079 ;
  assign n7205 = ( n5979 & n7079 ) | ( n5979 & n7204 ) | ( n7079 & n7204 ) ;
  assign n7206 = n7203 | n7205 ;
  assign n7207 = n7202 | n7206 ;
  assign n7208 = n7078 | n7207 ;
  assign n7209 = n7207 & n7208 ;
  assign n7210 = ( n6181 & n7208 ) | ( n6181 & n7209 ) | ( n7208 & n7209 ) ;
  assign n7211 = x8 & n7209 ;
  assign n7212 = x8 & n7208 ;
  assign n7213 = ( n6181 & n7211 ) | ( n6181 & n7212 ) | ( n7211 & n7212 ) ;
  assign n7214 = x8 & ~n7211 ;
  assign n7215 = x8 & ~n7212 ;
  assign n7216 = ( ~n6181 & n7214 ) | ( ~n6181 & n7215 ) | ( n7214 & n7215 ) ;
  assign n7217 = ( n7210 & ~n7213 ) | ( n7210 & n7216 ) | ( ~n7213 & n7216 ) ;
  assign n7218 = n7200 & n7217 ;
  assign n7219 = n7200 & ~n7218 ;
  assign n7220 = ~n7200 & n7217 ;
  assign n7221 = n7219 | n7220 ;
  assign n7222 = n6290 | n6310 ;
  assign n7223 = n6780 | n7222 ;
  assign n7224 = ~n6782 & n7223 ;
  assign n7225 = n5117 & n7068 ;
  assign n7226 = ( ~n5037 & n7068 ) | ( ~n5037 & n7225 ) | ( n7068 & n7225 ) ;
  assign n7227 = n5108 & n7079 ;
  assign n7228 = n5192 & n7074 ;
  assign n7229 = ( n5179 & n7074 ) | ( n5179 & n7228 ) | ( n7074 & n7228 ) ;
  assign n7230 = n7227 | n7229 ;
  assign n7231 = n7226 | n7230 ;
  assign n7232 = n7078 | n7231 ;
  assign n7233 = ( ~n5220 & n7231 ) | ( ~n5220 & n7232 ) | ( n7231 & n7232 ) ;
  assign n7234 = ~x8 & n7232 ;
  assign n7235 = ~x8 & n7231 ;
  assign n7236 = ( ~n5220 & n7234 ) | ( ~n5220 & n7235 ) | ( n7234 & n7235 ) ;
  assign n7237 = x8 | n7234 ;
  assign n7238 = x8 | n7235 ;
  assign n7239 = ( ~n5220 & n7237 ) | ( ~n5220 & n7238 ) | ( n7237 & n7238 ) ;
  assign n7240 = ( ~n7233 & n7236 ) | ( ~n7233 & n7239 ) | ( n7236 & n7239 ) ;
  assign n7241 = n7224 & n7240 ;
  assign n7242 = ~n6313 & n6779 ;
  assign n7243 = n6313 & ~n6779 ;
  assign n7244 = n7242 | n7243 ;
  assign n7245 = n4245 & n7074 ;
  assign n7246 = ( n4303 & n7074 ) | ( n4303 & n7245 ) | ( n7074 & n7245 ) ;
  assign n7247 = n5192 & n7068 ;
  assign n7248 = ( n5179 & n7068 ) | ( n5179 & n7247 ) | ( n7068 & n7247 ) ;
  assign n7249 = n7246 | n7248 ;
  assign n7250 = n5117 & n7079 ;
  assign n7251 = ( ~n5037 & n7079 ) | ( ~n5037 & n7250 ) | ( n7079 & n7250 ) ;
  assign n7252 = n7249 | n7251 ;
  assign n7253 = n7078 | n7251 ;
  assign n7254 = n7249 | n7253 ;
  assign n7255 = ( ~n5270 & n7252 ) | ( ~n5270 & n7254 ) | ( n7252 & n7254 ) ;
  assign n7256 = ~x8 & n7254 ;
  assign n7257 = ~x8 & n7252 ;
  assign n7258 = ( ~n5270 & n7256 ) | ( ~n5270 & n7257 ) | ( n7256 & n7257 ) ;
  assign n7259 = x8 | n7257 ;
  assign n7260 = x8 | n7256 ;
  assign n7261 = ( ~n5270 & n7259 ) | ( ~n5270 & n7260 ) | ( n7259 & n7260 ) ;
  assign n7262 = ( ~n7255 & n7258 ) | ( ~n7255 & n7261 ) | ( n7258 & n7261 ) ;
  assign n7263 = n7244 & n7262 ;
  assign n7264 = n6354 | n6776 ;
  assign n7265 = n6774 | n7264 ;
  assign n7266 = ~n6778 & n7265 ;
  assign n7267 = n4396 & n7074 ;
  assign n7268 = n4245 & n7068 ;
  assign n7269 = ( n4303 & n7068 ) | ( n4303 & n7268 ) | ( n7068 & n7268 ) ;
  assign n7270 = n7267 | n7269 ;
  assign n7271 = n5192 & n7079 ;
  assign n7272 = ( n5179 & n7079 ) | ( n5179 & n7271 ) | ( n7079 & n7271 ) ;
  assign n7274 = n7078 | n7272 ;
  assign n7275 = n7270 | n7274 ;
  assign n7273 = n7270 | n7272 ;
  assign n7276 = n7273 & n7275 ;
  assign n7277 = ( n5306 & n7275 ) | ( n5306 & n7276 ) | ( n7275 & n7276 ) ;
  assign n7278 = x8 & n7276 ;
  assign n7279 = x8 & n7275 ;
  assign n7280 = ( n5306 & n7278 ) | ( n5306 & n7279 ) | ( n7278 & n7279 ) ;
  assign n7281 = x8 & ~n7278 ;
  assign n7282 = x8 & ~n7279 ;
  assign n7283 = ( ~n5306 & n7281 ) | ( ~n5306 & n7282 ) | ( n7281 & n7282 ) ;
  assign n7284 = ( n7277 & ~n7280 ) | ( n7277 & n7283 ) | ( ~n7280 & n7283 ) ;
  assign n7285 = n7266 & n7284 ;
  assign n7286 = n7266 | n7284 ;
  assign n7287 = ~n7285 & n7286 ;
  assign n7288 = n6358 | n6773 ;
  assign n7289 = ~n6774 & n7288 ;
  assign n7290 = ~n4429 & n7074 ;
  assign n7291 = n4396 & n7068 ;
  assign n7292 = n7290 | n7291 ;
  assign n7293 = n4245 & n7079 ;
  assign n7294 = ( n4303 & n7079 ) | ( n4303 & n7293 ) | ( n7079 & n7293 ) ;
  assign n7296 = n7078 | n7294 ;
  assign n7297 = n7292 | n7296 ;
  assign n7295 = n7292 | n7294 ;
  assign n7298 = n7295 & n7297 ;
  assign n7299 = ( n4455 & n7297 ) | ( n4455 & n7298 ) | ( n7297 & n7298 ) ;
  assign n7300 = x8 & n7298 ;
  assign n7301 = x8 & n7297 ;
  assign n7302 = ( n4455 & n7300 ) | ( n4455 & n7301 ) | ( n7300 & n7301 ) ;
  assign n7303 = x8 & ~n7300 ;
  assign n7304 = x8 & ~n7301 ;
  assign n7305 = ( ~n4455 & n7303 ) | ( ~n4455 & n7304 ) | ( n7303 & n7304 ) ;
  assign n7306 = ( n7299 & ~n7302 ) | ( n7299 & n7305 ) | ( ~n7302 & n7305 ) ;
  assign n7307 = n7289 & n7306 ;
  assign n7308 = n7289 & ~n7307 ;
  assign n7309 = ~n7289 & n7306 ;
  assign n7310 = n7308 | n7309 ;
  assign n7311 = n6381 | n6771 ;
  assign n7312 = ~n6772 & n7311 ;
  assign n7313 = ~n4429 & n7068 ;
  assign n7314 = n7068 | n7074 ;
  assign n7315 = ( ~n4429 & n7074 ) | ( ~n4429 & n7314 ) | ( n7074 & n7314 ) ;
  assign n7316 = ( n4206 & n7313 ) | ( n4206 & n7315 ) | ( n7313 & n7315 ) ;
  assign n7317 = n4396 & n7079 ;
  assign n7319 = n7078 | n7317 ;
  assign n7320 = n7316 | n7319 ;
  assign n7318 = n7316 | n7317 ;
  assign n7321 = n7318 & n7320 ;
  assign n7322 = ( ~n4501 & n7320 ) | ( ~n4501 & n7321 ) | ( n7320 & n7321 ) ;
  assign n7323 = ~x8 & n7321 ;
  assign n7324 = ~x8 & n7320 ;
  assign n7325 = ( ~n4501 & n7323 ) | ( ~n4501 & n7324 ) | ( n7323 & n7324 ) ;
  assign n7326 = x8 | n7323 ;
  assign n7327 = x8 | n7324 ;
  assign n7328 = ( ~n4501 & n7326 ) | ( ~n4501 & n7327 ) | ( n7326 & n7327 ) ;
  assign n7329 = ( ~n7322 & n7325 ) | ( ~n7322 & n7328 ) | ( n7325 & n7328 ) ;
  assign n7330 = n7312 & n7329 ;
  assign n7331 = n7312 & ~n7330 ;
  assign n7332 = ~n7312 & n7329 ;
  assign n7333 = n7331 | n7332 ;
  assign n7334 = n6762 | n6768 ;
  assign n7335 = n6766 | n7334 ;
  assign n7336 = ~n6770 & n7335 ;
  assign n7337 = n4206 & n7068 ;
  assign n7338 = ~n4429 & n7079 ;
  assign n7339 = n3439 & n7074 ;
  assign n7340 = ( ~n3420 & n7074 ) | ( ~n3420 & n7339 ) | ( n7074 & n7339 ) ;
  assign n7341 = n7338 | n7340 ;
  assign n7342 = n7337 | n7341 ;
  assign n7343 = n7078 | n7337 ;
  assign n7344 = n7341 | n7343 ;
  assign n7345 = ( ~n4527 & n7342 ) | ( ~n4527 & n7344 ) | ( n7342 & n7344 ) ;
  assign n7346 = ~x8 & n7344 ;
  assign n7347 = ~x8 & n7342 ;
  assign n7348 = ( ~n4527 & n7346 ) | ( ~n4527 & n7347 ) | ( n7346 & n7347 ) ;
  assign n7349 = x8 | n7347 ;
  assign n7350 = x8 | n7346 ;
  assign n7351 = ( ~n4527 & n7349 ) | ( ~n4527 & n7350 ) | ( n7349 & n7350 ) ;
  assign n7352 = ( ~n7345 & n7348 ) | ( ~n7345 & n7351 ) | ( n7348 & n7351 ) ;
  assign n7353 = n7336 & n7352 ;
  assign n7354 = n6765 & ~n6766 ;
  assign n7355 = n6740 & ~n6765 ;
  assign n7356 = n7354 | n7355 ;
  assign n7357 = n4206 & n7079 ;
  assign n7358 = n3386 & n7074 ;
  assign n7359 = n3439 & n7068 ;
  assign n7360 = ( ~n3420 & n7068 ) | ( ~n3420 & n7359 ) | ( n7068 & n7359 ) ;
  assign n7361 = n7358 | n7360 ;
  assign n7362 = n7357 | n7361 ;
  assign n7363 = n7078 | n7357 ;
  assign n7364 = n7361 | n7363 ;
  assign n7365 = ( ~n4220 & n7362 ) | ( ~n4220 & n7364 ) | ( n7362 & n7364 ) ;
  assign n7366 = ~x8 & n7364 ;
  assign n7367 = ~x8 & n7362 ;
  assign n7368 = ( ~n4220 & n7366 ) | ( ~n4220 & n7367 ) | ( n7366 & n7367 ) ;
  assign n7369 = x8 | n7367 ;
  assign n7370 = x8 | n7366 ;
  assign n7371 = ( ~n4220 & n7369 ) | ( ~n4220 & n7370 ) | ( n7369 & n7370 ) ;
  assign n7372 = ( ~n7365 & n7368 ) | ( ~n7365 & n7371 ) | ( n7368 & n7371 ) ;
  assign n7373 = n7355 & n7372 ;
  assign n7374 = ( n7354 & n7372 ) | ( n7354 & n7373 ) | ( n7372 & n7373 ) ;
  assign n7375 = n7356 & ~n7374 ;
  assign n7376 = ~n7355 & n7372 ;
  assign n7377 = ~n7354 & n7376 ;
  assign n7378 = n7375 | n7377 ;
  assign n7379 = n6738 & ~n6739 ;
  assign n7380 = n6427 & ~n6739 ;
  assign n7381 = n7379 | n7380 ;
  assign n7382 = n3386 & n7068 ;
  assign n7383 = n3507 & n7074 ;
  assign n7384 = ( n3483 & n7074 ) | ( n3483 & n7383 ) | ( n7074 & n7383 ) ;
  assign n7385 = n3439 & n7079 ;
  assign n7386 = ( ~n3420 & n7079 ) | ( ~n3420 & n7385 ) | ( n7079 & n7385 ) ;
  assign n7387 = n7384 | n7386 ;
  assign n7388 = n7382 | n7387 ;
  assign n7389 = n7078 | n7388 ;
  assign n7390 = ( ~n3530 & n7388 ) | ( ~n3530 & n7389 ) | ( n7388 & n7389 ) ;
  assign n7391 = ~x8 & n7389 ;
  assign n7392 = ~x8 & n7388 ;
  assign n7393 = ( ~n3530 & n7391 ) | ( ~n3530 & n7392 ) | ( n7391 & n7392 ) ;
  assign n7394 = x8 | n7391 ;
  assign n7395 = x8 | n7392 ;
  assign n7396 = ( ~n3530 & n7394 ) | ( ~n3530 & n7395 ) | ( n7394 & n7395 ) ;
  assign n7397 = ( ~n7390 & n7393 ) | ( ~n7390 & n7396 ) | ( n7393 & n7396 ) ;
  assign n7398 = n7381 & n7397 ;
  assign n7399 = n7381 & ~n7398 ;
  assign n7400 = ~n7381 & n7397 ;
  assign n7401 = n7399 | n7400 ;
  assign n7402 = n6734 & n6736 ;
  assign n7403 = n6734 | n6736 ;
  assign n7404 = ~n7402 & n7403 ;
  assign n7405 = n2893 & n7074 ;
  assign n7406 = ( ~n2886 & n7074 ) | ( ~n2886 & n7405 ) | ( n7074 & n7405 ) ;
  assign n7407 = n3507 & n7068 ;
  assign n7408 = ( n3483 & n7068 ) | ( n3483 & n7407 ) | ( n7068 & n7407 ) ;
  assign n7409 = n7406 | n7408 ;
  assign n7410 = n3386 & n7079 ;
  assign n7412 = n7078 | n7410 ;
  assign n7413 = n7409 | n7412 ;
  assign n7411 = n7409 | n7410 ;
  assign n7414 = n7411 & n7413 ;
  assign n7415 = ( ~n3568 & n7413 ) | ( ~n3568 & n7414 ) | ( n7413 & n7414 ) ;
  assign n7416 = ~x8 & n7414 ;
  assign n7417 = ~x8 & n7413 ;
  assign n7418 = ( ~n3568 & n7416 ) | ( ~n3568 & n7417 ) | ( n7416 & n7417 ) ;
  assign n7419 = x8 | n7416 ;
  assign n7420 = x8 | n7417 ;
  assign n7421 = ( ~n3568 & n7419 ) | ( ~n3568 & n7420 ) | ( n7419 & n7420 ) ;
  assign n7422 = ( ~n7415 & n7418 ) | ( ~n7415 & n7421 ) | ( n7418 & n7421 ) ;
  assign n7423 = n7404 & n7422 ;
  assign n7424 = n6497 | n6730 ;
  assign n7425 = ~n6731 & n7424 ;
  assign n7426 = n2691 & n7074 ;
  assign n7427 = ( n2678 & n7074 ) | ( n2678 & n7426 ) | ( n7074 & n7426 ) ;
  assign n7428 = n2701 & n7068 ;
  assign n7429 = ( ~n2784 & n7068 ) | ( ~n2784 & n7428 ) | ( n7068 & n7428 ) ;
  assign n7430 = n7427 | n7429 ;
  assign n7431 = n2893 & n7079 ;
  assign n7432 = ( ~n2886 & n7079 ) | ( ~n2886 & n7431 ) | ( n7079 & n7431 ) ;
  assign n7433 = n7430 | n7432 ;
  assign n7434 = n7078 | n7433 ;
  assign n7435 = n7433 & n7434 ;
  assign n7436 = ( ~n2914 & n7434 ) | ( ~n2914 & n7435 ) | ( n7434 & n7435 ) ;
  assign n7437 = ~x8 & n7435 ;
  assign n7438 = ~x8 & n7434 ;
  assign n7439 = ( ~n2914 & n7437 ) | ( ~n2914 & n7438 ) | ( n7437 & n7438 ) ;
  assign n7440 = x8 | n7437 ;
  assign n7441 = x8 | n7438 ;
  assign n7442 = ( ~n2914 & n7440 ) | ( ~n2914 & n7441 ) | ( n7440 & n7441 ) ;
  assign n7443 = ( ~n7436 & n7439 ) | ( ~n7436 & n7442 ) | ( n7439 & n7442 ) ;
  assign n7444 = n7425 & n7443 ;
  assign n7445 = n7425 & ~n7444 ;
  assign n7446 = ~n7425 & n7443 ;
  assign n7447 = n7445 | n7446 ;
  assign n7448 = n6726 & n6728 ;
  assign n7449 = n6726 | n6728 ;
  assign n7450 = ~n7448 & n7449 ;
  assign n7451 = n2701 & n7079 ;
  assign n7452 = ( ~n2784 & n7079 ) | ( ~n2784 & n7451 ) | ( n7079 & n7451 ) ;
  assign n7453 = n2691 & n7068 ;
  assign n7454 = ( n2678 & n7068 ) | ( n2678 & n7453 ) | ( n7068 & n7453 ) ;
  assign n7455 = n7452 | n7454 ;
  assign n7456 = n2199 & n7074 ;
  assign n7457 = ( ~n2185 & n7074 ) | ( ~n2185 & n7456 ) | ( n7074 & n7456 ) ;
  assign n7458 = n7455 | n7457 ;
  assign n7459 = n7078 | n7457 ;
  assign n7460 = n7455 | n7459 ;
  assign n7461 = ( n2960 & n7458 ) | ( n2960 & n7460 ) | ( n7458 & n7460 ) ;
  assign n7462 = x8 & n7460 ;
  assign n7463 = x8 & n7458 ;
  assign n7464 = ( n2960 & n7462 ) | ( n2960 & n7463 ) | ( n7462 & n7463 ) ;
  assign n7465 = x8 & ~n7463 ;
  assign n7466 = x8 & ~n7462 ;
  assign n7467 = ( ~n2960 & n7465 ) | ( ~n2960 & n7466 ) | ( n7465 & n7466 ) ;
  assign n7468 = ( n7461 & ~n7464 ) | ( n7461 & n7467 ) | ( ~n7464 & n7467 ) ;
  assign n7469 = n7450 & n7468 ;
  assign n7470 = n6721 & n6724 ;
  assign n7471 = n6721 & ~n7470 ;
  assign n7474 = n2090 & n7074 ;
  assign n7475 = ( ~n2082 & n7074 ) | ( ~n2082 & n7474 ) | ( n7074 & n7474 ) ;
  assign n7476 = n2691 & n7079 ;
  assign n7477 = ( n2678 & n7079 ) | ( n2678 & n7476 ) | ( n7079 & n7476 ) ;
  assign n7478 = n2199 & n7068 ;
  assign n7479 = ( ~n2185 & n7068 ) | ( ~n2185 & n7478 ) | ( n7068 & n7478 ) ;
  assign n7480 = n7477 | n7479 ;
  assign n7481 = n7475 | n7480 ;
  assign n7482 = n7078 | n7481 ;
  assign n7483 = ( n2985 & n7481 ) | ( n2985 & n7482 ) | ( n7481 & n7482 ) ;
  assign n7484 = x8 & n7482 ;
  assign n7485 = x8 & n7481 ;
  assign n7486 = ( n2985 & n7484 ) | ( n2985 & n7485 ) | ( n7484 & n7485 ) ;
  assign n7487 = x8 & ~n7484 ;
  assign n7488 = x8 & ~n7485 ;
  assign n7489 = ( ~n2985 & n7487 ) | ( ~n2985 & n7488 ) | ( n7487 & n7488 ) ;
  assign n7490 = ( n7483 & ~n7486 ) | ( n7483 & n7489 ) | ( ~n7486 & n7489 ) ;
  assign n7472 = ~n6721 & n6724 ;
  assign n7491 = n7472 & n7490 ;
  assign n7492 = ( n7471 & n7490 ) | ( n7471 & n7491 ) | ( n7490 & n7491 ) ;
  assign n7473 = n7471 | n7472 ;
  assign n7493 = n7473 & ~n7492 ;
  assign n7494 = ~n7472 & n7490 ;
  assign n7495 = ~n7471 & n7494 ;
  assign n7496 = n7493 | n7495 ;
  assign n7497 = ~n6716 & n6719 ;
  assign n7498 = n6716 & ~n6719 ;
  assign n7499 = n7497 | n7498 ;
  assign n7500 = n2090 & n7068 ;
  assign n7501 = ( ~n2082 & n7068 ) | ( ~n2082 & n7500 ) | ( n7068 & n7500 ) ;
  assign n7502 = n2279 & n7074 ;
  assign n7503 = ( ~n2269 & n7074 ) | ( ~n2269 & n7502 ) | ( n7074 & n7502 ) ;
  assign n7504 = n2199 & n7079 ;
  assign n7505 = ( ~n2185 & n7079 ) | ( ~n2185 & n7504 ) | ( n7079 & n7504 ) ;
  assign n7506 = n7503 | n7505 ;
  assign n7507 = n7501 | n7506 ;
  assign n7508 = n7078 | n7507 ;
  assign n7509 = ( ~n2325 & n7507 ) | ( ~n2325 & n7508 ) | ( n7507 & n7508 ) ;
  assign n7510 = n7507 & n7508 ;
  assign n7511 = ( ~n2299 & n7509 ) | ( ~n2299 & n7510 ) | ( n7509 & n7510 ) ;
  assign n7512 = ~x8 & n7511 ;
  assign n7513 = x8 | n7511 ;
  assign n7514 = ( ~n7511 & n7512 ) | ( ~n7511 & n7513 ) | ( n7512 & n7513 ) ;
  assign n7515 = n7499 & n7514 ;
  assign n7516 = n7499 | n7514 ;
  assign n7517 = ~n7515 & n7516 ;
  assign n7518 = n6712 | n6714 ;
  assign n7519 = ~n6715 & n7518 ;
  assign n7520 = n1634 & n7074 ;
  assign n7521 = ( n1630 & n7074 ) | ( n1630 & n7520 ) | ( n7074 & n7520 ) ;
  assign n7522 = n2279 & n7068 ;
  assign n7523 = ( ~n2269 & n7068 ) | ( ~n2269 & n7522 ) | ( n7068 & n7522 ) ;
  assign n7524 = n7521 | n7523 ;
  assign n7525 = n2090 & n7079 ;
  assign n7526 = ( ~n2082 & n7079 ) | ( ~n2082 & n7525 ) | ( n7079 & n7525 ) ;
  assign n7527 = n7524 | n7526 ;
  assign n7528 = n7078 | n7527 ;
  assign n7529 = n7527 & n7528 ;
  assign n7530 = ( n2568 & n7528 ) | ( n2568 & n7529 ) | ( n7528 & n7529 ) ;
  assign n7531 = x8 & n7529 ;
  assign n7532 = x8 & n7528 ;
  assign n7533 = ( n2568 & n7531 ) | ( n2568 & n7532 ) | ( n7531 & n7532 ) ;
  assign n7534 = x8 & ~n7531 ;
  assign n7535 = x8 & ~n7532 ;
  assign n7536 = ( ~n2568 & n7534 ) | ( ~n2568 & n7535 ) | ( n7534 & n7535 ) ;
  assign n7537 = ( n7530 & ~n7533 ) | ( n7530 & n7536 ) | ( ~n7533 & n7536 ) ;
  assign n7538 = n7519 & n7537 ;
  assign n7539 = n6602 | n6710 ;
  assign n7540 = ~n6711 & n7539 ;
  assign n7541 = n1708 & n7074 ;
  assign n7542 = n1634 & n7068 ;
  assign n7543 = ( n1630 & n7068 ) | ( n1630 & n7542 ) | ( n7068 & n7542 ) ;
  assign n7544 = n2279 & n7079 ;
  assign n7545 = ( ~n2269 & n7079 ) | ( ~n2269 & n7544 ) | ( n7079 & n7544 ) ;
  assign n7546 = n7543 | n7545 ;
  assign n7547 = n7541 | n7546 ;
  assign n7548 = n7078 | n7547 ;
  assign n7549 = n7547 & n7548 ;
  assign n7550 = ( ~n2343 & n7548 ) | ( ~n2343 & n7549 ) | ( n7548 & n7549 ) ;
  assign n7551 = ~x8 & n7549 ;
  assign n7552 = ~x8 & n7548 ;
  assign n7553 = ( ~n2343 & n7551 ) | ( ~n2343 & n7552 ) | ( n7551 & n7552 ) ;
  assign n7554 = x8 | n7551 ;
  assign n7555 = x8 | n7552 ;
  assign n7556 = ( ~n2343 & n7554 ) | ( ~n2343 & n7555 ) | ( n7554 & n7555 ) ;
  assign n7557 = ( ~n7550 & n7553 ) | ( ~n7550 & n7556 ) | ( n7553 & n7556 ) ;
  assign n7558 = n7540 & n7557 ;
  assign n7559 = n6706 & n6708 ;
  assign n7560 = n6706 | n6708 ;
  assign n7561 = ~n7559 & n7560 ;
  assign n7562 = n1708 & n7068 ;
  assign n7563 = n1793 & n7074 ;
  assign n7564 = ( n1783 & n7074 ) | ( n1783 & n7563 ) | ( n7074 & n7563 ) ;
  assign n7565 = n1634 & n7079 ;
  assign n7566 = ( n1630 & n7079 ) | ( n1630 & n7565 ) | ( n7079 & n7565 ) ;
  assign n7567 = n7564 | n7566 ;
  assign n7568 = n7562 | n7567 ;
  assign n7569 = n7078 | n7568 ;
  assign n7570 = n7568 & n7569 ;
  assign n7571 = ( n1814 & n7569 ) | ( n1814 & n7570 ) | ( n7569 & n7570 ) ;
  assign n7572 = x8 & n7570 ;
  assign n7573 = x8 & n7569 ;
  assign n7574 = ( n1814 & n7572 ) | ( n1814 & n7573 ) | ( n7572 & n7573 ) ;
  assign n7575 = x8 & ~n7572 ;
  assign n7576 = x8 & ~n7573 ;
  assign n7577 = ( ~n1814 & n7575 ) | ( ~n1814 & n7576 ) | ( n7575 & n7576 ) ;
  assign n7578 = ( n7571 & ~n7574 ) | ( n7571 & n7577 ) | ( ~n7574 & n7577 ) ;
  assign n7579 = n7561 & n7578 ;
  assign n7580 = n6702 & n6704 ;
  assign n7581 = n6702 | n6704 ;
  assign n7582 = ~n7580 & n7581 ;
  assign n7583 = ~n523 & n7074 ;
  assign n7584 = n1793 & n7068 ;
  assign n7585 = ( n1783 & n7068 ) | ( n1783 & n7584 ) | ( n7068 & n7584 ) ;
  assign n7586 = n7583 | n7585 ;
  assign n7587 = n1708 & n7079 ;
  assign n7588 = n7586 | n7587 ;
  assign n7589 = n7078 | n7587 ;
  assign n7590 = n7586 | n7589 ;
  assign n7591 = ( ~n1852 & n7588 ) | ( ~n1852 & n7590 ) | ( n7588 & n7590 ) ;
  assign n7592 = ~x8 & n7590 ;
  assign n7593 = ~x8 & n7588 ;
  assign n7594 = ( ~n1852 & n7592 ) | ( ~n1852 & n7593 ) | ( n7592 & n7593 ) ;
  assign n7595 = x8 | n7593 ;
  assign n7596 = x8 | n7592 ;
  assign n7597 = ( ~n1852 & n7595 ) | ( ~n1852 & n7596 ) | ( n7595 & n7596 ) ;
  assign n7598 = ( ~n7591 & n7594 ) | ( ~n7591 & n7597 ) | ( n7594 & n7597 ) ;
  assign n7599 = n7582 & n7598 ;
  assign n7600 = n6698 | n6699 ;
  assign n7601 = n6682 | n7600 ;
  assign n7602 = ~n6701 & n7601 ;
  assign n7603 = ~n523 & n7068 ;
  assign n7604 = n352 & n7074 ;
  assign n7605 = ( ~n339 & n7074 ) | ( ~n339 & n7604 ) | ( n7074 & n7604 ) ;
  assign n7606 = n1793 & n7079 ;
  assign n7607 = ( n1783 & n7079 ) | ( n1783 & n7606 ) | ( n7079 & n7606 ) ;
  assign n7608 = n7605 | n7607 ;
  assign n7609 = n7603 | n7608 ;
  assign n7610 = n7078 | n7609 ;
  assign n7611 = n7609 & n7610 ;
  assign n7612 = ( n1884 & n7610 ) | ( n1884 & n7611 ) | ( n7610 & n7611 ) ;
  assign n7613 = x8 & n7611 ;
  assign n7614 = x8 & n7610 ;
  assign n7615 = ( n1884 & n7613 ) | ( n1884 & n7614 ) | ( n7613 & n7614 ) ;
  assign n7616 = x8 & ~n7613 ;
  assign n7617 = x8 & ~n7614 ;
  assign n7618 = ( ~n1884 & n7616 ) | ( ~n1884 & n7617 ) | ( n7616 & n7617 ) ;
  assign n7619 = ( n7612 & ~n7615 ) | ( n7612 & n7618 ) | ( ~n7615 & n7618 ) ;
  assign n7620 = n7602 & n7619 ;
  assign n7621 = n7602 | n7619 ;
  assign n7622 = ~n7620 & n7621 ;
  assign n7623 = ~n829 & n7074 ;
  assign n7624 = n352 & n7068 ;
  assign n7625 = ( ~n339 & n7068 ) | ( ~n339 & n7624 ) | ( n7068 & n7624 ) ;
  assign n7626 = n7623 | n7625 ;
  assign n7627 = ~n523 & n7079 ;
  assign n7628 = n7078 | n7627 ;
  assign n7629 = n7626 | n7628 ;
  assign n7630 = ~x8 & n7629 ;
  assign n7631 = n7626 | n7627 ;
  assign n7632 = ~x8 & n7631 ;
  assign n7633 = ( ~n1055 & n7630 ) | ( ~n1055 & n7632 ) | ( n7630 & n7632 ) ;
  assign n7634 = x8 & n7629 ;
  assign n7635 = x8 & ~n7634 ;
  assign n7636 = x8 & n7627 ;
  assign n7637 = ( x8 & n7626 ) | ( x8 & n7636 ) | ( n7626 & n7636 ) ;
  assign n7638 = x8 & ~n7637 ;
  assign n7639 = ( n1055 & n7635 ) | ( n1055 & n7638 ) | ( n7635 & n7638 ) ;
  assign n7640 = n7633 | n7639 ;
  assign n7641 = n6675 | n6677 ;
  assign n7642 = x11 & ~n6675 ;
  assign n7643 = ( n6658 & n7641 ) | ( n6658 & ~n7642 ) | ( n7641 & ~n7642 ) ;
  assign n7644 = ~n6680 & n7643 ;
  assign n7645 = n7640 & n7644 ;
  assign n7646 = x11 | n6672 ;
  assign n7647 = ( ~n6665 & n6672 ) | ( ~n6665 & n7646 ) | ( n6672 & n7646 ) ;
  assign n7648 = n6666 | n7647 ;
  assign n7649 = ~n6675 & n7648 ;
  assign n7650 = ~n829 & n7068 ;
  assign n7651 = n352 & n7079 ;
  assign n7652 = ( ~n339 & n7079 ) | ( ~n339 & n7651 ) | ( n7079 & n7651 ) ;
  assign n7653 = n7650 | n7652 ;
  assign n7654 = n692 & n7074 ;
  assign n7655 = ( n674 & n7074 ) | ( n674 & n7654 ) | ( n7074 & n7654 ) ;
  assign n7656 = n7653 | n7655 ;
  assign n7657 = n7078 | n7655 ;
  assign n7658 = n7653 | n7657 ;
  assign n7659 = ( ~n1209 & n7656 ) | ( ~n1209 & n7658 ) | ( n7656 & n7658 ) ;
  assign n7660 = ~x8 & n7658 ;
  assign n7661 = ~x8 & n7656 ;
  assign n7662 = ( ~n1209 & n7660 ) | ( ~n1209 & n7661 ) | ( n7660 & n7661 ) ;
  assign n7663 = x8 | n7661 ;
  assign n7664 = x8 | n7660 ;
  assign n7665 = ( ~n1209 & n7663 ) | ( ~n1209 & n7664 ) | ( n7663 & n7664 ) ;
  assign n7666 = ( ~n7659 & n7662 ) | ( ~n7659 & n7665 ) | ( n7662 & n7665 ) ;
  assign n7667 = n7649 & n7666 ;
  assign n7668 = ( ~n1027 & n6668 ) | ( ~n1027 & n6670 ) | ( n6668 & n6670 ) ;
  assign n7669 = ~n922 & n7068 ;
  assign n7670 = n1042 & n7074 ;
  assign n7671 = ( ~n1027 & n7074 ) | ( ~n1027 & n7670 ) | ( n7074 & n7670 ) ;
  assign n7672 = n7669 | n7671 ;
  assign n7673 = n692 & n7079 ;
  assign n7674 = ( n674 & n7079 ) | ( n674 & n7673 ) | ( n7079 & n7673 ) ;
  assign n7675 = n7672 | n7674 ;
  assign n7676 = ( n1538 & n7078 ) | ( n1538 & n7675 ) | ( n7078 & n7675 ) ;
  assign n7677 = ( x8 & ~n7675 ) | ( x8 & n7676 ) | ( ~n7675 & n7676 ) ;
  assign n7678 = ~n7676 & n7677 ;
  assign n7679 = ~n922 & n7079 ;
  assign n7680 = n1042 & n7068 ;
  assign n7681 = ( ~n1027 & n7068 ) | ( ~n1027 & n7680 ) | ( n7068 & n7680 ) ;
  assign n7682 = n7679 | n7681 ;
  assign n7683 = n7078 | n7681 ;
  assign n7684 = n7679 | n7683 ;
  assign n7685 = ( n1946 & n7682 ) | ( n1946 & n7684 ) | ( n7682 & n7684 ) ;
  assign n7686 = ~x8 & n7685 ;
  assign n7687 = n139 & n7067 ;
  assign n7688 = ( n1041 & n7067 ) | ( n1041 & n7687 ) | ( n7067 & n7687 ) ;
  assign n7689 = x8 & ~n7688 ;
  assign n7690 = n7067 | n7687 ;
  assign n7691 = x8 & ~n7690 ;
  assign n7692 = ( n1027 & n7689 ) | ( n1027 & n7691 ) | ( n7689 & n7691 ) ;
  assign n7693 = x8 & n7692 ;
  assign n7694 = ~n7685 & n7693 ;
  assign n7695 = ( n7686 & n7692 ) | ( n7686 & n7694 ) | ( n7692 & n7694 ) ;
  assign n7696 = x8 | n7675 ;
  assign n7697 = n7676 | n7696 ;
  assign n7698 = n7695 & n7697 ;
  assign n7699 = ~x8 & n7695 ;
  assign n7700 = ( n7678 & n7698 ) | ( n7678 & n7699 ) | ( n7698 & n7699 ) ;
  assign n7701 = n7668 & n7700 ;
  assign n7702 = n7700 & ~n7701 ;
  assign n7703 = ~n829 & n7079 ;
  assign n7704 = ~n922 & n7074 ;
  assign n7705 = n7703 | n7704 ;
  assign n7706 = n692 & n7068 ;
  assign n7707 = ( n674 & n7068 ) | ( n674 & n7706 ) | ( n7068 & n7706 ) ;
  assign n7708 = n7705 | n7707 ;
  assign n7709 = n7078 | n7707 ;
  assign n7710 = n7705 | n7709 ;
  assign n7711 = ( n1554 & n7708 ) | ( n1554 & n7710 ) | ( n7708 & n7710 ) ;
  assign n7712 = x8 & n7710 ;
  assign n7713 = x8 & n7708 ;
  assign n7714 = ( n1554 & n7712 ) | ( n1554 & n7713 ) | ( n7712 & n7713 ) ;
  assign n7715 = x8 & ~n7713 ;
  assign n7716 = x8 & ~n7712 ;
  assign n7717 = ( ~n1554 & n7715 ) | ( ~n1554 & n7716 ) | ( n7715 & n7716 ) ;
  assign n7718 = ( n7711 & ~n7714 ) | ( n7711 & n7717 ) | ( ~n7714 & n7717 ) ;
  assign n7719 = n7668 & ~n7700 ;
  assign n7720 = n7718 & n7719 ;
  assign n7721 = ( n7702 & n7718 ) | ( n7702 & n7720 ) | ( n7718 & n7720 ) ;
  assign n7722 = n7701 | n7721 ;
  assign n7723 = n7649 | n7666 ;
  assign n7724 = ~n7667 & n7723 ;
  assign n7725 = n7667 | n7724 ;
  assign n7726 = ( n7667 & n7722 ) | ( n7667 & n7725 ) | ( n7722 & n7725 ) ;
  assign n7727 = n7640 | n7644 ;
  assign n7728 = ~n7645 & n7727 ;
  assign n7729 = n7645 | n7728 ;
  assign n7730 = ( n7645 & n7726 ) | ( n7645 & n7729 ) | ( n7726 & n7729 ) ;
  assign n7731 = n7622 & n7730 ;
  assign n7732 = n7620 | n7731 ;
  assign n7733 = ~n7582 & n7598 ;
  assign n7734 = ( n7582 & ~n7599 ) | ( n7582 & n7733 ) | ( ~n7599 & n7733 ) ;
  assign n7735 = n7732 & n7734 ;
  assign n7736 = n7599 | n7735 ;
  assign n7737 = n7561 & ~n7579 ;
  assign n7738 = ~n7561 & n7578 ;
  assign n7739 = n7737 | n7738 ;
  assign n7740 = n7736 & n7739 ;
  assign n7741 = n7579 | n7740 ;
  assign n7742 = n7540 & ~n7558 ;
  assign n7743 = ~n7540 & n7557 ;
  assign n7744 = n7742 | n7743 ;
  assign n7745 = n7558 | n7744 ;
  assign n7746 = ( n7558 & n7741 ) | ( n7558 & n7745 ) | ( n7741 & n7745 ) ;
  assign n7747 = n7519 | n7537 ;
  assign n7748 = ~n7538 & n7747 ;
  assign n7749 = n7538 | n7748 ;
  assign n7750 = ( n7538 & n7746 ) | ( n7538 & n7749 ) | ( n7746 & n7749 ) ;
  assign n7751 = n7517 & n7750 ;
  assign n7752 = n7515 | n7751 ;
  assign n7753 = n7492 | n7752 ;
  assign n7754 = ( n7492 & n7496 ) | ( n7492 & n7753 ) | ( n7496 & n7753 ) ;
  assign n7755 = ~n7450 & n7468 ;
  assign n7756 = ( n7450 & ~n7469 ) | ( n7450 & n7755 ) | ( ~n7469 & n7755 ) ;
  assign n7757 = n7469 | n7756 ;
  assign n7758 = ( n7469 & n7754 ) | ( n7469 & n7757 ) | ( n7754 & n7757 ) ;
  assign n7759 = n7447 & n7758 ;
  assign n7760 = n7444 | n7759 ;
  assign n7761 = n6476 & n6732 ;
  assign n7762 = n6476 | n6732 ;
  assign n7763 = ~n7761 & n7762 ;
  assign n7764 = n2893 & n7068 ;
  assign n7765 = ( ~n2886 & n7068 ) | ( ~n2886 & n7764 ) | ( n7068 & n7764 ) ;
  assign n7766 = n2701 & n7074 ;
  assign n7767 = ( ~n2784 & n7074 ) | ( ~n2784 & n7766 ) | ( n7074 & n7766 ) ;
  assign n7768 = n3507 & n7079 ;
  assign n7769 = ( n3483 & n7079 ) | ( n3483 & n7768 ) | ( n7079 & n7768 ) ;
  assign n7770 = n7767 | n7769 ;
  assign n7771 = n7765 | n7770 ;
  assign n7772 = n7078 | n7771 ;
  assign n7773 = n7771 & n7772 ;
  assign n7774 = ( n3603 & n7772 ) | ( n3603 & n7773 ) | ( n7772 & n7773 ) ;
  assign n7775 = x8 & n7773 ;
  assign n7776 = x8 & n7772 ;
  assign n7777 = ( n3603 & n7775 ) | ( n3603 & n7776 ) | ( n7775 & n7776 ) ;
  assign n7778 = x8 & ~n7775 ;
  assign n7779 = x8 & ~n7776 ;
  assign n7780 = ( ~n3603 & n7778 ) | ( ~n3603 & n7779 ) | ( n7778 & n7779 ) ;
  assign n7781 = ( n7774 & ~n7777 ) | ( n7774 & n7780 ) | ( ~n7777 & n7780 ) ;
  assign n7782 = n7763 & n7781 ;
  assign n7783 = n7763 & ~n7782 ;
  assign n7784 = ~n7763 & n7781 ;
  assign n7785 = n7783 | n7784 ;
  assign n7786 = n7760 & n7785 ;
  assign n7787 = n7404 | n7422 ;
  assign n7788 = ~n7423 & n7787 ;
  assign n7789 = n7782 & n7788 ;
  assign n7790 = ( n7786 & n7788 ) | ( n7786 & n7789 ) | ( n7788 & n7789 ) ;
  assign n7791 = n7423 | n7790 ;
  assign n7792 = n7401 & n7791 ;
  assign n7793 = n7398 | n7792 ;
  assign n7794 = n7378 & n7793 ;
  assign n7795 = ~n7336 & n7352 ;
  assign n7796 = ( n7336 & ~n7353 ) | ( n7336 & n7795 ) | ( ~n7353 & n7795 ) ;
  assign n7797 = n7374 & n7796 ;
  assign n7798 = ( n7794 & n7796 ) | ( n7794 & n7797 ) | ( n7796 & n7797 ) ;
  assign n7799 = n7353 | n7798 ;
  assign n7800 = n7333 & n7799 ;
  assign n7801 = n7330 | n7800 ;
  assign n7802 = n7310 & n7801 ;
  assign n7803 = n7287 & n7307 ;
  assign n7804 = ( n7287 & n7802 ) | ( n7287 & n7803 ) | ( n7802 & n7803 ) ;
  assign n7805 = n7285 | n7804 ;
  assign n7806 = n7244 | n7262 ;
  assign n7807 = ~n7263 & n7806 ;
  assign n7808 = n7263 | n7807 ;
  assign n7809 = ( n7263 & n7805 ) | ( n7263 & n7808 ) | ( n7805 & n7808 ) ;
  assign n7810 = ~n7224 & n7240 ;
  assign n7811 = ( n7224 & ~n7241 ) | ( n7224 & n7810 ) | ( ~n7241 & n7810 ) ;
  assign n7812 = n7241 | n7811 ;
  assign n7813 = ( n7241 & n7809 ) | ( n7241 & n7812 ) | ( n7809 & n7812 ) ;
  assign n7814 = n7218 | n7813 ;
  assign n7815 = ( n7218 & n7221 ) | ( n7218 & n7814 ) | ( n7221 & n7814 ) ;
  assign n7816 = ~n7197 & n7815 ;
  assign n7817 = n7194 | n7816 ;
  assign n7818 = n7156 | n7174 ;
  assign n7819 = n7156 & n7173 ;
  assign n7820 = n7818 & ~n7819 ;
  assign n7821 = n7817 & ~n7820 ;
  assign n7822 = n7174 | n7821 ;
  assign n7823 = n7129 & ~n7154 ;
  assign n7824 = ~n7129 & n7153 ;
  assign n7825 = n7823 | n7824 ;
  assign n7826 = n7822 & n7825 ;
  assign n7827 = n7154 | n7826 ;
  assign n7828 = n7124 | n7827 ;
  assign n7829 = ( n7124 & ~n7127 ) | ( n7124 & n7828 ) | ( ~n7127 & n7828 ) ;
  assign n7830 = n7099 & n7829 ;
  assign n7831 = n7099 & ~n7830 ;
  assign n7832 = ~n7099 & n7829 ;
  assign n7833 = n7831 | n7832 ;
  assign n7834 = n182 | n460 ;
  assign n7835 = ( n418 & n5038 ) | ( n418 & ~n7834 ) | ( n5038 & ~n7834 ) ;
  assign n7836 = n7834 | n7835 ;
  assign n7837 = n5164 | n7836 ;
  assign n7838 = n608 | n648 ;
  assign n7839 = n562 | n7838 ;
  assign n7840 = n85 | n457 ;
  assign n7841 = n77 | n7840 ;
  assign n7842 = n7839 | n7841 ;
  assign n7843 = n777 | n5983 ;
  assign n7844 = n513 | n7843 ;
  assign n7845 = n7842 | n7844 ;
  assign n7846 = n176 | n331 ;
  assign n7847 = n384 | n399 ;
  assign n7848 = n7846 | n7847 ;
  assign n7849 = n237 | n388 ;
  assign n7850 = n381 | n7849 ;
  assign n7851 = n7848 | n7850 ;
  assign n7852 = n274 | n578 ;
  assign n7853 = n1303 | n7852 ;
  assign n7854 = n7851 | n7853 ;
  assign n7855 = n7845 | n7854 ;
  assign n7856 = n7837 | n7855 ;
  assign n7857 = n979 | n3425 ;
  assign n7858 = n461 | n590 ;
  assign n7859 = n631 | n7858 ;
  assign n7860 = n7857 | n7859 ;
  assign n7861 = n128 | n255 ;
  assign n7862 = n7860 | n7861 ;
  assign n7863 = n7856 | n7862 ;
  assign n7864 = n250 | n395 ;
  assign n7865 = n697 | n7864 ;
  assign n7866 = n225 | n7865 ;
  assign n7867 = n2244 | n7866 ;
  assign n7868 = n1131 | n7867 ;
  assign n7869 = n938 | n5183 ;
  assign n7870 = n217 | n7869 ;
  assign n7871 = n7868 | n7870 ;
  assign n7872 = n1028 | n3393 ;
  assign n7873 = n344 | n501 ;
  assign n7874 = n566 | n7873 ;
  assign n7875 = n7872 | n7874 ;
  assign n7876 = n234 | n895 ;
  assign n7877 = ( n197 & n263 ) | ( n197 & ~n7876 ) | ( n263 & ~n7876 ) ;
  assign n7878 = n7876 | n7877 ;
  assign n7879 = n7875 | n7878 ;
  assign n7880 = n356 | n858 ;
  assign n7881 = n278 | n491 ;
  assign n7882 = n309 | n7881 ;
  assign n7883 = n7880 | n7882 ;
  assign n7884 = n387 | n735 ;
  assign n7885 = n184 | n560 ;
  assign n7886 = n7884 | n7885 ;
  assign n7887 = n126 | n375 ;
  assign n7888 = n7886 | n7887 ;
  assign n7889 = n7883 | n7888 ;
  assign n7890 = n7879 | n7889 ;
  assign n7891 = n99 | n258 ;
  assign n7892 = n1763 | n7891 ;
  assign n7893 = n198 | n437 ;
  assign n7894 = n151 | n7893 ;
  assign n7895 = n7892 | n7894 ;
  assign n7896 = n424 | n448 ;
  assign n7897 = n1002 | n7896 ;
  assign n7898 = n702 | n7897 ;
  assign n7899 = n7895 | n7898 ;
  assign n7900 = n7890 | n7899 ;
  assign n7901 = n7871 | n7900 ;
  assign n7902 = n7863 | n7901 ;
  assign n7903 = n433 | n2156 ;
  assign n7904 = n292 | n720 ;
  assign n7905 = n689 | n7904 ;
  assign n7906 = n7903 | n7905 ;
  assign n7907 = n347 | n7906 ;
  assign n7908 = n7902 | n7907 ;
  assign n7909 = ~n6890 & n7908 ;
  assign n7910 = n6951 | n7038 ;
  assign n7911 = ( n6951 & ~n6953 ) | ( n6951 & n7910 ) | ( ~n6953 & n7910 ) ;
  assign n7912 = n6890 & ~n7908 ;
  assign n7913 = n7909 | n7912 ;
  assign n7914 = ~n7909 & n7913 ;
  assign n7915 = ( n7909 & n7911 ) | ( n7909 & ~n7914 ) | ( n7911 & ~n7914 ) ;
  assign n7916 = n341 | n901 ;
  assign n7917 = n6029 | n7916 ;
  assign n7918 = n6807 | n7917 ;
  assign n7919 = n868 | n870 ;
  assign n7920 = n1001 | n2117 ;
  assign n7921 = n821 | n7920 ;
  assign n7922 = ( n880 & ~n7919 ) | ( n880 & n7921 ) | ( ~n7919 & n7921 ) ;
  assign n7923 = n83 | n643 ;
  assign n7924 = n7919 | n7923 ;
  assign n7925 = n7922 | n7924 ;
  assign n7926 = n7918 | n7925 ;
  assign n7927 = n320 | n735 ;
  assign n7928 = n128 | n369 ;
  assign n7929 = n7927 | n7928 ;
  assign n7930 = n46 | n4145 ;
  assign n7931 = n7929 | n7930 ;
  assign n7932 = n321 | n7931 ;
  assign n7933 = n1080 | n2188 ;
  assign n7934 = n189 | n388 ;
  assign n7935 = n77 | n7934 ;
  assign n7936 = n7933 | n7935 ;
  assign n7937 = n340 | n974 ;
  assign n7938 = n7936 | n7937 ;
  assign n7939 = n7932 | n7938 ;
  assign n7940 = n215 | n2156 ;
  assign n7941 = n143 & ~n325 ;
  assign n7942 = ~n7940 & n7941 ;
  assign n7943 = ~n7939 & n7942 ;
  assign n7944 = ~n7926 & n7943 ;
  assign n7945 = n1035 | n2243 ;
  assign n7946 = n858 | n7945 ;
  assign n7947 = n7944 & ~n7946 ;
  assign n7948 = n412 | n1662 ;
  assign n7949 = n114 | n364 ;
  assign n7950 = n138 | n289 ;
  assign n7951 = n7949 | n7950 ;
  assign n7952 = n667 | n806 ;
  assign n7953 = n503 | n7952 ;
  assign n7954 = n7951 | n7953 ;
  assign n7955 = n261 | n722 ;
  assign n7956 = n112 | n168 ;
  assign n7957 = n1014 | n7956 ;
  assign n7958 = n7955 | n7957 ;
  assign n7959 = n7954 | n7958 ;
  assign n7960 = n7948 | n7959 ;
  assign n7961 = n384 | n7846 ;
  assign n7962 = n1332 | n7961 ;
  assign n7963 = n1282 | n4142 ;
  assign n7964 = n938 | n7963 ;
  assign n7965 = n7962 | n7964 ;
  assign n7966 = n581 | n959 ;
  assign n7967 = n94 | n461 ;
  assign n7968 = n7966 | n7967 ;
  assign n7969 = n7965 | n7968 ;
  assign n7970 = n7960 | n7969 ;
  assign n7971 = n124 | n479 ;
  assign n7972 = n88 | n7971 ;
  assign n7973 = n460 | n483 ;
  assign n7974 = n246 | n406 ;
  assign n7975 = n7973 | n7974 ;
  assign n7976 = n292 | n574 ;
  assign n7977 = n839 | n7976 ;
  assign n7978 = n7975 | n7977 ;
  assign n7979 = n7972 | n7978 ;
  assign n7980 = n7970 | n7979 ;
  assign n7981 = n7947 & ~n7980 ;
  assign n7982 = n223 | n303 ;
  assign n7983 = n257 | n7982 ;
  assign n7984 = n286 | n7983 ;
  assign n7985 = n363 | n623 ;
  assign n7986 = n104 | n312 ;
  assign n7987 = n7985 | n7986 ;
  assign n7988 = n7984 | n7987 ;
  assign n7989 = n496 | n7879 ;
  assign n7990 = n680 | n1690 ;
  assign n7991 = n888 | n7990 ;
  assign n7992 = n1689 | n7991 ;
  assign n7993 = n75 | n254 ;
  assign n7994 = n227 | n7993 ;
  assign n7995 = n7992 | n7994 ;
  assign n7996 = n7989 | n7995 ;
  assign n7997 = n679 | n4246 ;
  assign n7998 = n118 | n7997 ;
  assign n7999 = n171 | n2856 ;
  assign n8000 = n3375 | n7999 ;
  assign n8001 = n644 | n666 ;
  assign n8002 = ( n355 & n416 ) | ( n355 & ~n8001 ) | ( n416 & ~n8001 ) ;
  assign n8003 = n8001 | n8002 ;
  assign n8004 = n8000 | n8003 ;
  assign n8005 = n133 | n497 ;
  assign n8006 = n8004 | n8005 ;
  assign n8007 = n7998 | n8006 ;
  assign n8008 = n7996 | n8007 ;
  assign n8009 = n7988 | n8008 ;
  assign n8010 = n206 | n489 ;
  assign n8011 = n270 | n616 ;
  assign n8012 = n8010 | n8011 ;
  assign n8013 = n255 | n5946 ;
  assign n8014 = n8012 | n8013 ;
  assign n8015 = n141 | n8014 ;
  assign n8016 = n8009 | n8015 ;
  assign n8017 = n7981 & ~n8016 ;
  assign n8018 = ~n110 & n143 ;
  assign n8019 = ~n2047 & n8018 ;
  assign n8020 = ~n695 & n8019 ;
  assign n8021 = ~n7968 & n8020 ;
  assign n8022 = ~n7965 & n8021 ;
  assign n8023 = n208 | n869 ;
  assign n8024 = n7957 | n8023 ;
  assign n8025 = n126 | n245 ;
  assign n8026 = n71 | n555 ;
  assign n8027 = n349 | n381 ;
  assign n8028 = n8026 | n8027 ;
  assign n8029 = n8025 | n8028 ;
  assign n8030 = n8024 | n8029 ;
  assign n8031 = n1002 | n8030 ;
  assign n8032 = n8022 & ~n8031 ;
  assign n8033 = ~n225 & n8032 ;
  assign n8034 = n5929 | n7955 ;
  assign n8035 = n7954 | n8034 ;
  assign n8036 = n246 | n616 ;
  assign n8037 = n560 | n600 ;
  assign n8038 = n8036 | n8037 ;
  assign n8039 = n374 | n8038 ;
  assign n8040 = n697 | n1304 ;
  assign n8041 = n1637 | n8040 ;
  assign n8042 = n8039 | n8041 ;
  assign n8043 = n8035 | n8042 ;
  assign n8044 = n2853 | n8043 ;
  assign n8045 = n237 | n317 ;
  assign n8046 = n255 | n302 ;
  assign n8047 = n8045 | n8046 ;
  assign n8048 = n348 | n372 ;
  assign n8049 = n518 | n8048 ;
  assign n8050 = n8047 | n8049 ;
  assign n8051 = n413 | n8050 ;
  assign n8052 = n184 | n431 ;
  assign n8053 = n449 | n8052 ;
  assign n8054 = n661 | n3376 ;
  assign n8055 = n8053 | n8054 ;
  assign n8056 = n1146 | n1398 ;
  assign n8057 = n479 | n8056 ;
  assign n8058 = n8055 | n8057 ;
  assign n8059 = n412 | n465 ;
  assign n8060 = n203 | n206 ;
  assign n8061 = n8059 | n8060 ;
  assign n8062 = n1114 | n8061 ;
  assign n8063 = n151 | n196 ;
  assign n8064 = n424 | n443 ;
  assign n8065 = n8063 | n8064 ;
  assign n8066 = n8062 | n8065 ;
  assign n8067 = n8058 | n8066 ;
  assign n8068 = n8051 | n8067 ;
  assign n8069 = n8044 | n8068 ;
  assign n8070 = n8033 & ~n8069 ;
  assign n8071 = n987 | n4246 ;
  assign n8072 = n274 | n575 ;
  assign n8073 = n8071 | n8072 ;
  assign n8074 = n226 | n839 ;
  assign n8075 = n434 | n8074 ;
  assign n8076 = n476 | n8075 ;
  assign n8077 = n8073 | n8076 ;
  assign n8078 = n325 | n8077 ;
  assign n8079 = n155 | n8078 ;
  assign n8080 = n8070 & ~n8079 ;
  assign n8081 = n8017 | n8080 ;
  assign n8082 = n8017 & n8080 ;
  assign n8083 = n8081 & ~n8082 ;
  assign n8084 = n7908 & ~n8080 ;
  assign n8085 = ~n7908 & n8080 ;
  assign n8086 = n8084 | n8085 ;
  assign n8087 = ~n8084 & n8086 ;
  assign n8088 = n8083 & ~n8087 ;
  assign n8089 = n8083 & n8084 ;
  assign n8090 = ( n7915 & n8088 ) | ( n7915 & n8089 ) | ( n8088 & n8089 ) ;
  assign n8091 = ~n6951 & n6953 ;
  assign n8092 = ( ~n7909 & n7914 ) | ( ~n7909 & n8091 ) | ( n7914 & n8091 ) ;
  assign n8093 = ( n8088 & n8089 ) | ( n8088 & ~n8092 ) | ( n8089 & ~n8092 ) ;
  assign n8094 = ( n7050 & n8090 ) | ( n7050 & n8093 ) | ( n8090 & n8093 ) ;
  assign n8095 = ( n7054 & n8090 ) | ( n7054 & n8093 ) | ( n8090 & n8093 ) ;
  assign n8096 = ( n5216 & n8094 ) | ( n5216 & n8095 ) | ( n8094 & n8095 ) ;
  assign n8097 = ( n7915 & n8084 ) | ( n7915 & ~n8087 ) | ( n8084 & ~n8087 ) ;
  assign n8098 = ( ~n8084 & n8087 ) | ( ~n8084 & n8092 ) | ( n8087 & n8092 ) ;
  assign n8099 = ( n7054 & n8097 ) | ( n7054 & ~n8098 ) | ( n8097 & ~n8098 ) ;
  assign n8100 = n8083 | n8099 ;
  assign n8101 = ( n7050 & n8097 ) | ( n7050 & ~n8098 ) | ( n8097 & ~n8098 ) ;
  assign n8102 = n8083 | n8101 ;
  assign n8103 = ( n5216 & n8100 ) | ( n5216 & n8102 ) | ( n8100 & n8102 ) ;
  assign n8104 = ~n8096 & n8103 ;
  assign n8105 = ~x3 & x4 ;
  assign n8106 = x3 & ~x4 ;
  assign n8107 = n8105 | n8106 ;
  assign n8108 = x4 & ~x5 ;
  assign n8109 = ~x4 & x5 ;
  assign n8110 = n8108 | n8109 ;
  assign n8111 = x2 & ~x3 ;
  assign n8112 = ~x2 & x3 ;
  assign n8113 = n8111 | n8112 ;
  assign n8114 = n8110 & ~n8113 ;
  assign n8115 = ~n8107 & n8114 ;
  assign n8116 = n7907 & n8115 ;
  assign n8117 = ( n7902 & n8115 ) | ( n7902 & n8116 ) | ( n8115 & n8116 ) ;
  assign n8118 = n8107 & ~n8113 ;
  assign n8119 = n8079 & n8118 ;
  assign n8120 = ( ~n8070 & n8118 ) | ( ~n8070 & n8119 ) | ( n8118 & n8119 ) ;
  assign n8121 = n8117 | n8120 ;
  assign n8122 = ~n8110 & n8113 ;
  assign n8123 = ~n8017 & n8122 ;
  assign n8124 = n8121 | n8123 ;
  assign n8125 = n8110 & n8113 ;
  assign n8126 = n8121 | n8125 ;
  assign n8127 = n8123 | n8126 ;
  assign n8128 = ( n8104 & n8124 ) | ( n8104 & n8127 ) | ( n8124 & n8127 ) ;
  assign n8129 = x5 & n8127 ;
  assign n8130 = x5 & n8124 ;
  assign n8131 = ( n8104 & n8129 ) | ( n8104 & n8130 ) | ( n8129 & n8130 ) ;
  assign n8132 = x5 & ~n8130 ;
  assign n8133 = x5 & ~n8129 ;
  assign n8134 = ( ~n8104 & n8132 ) | ( ~n8104 & n8133 ) | ( n8132 & n8133 ) ;
  assign n8135 = ( n8128 & ~n8131 ) | ( n8128 & n8134 ) | ( ~n8131 & n8134 ) ;
  assign n8136 = n7832 & n8135 ;
  assign n8137 = ( n7831 & n8135 ) | ( n7831 & n8136 ) | ( n8135 & n8136 ) ;
  assign n8138 = n7833 & ~n8137 ;
  assign n8139 = ~n7832 & n8135 ;
  assign n8140 = ~n7831 & n8139 ;
  assign n8141 = n8138 | n8140 ;
  assign n8142 = ~n7127 & n7827 ;
  assign n8143 = n7127 | n8142 ;
  assign n8146 = n7915 & ~n8086 ;
  assign n8147 = n8086 | n8092 ;
  assign n8148 = ( n7050 & n8146 ) | ( n7050 & ~n8147 ) | ( n8146 & ~n8147 ) ;
  assign n8149 = ( n7054 & n8146 ) | ( n7054 & ~n8147 ) | ( n8146 & ~n8147 ) ;
  assign n8150 = ( n5216 & n8148 ) | ( n5216 & n8149 ) | ( n8148 & n8149 ) ;
  assign n8151 = ( n7054 & n7915 ) | ( n7054 & ~n8092 ) | ( n7915 & ~n8092 ) ;
  assign n8152 = n8086 & ~n8151 ;
  assign n8153 = ( n7050 & n7915 ) | ( n7050 & ~n8092 ) | ( n7915 & ~n8092 ) ;
  assign n8154 = n8086 & ~n8153 ;
  assign n8155 = ( ~n5216 & n8152 ) | ( ~n5216 & n8154 ) | ( n8152 & n8154 ) ;
  assign n8156 = n8150 | n8155 ;
  assign n8157 = n6889 & n8115 ;
  assign n8158 = ( ~n6884 & n8115 ) | ( ~n6884 & n8157 ) | ( n8115 & n8157 ) ;
  assign n8159 = n7907 & n8118 ;
  assign n8160 = ( n7902 & n8118 ) | ( n7902 & n8159 ) | ( n8118 & n8159 ) ;
  assign n8161 = n8079 & n8122 ;
  assign n8162 = ( ~n8070 & n8122 ) | ( ~n8070 & n8161 ) | ( n8122 & n8161 ) ;
  assign n8163 = n8160 | n8162 ;
  assign n8164 = n8158 | n8163 ;
  assign n8165 = n8125 | n8164 ;
  assign n8166 = ( ~n8156 & n8164 ) | ( ~n8156 & n8165 ) | ( n8164 & n8165 ) ;
  assign n8167 = ~x5 & n8165 ;
  assign n8168 = ~x5 & n8164 ;
  assign n8169 = ( ~n8156 & n8167 ) | ( ~n8156 & n8168 ) | ( n8167 & n8168 ) ;
  assign n8170 = x5 | n8167 ;
  assign n8171 = x5 | n8168 ;
  assign n8172 = ( ~n8156 & n8170 ) | ( ~n8156 & n8171 ) | ( n8170 & n8171 ) ;
  assign n8173 = ( ~n8166 & n8169 ) | ( ~n8166 & n8172 ) | ( n8169 & n8172 ) ;
  assign n8144 = n7127 & n7827 ;
  assign n8174 = n8144 & n8173 ;
  assign n8175 = ( ~n8143 & n8173 ) | ( ~n8143 & n8174 ) | ( n8173 & n8174 ) ;
  assign n8145 = n8143 & ~n8144 ;
  assign n8176 = n8145 | n8175 ;
  assign n8177 = ~n8144 & n8173 ;
  assign n8178 = n8143 & n8177 ;
  assign n8179 = n8176 & ~n8178 ;
  assign n8180 = n7822 & ~n7826 ;
  assign n8181 = n7825 & ~n7826 ;
  assign n8182 = n8180 | n8181 ;
  assign n8183 = n7911 & ~n7913 ;
  assign n8184 = n7913 | n8091 ;
  assign n8185 = ( n7050 & n8183 ) | ( n7050 & ~n8184 ) | ( n8183 & ~n8184 ) ;
  assign n8186 = ( n7054 & n8183 ) | ( n7054 & ~n8184 ) | ( n8183 & ~n8184 ) ;
  assign n8187 = ( n5216 & n8185 ) | ( n5216 & n8186 ) | ( n8185 & n8186 ) ;
  assign n8188 = ( n7054 & n7911 ) | ( n7054 & ~n8091 ) | ( n7911 & ~n8091 ) ;
  assign n8189 = n7913 & ~n8188 ;
  assign n8190 = ( n7050 & n7911 ) | ( n7050 & ~n8091 ) | ( n7911 & ~n8091 ) ;
  assign n8191 = n7913 & ~n8190 ;
  assign n8192 = ( ~n5216 & n8189 ) | ( ~n5216 & n8191 ) | ( n8189 & n8191 ) ;
  assign n8193 = n8187 | n8192 ;
  assign n8194 = n6950 & n8115 ;
  assign n8195 = n6889 & n8118 ;
  assign n8196 = ( ~n6884 & n8118 ) | ( ~n6884 & n8195 ) | ( n8118 & n8195 ) ;
  assign n8197 = n8194 | n8196 ;
  assign n8198 = n7907 & n8122 ;
  assign n8199 = ( n7902 & n8122 ) | ( n7902 & n8198 ) | ( n8122 & n8198 ) ;
  assign n8200 = n8197 | n8199 ;
  assign n8201 = n8125 | n8199 ;
  assign n8202 = n8197 | n8201 ;
  assign n8203 = ( ~n8193 & n8200 ) | ( ~n8193 & n8202 ) | ( n8200 & n8202 ) ;
  assign n8204 = ~x5 & n8202 ;
  assign n8205 = ~x5 & n8200 ;
  assign n8206 = ( ~n8193 & n8204 ) | ( ~n8193 & n8205 ) | ( n8204 & n8205 ) ;
  assign n8207 = x5 | n8205 ;
  assign n8208 = x5 | n8204 ;
  assign n8209 = ( ~n8193 & n8207 ) | ( ~n8193 & n8208 ) | ( n8207 & n8208 ) ;
  assign n8210 = ( ~n8203 & n8206 ) | ( ~n8203 & n8209 ) | ( n8206 & n8209 ) ;
  assign n8211 = n8182 & n8210 ;
  assign n8212 = n8182 & ~n8211 ;
  assign n8213 = ~n8182 & n8210 ;
  assign n8214 = n8212 | n8213 ;
  assign n8215 = n7817 & ~n7821 ;
  assign n8216 = n7820 | n7821 ;
  assign n8217 = ~n8215 & n8216 ;
  assign n8218 = n6950 & n8118 ;
  assign n8219 = n7036 & n8115 ;
  assign n8220 = ( n7023 & n8115 ) | ( n7023 & n8219 ) | ( n8115 & n8219 ) ;
  assign n8221 = n8218 | n8220 ;
  assign n8222 = n6889 & n8122 ;
  assign n8223 = ( ~n6884 & n8122 ) | ( ~n6884 & n8222 ) | ( n8122 & n8222 ) ;
  assign n8224 = n8221 | n8223 ;
  assign n8225 = n8125 | n8223 ;
  assign n8226 = n8221 | n8225 ;
  assign n8227 = ( ~n7061 & n8224 ) | ( ~n7061 & n8226 ) | ( n8224 & n8226 ) ;
  assign n8228 = ~x5 & n8226 ;
  assign n8229 = ~x5 & n8224 ;
  assign n8230 = ( ~n7061 & n8228 ) | ( ~n7061 & n8229 ) | ( n8228 & n8229 ) ;
  assign n8231 = x5 | n8229 ;
  assign n8232 = x5 | n8228 ;
  assign n8233 = ( ~n7061 & n8231 ) | ( ~n7061 & n8232 ) | ( n8231 & n8232 ) ;
  assign n8234 = ( ~n8227 & n8230 ) | ( ~n8227 & n8233 ) | ( n8230 & n8233 ) ;
  assign n8235 = ~n8217 & n8234 ;
  assign n8236 = n8217 | n8235 ;
  assign n8237 = n8217 & n8234 ;
  assign n8238 = n8236 & ~n8237 ;
  assign n8239 = n7815 & ~n7816 ;
  assign n8240 = n7197 | n7816 ;
  assign n8241 = ~n8239 & n8240 ;
  assign n8242 = ~n6091 & n8115 ;
  assign n8243 = n7036 & n8118 ;
  assign n8244 = ( n7023 & n8118 ) | ( n7023 & n8243 ) | ( n8118 & n8243 ) ;
  assign n8245 = n8242 | n8244 ;
  assign n8246 = n6950 & n8122 ;
  assign n8247 = n8245 | n8246 ;
  assign n8248 = n8125 | n8247 ;
  assign n8249 = ( ~n7107 & n8247 ) | ( ~n7107 & n8248 ) | ( n8247 & n8248 ) ;
  assign n8250 = ~x5 & n8248 ;
  assign n8251 = ~x5 & n8247 ;
  assign n8252 = ( ~n7107 & n8250 ) | ( ~n7107 & n8251 ) | ( n8250 & n8251 ) ;
  assign n8253 = x5 | n8250 ;
  assign n8254 = x5 | n8251 ;
  assign n8255 = ( ~n7107 & n8253 ) | ( ~n7107 & n8254 ) | ( n8253 & n8254 ) ;
  assign n8256 = ( ~n8249 & n8252 ) | ( ~n8249 & n8255 ) | ( n8252 & n8255 ) ;
  assign n8257 = ~n8241 & n8256 ;
  assign n8258 = n8241 | n8257 ;
  assign n8259 = n8241 & n8256 ;
  assign n8260 = n8258 & ~n8259 ;
  assign n8261 = n7221 & n7813 ;
  assign n8262 = n7221 & ~n8261 ;
  assign n8265 = n5857 & n8115 ;
  assign n8266 = ( ~n5899 & n8115 ) | ( ~n5899 & n8265 ) | ( n8115 & n8265 ) ;
  assign n8267 = ~n6091 & n8118 ;
  assign n8268 = n7036 & n8122 ;
  assign n8269 = ( n7023 & n8122 ) | ( n7023 & n8268 ) | ( n8122 & n8268 ) ;
  assign n8270 = n8267 | n8269 ;
  assign n8271 = n8266 | n8270 ;
  assign n8272 = n8125 | n8271 ;
  assign n8273 = ( n7136 & n8271 ) | ( n7136 & n8272 ) | ( n8271 & n8272 ) ;
  assign n8274 = x5 & n8272 ;
  assign n8275 = x5 & n8271 ;
  assign n8276 = ( n7136 & n8274 ) | ( n7136 & n8275 ) | ( n8274 & n8275 ) ;
  assign n8277 = x5 & ~n8274 ;
  assign n8278 = x5 & ~n8275 ;
  assign n8279 = ( ~n7136 & n8277 ) | ( ~n7136 & n8278 ) | ( n8277 & n8278 ) ;
  assign n8280 = ( n8273 & ~n8276 ) | ( n8273 & n8279 ) | ( ~n8276 & n8279 ) ;
  assign n8263 = ~n7221 & n7813 ;
  assign n8281 = n8263 & n8280 ;
  assign n8282 = ( n8262 & n8280 ) | ( n8262 & n8281 ) | ( n8280 & n8281 ) ;
  assign n8264 = n8262 | n8263 ;
  assign n8283 = n8264 & ~n8282 ;
  assign n8284 = ~n8263 & n8280 ;
  assign n8285 = ~n8262 & n8284 ;
  assign n8286 = n8283 | n8285 ;
  assign n8287 = n7809 & n7811 ;
  assign n8288 = n7809 | n7811 ;
  assign n8289 = ~n8287 & n8288 ;
  assign n8290 = n5857 & n8118 ;
  assign n8291 = ( ~n5899 & n8118 ) | ( ~n5899 & n8290 ) | ( n8118 & n8290 ) ;
  assign n8292 = ~n6091 & n8122 ;
  assign n8293 = n5997 & n8115 ;
  assign n8294 = ( n5979 & n8115 ) | ( n5979 & n8293 ) | ( n8115 & n8293 ) ;
  assign n8295 = n8292 | n8294 ;
  assign n8296 = n8291 | n8295 ;
  assign n8297 = n8125 | n8296 ;
  assign n8298 = n8296 & n8297 ;
  assign n8299 = ( n6108 & n8297 ) | ( n6108 & n8298 ) | ( n8297 & n8298 ) ;
  assign n8300 = x5 & n8298 ;
  assign n8301 = x5 & n8297 ;
  assign n8302 = ( n6108 & n8300 ) | ( n6108 & n8301 ) | ( n8300 & n8301 ) ;
  assign n8303 = x5 & ~n8300 ;
  assign n8304 = x5 & ~n8301 ;
  assign n8305 = ( ~n6108 & n8303 ) | ( ~n6108 & n8304 ) | ( n8303 & n8304 ) ;
  assign n8306 = ( n8299 & ~n8302 ) | ( n8299 & n8305 ) | ( ~n8302 & n8305 ) ;
  assign n8307 = n8289 & n8306 ;
  assign n8308 = n7805 & n7807 ;
  assign n8309 = n7805 | n7807 ;
  assign n8310 = ~n8308 & n8309 ;
  assign n8311 = n5108 & n8115 ;
  assign n8312 = n5997 & n8118 ;
  assign n8313 = ( n5979 & n8118 ) | ( n5979 & n8312 ) | ( n8118 & n8312 ) ;
  assign n8314 = n8311 | n8313 ;
  assign n8315 = n5857 & n8122 ;
  assign n8316 = ( ~n5899 & n8122 ) | ( ~n5899 & n8315 ) | ( n8122 & n8315 ) ;
  assign n8317 = n8314 | n8316 ;
  assign n8318 = n8125 | n8317 ;
  assign n8319 = n8317 & n8318 ;
  assign n8320 = ( ~n6151 & n8318 ) | ( ~n6151 & n8319 ) | ( n8318 & n8319 ) ;
  assign n8321 = ~x5 & n8319 ;
  assign n8322 = ~x5 & n8318 ;
  assign n8323 = ( ~n6151 & n8321 ) | ( ~n6151 & n8322 ) | ( n8321 & n8322 ) ;
  assign n8324 = x5 | n8321 ;
  assign n8325 = x5 | n8322 ;
  assign n8326 = ( ~n6151 & n8324 ) | ( ~n6151 & n8325 ) | ( n8324 & n8325 ) ;
  assign n8327 = ( ~n8320 & n8323 ) | ( ~n8320 & n8326 ) | ( n8323 & n8326 ) ;
  assign n8328 = n8310 & n8327 ;
  assign n8329 = n8310 & ~n8328 ;
  assign n8330 = ~n8310 & n8327 ;
  assign n8331 = n8329 | n8330 ;
  assign n8332 = n7287 | n7307 ;
  assign n8333 = n7802 | n8332 ;
  assign n8334 = ~n7804 & n8333 ;
  assign n8335 = n5117 & n8115 ;
  assign n8336 = ( ~n5037 & n8115 ) | ( ~n5037 & n8335 ) | ( n8115 & n8335 ) ;
  assign n8337 = n5108 & n8118 ;
  assign n8338 = n5997 & n8122 ;
  assign n8339 = ( n5979 & n8122 ) | ( n5979 & n8338 ) | ( n8122 & n8338 ) ;
  assign n8340 = n8337 | n8339 ;
  assign n8341 = n8336 | n8340 ;
  assign n8342 = n8125 | n8341 ;
  assign n8343 = ( n6181 & n8341 ) | ( n6181 & n8342 ) | ( n8341 & n8342 ) ;
  assign n8344 = x5 & n8342 ;
  assign n8345 = x5 & n8341 ;
  assign n8346 = ( n6181 & n8344 ) | ( n6181 & n8345 ) | ( n8344 & n8345 ) ;
  assign n8347 = x5 & ~n8344 ;
  assign n8348 = x5 & ~n8345 ;
  assign n8349 = ( ~n6181 & n8347 ) | ( ~n6181 & n8348 ) | ( n8347 & n8348 ) ;
  assign n8350 = ( n8343 & ~n8346 ) | ( n8343 & n8349 ) | ( ~n8346 & n8349 ) ;
  assign n8351 = n8334 & n8350 ;
  assign n8352 = ~n7310 & n7801 ;
  assign n8353 = n7310 & ~n7801 ;
  assign n8354 = n8352 | n8353 ;
  assign n8355 = n5117 & n8118 ;
  assign n8356 = ( ~n5037 & n8118 ) | ( ~n5037 & n8355 ) | ( n8118 & n8355 ) ;
  assign n8357 = n5108 & n8122 ;
  assign n8358 = n5192 & n8115 ;
  assign n8359 = ( n5179 & n8115 ) | ( n5179 & n8358 ) | ( n8115 & n8358 ) ;
  assign n8360 = n8357 | n8359 ;
  assign n8361 = n8356 | n8360 ;
  assign n8362 = n8125 | n8361 ;
  assign n8363 = ( ~n5220 & n8361 ) | ( ~n5220 & n8362 ) | ( n8361 & n8362 ) ;
  assign n8364 = ~x5 & n8362 ;
  assign n8365 = ~x5 & n8361 ;
  assign n8366 = ( ~n5220 & n8364 ) | ( ~n5220 & n8365 ) | ( n8364 & n8365 ) ;
  assign n8367 = x5 | n8364 ;
  assign n8368 = x5 | n8365 ;
  assign n8369 = ( ~n5220 & n8367 ) | ( ~n5220 & n8368 ) | ( n8367 & n8368 ) ;
  assign n8370 = ( ~n8363 & n8366 ) | ( ~n8363 & n8369 ) | ( n8366 & n8369 ) ;
  assign n8371 = n8354 & n8370 ;
  assign n8372 = n8354 | n8370 ;
  assign n8373 = ~n8371 & n8372 ;
  assign n8374 = ~n7333 & n7799 ;
  assign n8375 = n7333 & ~n7799 ;
  assign n8376 = n8374 | n8375 ;
  assign n8377 = n4245 & n8115 ;
  assign n8378 = ( n4303 & n8115 ) | ( n4303 & n8377 ) | ( n8115 & n8377 ) ;
  assign n8379 = n5192 & n8118 ;
  assign n8380 = ( n5179 & n8118 ) | ( n5179 & n8379 ) | ( n8118 & n8379 ) ;
  assign n8381 = n8378 | n8380 ;
  assign n8382 = n5117 & n8122 ;
  assign n8383 = ( ~n5037 & n8122 ) | ( ~n5037 & n8382 ) | ( n8122 & n8382 ) ;
  assign n8384 = n8381 | n8383 ;
  assign n8385 = n8125 | n8383 ;
  assign n8386 = n8381 | n8385 ;
  assign n8387 = ( ~n5270 & n8384 ) | ( ~n5270 & n8386 ) | ( n8384 & n8386 ) ;
  assign n8388 = ~x5 & n8386 ;
  assign n8389 = ~x5 & n8384 ;
  assign n8390 = ( ~n5270 & n8388 ) | ( ~n5270 & n8389 ) | ( n8388 & n8389 ) ;
  assign n8391 = x5 | n8389 ;
  assign n8392 = x5 | n8388 ;
  assign n8393 = ( ~n5270 & n8391 ) | ( ~n5270 & n8392 ) | ( n8391 & n8392 ) ;
  assign n8394 = ( ~n8387 & n8390 ) | ( ~n8387 & n8393 ) | ( n8390 & n8393 ) ;
  assign n8395 = n8376 & n8394 ;
  assign n8396 = n7374 | n7796 ;
  assign n8397 = n7794 | n8396 ;
  assign n8398 = ~n7798 & n8397 ;
  assign n8399 = n4396 & n8115 ;
  assign n8400 = n4245 & n8118 ;
  assign n8401 = ( n4303 & n8118 ) | ( n4303 & n8400 ) | ( n8118 & n8400 ) ;
  assign n8402 = n8399 | n8401 ;
  assign n8403 = n5192 & n8122 ;
  assign n8404 = ( n5179 & n8122 ) | ( n5179 & n8403 ) | ( n8122 & n8403 ) ;
  assign n8406 = n8125 | n8404 ;
  assign n8407 = n8402 | n8406 ;
  assign n8405 = n8402 | n8404 ;
  assign n8408 = n8405 & n8407 ;
  assign n8409 = ( n5306 & n8407 ) | ( n5306 & n8408 ) | ( n8407 & n8408 ) ;
  assign n8410 = x5 & n8408 ;
  assign n8411 = x5 & n8407 ;
  assign n8412 = ( n5306 & n8410 ) | ( n5306 & n8411 ) | ( n8410 & n8411 ) ;
  assign n8413 = x5 & ~n8410 ;
  assign n8414 = x5 & ~n8411 ;
  assign n8415 = ( ~n5306 & n8413 ) | ( ~n5306 & n8414 ) | ( n8413 & n8414 ) ;
  assign n8416 = ( n8409 & ~n8412 ) | ( n8409 & n8415 ) | ( ~n8412 & n8415 ) ;
  assign n8417 = n8398 & n8416 ;
  assign n8418 = n8398 | n8416 ;
  assign n8419 = ~n8417 & n8418 ;
  assign n8420 = n7378 | n7793 ;
  assign n8421 = ~n7794 & n8420 ;
  assign n8422 = ~n4429 & n8115 ;
  assign n8423 = n4396 & n8118 ;
  assign n8424 = n8422 | n8423 ;
  assign n8425 = n4245 & n8122 ;
  assign n8426 = ( n4303 & n8122 ) | ( n4303 & n8425 ) | ( n8122 & n8425 ) ;
  assign n8428 = n8125 | n8426 ;
  assign n8429 = n8424 | n8428 ;
  assign n8427 = n8424 | n8426 ;
  assign n8430 = n8427 & n8429 ;
  assign n8431 = ( n4455 & n8429 ) | ( n4455 & n8430 ) | ( n8429 & n8430 ) ;
  assign n8432 = x5 & n8430 ;
  assign n8433 = x5 & n8429 ;
  assign n8434 = ( n4455 & n8432 ) | ( n4455 & n8433 ) | ( n8432 & n8433 ) ;
  assign n8435 = x5 & ~n8432 ;
  assign n8436 = x5 & ~n8433 ;
  assign n8437 = ( ~n4455 & n8435 ) | ( ~n4455 & n8436 ) | ( n8435 & n8436 ) ;
  assign n8438 = ( n8431 & ~n8434 ) | ( n8431 & n8437 ) | ( ~n8434 & n8437 ) ;
  assign n8439 = n8421 & n8438 ;
  assign n8440 = n8421 & ~n8439 ;
  assign n8441 = ~n8421 & n8438 ;
  assign n8442 = n8440 | n8441 ;
  assign n8443 = n7401 | n7791 ;
  assign n8444 = ~n7792 & n8443 ;
  assign n8445 = ~n4429 & n8118 ;
  assign n8446 = n8115 | n8118 ;
  assign n8447 = ( ~n4429 & n8115 ) | ( ~n4429 & n8446 ) | ( n8115 & n8446 ) ;
  assign n8448 = ( n4206 & n8445 ) | ( n4206 & n8447 ) | ( n8445 & n8447 ) ;
  assign n8449 = n4396 & n8122 ;
  assign n8451 = n8125 | n8449 ;
  assign n8452 = n8448 | n8451 ;
  assign n8450 = n8448 | n8449 ;
  assign n8453 = n8450 & n8452 ;
  assign n8454 = ( ~n4501 & n8452 ) | ( ~n4501 & n8453 ) | ( n8452 & n8453 ) ;
  assign n8455 = ~x5 & n8453 ;
  assign n8456 = ~x5 & n8452 ;
  assign n8457 = ( ~n4501 & n8455 ) | ( ~n4501 & n8456 ) | ( n8455 & n8456 ) ;
  assign n8458 = x5 | n8455 ;
  assign n8459 = x5 | n8456 ;
  assign n8460 = ( ~n4501 & n8458 ) | ( ~n4501 & n8459 ) | ( n8458 & n8459 ) ;
  assign n8461 = ( ~n8454 & n8457 ) | ( ~n8454 & n8460 ) | ( n8457 & n8460 ) ;
  assign n8462 = n8444 & n8461 ;
  assign n8463 = n8444 & ~n8462 ;
  assign n8464 = ~n8444 & n8461 ;
  assign n8465 = n8463 | n8464 ;
  assign n8466 = n7782 | n7788 ;
  assign n8467 = n7786 | n8466 ;
  assign n8468 = ~n7790 & n8467 ;
  assign n8469 = n4206 & n8118 ;
  assign n8470 = ~n4429 & n8122 ;
  assign n8471 = n3439 & n8115 ;
  assign n8472 = ( ~n3420 & n8115 ) | ( ~n3420 & n8471 ) | ( n8115 & n8471 ) ;
  assign n8473 = n8470 | n8472 ;
  assign n8474 = n8469 | n8473 ;
  assign n8475 = n8125 | n8469 ;
  assign n8476 = n8473 | n8475 ;
  assign n8477 = ( ~n4527 & n8474 ) | ( ~n4527 & n8476 ) | ( n8474 & n8476 ) ;
  assign n8478 = ~x5 & n8476 ;
  assign n8479 = ~x5 & n8474 ;
  assign n8480 = ( ~n4527 & n8478 ) | ( ~n4527 & n8479 ) | ( n8478 & n8479 ) ;
  assign n8481 = x5 | n8479 ;
  assign n8482 = x5 | n8478 ;
  assign n8483 = ( ~n4527 & n8481 ) | ( ~n4527 & n8482 ) | ( n8481 & n8482 ) ;
  assign n8484 = ( ~n8477 & n8480 ) | ( ~n8477 & n8483 ) | ( n8480 & n8483 ) ;
  assign n8485 = n8468 & n8484 ;
  assign n8486 = n7785 & ~n7786 ;
  assign n8487 = n7760 & ~n7785 ;
  assign n8488 = n8486 | n8487 ;
  assign n8489 = n4206 & n8122 ;
  assign n8490 = n3386 & n8115 ;
  assign n8491 = n3439 & n8118 ;
  assign n8492 = ( ~n3420 & n8118 ) | ( ~n3420 & n8491 ) | ( n8118 & n8491 ) ;
  assign n8493 = n8490 | n8492 ;
  assign n8494 = n8489 | n8493 ;
  assign n8495 = n8125 | n8489 ;
  assign n8496 = n8493 | n8495 ;
  assign n8497 = ( ~n4220 & n8494 ) | ( ~n4220 & n8496 ) | ( n8494 & n8496 ) ;
  assign n8498 = ~x5 & n8496 ;
  assign n8499 = ~x5 & n8494 ;
  assign n8500 = ( ~n4220 & n8498 ) | ( ~n4220 & n8499 ) | ( n8498 & n8499 ) ;
  assign n8501 = x5 | n8499 ;
  assign n8502 = x5 | n8498 ;
  assign n8503 = ( ~n4220 & n8501 ) | ( ~n4220 & n8502 ) | ( n8501 & n8502 ) ;
  assign n8504 = ( ~n8497 & n8500 ) | ( ~n8497 & n8503 ) | ( n8500 & n8503 ) ;
  assign n8505 = n8487 & n8504 ;
  assign n8506 = ( n8486 & n8504 ) | ( n8486 & n8505 ) | ( n8504 & n8505 ) ;
  assign n8507 = n8488 & ~n8506 ;
  assign n8508 = ~n8487 & n8504 ;
  assign n8509 = ~n8486 & n8508 ;
  assign n8510 = n8507 | n8509 ;
  assign n8511 = n7758 & ~n7759 ;
  assign n8512 = n7447 & ~n7759 ;
  assign n8513 = n8511 | n8512 ;
  assign n8514 = n3386 & n8118 ;
  assign n8515 = n3507 & n8115 ;
  assign n8516 = ( n3483 & n8115 ) | ( n3483 & n8515 ) | ( n8115 & n8515 ) ;
  assign n8517 = n3439 & n8122 ;
  assign n8518 = ( ~n3420 & n8122 ) | ( ~n3420 & n8517 ) | ( n8122 & n8517 ) ;
  assign n8519 = n8516 | n8518 ;
  assign n8520 = n8514 | n8519 ;
  assign n8521 = n8125 | n8520 ;
  assign n8522 = ( ~n3530 & n8520 ) | ( ~n3530 & n8521 ) | ( n8520 & n8521 ) ;
  assign n8523 = ~x5 & n8521 ;
  assign n8524 = ~x5 & n8520 ;
  assign n8525 = ( ~n3530 & n8523 ) | ( ~n3530 & n8524 ) | ( n8523 & n8524 ) ;
  assign n8526 = x5 | n8523 ;
  assign n8527 = x5 | n8524 ;
  assign n8528 = ( ~n3530 & n8526 ) | ( ~n3530 & n8527 ) | ( n8526 & n8527 ) ;
  assign n8529 = ( ~n8522 & n8525 ) | ( ~n8522 & n8528 ) | ( n8525 & n8528 ) ;
  assign n8530 = n8513 & n8529 ;
  assign n8531 = n8513 & ~n8530 ;
  assign n8532 = ~n8513 & n8529 ;
  assign n8533 = n8531 | n8532 ;
  assign n8534 = n7754 & n7756 ;
  assign n8535 = n7754 | n7756 ;
  assign n8536 = ~n8534 & n8535 ;
  assign n8537 = n2893 & n8115 ;
  assign n8538 = ( ~n2886 & n8115 ) | ( ~n2886 & n8537 ) | ( n8115 & n8537 ) ;
  assign n8539 = n3507 & n8118 ;
  assign n8540 = ( n3483 & n8118 ) | ( n3483 & n8539 ) | ( n8118 & n8539 ) ;
  assign n8541 = n8538 | n8540 ;
  assign n8542 = n3386 & n8122 ;
  assign n8544 = n8125 | n8542 ;
  assign n8545 = n8541 | n8544 ;
  assign n8543 = n8541 | n8542 ;
  assign n8546 = n8543 & n8545 ;
  assign n8547 = ( ~n3568 & n8545 ) | ( ~n3568 & n8546 ) | ( n8545 & n8546 ) ;
  assign n8548 = ~x5 & n8546 ;
  assign n8549 = ~x5 & n8545 ;
  assign n8550 = ( ~n3568 & n8548 ) | ( ~n3568 & n8549 ) | ( n8548 & n8549 ) ;
  assign n8551 = x5 | n8548 ;
  assign n8552 = x5 | n8549 ;
  assign n8553 = ( ~n3568 & n8551 ) | ( ~n3568 & n8552 ) | ( n8551 & n8552 ) ;
  assign n8554 = ( ~n8547 & n8550 ) | ( ~n8547 & n8553 ) | ( n8550 & n8553 ) ;
  assign n8555 = n8536 & n8554 ;
  assign n8556 = n7517 | n7750 ;
  assign n8557 = ~n7751 & n8556 ;
  assign n8558 = n2691 & n8115 ;
  assign n8559 = ( n2678 & n8115 ) | ( n2678 & n8558 ) | ( n8115 & n8558 ) ;
  assign n8560 = n2701 & n8118 ;
  assign n8561 = ( ~n2784 & n8118 ) | ( ~n2784 & n8560 ) | ( n8118 & n8560 ) ;
  assign n8562 = n8559 | n8561 ;
  assign n8563 = n2893 & n8122 ;
  assign n8564 = ( ~n2886 & n8122 ) | ( ~n2886 & n8563 ) | ( n8122 & n8563 ) ;
  assign n8565 = n8562 | n8564 ;
  assign n8566 = n8125 | n8565 ;
  assign n8567 = n8565 & n8566 ;
  assign n8568 = ( ~n2914 & n8566 ) | ( ~n2914 & n8567 ) | ( n8566 & n8567 ) ;
  assign n8569 = ~x5 & n8567 ;
  assign n8570 = ~x5 & n8566 ;
  assign n8571 = ( ~n2914 & n8569 ) | ( ~n2914 & n8570 ) | ( n8569 & n8570 ) ;
  assign n8572 = x5 | n8569 ;
  assign n8573 = x5 | n8570 ;
  assign n8574 = ( ~n2914 & n8572 ) | ( ~n2914 & n8573 ) | ( n8572 & n8573 ) ;
  assign n8575 = ( ~n8568 & n8571 ) | ( ~n8568 & n8574 ) | ( n8571 & n8574 ) ;
  assign n8576 = n8557 & n8575 ;
  assign n8577 = n8557 & ~n8576 ;
  assign n8578 = ~n8557 & n8575 ;
  assign n8579 = n8577 | n8578 ;
  assign n8580 = n7746 & n7748 ;
  assign n8581 = n7746 | n7748 ;
  assign n8582 = ~n8580 & n8581 ;
  assign n8583 = n2701 & n8122 ;
  assign n8584 = ( ~n2784 & n8122 ) | ( ~n2784 & n8583 ) | ( n8122 & n8583 ) ;
  assign n8585 = n2691 & n8118 ;
  assign n8586 = ( n2678 & n8118 ) | ( n2678 & n8585 ) | ( n8118 & n8585 ) ;
  assign n8587 = n8584 | n8586 ;
  assign n8588 = n2199 & n8115 ;
  assign n8589 = ( ~n2185 & n8115 ) | ( ~n2185 & n8588 ) | ( n8115 & n8588 ) ;
  assign n8590 = n8587 | n8589 ;
  assign n8591 = n8125 | n8589 ;
  assign n8592 = n8587 | n8591 ;
  assign n8593 = ( n2960 & n8590 ) | ( n2960 & n8592 ) | ( n8590 & n8592 ) ;
  assign n8594 = x5 & n8592 ;
  assign n8595 = x5 & n8590 ;
  assign n8596 = ( n2960 & n8594 ) | ( n2960 & n8595 ) | ( n8594 & n8595 ) ;
  assign n8597 = x5 & ~n8595 ;
  assign n8598 = x5 & ~n8594 ;
  assign n8599 = ( ~n2960 & n8597 ) | ( ~n2960 & n8598 ) | ( n8597 & n8598 ) ;
  assign n8600 = ( n8593 & ~n8596 ) | ( n8593 & n8599 ) | ( ~n8596 & n8599 ) ;
  assign n8601 = n8582 & n8600 ;
  assign n8602 = n7741 & n7744 ;
  assign n8603 = n7741 & ~n8602 ;
  assign n8606 = n2090 & n8115 ;
  assign n8607 = ( ~n2082 & n8115 ) | ( ~n2082 & n8606 ) | ( n8115 & n8606 ) ;
  assign n8608 = n2691 & n8122 ;
  assign n8609 = ( n2678 & n8122 ) | ( n2678 & n8608 ) | ( n8122 & n8608 ) ;
  assign n8610 = n2199 & n8118 ;
  assign n8611 = ( ~n2185 & n8118 ) | ( ~n2185 & n8610 ) | ( n8118 & n8610 ) ;
  assign n8612 = n8609 | n8611 ;
  assign n8613 = n8607 | n8612 ;
  assign n8614 = n8125 | n8613 ;
  assign n8615 = ( n2985 & n8613 ) | ( n2985 & n8614 ) | ( n8613 & n8614 ) ;
  assign n8616 = x5 & n8614 ;
  assign n8617 = x5 & n8613 ;
  assign n8618 = ( n2985 & n8616 ) | ( n2985 & n8617 ) | ( n8616 & n8617 ) ;
  assign n8619 = x5 & ~n8616 ;
  assign n8620 = x5 & ~n8617 ;
  assign n8621 = ( ~n2985 & n8619 ) | ( ~n2985 & n8620 ) | ( n8619 & n8620 ) ;
  assign n8622 = ( n8615 & ~n8618 ) | ( n8615 & n8621 ) | ( ~n8618 & n8621 ) ;
  assign n8604 = ~n7741 & n7744 ;
  assign n8623 = n8604 & n8622 ;
  assign n8624 = ( n8603 & n8622 ) | ( n8603 & n8623 ) | ( n8622 & n8623 ) ;
  assign n8605 = n8603 | n8604 ;
  assign n8625 = n8605 & ~n8624 ;
  assign n8626 = ~n8604 & n8622 ;
  assign n8627 = ~n8603 & n8626 ;
  assign n8628 = n8625 | n8627 ;
  assign n8629 = ~n7736 & n7739 ;
  assign n8630 = n7736 & ~n7739 ;
  assign n8631 = n8629 | n8630 ;
  assign n8632 = n2090 & n8118 ;
  assign n8633 = ( ~n2082 & n8118 ) | ( ~n2082 & n8632 ) | ( n8118 & n8632 ) ;
  assign n8634 = n2279 & n8115 ;
  assign n8635 = ( ~n2269 & n8115 ) | ( ~n2269 & n8634 ) | ( n8115 & n8634 ) ;
  assign n8636 = n2199 & n8122 ;
  assign n8637 = ( ~n2185 & n8122 ) | ( ~n2185 & n8636 ) | ( n8122 & n8636 ) ;
  assign n8638 = n8635 | n8637 ;
  assign n8639 = n8633 | n8638 ;
  assign n8640 = n8125 | n8639 ;
  assign n8641 = ( ~n2325 & n8639 ) | ( ~n2325 & n8640 ) | ( n8639 & n8640 ) ;
  assign n8642 = n8639 & n8640 ;
  assign n8643 = ( ~n2299 & n8641 ) | ( ~n2299 & n8642 ) | ( n8641 & n8642 ) ;
  assign n8644 = ~x5 & n8643 ;
  assign n8645 = x5 | n8643 ;
  assign n8646 = ( ~n8643 & n8644 ) | ( ~n8643 & n8645 ) | ( n8644 & n8645 ) ;
  assign n8647 = n8631 & n8646 ;
  assign n8648 = n8631 | n8646 ;
  assign n8649 = ~n8647 & n8648 ;
  assign n8650 = n7732 | n7734 ;
  assign n8651 = ~n7735 & n8650 ;
  assign n8652 = n1634 & n8115 ;
  assign n8653 = ( n1630 & n8115 ) | ( n1630 & n8652 ) | ( n8115 & n8652 ) ;
  assign n8654 = n2279 & n8118 ;
  assign n8655 = ( ~n2269 & n8118 ) | ( ~n2269 & n8654 ) | ( n8118 & n8654 ) ;
  assign n8656 = n8653 | n8655 ;
  assign n8657 = n2090 & n8122 ;
  assign n8658 = ( ~n2082 & n8122 ) | ( ~n2082 & n8657 ) | ( n8122 & n8657 ) ;
  assign n8659 = n8656 | n8658 ;
  assign n8660 = n8125 | n8659 ;
  assign n8661 = n8659 & n8660 ;
  assign n8662 = ( n2568 & n8660 ) | ( n2568 & n8661 ) | ( n8660 & n8661 ) ;
  assign n8663 = x5 & n8661 ;
  assign n8664 = x5 & n8660 ;
  assign n8665 = ( n2568 & n8663 ) | ( n2568 & n8664 ) | ( n8663 & n8664 ) ;
  assign n8666 = x5 & ~n8663 ;
  assign n8667 = x5 & ~n8664 ;
  assign n8668 = ( ~n2568 & n8666 ) | ( ~n2568 & n8667 ) | ( n8666 & n8667 ) ;
  assign n8669 = ( n8662 & ~n8665 ) | ( n8662 & n8668 ) | ( ~n8665 & n8668 ) ;
  assign n8670 = n8651 & n8669 ;
  assign n8671 = n7622 | n7730 ;
  assign n8672 = ~n7731 & n8671 ;
  assign n8673 = n1708 & n8115 ;
  assign n8674 = n1634 & n8118 ;
  assign n8675 = ( n1630 & n8118 ) | ( n1630 & n8674 ) | ( n8118 & n8674 ) ;
  assign n8676 = n2279 & n8122 ;
  assign n8677 = ( ~n2269 & n8122 ) | ( ~n2269 & n8676 ) | ( n8122 & n8676 ) ;
  assign n8678 = n8675 | n8677 ;
  assign n8679 = n8673 | n8678 ;
  assign n8680 = n8125 | n8679 ;
  assign n8681 = n8679 & n8680 ;
  assign n8682 = ( ~n2343 & n8680 ) | ( ~n2343 & n8681 ) | ( n8680 & n8681 ) ;
  assign n8683 = ~x5 & n8681 ;
  assign n8684 = ~x5 & n8680 ;
  assign n8685 = ( ~n2343 & n8683 ) | ( ~n2343 & n8684 ) | ( n8683 & n8684 ) ;
  assign n8686 = x5 | n8683 ;
  assign n8687 = x5 | n8684 ;
  assign n8688 = ( ~n2343 & n8686 ) | ( ~n2343 & n8687 ) | ( n8686 & n8687 ) ;
  assign n8689 = ( ~n8682 & n8685 ) | ( ~n8682 & n8688 ) | ( n8685 & n8688 ) ;
  assign n8690 = n8672 & n8689 ;
  assign n8691 = n7726 & n7728 ;
  assign n8692 = n7726 | n7728 ;
  assign n8693 = ~n8691 & n8692 ;
  assign n8694 = n1708 & n8118 ;
  assign n8695 = n1793 & n8115 ;
  assign n8696 = ( n1783 & n8115 ) | ( n1783 & n8695 ) | ( n8115 & n8695 ) ;
  assign n8697 = n1634 & n8122 ;
  assign n8698 = ( n1630 & n8122 ) | ( n1630 & n8697 ) | ( n8122 & n8697 ) ;
  assign n8699 = n8696 | n8698 ;
  assign n8700 = n8694 | n8699 ;
  assign n8701 = n8125 | n8700 ;
  assign n8702 = n8700 & n8701 ;
  assign n8703 = ( n1814 & n8701 ) | ( n1814 & n8702 ) | ( n8701 & n8702 ) ;
  assign n8704 = x5 & n8702 ;
  assign n8705 = x5 & n8701 ;
  assign n8706 = ( n1814 & n8704 ) | ( n1814 & n8705 ) | ( n8704 & n8705 ) ;
  assign n8707 = x5 & ~n8704 ;
  assign n8708 = x5 & ~n8705 ;
  assign n8709 = ( ~n1814 & n8707 ) | ( ~n1814 & n8708 ) | ( n8707 & n8708 ) ;
  assign n8710 = ( n8703 & ~n8706 ) | ( n8703 & n8709 ) | ( ~n8706 & n8709 ) ;
  assign n8711 = n8693 & n8710 ;
  assign n8712 = n7722 & n7724 ;
  assign n8713 = n7722 | n7724 ;
  assign n8714 = ~n8712 & n8713 ;
  assign n8715 = ~n523 & n8115 ;
  assign n8716 = n1793 & n8118 ;
  assign n8717 = ( n1783 & n8118 ) | ( n1783 & n8716 ) | ( n8118 & n8716 ) ;
  assign n8718 = n8715 | n8717 ;
  assign n8719 = n1708 & n8122 ;
  assign n8720 = n8718 | n8719 ;
  assign n8721 = n8125 | n8719 ;
  assign n8722 = n8718 | n8721 ;
  assign n8723 = ( ~n1852 & n8720 ) | ( ~n1852 & n8722 ) | ( n8720 & n8722 ) ;
  assign n8724 = ~x5 & n8722 ;
  assign n8725 = ~x5 & n8720 ;
  assign n8726 = ( ~n1852 & n8724 ) | ( ~n1852 & n8725 ) | ( n8724 & n8725 ) ;
  assign n8727 = x5 | n8725 ;
  assign n8728 = x5 | n8724 ;
  assign n8729 = ( ~n1852 & n8727 ) | ( ~n1852 & n8728 ) | ( n8727 & n8728 ) ;
  assign n8730 = ( ~n8723 & n8726 ) | ( ~n8723 & n8729 ) | ( n8726 & n8729 ) ;
  assign n8731 = n8714 & n8730 ;
  assign n8732 = n7718 | n7719 ;
  assign n8733 = n7702 | n8732 ;
  assign n8734 = ~n7721 & n8733 ;
  assign n8735 = ~n523 & n8118 ;
  assign n8736 = n352 & n8115 ;
  assign n8737 = ( ~n339 & n8115 ) | ( ~n339 & n8736 ) | ( n8115 & n8736 ) ;
  assign n8738 = n1793 & n8122 ;
  assign n8739 = ( n1783 & n8122 ) | ( n1783 & n8738 ) | ( n8122 & n8738 ) ;
  assign n8740 = n8737 | n8739 ;
  assign n8741 = n8735 | n8740 ;
  assign n8742 = n8125 | n8741 ;
  assign n8743 = n8741 & n8742 ;
  assign n8744 = ( n1884 & n8742 ) | ( n1884 & n8743 ) | ( n8742 & n8743 ) ;
  assign n8745 = x5 & n8743 ;
  assign n8746 = x5 & n8742 ;
  assign n8747 = ( n1884 & n8745 ) | ( n1884 & n8746 ) | ( n8745 & n8746 ) ;
  assign n8748 = x5 & ~n8745 ;
  assign n8749 = x5 & ~n8746 ;
  assign n8750 = ( ~n1884 & n8748 ) | ( ~n1884 & n8749 ) | ( n8748 & n8749 ) ;
  assign n8751 = ( n8744 & ~n8747 ) | ( n8744 & n8750 ) | ( ~n8747 & n8750 ) ;
  assign n8752 = n8734 & n8751 ;
  assign n8753 = n8734 | n8751 ;
  assign n8754 = ~n8752 & n8753 ;
  assign n8755 = ~n829 & n8115 ;
  assign n8756 = n352 & n8118 ;
  assign n8757 = ( ~n339 & n8118 ) | ( ~n339 & n8756 ) | ( n8118 & n8756 ) ;
  assign n8758 = n8755 | n8757 ;
  assign n8759 = ~n523 & n8122 ;
  assign n8760 = n8125 | n8759 ;
  assign n8761 = n8758 | n8760 ;
  assign n8762 = ~x5 & n8761 ;
  assign n8763 = n8758 | n8759 ;
  assign n8764 = ~x5 & n8763 ;
  assign n8765 = ( ~n1055 & n8762 ) | ( ~n1055 & n8764 ) | ( n8762 & n8764 ) ;
  assign n8766 = x5 & n8761 ;
  assign n8767 = x5 & ~n8766 ;
  assign n8768 = x5 & n8759 ;
  assign n8769 = ( x5 & n8758 ) | ( x5 & n8768 ) | ( n8758 & n8768 ) ;
  assign n8770 = x5 & ~n8769 ;
  assign n8771 = ( n1055 & n8767 ) | ( n1055 & n8770 ) | ( n8767 & n8770 ) ;
  assign n8772 = n8765 | n8771 ;
  assign n8773 = n7695 | n7697 ;
  assign n8774 = x8 & ~n7695 ;
  assign n8775 = ( n7678 & n8773 ) | ( n7678 & ~n8774 ) | ( n8773 & ~n8774 ) ;
  assign n8776 = ~n7700 & n8775 ;
  assign n8777 = n8772 & n8776 ;
  assign n8778 = x8 | n7692 ;
  assign n8779 = ( ~n7685 & n7692 ) | ( ~n7685 & n8778 ) | ( n7692 & n8778 ) ;
  assign n8780 = n7686 | n8779 ;
  assign n8781 = ~n7695 & n8780 ;
  assign n8782 = ~n829 & n8118 ;
  assign n8783 = n352 & n8122 ;
  assign n8784 = ( ~n339 & n8122 ) | ( ~n339 & n8783 ) | ( n8122 & n8783 ) ;
  assign n8785 = n8782 | n8784 ;
  assign n8786 = n692 & n8115 ;
  assign n8787 = ( n674 & n8115 ) | ( n674 & n8786 ) | ( n8115 & n8786 ) ;
  assign n8788 = n8785 | n8787 ;
  assign n8789 = n8125 | n8787 ;
  assign n8790 = n8785 | n8789 ;
  assign n8791 = ( ~n1209 & n8788 ) | ( ~n1209 & n8790 ) | ( n8788 & n8790 ) ;
  assign n8792 = ~x5 & n8790 ;
  assign n8793 = ~x5 & n8788 ;
  assign n8794 = ( ~n1209 & n8792 ) | ( ~n1209 & n8793 ) | ( n8792 & n8793 ) ;
  assign n8795 = x5 | n8793 ;
  assign n8796 = x5 | n8792 ;
  assign n8797 = ( ~n1209 & n8795 ) | ( ~n1209 & n8796 ) | ( n8795 & n8796 ) ;
  assign n8798 = ( ~n8791 & n8794 ) | ( ~n8791 & n8797 ) | ( n8794 & n8797 ) ;
  assign n8799 = n8781 & n8798 ;
  assign n8800 = ( ~n1027 & n7688 ) | ( ~n1027 & n7690 ) | ( n7688 & n7690 ) ;
  assign n8801 = ~n922 & n8118 ;
  assign n8802 = n1042 & n8115 ;
  assign n8803 = ( ~n1027 & n8115 ) | ( ~n1027 & n8802 ) | ( n8115 & n8802 ) ;
  assign n8804 = n8801 | n8803 ;
  assign n8805 = n692 & n8122 ;
  assign n8806 = ( n674 & n8122 ) | ( n674 & n8805 ) | ( n8122 & n8805 ) ;
  assign n8807 = n8804 | n8806 ;
  assign n8808 = ( n1538 & n8125 ) | ( n1538 & n8807 ) | ( n8125 & n8807 ) ;
  assign n8809 = ( x5 & ~n8807 ) | ( x5 & n8808 ) | ( ~n8807 & n8808 ) ;
  assign n8810 = ~n8808 & n8809 ;
  assign n8811 = ~n922 & n8122 ;
  assign n8812 = n1042 & n8118 ;
  assign n8813 = ( ~n1027 & n8118 ) | ( ~n1027 & n8812 ) | ( n8118 & n8812 ) ;
  assign n8814 = n8811 | n8813 ;
  assign n8815 = n8125 | n8813 ;
  assign n8816 = n8811 | n8815 ;
  assign n8817 = ( n1946 & n8814 ) | ( n1946 & n8816 ) | ( n8814 & n8816 ) ;
  assign n8818 = ~x5 & n8817 ;
  assign n8819 = n139 & n8113 ;
  assign n8820 = ( n1041 & n8113 ) | ( n1041 & n8819 ) | ( n8113 & n8819 ) ;
  assign n8821 = x5 & ~n8820 ;
  assign n8822 = n8113 | n8819 ;
  assign n8823 = x5 & ~n8822 ;
  assign n8824 = ( n1027 & n8821 ) | ( n1027 & n8823 ) | ( n8821 & n8823 ) ;
  assign n8825 = x5 & n8824 ;
  assign n8826 = ~n8817 & n8825 ;
  assign n8827 = ( n8818 & n8824 ) | ( n8818 & n8826 ) | ( n8824 & n8826 ) ;
  assign n8828 = x5 | n8807 ;
  assign n8829 = n8808 | n8828 ;
  assign n8830 = n8827 & n8829 ;
  assign n8831 = ~x5 & n8827 ;
  assign n8832 = ( n8810 & n8830 ) | ( n8810 & n8831 ) | ( n8830 & n8831 ) ;
  assign n8833 = n8800 & n8832 ;
  assign n8834 = n8832 & ~n8833 ;
  assign n8835 = ~n829 & n8122 ;
  assign n8836 = ~n922 & n8115 ;
  assign n8837 = n8835 | n8836 ;
  assign n8838 = n692 & n8118 ;
  assign n8839 = ( n674 & n8118 ) | ( n674 & n8838 ) | ( n8118 & n8838 ) ;
  assign n8840 = n8837 | n8839 ;
  assign n8841 = n8125 | n8839 ;
  assign n8842 = n8837 | n8841 ;
  assign n8843 = ( n1554 & n8840 ) | ( n1554 & n8842 ) | ( n8840 & n8842 ) ;
  assign n8844 = x5 & n8842 ;
  assign n8845 = x5 & n8840 ;
  assign n8846 = ( n1554 & n8844 ) | ( n1554 & n8845 ) | ( n8844 & n8845 ) ;
  assign n8847 = x5 & ~n8845 ;
  assign n8848 = x5 & ~n8844 ;
  assign n8849 = ( ~n1554 & n8847 ) | ( ~n1554 & n8848 ) | ( n8847 & n8848 ) ;
  assign n8850 = ( n8843 & ~n8846 ) | ( n8843 & n8849 ) | ( ~n8846 & n8849 ) ;
  assign n8851 = n8800 & ~n8832 ;
  assign n8852 = n8850 & n8851 ;
  assign n8853 = ( n8834 & n8850 ) | ( n8834 & n8852 ) | ( n8850 & n8852 ) ;
  assign n8854 = n8833 | n8853 ;
  assign n8855 = n8781 | n8798 ;
  assign n8856 = ~n8799 & n8855 ;
  assign n8857 = n8799 | n8856 ;
  assign n8858 = ( n8799 & n8854 ) | ( n8799 & n8857 ) | ( n8854 & n8857 ) ;
  assign n8859 = n8772 | n8776 ;
  assign n8860 = ~n8777 & n8859 ;
  assign n8861 = n8777 | n8860 ;
  assign n8862 = ( n8777 & n8858 ) | ( n8777 & n8861 ) | ( n8858 & n8861 ) ;
  assign n8863 = n8754 & n8862 ;
  assign n8864 = n8752 | n8863 ;
  assign n8865 = ~n8714 & n8730 ;
  assign n8866 = ( n8714 & ~n8731 ) | ( n8714 & n8865 ) | ( ~n8731 & n8865 ) ;
  assign n8867 = n8864 & n8866 ;
  assign n8868 = n8731 | n8867 ;
  assign n8869 = n8693 & ~n8711 ;
  assign n8870 = ~n8693 & n8710 ;
  assign n8871 = n8869 | n8870 ;
  assign n8872 = n8868 & n8871 ;
  assign n8873 = n8711 | n8872 ;
  assign n8874 = n8672 & ~n8690 ;
  assign n8875 = ~n8672 & n8689 ;
  assign n8876 = n8874 | n8875 ;
  assign n8877 = n8690 | n8876 ;
  assign n8878 = ( n8690 & n8873 ) | ( n8690 & n8877 ) | ( n8873 & n8877 ) ;
  assign n8879 = n8651 | n8669 ;
  assign n8880 = ~n8670 & n8879 ;
  assign n8881 = n8670 | n8880 ;
  assign n8882 = ( n8670 & n8878 ) | ( n8670 & n8881 ) | ( n8878 & n8881 ) ;
  assign n8883 = n8649 & n8882 ;
  assign n8884 = n8647 | n8883 ;
  assign n8885 = n8624 | n8884 ;
  assign n8886 = ( n8624 & n8628 ) | ( n8624 & n8885 ) | ( n8628 & n8885 ) ;
  assign n8887 = ~n8582 & n8600 ;
  assign n8888 = ( n8582 & ~n8601 ) | ( n8582 & n8887 ) | ( ~n8601 & n8887 ) ;
  assign n8889 = n8601 | n8888 ;
  assign n8890 = ( n8601 & n8886 ) | ( n8601 & n8889 ) | ( n8886 & n8889 ) ;
  assign n8891 = n8579 & n8890 ;
  assign n8892 = n8576 | n8891 ;
  assign n8893 = n7496 & n7752 ;
  assign n8894 = n7496 | n7752 ;
  assign n8895 = ~n8893 & n8894 ;
  assign n8896 = n2893 & n8118 ;
  assign n8897 = ( ~n2886 & n8118 ) | ( ~n2886 & n8896 ) | ( n8118 & n8896 ) ;
  assign n8898 = n2701 & n8115 ;
  assign n8899 = ( ~n2784 & n8115 ) | ( ~n2784 & n8898 ) | ( n8115 & n8898 ) ;
  assign n8900 = n3507 & n8122 ;
  assign n8901 = ( n3483 & n8122 ) | ( n3483 & n8900 ) | ( n8122 & n8900 ) ;
  assign n8902 = n8899 | n8901 ;
  assign n8903 = n8897 | n8902 ;
  assign n8904 = n8125 | n8903 ;
  assign n8905 = n8903 & n8904 ;
  assign n8906 = ( n3603 & n8904 ) | ( n3603 & n8905 ) | ( n8904 & n8905 ) ;
  assign n8907 = x5 & n8905 ;
  assign n8908 = x5 & n8904 ;
  assign n8909 = ( n3603 & n8907 ) | ( n3603 & n8908 ) | ( n8907 & n8908 ) ;
  assign n8910 = x5 & ~n8907 ;
  assign n8911 = x5 & ~n8908 ;
  assign n8912 = ( ~n3603 & n8910 ) | ( ~n3603 & n8911 ) | ( n8910 & n8911 ) ;
  assign n8913 = ( n8906 & ~n8909 ) | ( n8906 & n8912 ) | ( ~n8909 & n8912 ) ;
  assign n8914 = n8895 & n8913 ;
  assign n8915 = n8895 & ~n8914 ;
  assign n8916 = ~n8895 & n8913 ;
  assign n8917 = n8915 | n8916 ;
  assign n8918 = n8892 & n8917 ;
  assign n8919 = n8536 | n8554 ;
  assign n8920 = ~n8555 & n8919 ;
  assign n8921 = n8914 & n8920 ;
  assign n8922 = ( n8918 & n8920 ) | ( n8918 & n8921 ) | ( n8920 & n8921 ) ;
  assign n8923 = n8555 | n8922 ;
  assign n8924 = n8533 & n8923 ;
  assign n8925 = n8530 | n8924 ;
  assign n8926 = n8510 & n8925 ;
  assign n8927 = ~n8468 & n8484 ;
  assign n8928 = ( n8468 & ~n8485 ) | ( n8468 & n8927 ) | ( ~n8485 & n8927 ) ;
  assign n8929 = n8506 & n8928 ;
  assign n8930 = ( n8926 & n8928 ) | ( n8926 & n8929 ) | ( n8928 & n8929 ) ;
  assign n8931 = n8485 | n8930 ;
  assign n8932 = n8465 & n8931 ;
  assign n8933 = n8462 | n8932 ;
  assign n8934 = n8442 & n8933 ;
  assign n8935 = n8419 & n8439 ;
  assign n8936 = ( n8419 & n8934 ) | ( n8419 & n8935 ) | ( n8934 & n8935 ) ;
  assign n8937 = n8417 | n8936 ;
  assign n8938 = n8376 | n8394 ;
  assign n8939 = ~n8395 & n8938 ;
  assign n8940 = n8395 | n8939 ;
  assign n8941 = ( n8395 & n8937 ) | ( n8395 & n8940 ) | ( n8937 & n8940 ) ;
  assign n8942 = n8373 & n8941 ;
  assign n8943 = n8371 | n8942 ;
  assign n8944 = ~n8334 & n8350 ;
  assign n8945 = ( n8334 & ~n8351 ) | ( n8334 & n8944 ) | ( ~n8351 & n8944 ) ;
  assign n8946 = n8351 | n8945 ;
  assign n8947 = ( n8351 & n8943 ) | ( n8351 & n8946 ) | ( n8943 & n8946 ) ;
  assign n8948 = n8331 & n8947 ;
  assign n8949 = n8289 | n8306 ;
  assign n8950 = ~n8307 & n8949 ;
  assign n8951 = n8328 & n8950 ;
  assign n8952 = ( n8948 & n8950 ) | ( n8948 & n8951 ) | ( n8950 & n8951 ) ;
  assign n8953 = n8307 | n8952 ;
  assign n8954 = n8286 & n8953 ;
  assign n8955 = n8282 | n8954 ;
  assign n8956 = ~n8260 & n8955 ;
  assign n8957 = n8257 | n8956 ;
  assign n8958 = ~n8238 & n8957 ;
  assign n8959 = n8235 | n8958 ;
  assign n8960 = n8214 & n8959 ;
  assign n8961 = n8211 | n8960 ;
  assign n8962 = ~n8179 & n8961 ;
  assign n8963 = n8175 | n8962 ;
  assign n8964 = n8141 & n8963 ;
  assign n8965 = n8141 | n8963 ;
  assign n8966 = ~n8964 & n8965 ;
  assign n8971 = n343 | n356 ;
  assign n8972 = n555 | n8971 ;
  assign n8973 = n6826 | n8972 ;
  assign n8974 = n349 | n395 ;
  assign n8975 = n7982 | n8974 ;
  assign n8976 = n382 | n8975 ;
  assign n8977 = n8973 | n8976 ;
  assign n8978 = n143 & ~n497 ;
  assign n8979 = n311 | n1615 ;
  assign n8980 = n5154 | n8979 ;
  assign n8981 = n8978 & ~n8980 ;
  assign n8982 = ~n8977 & n8981 ;
  assign n8983 = n167 | n233 ;
  assign n8984 = n811 | n8983 ;
  assign n8985 = n6009 | n8984 ;
  assign n8986 = n682 | n3445 ;
  assign n8987 = n442 | n8986 ;
  assign n8988 = n8985 | n8987 ;
  assign n8989 = n182 | n354 ;
  assign n8990 = n1126 | n8989 ;
  assign n8991 = n117 | n1172 ;
  assign n8992 = n85 | n8991 ;
  assign n8993 = n8990 | n8992 ;
  assign n8994 = n487 | n8993 ;
  assign n8995 = n8988 | n8994 ;
  assign n8996 = n375 | n758 ;
  assign n8997 = n578 | n8996 ;
  assign n8998 = n1124 | n2047 ;
  assign n8999 = n8997 | n8998 ;
  assign n9000 = n110 | n8999 ;
  assign n9001 = n8995 | n9000 ;
  assign n9002 = n8982 & ~n9001 ;
  assign n9003 = n7992 | n7993 ;
  assign n9004 = n636 | n1286 ;
  assign n9005 = n764 | n5946 ;
  assign n9006 = n9004 | n9005 ;
  assign n9007 = n159 | n431 ;
  assign n9008 = n197 | n283 ;
  assign n9009 = n104 | n689 ;
  assign n9010 = n9008 | n9009 ;
  assign n9011 = n9007 | n9010 ;
  assign n9012 = n9006 | n9011 ;
  assign n9013 = n9003 | n9012 ;
  assign n9014 = n225 | n263 ;
  assign n9015 = n1648 | n1653 ;
  assign n9016 = n1645 | n9015 ;
  assign n9017 = n9014 | n9016 ;
  assign n9018 = n9013 | n9017 ;
  assign n9019 = n9002 & ~n9018 ;
  assign n8967 = x1 & ~x2 ;
  assign n8968 = ~x1 & x2 ;
  assign n8969 = n8967 | n8968 ;
  assign n9020 = x0 | x1 ;
  assign n9021 = n8969 & ~n9020 ;
  assign n9022 = n170 | n262 ;
  assign n9023 = n9021 & ~n9022 ;
  assign n9024 = ~x0 & x1 ;
  assign n9025 = n2768 | n3393 ;
  assign n9026 = n496 | n796 ;
  assign n9027 = n9025 | n9026 ;
  assign n9028 = n447 | n491 ;
  assign n9029 = n560 | n801 ;
  assign n9030 = n9028 | n9029 ;
  assign n9031 = n9027 | n9030 ;
  assign n9032 = n192 | n607 ;
  assign n9033 = n2024 | n9032 ;
  assign n9034 = n131 | n278 ;
  assign n9035 = n99 | n9034 ;
  assign n9036 = n9033 | n9035 ;
  assign n9037 = n514 | n600 ;
  assign n9038 = n1240 | n9037 ;
  assign n9039 = n9036 | n9038 ;
  assign n9040 = n9031 | n9039 ;
  assign n9041 = n1723 | n4246 ;
  assign n9042 = n433 | n3425 ;
  assign n9043 = n9041 | n9042 ;
  assign n9044 = n139 | n9043 ;
  assign n9045 = n141 | n302 ;
  assign n9046 = n255 | n9045 ;
  assign n9047 = n8012 | n9046 ;
  assign n9048 = n262 | n401 ;
  assign n9049 = n9047 | n9048 ;
  assign n9050 = n9044 | n9049 ;
  assign n9051 = n9040 | n9050 ;
  assign n9052 = ~n8982 & n9024 ;
  assign n9053 = ( n9024 & n9051 ) | ( n9024 & n9052 ) | ( n9051 & n9052 ) ;
  assign n9054 = ( n9021 & ~n9023 ) | ( n9021 & n9053 ) | ( ~n9023 & n9053 ) ;
  assign n9055 = n9021 | n9053 ;
  assign n9056 = ( ~n9019 & n9054 ) | ( ~n9019 & n9055 ) | ( n9054 & n9055 ) ;
  assign n8970 = x0 & n8969 ;
  assign n9057 = n8970 | n9056 ;
  assign n9058 = n9019 & ~n9022 ;
  assign n9059 = n8017 | n9058 ;
  assign n9060 = n8017 & n9058 ;
  assign n9061 = n9059 & ~n9060 ;
  assign n9062 = n8081 & ~n8089 ;
  assign n9063 = n8081 & ~n8088 ;
  assign n9064 = ( ~n7915 & n9062 ) | ( ~n7915 & n9063 ) | ( n9062 & n9063 ) ;
  assign n9065 = n9061 & ~n9064 ;
  assign n9066 = ( n8092 & n9062 ) | ( n8092 & n9063 ) | ( n9062 & n9063 ) ;
  assign n9067 = n9061 & ~n9066 ;
  assign n9068 = ( n7054 & n9065 ) | ( n7054 & n9067 ) | ( n9065 & n9067 ) ;
  assign n9069 = n9059 & ~n9068 ;
  assign n9070 = ( n7050 & n9065 ) | ( n7050 & n9067 ) | ( n9065 & n9067 ) ;
  assign n9071 = n9059 & ~n9070 ;
  assign n9072 = ( ~n5216 & n9069 ) | ( ~n5216 & n9071 ) | ( n9069 & n9071 ) ;
  assign n9073 = n9058 | n9072 ;
  assign n9074 = n8982 & ~n9051 ;
  assign n9075 = n9072 | n9074 ;
  assign n9076 = n9022 | n9074 ;
  assign n9077 = n9019 & ~n9076 ;
  assign n9078 = ( ~n9073 & n9075 ) | ( ~n9073 & n9077 ) | ( n9075 & n9077 ) ;
  assign n9079 = ( n9056 & n9057 ) | ( n9056 & n9078 ) | ( n9057 & n9078 ) ;
  assign n9080 = x2 & n9057 ;
  assign n9081 = x2 & n9056 ;
  assign n9082 = ( n9078 & n9080 ) | ( n9078 & n9081 ) | ( n9080 & n9081 ) ;
  assign n9083 = x2 & ~n9080 ;
  assign n9084 = x2 & ~n9081 ;
  assign n9085 = ( ~n9078 & n9083 ) | ( ~n9078 & n9084 ) | ( n9083 & n9084 ) ;
  assign n9086 = ( n9079 & ~n9082 ) | ( n9079 & n9085 ) | ( ~n9082 & n9085 ) ;
  assign n9087 = n8966 & n9086 ;
  assign n9404 = n7096 | n7829 ;
  assign n9405 = ( n7096 & n7099 ) | ( n7096 & n9404 ) | ( n7099 & n9404 ) ;
  assign n9088 = n5252 | n5853 ;
  assign n9248 = n4110 | n4113 ;
  assign n9249 = ( n3971 & n4110 ) | ( n3971 & n9248 ) | ( n4110 & n9248 ) ;
  assign n9089 = n1057 & n1708 ;
  assign n9090 = ~n523 & n1060 ;
  assign n9091 = n1065 & n1793 ;
  assign n9092 = ( n1065 & n1783 ) | ( n1065 & n9091 ) | ( n1783 & n9091 ) ;
  assign n9093 = n1062 | n9092 ;
  assign n9094 = n9090 | n9093 ;
  assign n9095 = n9089 | n9094 ;
  assign n9096 = n9090 | n9092 ;
  assign n9097 = n9089 | n9096 ;
  assign n9098 = ( ~n1852 & n9095 ) | ( ~n1852 & n9097 ) | ( n9095 & n9097 ) ;
  assign n9099 = n1693 | n5123 ;
  assign n9100 = n141 | n560 ;
  assign n9101 = n1166 | n9100 ;
  assign n9102 = n9099 | n9101 ;
  assign n9103 = n930 | n2023 ;
  assign n9104 = n3983 | n9103 ;
  assign n9105 = n9102 | n9104 ;
  assign n9106 = n399 | n479 ;
  assign n9107 = n213 | n9106 ;
  assign n9108 = n9105 | n9107 ;
  assign n9109 = n124 | n460 ;
  assign n9110 = n514 | n758 ;
  assign n9111 = n9109 | n9110 ;
  assign n9112 = n228 | n270 ;
  assign n9113 = n887 | n9112 ;
  assign n9114 = n5069 | n7011 ;
  assign n9115 = n9113 | n9114 ;
  assign n9116 = n9111 | n9115 ;
  assign n9117 = n155 | n240 ;
  assign n9118 = n178 | n638 ;
  assign n9119 = n193 | n542 ;
  assign n9120 = n9118 | n9119 ;
  assign n9121 = n332 | n929 ;
  assign n9122 = n9120 | n9121 ;
  assign n9123 = n9117 | n9122 ;
  assign n9124 = n9116 | n9123 ;
  assign n9125 = n9108 | n9124 ;
  assign n9126 = n176 | n644 ;
  assign n9127 = n274 | n9126 ;
  assign n9128 = n71 | n303 ;
  assign n9129 = n39 | n9128 ;
  assign n9130 = n9127 | n9129 ;
  assign n9131 = n234 | n1714 ;
  assign n9132 = n9130 | n9131 ;
  assign n9133 = n103 | n5092 ;
  assign n9134 = n1765 | n9133 ;
  assign n9135 = n9132 | n9134 ;
  assign n9136 = n414 | n764 ;
  assign n9137 = n1126 | n1304 ;
  assign n9138 = n9136 | n9137 ;
  assign n9139 = n648 | n9138 ;
  assign n9140 = n441 | n480 ;
  assign n9141 = n189 | n461 ;
  assign n9142 = n9140 | n9141 ;
  assign n9143 = n92 | n643 ;
  assign n9144 = n401 | n9143 ;
  assign n9145 = n9142 | n9144 ;
  assign n9146 = n9139 | n9145 ;
  assign n9147 = n9135 | n9146 ;
  assign n9148 = n9125 | n9147 ;
  assign n9149 = n2774 | n2777 ;
  assign n9150 = n489 | n735 ;
  assign n9151 = n527 | n806 ;
  assign n9152 = n531 | n9151 ;
  assign n9153 = n9150 | n9152 ;
  assign n9154 = n79 | n938 ;
  assign n9155 = n369 | n432 ;
  assign n9156 = n9154 | n9155 ;
  assign n9157 = n374 | n1114 ;
  assign n9158 = n9156 | n9157 ;
  assign n9159 = n9153 | n9158 ;
  assign n9160 = n4142 | n9159 ;
  assign n9161 = n9149 | n9160 ;
  assign n9162 = n59 | n247 ;
  assign n9163 = n349 | n9162 ;
  assign n9164 = n1355 | n2147 ;
  assign n9165 = n1251 | n6029 ;
  assign n9166 = n9164 | n9165 ;
  assign n9167 = n317 | n591 ;
  assign n9168 = n9166 | n9167 ;
  assign n9169 = n9163 | n9168 ;
  assign n9170 = n9161 | n9169 ;
  assign n9171 = n9148 | n9170 ;
  assign n9172 = n1615 | n2053 ;
  assign n9173 = n3375 | n9172 ;
  assign n9174 = n64 | n289 ;
  assign n9175 = n223 | n9174 ;
  assign n9176 = n372 | n9175 ;
  assign n9177 = n9173 | n9176 ;
  assign n9178 = n424 | n9177 ;
  assign n9179 = n9171 | n9178 ;
  assign n9180 = n9089 & n9179 ;
  assign n9181 = ( n9094 & n9179 ) | ( n9094 & n9180 ) | ( n9179 & n9180 ) ;
  assign n9182 = ( n9096 & n9179 ) | ( n9096 & n9180 ) | ( n9179 & n9180 ) ;
  assign n9183 = ( ~n1852 & n9181 ) | ( ~n1852 & n9182 ) | ( n9181 & n9182 ) ;
  assign n9184 = n9098 & ~n9183 ;
  assign n9185 = ~n9097 & n9179 ;
  assign n9186 = ~n9095 & n9179 ;
  assign n9187 = ( n1852 & n9185 ) | ( n1852 & n9186 ) | ( n9185 & n9186 ) ;
  assign n9188 = n9184 | n9187 ;
  assign n9189 = n4057 & n9188 ;
  assign n9190 = ( n4064 & n9188 ) | ( n4064 & n9189 ) | ( n9188 & n9189 ) ;
  assign n9191 = n4057 | n9188 ;
  assign n9192 = n4064 | n9191 ;
  assign n9193 = ~n9190 & n9192 ;
  assign n9194 = n1634 & n1826 ;
  assign n9195 = ( n1630 & n1826 ) | ( n1630 & n9194 ) | ( n1826 & n9194 ) ;
  assign n9196 = n1823 & n2279 ;
  assign n9197 = ( n1823 & ~n2269 ) | ( n1823 & n9196 ) | ( ~n2269 & n9196 ) ;
  assign n9198 = n9195 | n9197 ;
  assign n9199 = n1829 & n2090 ;
  assign n9200 = ( n1829 & ~n2082 ) | ( n1829 & n9199 ) | ( ~n2082 & n9199 ) ;
  assign n9201 = n9198 | n9200 ;
  assign n9202 = n1821 | n9201 ;
  assign n9203 = n9201 & n9202 ;
  assign n9204 = ( n2568 & n9202 ) | ( n2568 & n9203 ) | ( n9202 & n9203 ) ;
  assign n9205 = x29 & n9203 ;
  assign n9206 = x29 & n9202 ;
  assign n9207 = ( n2568 & n9205 ) | ( n2568 & n9206 ) | ( n9205 & n9206 ) ;
  assign n9208 = x29 & ~n9205 ;
  assign n9209 = x29 & ~n9206 ;
  assign n9210 = ( ~n2568 & n9208 ) | ( ~n2568 & n9209 ) | ( n9208 & n9209 ) ;
  assign n9211 = ( n9204 & ~n9207 ) | ( n9204 & n9210 ) | ( ~n9207 & n9210 ) ;
  assign n9212 = n9193 & n9211 ;
  assign n9213 = n9193 | n9211 ;
  assign n9214 = ~n9212 & n9213 ;
  assign n9215 = n4085 | n4087 ;
  assign n9216 = ( n1843 & n4085 ) | ( n1843 & n9215 ) | ( n4085 & n9215 ) ;
  assign n9217 = n4085 | n9215 ;
  assign n9218 = ( n2020 & n9216 ) | ( n2020 & n9217 ) | ( n9216 & n9217 ) ;
  assign n9219 = n9214 | n9218 ;
  assign n9220 = ( n4085 & n4088 ) | ( n4085 & n9214 ) | ( n4088 & n9214 ) ;
  assign n9221 = ( n4085 & n4087 ) | ( n4085 & n9214 ) | ( n4087 & n9214 ) ;
  assign n9222 = ( n2020 & n9220 ) | ( n2020 & n9221 ) | ( n9220 & n9221 ) ;
  assign n9223 = n9219 & ~n9222 ;
  assign n9224 = n2315 & n2701 ;
  assign n9225 = ( n2315 & ~n2784 ) | ( n2315 & n9224 ) | ( ~n2784 & n9224 ) ;
  assign n9226 = n2308 & n2691 ;
  assign n9227 = ( n2308 & n2678 ) | ( n2308 & n9226 ) | ( n2678 & n9226 ) ;
  assign n9228 = n9225 | n9227 ;
  assign n9229 = n2199 & n2312 ;
  assign n9230 = ( ~n2185 & n2312 ) | ( ~n2185 & n9229 ) | ( n2312 & n9229 ) ;
  assign n9231 = n9228 | n9230 ;
  assign n9232 = n2306 | n9230 ;
  assign n9233 = n9228 | n9232 ;
  assign n9234 = ( n2960 & n9231 ) | ( n2960 & n9233 ) | ( n9231 & n9233 ) ;
  assign n9235 = x26 & n9233 ;
  assign n9236 = x26 & n9231 ;
  assign n9237 = ( n2960 & n9235 ) | ( n2960 & n9236 ) | ( n9235 & n9236 ) ;
  assign n9238 = x26 & ~n9236 ;
  assign n9239 = x26 & ~n9235 ;
  assign n9240 = ( ~n2960 & n9238 ) | ( ~n2960 & n9239 ) | ( n9238 & n9239 ) ;
  assign n9241 = ( n9234 & ~n9237 ) | ( n9234 & n9240 ) | ( ~n9237 & n9240 ) ;
  assign n9242 = ~n9222 & n9241 ;
  assign n9243 = n9219 & n9242 ;
  assign n9244 = n9223 & ~n9243 ;
  assign n9245 = n9222 & n9241 ;
  assign n9246 = ( ~n9219 & n9241 ) | ( ~n9219 & n9245 ) | ( n9241 & n9245 ) ;
  assign n9247 = n9244 | n9246 ;
  assign n9250 = n9247 & n9249 ;
  assign n9251 = n9249 & ~n9250 ;
  assign n9252 = n2893 & n2925 ;
  assign n9253 = ( ~n2886 & n2925 ) | ( ~n2886 & n9252 ) | ( n2925 & n9252 ) ;
  assign n9254 = n2928 & n3507 ;
  assign n9255 = ( n2928 & n3483 ) | ( n2928 & n9254 ) | ( n3483 & n9254 ) ;
  assign n9256 = n9253 | n9255 ;
  assign n9257 = n2932 & n3386 ;
  assign n9258 = n9256 | n9257 ;
  assign n9259 = n2936 | n9257 ;
  assign n9260 = n9256 | n9259 ;
  assign n9261 = ( ~n3568 & n9258 ) | ( ~n3568 & n9260 ) | ( n9258 & n9260 ) ;
  assign n9262 = ~x23 & n9260 ;
  assign n9263 = ~x23 & n9258 ;
  assign n9264 = ( ~n3568 & n9262 ) | ( ~n3568 & n9263 ) | ( n9262 & n9263 ) ;
  assign n9265 = x23 | n9263 ;
  assign n9266 = x23 | n9262 ;
  assign n9267 = ( ~n3568 & n9265 ) | ( ~n3568 & n9266 ) | ( n9265 & n9266 ) ;
  assign n9268 = ( ~n9261 & n9264 ) | ( ~n9261 & n9267 ) | ( n9264 & n9267 ) ;
  assign n9269 = n9247 & ~n9249 ;
  assign n9270 = n9268 & n9269 ;
  assign n9271 = ( n9251 & n9268 ) | ( n9251 & n9270 ) | ( n9268 & n9270 ) ;
  assign n9272 = n9268 | n9269 ;
  assign n9273 = n9251 | n9272 ;
  assign n9274 = ~n9271 & n9273 ;
  assign n9275 = n4134 | n4136 ;
  assign n9276 = ( n4134 & n4138 ) | ( n4134 & n9275 ) | ( n4138 & n9275 ) ;
  assign n9277 = n9274 & n9276 ;
  assign n9278 = n9274 | n9276 ;
  assign n9279 = ~n9277 & n9278 ;
  assign n9280 = n3541 & n4206 ;
  assign n9281 = n3547 & ~n4429 ;
  assign n9282 = n3439 & n3544 ;
  assign n9283 = ( ~n3420 & n3544 ) | ( ~n3420 & n9282 ) | ( n3544 & n9282 ) ;
  assign n9284 = n9281 | n9283 ;
  assign n9285 = n9280 | n9284 ;
  assign n9286 = n3537 | n9280 ;
  assign n9287 = n9284 | n9286 ;
  assign n9288 = ( ~n4527 & n9285 ) | ( ~n4527 & n9287 ) | ( n9285 & n9287 ) ;
  assign n9289 = ~x20 & n9287 ;
  assign n9290 = ~x20 & n9285 ;
  assign n9291 = ( ~n4527 & n9289 ) | ( ~n4527 & n9290 ) | ( n9289 & n9290 ) ;
  assign n9292 = x20 | n9290 ;
  assign n9293 = x20 | n9289 ;
  assign n9294 = ( ~n4527 & n9292 ) | ( ~n4527 & n9293 ) | ( n9292 & n9293 ) ;
  assign n9295 = ( ~n9288 & n9291 ) | ( ~n9288 & n9294 ) | ( n9291 & n9294 ) ;
  assign n9296 = n9279 & n9295 ;
  assign n9297 = n9279 & ~n9296 ;
  assign n9298 = ~n9279 & n9295 ;
  assign n9299 = n9297 | n9298 ;
  assign n9300 = n4237 | n4240 ;
  assign n9301 = ( n3970 & n4237 ) | ( n3970 & n9300 ) | ( n4237 & n9300 ) ;
  assign n9302 = n9299 & ~n9301 ;
  assign n9303 = ~n9299 & n9301 ;
  assign n9304 = n9302 | n9303 ;
  assign n9305 = n4396 & n4466 ;
  assign n9306 = n4245 & n4468 ;
  assign n9307 = ( n4303 & n4468 ) | ( n4303 & n9306 ) | ( n4468 & n9306 ) ;
  assign n9308 = n9305 | n9307 ;
  assign n9309 = n4471 & n5192 ;
  assign n9310 = ( n4471 & n5179 ) | ( n4471 & n9309 ) | ( n5179 & n9309 ) ;
  assign n9311 = n9308 | n9310 ;
  assign n9312 = n4475 | n9310 ;
  assign n9313 = n9308 | n9312 ;
  assign n9314 = ( n5306 & n9311 ) | ( n5306 & n9313 ) | ( n9311 & n9313 ) ;
  assign n9315 = x17 & n9313 ;
  assign n9316 = x17 & n9311 ;
  assign n9317 = ( n5306 & n9315 ) | ( n5306 & n9316 ) | ( n9315 & n9316 ) ;
  assign n9318 = x17 & ~n9316 ;
  assign n9319 = x17 & ~n9315 ;
  assign n9320 = ( ~n5306 & n9318 ) | ( ~n5306 & n9319 ) | ( n9318 & n9319 ) ;
  assign n9321 = ( n9314 & ~n9317 ) | ( n9314 & n9320 ) | ( ~n9317 & n9320 ) ;
  assign n9322 = n9304 & n9321 ;
  assign n9323 = n9304 | n9321 ;
  assign n9324 = ~n9322 & n9323 ;
  assign n9325 = n4487 | n4999 ;
  assign n9326 = ( n4487 & n4491 ) | ( n4487 & n9325 ) | ( n4491 & n9325 ) ;
  assign n9327 = n9324 & n9326 ;
  assign n9328 = n9324 | n9326 ;
  assign n9329 = ~n9327 & n9328 ;
  assign n9330 = n5117 & n5237 ;
  assign n9331 = ( ~n5037 & n5237 ) | ( ~n5037 & n9330 ) | ( n5237 & n9330 ) ;
  assign n9332 = n5108 & n5231 ;
  assign n9333 = n5234 & n5997 ;
  assign n9334 = ( n5234 & n5979 ) | ( n5234 & n9333 ) | ( n5979 & n9333 ) ;
  assign n9335 = n9332 | n9334 ;
  assign n9336 = n9331 | n9335 ;
  assign n9337 = n5227 | n9336 ;
  assign n9338 = n9336 & n9337 ;
  assign n9339 = ( n6181 & n9337 ) | ( n6181 & n9338 ) | ( n9337 & n9338 ) ;
  assign n9340 = x14 & n9338 ;
  assign n9341 = x14 & n9337 ;
  assign n9342 = ( n6181 & n9340 ) | ( n6181 & n9341 ) | ( n9340 & n9341 ) ;
  assign n9343 = x14 & ~n9340 ;
  assign n9344 = x14 & ~n9341 ;
  assign n9345 = ( ~n6181 & n9343 ) | ( ~n6181 & n9344 ) | ( n9343 & n9344 ) ;
  assign n9346 = ( n9339 & ~n9342 ) | ( n9339 & n9345 ) | ( ~n9342 & n9345 ) ;
  assign n9347 = n9329 & n9346 ;
  assign n9348 = n9329 & ~n9347 ;
  assign n9349 = ~n9329 & n9346 ;
  assign n9350 = n9348 | n9349 ;
  assign n9351 = n9088 & n9350 ;
  assign n9352 = n9088 & ~n9351 ;
  assign n9353 = ~n9088 & n9350 ;
  assign n9354 = n9352 | n9353 ;
  assign n9355 = n5857 & n6125 ;
  assign n9356 = ( ~n5899 & n6125 ) | ( ~n5899 & n9355 ) | ( n6125 & n9355 ) ;
  assign n9357 = ~n6091 & n6119 ;
  assign n9358 = n6122 & n7036 ;
  assign n9359 = ( n6122 & n7023 ) | ( n6122 & n9358 ) | ( n7023 & n9358 ) ;
  assign n9360 = n9357 | n9359 ;
  assign n9361 = n9356 | n9360 ;
  assign n9362 = n6115 | n9361 ;
  assign n9363 = ( n7136 & n9361 ) | ( n7136 & n9362 ) | ( n9361 & n9362 ) ;
  assign n9364 = x11 & n9362 ;
  assign n9365 = x11 & n9361 ;
  assign n9366 = ( n7136 & n9364 ) | ( n7136 & n9365 ) | ( n9364 & n9365 ) ;
  assign n9367 = x11 & ~n9364 ;
  assign n9368 = x11 & ~n9365 ;
  assign n9369 = ( ~n7136 & n9367 ) | ( ~n7136 & n9368 ) | ( n9367 & n9368 ) ;
  assign n9370 = ( n9363 & ~n9366 ) | ( n9363 & n9369 ) | ( ~n9366 & n9369 ) ;
  assign n9371 = n9353 & n9370 ;
  assign n9372 = ( n9352 & n9370 ) | ( n9352 & n9371 ) | ( n9370 & n9371 ) ;
  assign n9373 = n9354 & ~n9372 ;
  assign n9374 = ~n9353 & n9370 ;
  assign n9375 = ~n9352 & n9374 ;
  assign n9376 = n9373 | n9375 ;
  assign n9377 = n6139 | n6795 ;
  assign n9378 = ( n6139 & n6142 ) | ( n6139 & n9377 ) | ( n6142 & n9377 ) ;
  assign n9379 = n9376 & n9378 ;
  assign n9380 = n9376 | n9378 ;
  assign n9381 = ~n9379 & n9380 ;
  assign n9382 = n6950 & n7074 ;
  assign n9383 = n6889 & n7068 ;
  assign n9384 = ( ~n6884 & n7068 ) | ( ~n6884 & n9383 ) | ( n7068 & n9383 ) ;
  assign n9385 = n9382 | n9384 ;
  assign n9386 = n7079 & n7907 ;
  assign n9387 = ( n7079 & n7902 ) | ( n7079 & n9386 ) | ( n7902 & n9386 ) ;
  assign n9389 = n7078 | n9387 ;
  assign n9390 = n9385 | n9389 ;
  assign n9388 = n9385 | n9387 ;
  assign n9391 = n9388 & n9390 ;
  assign n9392 = ( ~n8193 & n9390 ) | ( ~n8193 & n9391 ) | ( n9390 & n9391 ) ;
  assign n9393 = ~x8 & n9391 ;
  assign n9394 = ~x8 & n9390 ;
  assign n9395 = ( ~n8193 & n9393 ) | ( ~n8193 & n9394 ) | ( n9393 & n9394 ) ;
  assign n9396 = x8 | n9393 ;
  assign n9397 = x8 | n9394 ;
  assign n9398 = ( ~n8193 & n9396 ) | ( ~n8193 & n9397 ) | ( n9396 & n9397 ) ;
  assign n9399 = ( ~n9392 & n9395 ) | ( ~n9392 & n9398 ) | ( n9395 & n9398 ) ;
  assign n9400 = n9381 & n9399 ;
  assign n9401 = n9381 & ~n9400 ;
  assign n9402 = ~n9381 & n9399 ;
  assign n9403 = n9401 | n9402 ;
  assign n9406 = n9403 & n9405 ;
  assign n9407 = n9405 & ~n9406 ;
  assign n9408 = n9403 & ~n9406 ;
  assign n9409 = n9407 | n9408 ;
  assign n9410 = ( n5216 & n9068 ) | ( n5216 & n9070 ) | ( n9068 & n9070 ) ;
  assign n9411 = ( ~n7054 & n9064 ) | ( ~n7054 & n9066 ) | ( n9064 & n9066 ) ;
  assign n9412 = ~n9061 & n9411 ;
  assign n9413 = ( ~n7050 & n9064 ) | ( ~n7050 & n9066 ) | ( n9064 & n9066 ) ;
  assign n9414 = ~n9061 & n9413 ;
  assign n9415 = ( ~n5216 & n9412 ) | ( ~n5216 & n9414 ) | ( n9412 & n9414 ) ;
  assign n9416 = n9410 | n9415 ;
  assign n9417 = n8079 & n8115 ;
  assign n9418 = ( ~n8070 & n8115 ) | ( ~n8070 & n9417 ) | ( n8115 & n9417 ) ;
  assign n9419 = n8118 | n9418 ;
  assign n9420 = ( ~n8017 & n9418 ) | ( ~n8017 & n9419 ) | ( n9418 & n9419 ) ;
  assign n9421 = n8122 & n9022 ;
  assign n9422 = ( n8122 & ~n9019 ) | ( n8122 & n9421 ) | ( ~n9019 & n9421 ) ;
  assign n9423 = n9420 | n9422 ;
  assign n9424 = n8125 | n9422 ;
  assign n9425 = n9420 | n9424 ;
  assign n9426 = ( ~n9416 & n9423 ) | ( ~n9416 & n9425 ) | ( n9423 & n9425 ) ;
  assign n9427 = ~x5 & n9425 ;
  assign n9428 = ~x5 & n9423 ;
  assign n9429 = ( ~n9416 & n9427 ) | ( ~n9416 & n9428 ) | ( n9427 & n9428 ) ;
  assign n9430 = x5 | n9428 ;
  assign n9431 = x5 | n9427 ;
  assign n9432 = ( ~n9416 & n9430 ) | ( ~n9416 & n9431 ) | ( n9430 & n9431 ) ;
  assign n9433 = ( ~n9426 & n9429 ) | ( ~n9426 & n9432 ) | ( n9429 & n9432 ) ;
  assign n9434 = ~n8982 & n9022 ;
  assign n9435 = ( n9022 & n9051 ) | ( n9022 & n9434 ) | ( n9051 & n9434 ) ;
  assign n9436 = ( n9019 & n9074 ) | ( n9019 & ~n9435 ) | ( n9074 & ~n9435 ) ;
  assign n9437 = n8982 & ~n9022 ;
  assign n9438 = ~n9051 & n9437 ;
  assign n9439 = n9019 & n9438 ;
  assign n9440 = n9436 & ~n9439 ;
  assign n9441 = n9022 & ~n9074 ;
  assign n9442 = ( n9019 & n9074 ) | ( n9019 & ~n9441 ) | ( n9074 & ~n9441 ) ;
  assign n9443 = ( n9074 & ~n9440 ) | ( n9074 & n9442 ) | ( ~n9440 & n9442 ) ;
  assign n9444 = ~n8982 & n9021 ;
  assign n9445 = ( n9021 & n9051 ) | ( n9021 & n9444 ) | ( n9051 & n9444 ) ;
  assign n9446 = n8970 | n9445 ;
  assign n9447 = ( ~n9443 & n9445 ) | ( ~n9443 & n9446 ) | ( n9445 & n9446 ) ;
  assign n9448 = ( ~n9442 & n9445 ) | ( ~n9442 & n9446 ) | ( n9445 & n9446 ) ;
  assign n9449 = ( ~n9072 & n9447 ) | ( ~n9072 & n9448 ) | ( n9447 & n9448 ) ;
  assign n9450 = ~x2 & n9447 ;
  assign n9451 = ~x2 & n9448 ;
  assign n9452 = ( ~n9072 & n9450 ) | ( ~n9072 & n9451 ) | ( n9450 & n9451 ) ;
  assign n9453 = x2 | n9450 ;
  assign n9454 = x2 | n9451 ;
  assign n9455 = ( ~n9072 & n9453 ) | ( ~n9072 & n9454 ) | ( n9453 & n9454 ) ;
  assign n9456 = ( ~n9449 & n9452 ) | ( ~n9449 & n9455 ) | ( n9452 & n9455 ) ;
  assign n9457 = n9433 & n9456 ;
  assign n9458 = n9433 & ~n9457 ;
  assign n9459 = ~n9433 & n9456 ;
  assign n9460 = n9458 | n9459 ;
  assign n9461 = ~n9409 & n9460 ;
  assign n9462 = n9409 & ~n9460 ;
  assign n9463 = n9461 | n9462 ;
  assign n9464 = n8137 | n8964 ;
  assign n9465 = n9463 & n9464 ;
  assign n9466 = n9463 | n9464 ;
  assign n9467 = ~n9465 & n9466 ;
  assign n9468 = n9087 | n9467 ;
  assign n9469 = n8260 & ~n8955 ;
  assign n9470 = n8956 | n9469 ;
  assign n9471 = n6889 & n9021 ;
  assign n9472 = ( ~n6884 & n9021 ) | ( ~n6884 & n9471 ) | ( n9021 & n9471 ) ;
  assign n9473 = n7907 & n9024 ;
  assign n9474 = ( n7902 & n9024 ) | ( n7902 & n9473 ) | ( n9024 & n9473 ) ;
  assign n9475 = x0 & ~n8969 ;
  assign n9476 = n8079 & n9475 ;
  assign n9477 = ( ~n8070 & n9475 ) | ( ~n8070 & n9476 ) | ( n9475 & n9476 ) ;
  assign n9478 = n9474 | n9477 ;
  assign n9479 = n9472 | n9478 ;
  assign n9480 = n8970 | n9479 ;
  assign n9481 = n9479 & n9480 ;
  assign n9482 = ( ~n8156 & n9480 ) | ( ~n8156 & n9481 ) | ( n9480 & n9481 ) ;
  assign n9483 = ~x2 & n9481 ;
  assign n9484 = ~x2 & n9480 ;
  assign n9485 = ( ~n8156 & n9483 ) | ( ~n8156 & n9484 ) | ( n9483 & n9484 ) ;
  assign n9486 = x2 | n9483 ;
  assign n9487 = x2 | n9484 ;
  assign n9488 = ( ~n8156 & n9486 ) | ( ~n8156 & n9487 ) | ( n9486 & n9487 ) ;
  assign n9489 = ( ~n9482 & n9485 ) | ( ~n9482 & n9488 ) | ( n9485 & n9488 ) ;
  assign n9490 = ~n9470 & n9489 ;
  assign n9491 = n9470 | n9490 ;
  assign n9492 = n9470 & n9489 ;
  assign n9493 = n9491 & ~n9492 ;
  assign n9494 = n8286 & ~n8953 ;
  assign n9495 = n8943 & n8945 ;
  assign n9496 = n8943 | n8945 ;
  assign n9497 = ~n9495 & n9496 ;
  assign n9498 = n5857 & n9024 ;
  assign n9499 = ( ~n5899 & n9024 ) | ( ~n5899 & n9498 ) | ( n9024 & n9498 ) ;
  assign n9500 = ~n6091 & n9475 ;
  assign n9501 = n5997 & n9021 ;
  assign n9502 = ( n5979 & n9021 ) | ( n5979 & n9501 ) | ( n9021 & n9501 ) ;
  assign n9503 = n9500 | n9502 ;
  assign n9504 = n9499 | n9503 ;
  assign n9505 = n8970 | n9504 ;
  assign n9506 = n9504 & n9505 ;
  assign n9507 = ( n6108 & n9505 ) | ( n6108 & n9506 ) | ( n9505 & n9506 ) ;
  assign n9508 = x2 & n9506 ;
  assign n9509 = x2 & n9505 ;
  assign n9510 = ( n6108 & n9508 ) | ( n6108 & n9509 ) | ( n9508 & n9509 ) ;
  assign n9511 = x2 & ~n9508 ;
  assign n9512 = x2 & ~n9509 ;
  assign n9513 = ( ~n6108 & n9511 ) | ( ~n6108 & n9512 ) | ( n9511 & n9512 ) ;
  assign n9514 = ( n9507 & ~n9510 ) | ( n9507 & n9513 ) | ( ~n9510 & n9513 ) ;
  assign n9515 = n4396 & n9021 ;
  assign n9516 = n4245 & n9024 ;
  assign n9517 = ( n4303 & n9024 ) | ( n4303 & n9516 ) | ( n9024 & n9516 ) ;
  assign n9518 = n9515 | n9517 ;
  assign n9519 = n5192 & n9475 ;
  assign n9520 = ( n5179 & n9475 ) | ( n5179 & n9519 ) | ( n9475 & n9519 ) ;
  assign n9522 = n8970 | n9520 ;
  assign n9523 = n9518 | n9522 ;
  assign n9521 = n9518 | n9520 ;
  assign n9524 = n9521 & n9523 ;
  assign n9525 = ( n5306 & n9523 ) | ( n5306 & n9524 ) | ( n9523 & n9524 ) ;
  assign n9526 = x2 & n9524 ;
  assign n9527 = x2 & n9523 ;
  assign n9528 = ( n5306 & n9526 ) | ( n5306 & n9527 ) | ( n9526 & n9527 ) ;
  assign n9529 = x2 & ~n9526 ;
  assign n9530 = x2 & ~n9527 ;
  assign n9531 = ( ~n5306 & n9529 ) | ( ~n5306 & n9530 ) | ( n9529 & n9530 ) ;
  assign n9532 = ( n9525 & ~n9528 ) | ( n9525 & n9531 ) | ( ~n9528 & n9531 ) ;
  assign n9533 = ~n4429 & n9021 ;
  assign n9534 = n4396 & n9024 ;
  assign n9535 = n9533 | n9534 ;
  assign n9536 = n4245 & n9475 ;
  assign n9537 = ( n4303 & n9475 ) | ( n4303 & n9536 ) | ( n9475 & n9536 ) ;
  assign n9539 = n8970 | n9537 ;
  assign n9540 = n9535 | n9539 ;
  assign n9538 = n9535 | n9537 ;
  assign n9541 = n9538 & n9540 ;
  assign n9542 = ( n4455 & n9540 ) | ( n4455 & n9541 ) | ( n9540 & n9541 ) ;
  assign n9543 = x2 & n9541 ;
  assign n9544 = x2 & n9540 ;
  assign n9545 = ( n4455 & n9543 ) | ( n4455 & n9544 ) | ( n9543 & n9544 ) ;
  assign n9546 = x2 & ~n9543 ;
  assign n9547 = x2 & ~n9544 ;
  assign n9548 = ( ~n4455 & n9546 ) | ( ~n4455 & n9547 ) | ( n9546 & n9547 ) ;
  assign n9549 = ( n9542 & ~n9545 ) | ( n9542 & n9548 ) | ( ~n9545 & n9548 ) ;
  assign n9550 = n8886 & n8888 ;
  assign n9551 = n8886 | n8888 ;
  assign n9552 = ~n9550 & n9551 ;
  assign n9553 = n2893 & n9024 ;
  assign n9554 = ( ~n2886 & n9024 ) | ( ~n2886 & n9553 ) | ( n9024 & n9553 ) ;
  assign n9555 = n2701 & n9021 ;
  assign n9556 = ( ~n2784 & n9021 ) | ( ~n2784 & n9555 ) | ( n9021 & n9555 ) ;
  assign n9557 = n3507 & n9475 ;
  assign n9558 = ( n3483 & n9475 ) | ( n3483 & n9557 ) | ( n9475 & n9557 ) ;
  assign n9559 = n9556 | n9558 ;
  assign n9560 = n9554 | n9559 ;
  assign n9561 = n8970 | n9560 ;
  assign n9562 = n9560 & n9561 ;
  assign n9563 = ( n3603 & n9561 ) | ( n3603 & n9562 ) | ( n9561 & n9562 ) ;
  assign n9564 = x2 & n9562 ;
  assign n9565 = x2 & n9561 ;
  assign n9566 = ( n3603 & n9564 ) | ( n3603 & n9565 ) | ( n9564 & n9565 ) ;
  assign n9567 = x2 & ~n9564 ;
  assign n9568 = x2 & ~n9565 ;
  assign n9569 = ( ~n3603 & n9567 ) | ( ~n3603 & n9568 ) | ( n9567 & n9568 ) ;
  assign n9570 = ( n9563 & ~n9566 ) | ( n9563 & n9569 ) | ( ~n9566 & n9569 ) ;
  assign n9571 = n8731 | n8870 ;
  assign n9572 = n8869 | n9571 ;
  assign n9573 = n8867 | n9572 ;
  assign n9574 = ~n8872 & n9573 ;
  assign n9575 = n1634 & n9021 ;
  assign n9576 = ( n1630 & n9021 ) | ( n1630 & n9575 ) | ( n9021 & n9575 ) ;
  assign n9577 = n2279 & n9024 ;
  assign n9578 = ( ~n2269 & n9024 ) | ( ~n2269 & n9577 ) | ( n9024 & n9577 ) ;
  assign n9579 = n9576 | n9578 ;
  assign n9580 = n2090 & n9475 ;
  assign n9581 = ( ~n2082 & n9475 ) | ( ~n2082 & n9580 ) | ( n9475 & n9580 ) ;
  assign n9582 = n9579 | n9581 ;
  assign n9583 = n8970 | n9582 ;
  assign n9584 = n9582 & n9583 ;
  assign n9585 = ( n2568 & n9583 ) | ( n2568 & n9584 ) | ( n9583 & n9584 ) ;
  assign n9586 = x2 & n9584 ;
  assign n9587 = x2 & n9583 ;
  assign n9588 = ( n2568 & n9586 ) | ( n2568 & n9587 ) | ( n9586 & n9587 ) ;
  assign n9589 = x2 & ~n9586 ;
  assign n9590 = x2 & ~n9587 ;
  assign n9591 = ( ~n2568 & n9589 ) | ( ~n2568 & n9590 ) | ( n9589 & n9590 ) ;
  assign n9592 = ( n9585 & ~n9588 ) | ( n9585 & n9591 ) | ( ~n9588 & n9591 ) ;
  assign n9593 = n8858 & n8860 ;
  assign n9594 = n8858 | n8860 ;
  assign n9595 = ~n9593 & n9594 ;
  assign n9596 = n8850 | n8851 ;
  assign n9597 = n8834 | n9596 ;
  assign n9598 = ~n8853 & n9597 ;
  assign n9599 = ~n829 & n9024 ;
  assign n9600 = n352 & n9475 ;
  assign n9601 = ( ~n339 & n9475 ) | ( ~n339 & n9600 ) | ( n9475 & n9600 ) ;
  assign n9602 = n9599 | n9601 ;
  assign n9603 = n692 & n9021 ;
  assign n9604 = ( n674 & n9021 ) | ( n674 & n9603 ) | ( n9021 & n9603 ) ;
  assign n9605 = n9602 | n9604 ;
  assign n9606 = n8970 | n9604 ;
  assign n9607 = n9602 | n9606 ;
  assign n9608 = ( ~n1209 & n9605 ) | ( ~n1209 & n9607 ) | ( n9605 & n9607 ) ;
  assign n9609 = ~x2 & n9607 ;
  assign n9610 = ~x2 & n9605 ;
  assign n9611 = ( ~n1209 & n9609 ) | ( ~n1209 & n9610 ) | ( n9609 & n9610 ) ;
  assign n9612 = x2 | n9610 ;
  assign n9613 = x2 | n9609 ;
  assign n9614 = ( ~n1209 & n9612 ) | ( ~n1209 & n9613 ) | ( n9612 & n9613 ) ;
  assign n9615 = ( ~n9608 & n9611 ) | ( ~n9608 & n9614 ) | ( n9611 & n9614 ) ;
  assign n9616 = ~n829 & n9475 ;
  assign n9617 = ~n922 & n9021 ;
  assign n9618 = n9616 | n9617 ;
  assign n9619 = n692 & n9024 ;
  assign n9620 = ( n674 & n9024 ) | ( n674 & n9619 ) | ( n9024 & n9619 ) ;
  assign n9621 = n9618 | n9620 ;
  assign n9622 = n8970 | n9620 ;
  assign n9623 = n9618 | n9622 ;
  assign n9624 = ( n1554 & n9621 ) | ( n1554 & n9623 ) | ( n9621 & n9623 ) ;
  assign n9625 = x2 & n9623 ;
  assign n9626 = x2 & n9621 ;
  assign n9627 = ( n1554 & n9625 ) | ( n1554 & n9626 ) | ( n9625 & n9626 ) ;
  assign n9628 = x2 & ~n9626 ;
  assign n9629 = x2 & ~n9625 ;
  assign n9630 = ( ~n1554 & n9628 ) | ( ~n1554 & n9629 ) | ( n9628 & n9629 ) ;
  assign n9631 = ( n9624 & ~n9627 ) | ( n9624 & n9630 ) | ( ~n9627 & n9630 ) ;
  assign n9632 = x0 & x2 ;
  assign n9633 = n8969 & n9632 ;
  assign n9634 = n1538 & n9633 ;
  assign n9635 = ~n8969 & n9632 ;
  assign n9636 = n919 & n9635 ;
  assign n9637 = ( n918 & n9635 ) | ( n918 & n9636 ) | ( n9635 & n9636 ) ;
  assign n9638 = x2 & ~n9637 ;
  assign n9639 = x2 & ~n9632 ;
  assign n9640 = ( x2 & n8969 ) | ( x2 & n9639 ) | ( n8969 & n9639 ) ;
  assign n9641 = ( n916 & n9638 ) | ( n916 & n9640 ) | ( n9638 & n9640 ) ;
  assign n9642 = n9638 & n9640 ;
  assign n9643 = ( ~n874 & n9641 ) | ( ~n874 & n9642 ) | ( n9641 & n9642 ) ;
  assign n9644 = x2 & n9024 ;
  assign n9645 = n1042 & n9644 ;
  assign n9646 = ( ~n1027 & n9644 ) | ( ~n1027 & n9645 ) | ( n9644 & n9645 ) ;
  assign n9647 = n9643 & ~n9646 ;
  assign n9648 = ~n9633 & n9647 ;
  assign n9649 = ( ~n1946 & n9647 ) | ( ~n1946 & n9648 ) | ( n9647 & n9648 ) ;
  assign n9650 = ~n922 & n9024 ;
  assign n9651 = n1042 & n9021 ;
  assign n9652 = ( ~n1027 & n9021 ) | ( ~n1027 & n9651 ) | ( n9021 & n9651 ) ;
  assign n9653 = n9650 | n9652 ;
  assign n9654 = n692 & n9475 ;
  assign n9655 = ( n674 & n9475 ) | ( n674 & n9654 ) | ( n9475 & n9654 ) ;
  assign n9656 = x2 & n9655 ;
  assign n9657 = ( x2 & n9653 ) | ( x2 & n9656 ) | ( n9653 & n9656 ) ;
  assign n9658 = n9649 & ~n9657 ;
  assign n9659 = ~n9634 & n9658 ;
  assign n9660 = n8970 | n9475 ;
  assign n9661 = n1042 & n9660 ;
  assign n9662 = ( ~n1027 & n9660 ) | ( ~n1027 & n9661 ) | ( n9660 & n9661 ) ;
  assign n9663 = n9659 & ~n9662 ;
  assign n9664 = ( ~n1027 & n8820 ) | ( ~n1027 & n8822 ) | ( n8820 & n8822 ) ;
  assign n9665 = ( n9631 & n9663 ) | ( n9631 & n9664 ) | ( n9663 & n9664 ) ;
  assign n9666 = n9615 | n9665 ;
  assign n9667 = x5 | n8824 ;
  assign n9668 = ( ~n8817 & n8824 ) | ( ~n8817 & n9667 ) | ( n8824 & n9667 ) ;
  assign n9669 = n8818 | n9668 ;
  assign n9670 = ~n8827 & n9669 ;
  assign n9671 = n9666 & n9670 ;
  assign n9672 = n8827 | n8829 ;
  assign n9673 = x5 & ~n8827 ;
  assign n9674 = ( n8810 & n9672 ) | ( n8810 & ~n9673 ) | ( n9672 & ~n9673 ) ;
  assign n9675 = ~n8832 & n9674 ;
  assign n9676 = n9615 & n9665 ;
  assign n9677 = n9675 | n9676 ;
  assign n9678 = n9671 | n9677 ;
  assign n9679 = ~n829 & n9021 ;
  assign n9680 = n352 & n9024 ;
  assign n9681 = ( ~n339 & n9024 ) | ( ~n339 & n9680 ) | ( n9024 & n9680 ) ;
  assign n9682 = n9679 | n9681 ;
  assign n9683 = ~n523 & n9475 ;
  assign n9684 = n9682 | n9683 ;
  assign n9685 = n8970 | n9683 ;
  assign n9686 = n9682 | n9685 ;
  assign n9687 = ( ~n1055 & n9684 ) | ( ~n1055 & n9686 ) | ( n9684 & n9686 ) ;
  assign n9688 = ~x2 & n9686 ;
  assign n9689 = ~x2 & n9684 ;
  assign n9690 = ( ~n1055 & n9688 ) | ( ~n1055 & n9689 ) | ( n9688 & n9689 ) ;
  assign n9691 = x2 | n9689 ;
  assign n9692 = x2 | n9688 ;
  assign n9693 = ( ~n1055 & n9691 ) | ( ~n1055 & n9692 ) | ( n9691 & n9692 ) ;
  assign n9694 = ( ~n9687 & n9690 ) | ( ~n9687 & n9693 ) | ( n9690 & n9693 ) ;
  assign n9695 = n9678 & n9694 ;
  assign n9696 = n9675 & n9676 ;
  assign n9697 = ( n9671 & n9675 ) | ( n9671 & n9696 ) | ( n9675 & n9696 ) ;
  assign n9698 = ~n523 & n9024 ;
  assign n9699 = n352 & n9021 ;
  assign n9700 = ( ~n339 & n9021 ) | ( ~n339 & n9699 ) | ( n9021 & n9699 ) ;
  assign n9701 = n1793 & n9475 ;
  assign n9702 = ( n1783 & n9475 ) | ( n1783 & n9701 ) | ( n9475 & n9701 ) ;
  assign n9703 = n9700 | n9702 ;
  assign n9704 = n9698 | n9703 ;
  assign n9705 = n8970 | n9704 ;
  assign n9706 = n9704 & n9705 ;
  assign n9707 = ( n1884 & n9705 ) | ( n1884 & n9706 ) | ( n9705 & n9706 ) ;
  assign n9708 = x2 & n9706 ;
  assign n9709 = x2 & n9705 ;
  assign n9710 = ( n1884 & n9708 ) | ( n1884 & n9709 ) | ( n9708 & n9709 ) ;
  assign n9711 = x2 & ~n9708 ;
  assign n9712 = x2 & ~n9709 ;
  assign n9713 = ( ~n1884 & n9711 ) | ( ~n1884 & n9712 ) | ( n9711 & n9712 ) ;
  assign n9714 = ( n9707 & ~n9710 ) | ( n9707 & n9713 ) | ( ~n9710 & n9713 ) ;
  assign n9715 = n9697 | n9714 ;
  assign n9716 = n9695 | n9715 ;
  assign n9717 = n9598 & n9716 ;
  assign n9718 = n8854 & n8856 ;
  assign n9719 = n8854 | n8856 ;
  assign n9720 = ~n9718 & n9719 ;
  assign n9721 = n9697 & n9714 ;
  assign n9722 = ( n9695 & n9714 ) | ( n9695 & n9721 ) | ( n9714 & n9721 ) ;
  assign n9723 = n9720 | n9722 ;
  assign n9724 = n9717 | n9723 ;
  assign n9725 = ~n523 & n9021 ;
  assign n9726 = n1793 & n9024 ;
  assign n9727 = ( n1783 & n9024 ) | ( n1783 & n9726 ) | ( n9024 & n9726 ) ;
  assign n9728 = n9725 | n9727 ;
  assign n9729 = n1708 & n9475 ;
  assign n9730 = n9728 | n9729 ;
  assign n9731 = n8970 | n9729 ;
  assign n9732 = n9728 | n9731 ;
  assign n9733 = ( ~n1852 & n9730 ) | ( ~n1852 & n9732 ) | ( n9730 & n9732 ) ;
  assign n9734 = ~x2 & n9732 ;
  assign n9735 = ~x2 & n9730 ;
  assign n9736 = ( ~n1852 & n9734 ) | ( ~n1852 & n9735 ) | ( n9734 & n9735 ) ;
  assign n9737 = x2 | n9735 ;
  assign n9738 = x2 | n9734 ;
  assign n9739 = ( ~n1852 & n9737 ) | ( ~n1852 & n9738 ) | ( n9737 & n9738 ) ;
  assign n9740 = ( ~n9733 & n9736 ) | ( ~n9733 & n9739 ) | ( n9736 & n9739 ) ;
  assign n9741 = n9724 & n9740 ;
  assign n9742 = n9720 & n9722 ;
  assign n9743 = ( n9717 & n9720 ) | ( n9717 & n9742 ) | ( n9720 & n9742 ) ;
  assign n9744 = n1708 & n9024 ;
  assign n9745 = n1793 & n9021 ;
  assign n9746 = ( n1783 & n9021 ) | ( n1783 & n9745 ) | ( n9021 & n9745 ) ;
  assign n9747 = n1634 & n9475 ;
  assign n9748 = ( n1630 & n9475 ) | ( n1630 & n9747 ) | ( n9475 & n9747 ) ;
  assign n9749 = n9746 | n9748 ;
  assign n9750 = n9744 | n9749 ;
  assign n9751 = n8970 | n9750 ;
  assign n9752 = n9750 & n9751 ;
  assign n9753 = ( n1814 & n9751 ) | ( n1814 & n9752 ) | ( n9751 & n9752 ) ;
  assign n9754 = x2 & n9752 ;
  assign n9755 = x2 & n9751 ;
  assign n9756 = ( n1814 & n9754 ) | ( n1814 & n9755 ) | ( n9754 & n9755 ) ;
  assign n9757 = x2 & ~n9754 ;
  assign n9758 = x2 & ~n9755 ;
  assign n9759 = ( ~n1814 & n9757 ) | ( ~n1814 & n9758 ) | ( n9757 & n9758 ) ;
  assign n9760 = ( n9753 & ~n9756 ) | ( n9753 & n9759 ) | ( ~n9756 & n9759 ) ;
  assign n9761 = n9743 | n9760 ;
  assign n9762 = n9741 | n9761 ;
  assign n9763 = n9595 & n9762 ;
  assign n9764 = n1708 & n9021 ;
  assign n9765 = n1634 & n9024 ;
  assign n9766 = ( n1630 & n9024 ) | ( n1630 & n9765 ) | ( n9024 & n9765 ) ;
  assign n9767 = n2279 & n9475 ;
  assign n9768 = ( ~n2269 & n9475 ) | ( ~n2269 & n9767 ) | ( n9475 & n9767 ) ;
  assign n9769 = n9766 | n9768 ;
  assign n9770 = n9764 | n9769 ;
  assign n9771 = n8970 | n9770 ;
  assign n9772 = n9770 & n9771 ;
  assign n9773 = ( ~n2343 & n9771 ) | ( ~n2343 & n9772 ) | ( n9771 & n9772 ) ;
  assign n9774 = ~x2 & n9772 ;
  assign n9775 = ~x2 & n9771 ;
  assign n9776 = ( ~n2343 & n9774 ) | ( ~n2343 & n9775 ) | ( n9774 & n9775 ) ;
  assign n9777 = x2 | n9774 ;
  assign n9778 = x2 | n9775 ;
  assign n9779 = ( ~n2343 & n9777 ) | ( ~n2343 & n9778 ) | ( n9777 & n9778 ) ;
  assign n9780 = ( ~n9773 & n9776 ) | ( ~n9773 & n9779 ) | ( n9776 & n9779 ) ;
  assign n9781 = n9743 & n9760 ;
  assign n9782 = ( n9741 & n9760 ) | ( n9741 & n9781 ) | ( n9760 & n9781 ) ;
  assign n9783 = n9780 & n9782 ;
  assign n9784 = ( n9763 & n9780 ) | ( n9763 & n9783 ) | ( n9780 & n9783 ) ;
  assign n9785 = n9592 & n9784 ;
  assign n9786 = n9780 | n9782 ;
  assign n9787 = n9763 | n9786 ;
  assign n9788 = n8862 & ~n8863 ;
  assign n9789 = n8754 & ~n8863 ;
  assign n9790 = ( n9787 & n9788 ) | ( n9787 & n9789 ) | ( n9788 & n9789 ) ;
  assign n9791 = ( n9592 & n9785 ) | ( n9592 & n9790 ) | ( n9785 & n9790 ) ;
  assign n9792 = n9574 | n9791 ;
  assign n9793 = n9592 | n9784 ;
  assign n9794 = n9790 | n9793 ;
  assign n9795 = n8866 & ~n8867 ;
  assign n9796 = n8864 & ~n8867 ;
  assign n9797 = ( n9794 & n9795 ) | ( n9794 & n9796 ) | ( n9795 & n9796 ) ;
  assign n9798 = n9792 | n9797 ;
  assign n9799 = n2090 & n9024 ;
  assign n9800 = ( ~n2082 & n9024 ) | ( ~n2082 & n9799 ) | ( n9024 & n9799 ) ;
  assign n9801 = n2279 & n9021 ;
  assign n9802 = ( ~n2269 & n9021 ) | ( ~n2269 & n9801 ) | ( n9021 & n9801 ) ;
  assign n9803 = n2199 & n9475 ;
  assign n9804 = ( ~n2185 & n9475 ) | ( ~n2185 & n9803 ) | ( n9475 & n9803 ) ;
  assign n9805 = n9802 | n9804 ;
  assign n9806 = n9800 | n9805 ;
  assign n9807 = n8970 | n9806 ;
  assign n9808 = ( ~n2325 & n9806 ) | ( ~n2325 & n9807 ) | ( n9806 & n9807 ) ;
  assign n9809 = n9806 & n9807 ;
  assign n9810 = ( ~n2299 & n9808 ) | ( ~n2299 & n9809 ) | ( n9808 & n9809 ) ;
  assign n9811 = ~x2 & n9810 ;
  assign n9812 = x2 | n9810 ;
  assign n9813 = ( ~n9810 & n9811 ) | ( ~n9810 & n9812 ) | ( n9811 & n9812 ) ;
  assign n9814 = n9798 & n9813 ;
  assign n9815 = n8873 & n8876 ;
  assign n9816 = n8873 | n8876 ;
  assign n9817 = ~n9815 & n9816 ;
  assign n9818 = n9574 & n9791 ;
  assign n9819 = ( n9574 & n9797 ) | ( n9574 & n9818 ) | ( n9797 & n9818 ) ;
  assign n9820 = n9817 | n9819 ;
  assign n9821 = n9814 | n9820 ;
  assign n9822 = n2090 & n9021 ;
  assign n9823 = ( ~n2082 & n9021 ) | ( ~n2082 & n9822 ) | ( n9021 & n9822 ) ;
  assign n9824 = n2691 & n9475 ;
  assign n9825 = ( n2678 & n9475 ) | ( n2678 & n9824 ) | ( n9475 & n9824 ) ;
  assign n9826 = n2199 & n9024 ;
  assign n9827 = ( ~n2185 & n9024 ) | ( ~n2185 & n9826 ) | ( n9024 & n9826 ) ;
  assign n9828 = n9825 | n9827 ;
  assign n9829 = n9823 | n9828 ;
  assign n9830 = n8970 | n9829 ;
  assign n9831 = ( n2985 & n9829 ) | ( n2985 & n9830 ) | ( n9829 & n9830 ) ;
  assign n9832 = x2 & n9830 ;
  assign n9833 = x2 & n9829 ;
  assign n9834 = ( n2985 & n9832 ) | ( n2985 & n9833 ) | ( n9832 & n9833 ) ;
  assign n9835 = x2 & ~n9832 ;
  assign n9836 = x2 & ~n9833 ;
  assign n9837 = ( ~n2985 & n9835 ) | ( ~n2985 & n9836 ) | ( n9835 & n9836 ) ;
  assign n9838 = ( n9831 & ~n9834 ) | ( n9831 & n9837 ) | ( ~n9834 & n9837 ) ;
  assign n9839 = n9821 & n9838 ;
  assign n9840 = n8878 & n8880 ;
  assign n9841 = n8878 | n8880 ;
  assign n9842 = ~n9840 & n9841 ;
  assign n9843 = n9817 & n9819 ;
  assign n9844 = ( n9814 & n9817 ) | ( n9814 & n9843 ) | ( n9817 & n9843 ) ;
  assign n9845 = n9842 | n9844 ;
  assign n9846 = n9839 | n9845 ;
  assign n9847 = n2701 & n9475 ;
  assign n9848 = ( ~n2784 & n9475 ) | ( ~n2784 & n9847 ) | ( n9475 & n9847 ) ;
  assign n9849 = n2691 & n9024 ;
  assign n9850 = ( n2678 & n9024 ) | ( n2678 & n9849 ) | ( n9024 & n9849 ) ;
  assign n9851 = n9848 | n9850 ;
  assign n9852 = n2199 & n9021 ;
  assign n9853 = ( ~n2185 & n9021 ) | ( ~n2185 & n9852 ) | ( n9021 & n9852 ) ;
  assign n9854 = n9851 | n9853 ;
  assign n9855 = n8970 | n9853 ;
  assign n9856 = n9851 | n9855 ;
  assign n9857 = ( n2960 & n9854 ) | ( n2960 & n9856 ) | ( n9854 & n9856 ) ;
  assign n9858 = x2 & n9856 ;
  assign n9859 = x2 & n9854 ;
  assign n9860 = ( n2960 & n9858 ) | ( n2960 & n9859 ) | ( n9858 & n9859 ) ;
  assign n9861 = x2 & ~n9859 ;
  assign n9862 = x2 & ~n9858 ;
  assign n9863 = ( ~n2960 & n9861 ) | ( ~n2960 & n9862 ) | ( n9861 & n9862 ) ;
  assign n9864 = ( n9857 & ~n9860 ) | ( n9857 & n9863 ) | ( ~n9860 & n9863 ) ;
  assign n9865 = n9846 & n9864 ;
  assign n9866 = n2691 & n9021 ;
  assign n9867 = ( n2678 & n9021 ) | ( n2678 & n9866 ) | ( n9021 & n9866 ) ;
  assign n9868 = n2701 & n9024 ;
  assign n9869 = ( ~n2784 & n9024 ) | ( ~n2784 & n9868 ) | ( n9024 & n9868 ) ;
  assign n9870 = n9867 | n9869 ;
  assign n9871 = n2893 & n9475 ;
  assign n9872 = ( ~n2886 & n9475 ) | ( ~n2886 & n9871 ) | ( n9475 & n9871 ) ;
  assign n9873 = n9870 | n9872 ;
  assign n9874 = n8970 | n9873 ;
  assign n9875 = n9873 & n9874 ;
  assign n9876 = ( ~n2914 & n9874 ) | ( ~n2914 & n9875 ) | ( n9874 & n9875 ) ;
  assign n9877 = ~x2 & n9875 ;
  assign n9878 = ~x2 & n9874 ;
  assign n9879 = ( ~n2914 & n9877 ) | ( ~n2914 & n9878 ) | ( n9877 & n9878 ) ;
  assign n9880 = x2 | n9877 ;
  assign n9881 = x2 | n9878 ;
  assign n9882 = ( ~n2914 & n9880 ) | ( ~n2914 & n9881 ) | ( n9880 & n9881 ) ;
  assign n9883 = ( ~n9876 & n9879 ) | ( ~n9876 & n9882 ) | ( n9879 & n9882 ) ;
  assign n9884 = n9842 & n9844 ;
  assign n9885 = ( n9839 & n9842 ) | ( n9839 & n9884 ) | ( n9842 & n9884 ) ;
  assign n9886 = n9883 & n9885 ;
  assign n9887 = ( n9865 & n9883 ) | ( n9865 & n9886 ) | ( n9883 & n9886 ) ;
  assign n9888 = n9570 & n9887 ;
  assign n9889 = n8649 & ~n8882 ;
  assign n9890 = n9883 | n9885 ;
  assign n9891 = n9865 | n9890 ;
  assign n9892 = ( ~n8649 & n8882 ) | ( ~n8649 & n9889 ) | ( n8882 & n9889 ) ;
  assign n9893 = ( n9889 & n9891 ) | ( n9889 & n9892 ) | ( n9891 & n9892 ) ;
  assign n9894 = ( n9570 & n9888 ) | ( n9570 & n9893 ) | ( n9888 & n9893 ) ;
  assign n9895 = n2893 & n9021 ;
  assign n9896 = ( ~n2886 & n9021 ) | ( ~n2886 & n9895 ) | ( n9021 & n9895 ) ;
  assign n9897 = n3507 & n9024 ;
  assign n9898 = ( n3483 & n9024 ) | ( n3483 & n9897 ) | ( n9024 & n9897 ) ;
  assign n9899 = n9896 | n9898 ;
  assign n9900 = n3386 & n9475 ;
  assign n9902 = n8970 | n9900 ;
  assign n9903 = n9899 | n9902 ;
  assign n9901 = n9899 | n9900 ;
  assign n9904 = n9901 & n9903 ;
  assign n9905 = ( ~n3568 & n9903 ) | ( ~n3568 & n9904 ) | ( n9903 & n9904 ) ;
  assign n9906 = ~x2 & n9904 ;
  assign n9907 = ~x2 & n9903 ;
  assign n9908 = ( ~n3568 & n9906 ) | ( ~n3568 & n9907 ) | ( n9906 & n9907 ) ;
  assign n9909 = x2 | n9906 ;
  assign n9910 = x2 | n9907 ;
  assign n9911 = ( ~n3568 & n9909 ) | ( ~n3568 & n9910 ) | ( n9909 & n9910 ) ;
  assign n9912 = ( ~n9905 & n9908 ) | ( ~n9905 & n9911 ) | ( n9908 & n9911 ) ;
  assign n9913 = n9894 | n9912 ;
  assign n9914 = n8628 & ~n8884 ;
  assign n9915 = n9570 | n9887 ;
  assign n9916 = n9893 | n9915 ;
  assign n9917 = ( ~n8628 & n8884 ) | ( ~n8628 & n9914 ) | ( n8884 & n9914 ) ;
  assign n9918 = ( n9914 & n9916 ) | ( n9914 & n9917 ) | ( n9916 & n9917 ) ;
  assign n9919 = n9913 | n9918 ;
  assign n9920 = n9552 & n9919 ;
  assign n9921 = ( n8577 & n8578 ) | ( n8577 & ~n8890 ) | ( n8578 & ~n8890 ) ;
  assign n9922 = n8890 | n9921 ;
  assign n9923 = ~n8891 & n9922 ;
  assign n9924 = n9894 & n9912 ;
  assign n9925 = ( n9912 & n9918 ) | ( n9912 & n9924 ) | ( n9918 & n9924 ) ;
  assign n9926 = n9923 | n9925 ;
  assign n9927 = n9920 | n9926 ;
  assign n9928 = n3386 & n9024 ;
  assign n9929 = n3507 & n9021 ;
  assign n9930 = ( n3483 & n9021 ) | ( n3483 & n9929 ) | ( n9021 & n9929 ) ;
  assign n9931 = n3439 & n9475 ;
  assign n9932 = ( ~n3420 & n9475 ) | ( ~n3420 & n9931 ) | ( n9475 & n9931 ) ;
  assign n9933 = n9930 | n9932 ;
  assign n9934 = n9928 | n9933 ;
  assign n9935 = n8970 | n9934 ;
  assign n9936 = ( ~n3530 & n9934 ) | ( ~n3530 & n9935 ) | ( n9934 & n9935 ) ;
  assign n9937 = ~x2 & n9935 ;
  assign n9938 = ~x2 & n9934 ;
  assign n9939 = ( ~n3530 & n9937 ) | ( ~n3530 & n9938 ) | ( n9937 & n9938 ) ;
  assign n9940 = x2 | n9937 ;
  assign n9941 = x2 | n9938 ;
  assign n9942 = ( ~n3530 & n9940 ) | ( ~n3530 & n9941 ) | ( n9940 & n9941 ) ;
  assign n9943 = ( ~n9936 & n9939 ) | ( ~n9936 & n9942 ) | ( n9939 & n9942 ) ;
  assign n9944 = n9927 & n9943 ;
  assign n9945 = ( ~n8892 & n8915 ) | ( ~n8892 & n8916 ) | ( n8915 & n8916 ) ;
  assign n9946 = n8892 | n9945 ;
  assign n9947 = ~n8918 & n9946 ;
  assign n9948 = n9923 & n9925 ;
  assign n9949 = ( n9920 & n9923 ) | ( n9920 & n9948 ) | ( n9923 & n9948 ) ;
  assign n9950 = n9947 | n9949 ;
  assign n9951 = n9944 | n9950 ;
  assign n9952 = n4206 & n9475 ;
  assign n9953 = n3386 & n9021 ;
  assign n9954 = n3439 & n9024 ;
  assign n9955 = ( ~n3420 & n9024 ) | ( ~n3420 & n9954 ) | ( n9024 & n9954 ) ;
  assign n9956 = n9953 | n9955 ;
  assign n9957 = n9952 | n9956 ;
  assign n9958 = n8970 | n9952 ;
  assign n9959 = n9956 | n9958 ;
  assign n9960 = ( ~n4220 & n9957 ) | ( ~n4220 & n9959 ) | ( n9957 & n9959 ) ;
  assign n9961 = ~x2 & n9959 ;
  assign n9962 = ~x2 & n9957 ;
  assign n9963 = ( ~n4220 & n9961 ) | ( ~n4220 & n9962 ) | ( n9961 & n9962 ) ;
  assign n9964 = x2 | n9962 ;
  assign n9965 = x2 | n9961 ;
  assign n9966 = ( ~n4220 & n9964 ) | ( ~n4220 & n9965 ) | ( n9964 & n9965 ) ;
  assign n9967 = ( ~n9960 & n9963 ) | ( ~n9960 & n9966 ) | ( n9963 & n9966 ) ;
  assign n9968 = n9951 & n9967 ;
  assign n9969 = n8914 | n8920 ;
  assign n9970 = n8918 | n9969 ;
  assign n9971 = ~n8922 & n9970 ;
  assign n9972 = n9947 & n9949 ;
  assign n9973 = ( n9944 & n9947 ) | ( n9944 & n9972 ) | ( n9947 & n9972 ) ;
  assign n9974 = n9971 | n9973 ;
  assign n9975 = n9968 | n9974 ;
  assign n9976 = n4206 & n9024 ;
  assign n9977 = ~n4429 & n9475 ;
  assign n9978 = n3439 & n9021 ;
  assign n9979 = ( ~n3420 & n9021 ) | ( ~n3420 & n9978 ) | ( n9021 & n9978 ) ;
  assign n9980 = n9977 | n9979 ;
  assign n9981 = n9976 | n9980 ;
  assign n9982 = n8970 | n9976 ;
  assign n9983 = n9980 | n9982 ;
  assign n9984 = ( ~n4527 & n9981 ) | ( ~n4527 & n9983 ) | ( n9981 & n9983 ) ;
  assign n9985 = ~x2 & n9983 ;
  assign n9986 = ~x2 & n9981 ;
  assign n9987 = ( ~n4527 & n9985 ) | ( ~n4527 & n9986 ) | ( n9985 & n9986 ) ;
  assign n9988 = x2 | n9986 ;
  assign n9989 = x2 | n9985 ;
  assign n9990 = ( ~n4527 & n9988 ) | ( ~n4527 & n9989 ) | ( n9988 & n9989 ) ;
  assign n9991 = ( ~n9984 & n9987 ) | ( ~n9984 & n9990 ) | ( n9987 & n9990 ) ;
  assign n9992 = n9975 & n9991 ;
  assign n9993 = ~n4429 & n9024 ;
  assign n9994 = n9021 | n9024 ;
  assign n9995 = ( ~n4429 & n9021 ) | ( ~n4429 & n9994 ) | ( n9021 & n9994 ) ;
  assign n9996 = ( n4206 & n9993 ) | ( n4206 & n9995 ) | ( n9993 & n9995 ) ;
  assign n9997 = n4396 & n9475 ;
  assign n9999 = n8970 | n9997 ;
  assign n10000 = n9996 | n9999 ;
  assign n9998 = n9996 | n9997 ;
  assign n10001 = n9998 & n10000 ;
  assign n10002 = ( ~n4501 & n10000 ) | ( ~n4501 & n10001 ) | ( n10000 & n10001 ) ;
  assign n10003 = ~x2 & n10001 ;
  assign n10004 = ~x2 & n10000 ;
  assign n10005 = ( ~n4501 & n10003 ) | ( ~n4501 & n10004 ) | ( n10003 & n10004 ) ;
  assign n10006 = x2 | n10003 ;
  assign n10007 = x2 | n10004 ;
  assign n10008 = ( ~n4501 & n10006 ) | ( ~n4501 & n10007 ) | ( n10006 & n10007 ) ;
  assign n10009 = ( ~n10002 & n10005 ) | ( ~n10002 & n10008 ) | ( n10005 & n10008 ) ;
  assign n10010 = n9971 & n9973 ;
  assign n10011 = ( n9968 & n9971 ) | ( n9968 & n10010 ) | ( n9971 & n10010 ) ;
  assign n10012 = n10009 & n10011 ;
  assign n10013 = ( n9992 & n10009 ) | ( n9992 & n10012 ) | ( n10009 & n10012 ) ;
  assign n10014 = n9549 & n10013 ;
  assign n10015 = n8533 & ~n8923 ;
  assign n10016 = n10009 | n10011 ;
  assign n10017 = n9992 | n10016 ;
  assign n10018 = ( ~n8533 & n8923 ) | ( ~n8533 & n10015 ) | ( n8923 & n10015 ) ;
  assign n10019 = ( n10015 & n10017 ) | ( n10015 & n10018 ) | ( n10017 & n10018 ) ;
  assign n10020 = ( n9549 & n10014 ) | ( n9549 & n10019 ) | ( n10014 & n10019 ) ;
  assign n10021 = n9532 & n10020 ;
  assign n10022 = n8510 & ~n8925 ;
  assign n10023 = n9549 | n10013 ;
  assign n10024 = n10019 | n10023 ;
  assign n10025 = ( ~n8510 & n8925 ) | ( ~n8510 & n10022 ) | ( n8925 & n10022 ) ;
  assign n10026 = ( n10022 & n10024 ) | ( n10022 & n10025 ) | ( n10024 & n10025 ) ;
  assign n10027 = ( n9532 & n10021 ) | ( n9532 & n10026 ) | ( n10021 & n10026 ) ;
  assign n10028 = n8465 | n8931 ;
  assign n10029 = ~n8931 & n10028 ;
  assign n10030 = ( ~n8465 & n10028 ) | ( ~n8465 & n10029 ) | ( n10028 & n10029 ) ;
  assign n10031 = n10027 | n10030 ;
  assign n10032 = n9532 | n10020 ;
  assign n10033 = n10026 | n10032 ;
  assign n10034 = n8506 & ~n8928 ;
  assign n10035 = ( n8926 & ~n8928 ) | ( n8926 & n10034 ) | ( ~n8928 & n10034 ) ;
  assign n10036 = n8506 | n8926 ;
  assign n10037 = ( n8928 & n10035 ) | ( n8928 & ~n10036 ) | ( n10035 & ~n10036 ) ;
  assign n10038 = ( n10033 & n10035 ) | ( n10033 & n10037 ) | ( n10035 & n10037 ) ;
  assign n10039 = n10031 | n10038 ;
  assign n10040 = n4245 & n9021 ;
  assign n10041 = ( n4303 & n9021 ) | ( n4303 & n10040 ) | ( n9021 & n10040 ) ;
  assign n10042 = n5192 & n9024 ;
  assign n10043 = ( n5179 & n9024 ) | ( n5179 & n10042 ) | ( n9024 & n10042 ) ;
  assign n10044 = n10041 | n10043 ;
  assign n10045 = n5117 & n9475 ;
  assign n10046 = ( ~n5037 & n9475 ) | ( ~n5037 & n10045 ) | ( n9475 & n10045 ) ;
  assign n10047 = n10044 | n10046 ;
  assign n10048 = n8970 | n10046 ;
  assign n10049 = n10044 | n10048 ;
  assign n10050 = ( ~n5270 & n10047 ) | ( ~n5270 & n10049 ) | ( n10047 & n10049 ) ;
  assign n10051 = ~x2 & n10049 ;
  assign n10052 = ~x2 & n10047 ;
  assign n10053 = ( ~n5270 & n10051 ) | ( ~n5270 & n10052 ) | ( n10051 & n10052 ) ;
  assign n10054 = x2 | n10052 ;
  assign n10055 = x2 | n10051 ;
  assign n10056 = ( ~n5270 & n10054 ) | ( ~n5270 & n10055 ) | ( n10054 & n10055 ) ;
  assign n10057 = ( ~n10050 & n10053 ) | ( ~n10050 & n10056 ) | ( n10053 & n10056 ) ;
  assign n10058 = n10039 & n10057 ;
  assign n10059 = n10027 & n10030 ;
  assign n10060 = ( n10030 & n10038 ) | ( n10030 & n10059 ) | ( n10038 & n10059 ) ;
  assign n10061 = n8442 | n8933 ;
  assign n10062 = ~n8933 & n10061 ;
  assign n10063 = ( ~n8442 & n10061 ) | ( ~n8442 & n10062 ) | ( n10061 & n10062 ) ;
  assign n10064 = n10060 | n10063 ;
  assign n10065 = n10058 | n10064 ;
  assign n10066 = n5117 & n9024 ;
  assign n10067 = ( ~n5037 & n9024 ) | ( ~n5037 & n10066 ) | ( n9024 & n10066 ) ;
  assign n10068 = n5108 & n9475 ;
  assign n10069 = n5192 & n9021 ;
  assign n10070 = ( n5179 & n9021 ) | ( n5179 & n10069 ) | ( n9021 & n10069 ) ;
  assign n10071 = n10068 | n10070 ;
  assign n10072 = n10067 | n10071 ;
  assign n10073 = n8970 | n10072 ;
  assign n10074 = ( ~n5220 & n10072 ) | ( ~n5220 & n10073 ) | ( n10072 & n10073 ) ;
  assign n10075 = ~x2 & n10073 ;
  assign n10076 = ~x2 & n10072 ;
  assign n10077 = ( ~n5220 & n10075 ) | ( ~n5220 & n10076 ) | ( n10075 & n10076 ) ;
  assign n10078 = x2 | n10075 ;
  assign n10079 = x2 | n10076 ;
  assign n10080 = ( ~n5220 & n10078 ) | ( ~n5220 & n10079 ) | ( n10078 & n10079 ) ;
  assign n10081 = ( ~n10074 & n10077 ) | ( ~n10074 & n10080 ) | ( n10077 & n10080 ) ;
  assign n10082 = n10065 & n10081 ;
  assign n10083 = n8419 | n8439 ;
  assign n10084 = n8934 | n10083 ;
  assign n10085 = ~n8936 & n10084 ;
  assign n10086 = n10060 & n10063 ;
  assign n10087 = ( n10058 & n10063 ) | ( n10058 & n10086 ) | ( n10063 & n10086 ) ;
  assign n10088 = n10085 | n10087 ;
  assign n10089 = n10082 | n10088 ;
  assign n10090 = n5117 & n9021 ;
  assign n10091 = ( ~n5037 & n9021 ) | ( ~n5037 & n10090 ) | ( n9021 & n10090 ) ;
  assign n10092 = n5108 & n9024 ;
  assign n10093 = n5997 & n9475 ;
  assign n10094 = ( n5979 & n9475 ) | ( n5979 & n10093 ) | ( n9475 & n10093 ) ;
  assign n10095 = n10092 | n10094 ;
  assign n10096 = n10091 | n10095 ;
  assign n10097 = n8970 | n10096 ;
  assign n10098 = ( n6181 & n10096 ) | ( n6181 & n10097 ) | ( n10096 & n10097 ) ;
  assign n10099 = x2 & n10097 ;
  assign n10100 = x2 & n10096 ;
  assign n10101 = ( n6181 & n10099 ) | ( n6181 & n10100 ) | ( n10099 & n10100 ) ;
  assign n10102 = x2 & ~n10099 ;
  assign n10103 = x2 & ~n10100 ;
  assign n10104 = ( ~n6181 & n10102 ) | ( ~n6181 & n10103 ) | ( n10102 & n10103 ) ;
  assign n10105 = ( n10098 & ~n10101 ) | ( n10098 & n10104 ) | ( ~n10101 & n10104 ) ;
  assign n10106 = n10089 & n10105 ;
  assign n10107 = n5108 & n9021 ;
  assign n10108 = n5997 & n9024 ;
  assign n10109 = ( n5979 & n9024 ) | ( n5979 & n10108 ) | ( n9024 & n10108 ) ;
  assign n10110 = n10107 | n10109 ;
  assign n10111 = n5857 & n9475 ;
  assign n10112 = ( ~n5899 & n9475 ) | ( ~n5899 & n10111 ) | ( n9475 & n10111 ) ;
  assign n10113 = n10110 | n10112 ;
  assign n10114 = n8970 | n10113 ;
  assign n10115 = n10113 & n10114 ;
  assign n10116 = ( ~n6151 & n10114 ) | ( ~n6151 & n10115 ) | ( n10114 & n10115 ) ;
  assign n10117 = ~x2 & n10115 ;
  assign n10118 = ~x2 & n10114 ;
  assign n10119 = ( ~n6151 & n10117 ) | ( ~n6151 & n10118 ) | ( n10117 & n10118 ) ;
  assign n10120 = x2 | n10117 ;
  assign n10121 = x2 | n10118 ;
  assign n10122 = ( ~n6151 & n10120 ) | ( ~n6151 & n10121 ) | ( n10120 & n10121 ) ;
  assign n10123 = ( ~n10116 & n10119 ) | ( ~n10116 & n10122 ) | ( n10119 & n10122 ) ;
  assign n10124 = n10085 & n10087 ;
  assign n10125 = ( n10082 & n10085 ) | ( n10082 & n10124 ) | ( n10085 & n10124 ) ;
  assign n10126 = n10123 & n10125 ;
  assign n10127 = ( n10106 & n10123 ) | ( n10106 & n10126 ) | ( n10123 & n10126 ) ;
  assign n10128 = n9514 & n10127 ;
  assign n10129 = ~n8937 & n8939 ;
  assign n10130 = n10123 | n10125 ;
  assign n10131 = n10106 | n10130 ;
  assign n10132 = ( n8937 & ~n8939 ) | ( n8937 & n10129 ) | ( ~n8939 & n10129 ) ;
  assign n10133 = ( n10129 & n10131 ) | ( n10129 & n10132 ) | ( n10131 & n10132 ) ;
  assign n10134 = ( n9514 & n10128 ) | ( n9514 & n10133 ) | ( n10128 & n10133 ) ;
  assign n10135 = n5857 & n9021 ;
  assign n10136 = ( ~n5899 & n9021 ) | ( ~n5899 & n10135 ) | ( n9021 & n10135 ) ;
  assign n10137 = ~n6091 & n9024 ;
  assign n10138 = n7036 & n9475 ;
  assign n10139 = ( n7023 & n9475 ) | ( n7023 & n10138 ) | ( n9475 & n10138 ) ;
  assign n10140 = n10137 | n10139 ;
  assign n10141 = n10136 | n10140 ;
  assign n10142 = n8970 | n10141 ;
  assign n10143 = n10141 & n10142 ;
  assign n10144 = ( n7136 & n10142 ) | ( n7136 & n10143 ) | ( n10142 & n10143 ) ;
  assign n10145 = x2 & n10143 ;
  assign n10146 = x2 & n10142 ;
  assign n10147 = ( n7136 & n10145 ) | ( n7136 & n10146 ) | ( n10145 & n10146 ) ;
  assign n10148 = x2 & ~n10145 ;
  assign n10149 = x2 & ~n10146 ;
  assign n10150 = ( ~n7136 & n10148 ) | ( ~n7136 & n10149 ) | ( n10148 & n10149 ) ;
  assign n10151 = ( n10144 & ~n10147 ) | ( n10144 & n10150 ) | ( ~n10147 & n10150 ) ;
  assign n10152 = n10134 | n10151 ;
  assign n10153 = n8373 & ~n8941 ;
  assign n10154 = n9514 | n10127 ;
  assign n10155 = n10133 | n10154 ;
  assign n10156 = ( ~n8373 & n8941 ) | ( ~n8373 & n10153 ) | ( n8941 & n10153 ) ;
  assign n10157 = ( n10153 & n10155 ) | ( n10153 & n10156 ) | ( n10155 & n10156 ) ;
  assign n10158 = n10152 | n10157 ;
  assign n10159 = n9497 & n10158 ;
  assign n10160 = ( n8329 & n8330 ) | ( n8329 & ~n8947 ) | ( n8330 & ~n8947 ) ;
  assign n10161 = n8947 | n10160 ;
  assign n10162 = ~n8948 & n10161 ;
  assign n10163 = n10134 & n10151 ;
  assign n10164 = ( n10151 & n10157 ) | ( n10151 & n10163 ) | ( n10157 & n10163 ) ;
  assign n10165 = n10162 | n10164 ;
  assign n10166 = n10159 | n10165 ;
  assign n10167 = ~n6091 & n9021 ;
  assign n10168 = n7036 & n9024 ;
  assign n10169 = ( n7023 & n9024 ) | ( n7023 & n10168 ) | ( n9024 & n10168 ) ;
  assign n10170 = n10167 | n10169 ;
  assign n10171 = n6950 & n9475 ;
  assign n10172 = n10170 | n10171 ;
  assign n10173 = n8970 | n10172 ;
  assign n10174 = ( ~n7107 & n10172 ) | ( ~n7107 & n10173 ) | ( n10172 & n10173 ) ;
  assign n10175 = ~x2 & n10173 ;
  assign n10176 = ~x2 & n10172 ;
  assign n10177 = ( ~n7107 & n10175 ) | ( ~n7107 & n10176 ) | ( n10175 & n10176 ) ;
  assign n10178 = x2 | n10175 ;
  assign n10179 = x2 | n10176 ;
  assign n10180 = ( ~n7107 & n10178 ) | ( ~n7107 & n10179 ) | ( n10178 & n10179 ) ;
  assign n10181 = ( ~n10174 & n10177 ) | ( ~n10174 & n10180 ) | ( n10177 & n10180 ) ;
  assign n10182 = n10166 & n10181 ;
  assign n10183 = n8328 | n8950 ;
  assign n10184 = n8948 | n10183 ;
  assign n10185 = ~n8952 & n10184 ;
  assign n10186 = n10162 & n10164 ;
  assign n10187 = ( n10159 & n10162 ) | ( n10159 & n10186 ) | ( n10162 & n10186 ) ;
  assign n10188 = n10185 | n10187 ;
  assign n10189 = n10182 | n10188 ;
  assign n10190 = n6950 & n9024 ;
  assign n10191 = n7036 & n9021 ;
  assign n10192 = ( n7023 & n9021 ) | ( n7023 & n10191 ) | ( n9021 & n10191 ) ;
  assign n10193 = n10190 | n10192 ;
  assign n10194 = n6889 & n9475 ;
  assign n10195 = ( ~n6884 & n9475 ) | ( ~n6884 & n10194 ) | ( n9475 & n10194 ) ;
  assign n10196 = n10193 | n10195 ;
  assign n10197 = n8970 | n10195 ;
  assign n10198 = n10193 | n10197 ;
  assign n10199 = ( ~n7061 & n10196 ) | ( ~n7061 & n10198 ) | ( n10196 & n10198 ) ;
  assign n10200 = ~x2 & n10198 ;
  assign n10201 = ~x2 & n10196 ;
  assign n10202 = ( ~n7061 & n10200 ) | ( ~n7061 & n10201 ) | ( n10200 & n10201 ) ;
  assign n10203 = x2 | n10201 ;
  assign n10204 = x2 | n10200 ;
  assign n10205 = ( ~n7061 & n10203 ) | ( ~n7061 & n10204 ) | ( n10203 & n10204 ) ;
  assign n10206 = ( ~n10199 & n10202 ) | ( ~n10199 & n10205 ) | ( n10202 & n10205 ) ;
  assign n10207 = n10189 & n10206 ;
  assign n10208 = n10185 & n10187 ;
  assign n10209 = ( n10182 & n10185 ) | ( n10182 & n10208 ) | ( n10185 & n10208 ) ;
  assign n10210 = n6950 & n9021 ;
  assign n10211 = n6889 & n9024 ;
  assign n10212 = ( ~n6884 & n9024 ) | ( ~n6884 & n10211 ) | ( n9024 & n10211 ) ;
  assign n10213 = n10210 | n10212 ;
  assign n10214 = n7907 & n9475 ;
  assign n10215 = ( n7902 & n9475 ) | ( n7902 & n10214 ) | ( n9475 & n10214 ) ;
  assign n10217 = n8970 | n10215 ;
  assign n10218 = n10213 | n10217 ;
  assign n10216 = n10213 | n10215 ;
  assign n10219 = n10216 & n10218 ;
  assign n10220 = ( ~n8193 & n10218 ) | ( ~n8193 & n10219 ) | ( n10218 & n10219 ) ;
  assign n10221 = ~x2 & n10219 ;
  assign n10222 = ~x2 & n10218 ;
  assign n10223 = ( ~n8193 & n10221 ) | ( ~n8193 & n10222 ) | ( n10221 & n10222 ) ;
  assign n10224 = x2 | n10221 ;
  assign n10225 = x2 | n10222 ;
  assign n10226 = ( ~n8193 & n10224 ) | ( ~n8193 & n10225 ) | ( n10224 & n10225 ) ;
  assign n10227 = ( ~n10220 & n10223 ) | ( ~n10220 & n10226 ) | ( n10223 & n10226 ) ;
  assign n10228 = n10209 | n10227 ;
  assign n10229 = n10207 | n10228 ;
  assign n10230 = ( ~n8286 & n8953 ) | ( ~n8286 & n9494 ) | ( n8953 & n9494 ) ;
  assign n10231 = ( n9494 & n10229 ) | ( n9494 & n10230 ) | ( n10229 & n10230 ) ;
  assign n10232 = n10209 & n10227 ;
  assign n10233 = ( n10207 & n10227 ) | ( n10207 & n10232 ) | ( n10227 & n10232 ) ;
  assign n10234 = ~n9493 & n10233 ;
  assign n10235 = ( ~n9493 & n10231 ) | ( ~n9493 & n10234 ) | ( n10231 & n10234 ) ;
  assign n10236 = n8966 | n9086 ;
  assign n10237 = ~n9087 & n10236 ;
  assign n10238 = n8179 & ~n8961 ;
  assign n10239 = n8962 | n10238 ;
  assign n10240 = ~n9072 & n9440 ;
  assign n10241 = n9072 & ~n9440 ;
  assign n10242 = n10240 | n10241 ;
  assign n10243 = ~n8982 & n9475 ;
  assign n10244 = ( n9051 & n9475 ) | ( n9051 & n10243 ) | ( n9475 & n10243 ) ;
  assign n10245 = n9022 & n9024 ;
  assign n10246 = n10244 | n10245 ;
  assign n10247 = n9024 | n10244 ;
  assign n10248 = ( ~n9019 & n10246 ) | ( ~n9019 & n10247 ) | ( n10246 & n10247 ) ;
  assign n10249 = n9021 | n10248 ;
  assign n10250 = ( ~n8017 & n10248 ) | ( ~n8017 & n10249 ) | ( n10248 & n10249 ) ;
  assign n10251 = n8970 | n10250 ;
  assign n10252 = ( ~n10242 & n10250 ) | ( ~n10242 & n10251 ) | ( n10250 & n10251 ) ;
  assign n10253 = ~x2 & n10251 ;
  assign n10254 = ~x2 & n10250 ;
  assign n10255 = ( ~n10242 & n10253 ) | ( ~n10242 & n10254 ) | ( n10253 & n10254 ) ;
  assign n10256 = x2 | n10253 ;
  assign n10257 = x2 | n10254 ;
  assign n10258 = ( ~n10242 & n10256 ) | ( ~n10242 & n10257 ) | ( n10256 & n10257 ) ;
  assign n10259 = ( ~n10252 & n10255 ) | ( ~n10252 & n10258 ) | ( n10255 & n10258 ) ;
  assign n10260 = ~n10239 & n10259 ;
  assign n10261 = n10239 & ~n10259 ;
  assign n10262 = n10260 | n10261 ;
  assign n10263 = n8214 | n8959 ;
  assign n10264 = ~n8960 & n10263 ;
  assign n10265 = n8079 & n9021 ;
  assign n10266 = ( ~n8070 & n9021 ) | ( ~n8070 & n10265 ) | ( n9021 & n10265 ) ;
  assign n10267 = n9024 | n10266 ;
  assign n10268 = ( ~n8017 & n10266 ) | ( ~n8017 & n10267 ) | ( n10266 & n10267 ) ;
  assign n10269 = n9022 & n9475 ;
  assign n10270 = ( ~n9019 & n9475 ) | ( ~n9019 & n10269 ) | ( n9475 & n10269 ) ;
  assign n10272 = n8970 | n10270 ;
  assign n10273 = n10268 | n10272 ;
  assign n10271 = n10268 | n10270 ;
  assign n10274 = n10271 & n10273 ;
  assign n10275 = ( ~n9416 & n10273 ) | ( ~n9416 & n10274 ) | ( n10273 & n10274 ) ;
  assign n10276 = ~x2 & n10274 ;
  assign n10277 = ~x2 & n10273 ;
  assign n10278 = ( ~n9416 & n10276 ) | ( ~n9416 & n10277 ) | ( n10276 & n10277 ) ;
  assign n10279 = x2 | n10276 ;
  assign n10280 = x2 | n10277 ;
  assign n10281 = ( ~n9416 & n10279 ) | ( ~n9416 & n10280 ) | ( n10279 & n10280 ) ;
  assign n10282 = ( ~n10275 & n10278 ) | ( ~n10275 & n10281 ) | ( n10278 & n10281 ) ;
  assign n10283 = n10264 & n10282 ;
  assign n10284 = n10264 | n10282 ;
  assign n10285 = ~n10283 & n10284 ;
  assign n10286 = n8238 & ~n8957 ;
  assign n10287 = n8958 | n10286 ;
  assign n10293 = ~n8017 & n9475 ;
  assign n10288 = n7907 & n9021 ;
  assign n10289 = ( n7902 & n9021 ) | ( n7902 & n10288 ) | ( n9021 & n10288 ) ;
  assign n10290 = n8079 & n9024 ;
  assign n10291 = ( ~n8070 & n9024 ) | ( ~n8070 & n10290 ) | ( n9024 & n10290 ) ;
  assign n10292 = n10289 | n10291 ;
  assign n10295 = n8970 | n10292 ;
  assign n10296 = n10293 | n10295 ;
  assign n10294 = n10292 | n10293 ;
  assign n10297 = n10294 & n10296 ;
  assign n10298 = ( n8104 & n10296 ) | ( n8104 & n10297 ) | ( n10296 & n10297 ) ;
  assign n10299 = x2 & n10297 ;
  assign n10300 = x2 & n10296 ;
  assign n10301 = ( n8104 & n10299 ) | ( n8104 & n10300 ) | ( n10299 & n10300 ) ;
  assign n10302 = x2 & ~n10299 ;
  assign n10303 = x2 & ~n10300 ;
  assign n10304 = ( ~n8104 & n10302 ) | ( ~n8104 & n10303 ) | ( n10302 & n10303 ) ;
  assign n10305 = ( n10298 & ~n10301 ) | ( n10298 & n10304 ) | ( ~n10301 & n10304 ) ;
  assign n10306 = ~n10287 & n10305 ;
  assign n10307 = n10287 & ~n10305 ;
  assign n10308 = n10306 | n10307 ;
  assign n10309 = ~n10306 & n10308 ;
  assign n10310 = n10285 & ~n10309 ;
  assign n10311 = n10283 | n10310 ;
  assign n10312 = ~n10262 & n10311 ;
  assign n10313 = n10260 | n10312 ;
  assign n10314 = n10237 & n10313 ;
  assign n10315 = n9490 | n10306 ;
  assign n10316 = ( n10306 & ~n10308 ) | ( n10306 & n10315 ) | ( ~n10308 & n10315 ) ;
  assign n10317 = n10285 & n10316 ;
  assign n10318 = n10283 | n10317 ;
  assign n10319 = ~n10262 & n10318 ;
  assign n10320 = n10260 | n10319 ;
  assign n10321 = n10237 & n10320 ;
  assign n10322 = ( n10235 & n10314 ) | ( n10235 & n10321 ) | ( n10314 & n10321 ) ;
  assign n10323 = n9468 | n10322 ;
  assign n10324 = ( n9087 & n9467 ) | ( n9087 & n10322 ) | ( n9467 & n10322 ) ;
  assign n10325 = n10323 & ~n10324 ;
  assign n10326 = n9400 | n9406 ;
  assign n10327 = n9372 | n9379 ;
  assign n10328 = n1065 & n1708 ;
  assign n10329 = n1060 & n1793 ;
  assign n10330 = ( n1060 & n1783 ) | ( n1060 & n10329 ) | ( n1783 & n10329 ) ;
  assign n10331 = n1057 & n1634 ;
  assign n10332 = ( n1057 & n1630 ) | ( n1057 & n10331 ) | ( n1630 & n10331 ) ;
  assign n10333 = n10330 | n10332 ;
  assign n10334 = n10328 | n10333 ;
  assign n10335 = n1062 | n10334 ;
  assign n10336 = ( n1814 & n10334 ) | ( n1814 & n10335 ) | ( n10334 & n10335 ) ;
  assign n10337 = n292 | n399 ;
  assign n10338 = n356 | n10337 ;
  assign n10339 = n76 | n839 ;
  assign n10340 = n10338 | n10339 ;
  assign n10341 = n171 | n10340 ;
  assign n10342 = n1287 | n8996 ;
  assign n10343 = n557 | n10342 ;
  assign n10344 = n348 | n402 ;
  assign n10345 = n1336 | n10344 ;
  assign n10346 = n10343 | n10345 ;
  assign n10347 = n10341 | n10346 ;
  assign n10348 = n1615 | n2651 ;
  assign n10349 = n2666 | n10348 ;
  assign n10350 = n682 | n10349 ;
  assign n10351 = n233 | n457 ;
  assign n10352 = n340 | n901 ;
  assign n10353 = n10351 | n10352 ;
  assign n10354 = n312 | n10353 ;
  assign n10355 = n10350 | n10354 ;
  assign n10356 = n10347 | n10355 ;
  assign n10357 = n240 | n246 ;
  assign n10358 = n3983 | n10357 ;
  assign n10359 = n1232 | n1270 ;
  assign n10360 = n10358 | n10359 ;
  assign n10361 = n930 | n10360 ;
  assign n10362 = n193 | n261 ;
  assign n10363 = n1126 | n10362 ;
  assign n10364 = n306 | n607 ;
  assign n10365 = n437 | n10364 ;
  assign n10366 = n10363 | n10365 ;
  assign n10367 = n10361 | n10366 ;
  assign n10368 = n939 | n3444 ;
  assign n10369 = n330 | n479 ;
  assign n10370 = n92 | n10369 ;
  assign n10371 = n10368 | n10370 ;
  assign n10372 = n118 | n313 ;
  assign n10373 = n250 | n10372 ;
  assign n10374 = n10371 | n10373 ;
  assign n10375 = n1012 | n10374 ;
  assign n10376 = n10367 | n10375 ;
  assign n10377 = n10356 | n10376 ;
  assign n10378 = n161 | n10377 ;
  assign n10379 = n162 | n291 ;
  assign n10380 = n280 | n448 ;
  assign n10381 = n10379 | n10380 ;
  assign n10382 = n254 | n413 ;
  assign n10383 = x2 | n10382 ;
  assign n10384 = n10381 | n10383 ;
  assign n10385 = n4204 | n10384 ;
  assign n10386 = n10378 | n10385 ;
  assign n10387 = x2 & n10382 ;
  assign n10388 = ( x2 & n10381 ) | ( x2 & n10387 ) | ( n10381 & n10387 ) ;
  assign n10389 = ( x2 & n4204 ) | ( x2 & n10388 ) | ( n4204 & n10388 ) ;
  assign n10390 = x2 | n10388 ;
  assign n10391 = ( n10378 & n10389 ) | ( n10378 & n10390 ) | ( n10389 & n10390 ) ;
  assign n10392 = n1062 & ~n10391 ;
  assign n10393 = n10386 & n10392 ;
  assign n10394 = n10386 & ~n10391 ;
  assign n10395 = ( n10334 & n10393 ) | ( n10334 & n10394 ) | ( n10393 & n10394 ) ;
  assign n10396 = n10334 & n10394 ;
  assign n10397 = ( n1814 & n10395 ) | ( n1814 & n10396 ) | ( n10395 & n10396 ) ;
  assign n10398 = n10336 & ~n10397 ;
  assign n10399 = n10391 | n10395 ;
  assign n10400 = n10386 & ~n10399 ;
  assign n10401 = n10391 | n10394 ;
  assign n10402 = ( n10334 & n10391 ) | ( n10334 & n10401 ) | ( n10391 & n10401 ) ;
  assign n10403 = n10386 & ~n10402 ;
  assign n10404 = ( ~n1814 & n10400 ) | ( ~n1814 & n10403 ) | ( n10400 & n10403 ) ;
  assign n10405 = n10398 | n10404 ;
  assign n10406 = n9183 & n10404 ;
  assign n10407 = ( n9183 & n10398 ) | ( n9183 & n10406 ) | ( n10398 & n10406 ) ;
  assign n10408 = ( n9190 & n10405 ) | ( n9190 & n10407 ) | ( n10405 & n10407 ) ;
  assign n10409 = n9183 | n10404 ;
  assign n10410 = n10398 | n10409 ;
  assign n10411 = n9190 | n10410 ;
  assign n10412 = ~n10408 & n10411 ;
  assign n10413 = n1823 & n2090 ;
  assign n10414 = ( n1823 & ~n2082 ) | ( n1823 & n10413 ) | ( ~n2082 & n10413 ) ;
  assign n10415 = n1826 & n2279 ;
  assign n10416 = ( n1826 & ~n2269 ) | ( n1826 & n10415 ) | ( ~n2269 & n10415 ) ;
  assign n10417 = n1829 & n2199 ;
  assign n10418 = ( n1829 & ~n2185 ) | ( n1829 & n10417 ) | ( ~n2185 & n10417 ) ;
  assign n10419 = n10416 | n10418 ;
  assign n10420 = n10414 | n10419 ;
  assign n10421 = n1821 | n10420 ;
  assign n10422 = ( ~n2325 & n10420 ) | ( ~n2325 & n10421 ) | ( n10420 & n10421 ) ;
  assign n10423 = n10420 & n10421 ;
  assign n10424 = ( ~n2299 & n10422 ) | ( ~n2299 & n10423 ) | ( n10422 & n10423 ) ;
  assign n10425 = ~x29 & n10424 ;
  assign n10426 = x29 | n10424 ;
  assign n10427 = ( ~n10424 & n10425 ) | ( ~n10424 & n10426 ) | ( n10425 & n10426 ) ;
  assign n10428 = n10412 & n10427 ;
  assign n10429 = n10412 | n10427 ;
  assign n10430 = ~n10428 & n10429 ;
  assign n10431 = n9212 & n10430 ;
  assign n10432 = ( n9222 & n10430 ) | ( n9222 & n10431 ) | ( n10430 & n10431 ) ;
  assign n10433 = n9212 | n10430 ;
  assign n10434 = n9222 | n10433 ;
  assign n10435 = ~n10432 & n10434 ;
  assign n10436 = n2312 & n2691 ;
  assign n10437 = ( n2312 & n2678 ) | ( n2312 & n10436 ) | ( n2678 & n10436 ) ;
  assign n10438 = n2308 & n2701 ;
  assign n10439 = ( n2308 & ~n2784 ) | ( n2308 & n10438 ) | ( ~n2784 & n10438 ) ;
  assign n10440 = n10437 | n10439 ;
  assign n10441 = n2315 & n2893 ;
  assign n10442 = ( n2315 & ~n2886 ) | ( n2315 & n10441 ) | ( ~n2886 & n10441 ) ;
  assign n10443 = n10440 | n10442 ;
  assign n10444 = n2306 | n10443 ;
  assign n10445 = ( ~n2914 & n10443 ) | ( ~n2914 & n10444 ) | ( n10443 & n10444 ) ;
  assign n10446 = ~x26 & n10444 ;
  assign n10447 = ~x26 & n10443 ;
  assign n10448 = ( ~n2914 & n10446 ) | ( ~n2914 & n10447 ) | ( n10446 & n10447 ) ;
  assign n10449 = x26 | n10446 ;
  assign n10450 = x26 | n10447 ;
  assign n10451 = ( ~n2914 & n10449 ) | ( ~n2914 & n10450 ) | ( n10449 & n10450 ) ;
  assign n10452 = ( ~n10445 & n10448 ) | ( ~n10445 & n10451 ) | ( n10448 & n10451 ) ;
  assign n10453 = n10435 & n10452 ;
  assign n10454 = n10435 | n10452 ;
  assign n10455 = ~n10453 & n10454 ;
  assign n10456 = n9243 | n9246 ;
  assign n10457 = n9244 | n10456 ;
  assign n10458 = n10455 & n10457 ;
  assign n10459 = n9243 & n10455 ;
  assign n10460 = ( n9249 & n10458 ) | ( n9249 & n10459 ) | ( n10458 & n10459 ) ;
  assign n10461 = n10455 | n10457 ;
  assign n10462 = n9243 | n10455 ;
  assign n10463 = ( n9249 & n10461 ) | ( n9249 & n10462 ) | ( n10461 & n10462 ) ;
  assign n10464 = ~n10460 & n10463 ;
  assign n10465 = n2928 & n3386 ;
  assign n10466 = n2925 & n3507 ;
  assign n10467 = ( n2925 & n3483 ) | ( n2925 & n10466 ) | ( n3483 & n10466 ) ;
  assign n10468 = n2932 & n3439 ;
  assign n10469 = ( n2932 & ~n3420 ) | ( n2932 & n10468 ) | ( ~n3420 & n10468 ) ;
  assign n10470 = n10467 | n10469 ;
  assign n10471 = n10465 | n10470 ;
  assign n10472 = n2936 | n10471 ;
  assign n10473 = ( ~n3530 & n10471 ) | ( ~n3530 & n10472 ) | ( n10471 & n10472 ) ;
  assign n10474 = ~x23 & n10472 ;
  assign n10475 = ~x23 & n10471 ;
  assign n10476 = ( ~n3530 & n10474 ) | ( ~n3530 & n10475 ) | ( n10474 & n10475 ) ;
  assign n10477 = x23 | n10474 ;
  assign n10478 = x23 | n10475 ;
  assign n10479 = ( ~n3530 & n10477 ) | ( ~n3530 & n10478 ) | ( n10477 & n10478 ) ;
  assign n10480 = ( ~n10473 & n10476 ) | ( ~n10473 & n10479 ) | ( n10476 & n10479 ) ;
  assign n10481 = n10464 & n10480 ;
  assign n10482 = n10464 | n10480 ;
  assign n10483 = ~n10481 & n10482 ;
  assign n10484 = n9271 | n9274 ;
  assign n10485 = ( n9271 & n9276 ) | ( n9271 & n10484 ) | ( n9276 & n10484 ) ;
  assign n10486 = n10483 & n10485 ;
  assign n10487 = n10483 | n10485 ;
  assign n10488 = ~n10486 & n10487 ;
  assign n10489 = n3541 & ~n4429 ;
  assign n10490 = n3541 | n3544 ;
  assign n10491 = ( n3544 & ~n4429 ) | ( n3544 & n10490 ) | ( ~n4429 & n10490 ) ;
  assign n10492 = ( n4206 & n10489 ) | ( n4206 & n10491 ) | ( n10489 & n10491 ) ;
  assign n10493 = n3547 & n4396 ;
  assign n10494 = n10492 | n10493 ;
  assign n10495 = n3537 | n10493 ;
  assign n10496 = n10492 | n10495 ;
  assign n10497 = ( ~n4501 & n10494 ) | ( ~n4501 & n10496 ) | ( n10494 & n10496 ) ;
  assign n10498 = ~x20 & n10496 ;
  assign n10499 = ~x20 & n10494 ;
  assign n10500 = ( ~n4501 & n10498 ) | ( ~n4501 & n10499 ) | ( n10498 & n10499 ) ;
  assign n10501 = x20 | n10499 ;
  assign n10502 = x20 | n10498 ;
  assign n10503 = ( ~n4501 & n10501 ) | ( ~n4501 & n10502 ) | ( n10501 & n10502 ) ;
  assign n10504 = ( ~n10497 & n10500 ) | ( ~n10497 & n10503 ) | ( n10500 & n10503 ) ;
  assign n10505 = n10488 & n10504 ;
  assign n10506 = n10488 | n10504 ;
  assign n10507 = ~n10505 & n10506 ;
  assign n10508 = n9296 | n9299 ;
  assign n10509 = ( n9296 & n9301 ) | ( n9296 & n10508 ) | ( n9301 & n10508 ) ;
  assign n10510 = n10507 & n10509 ;
  assign n10511 = n10507 | n10509 ;
  assign n10512 = ~n10510 & n10511 ;
  assign n10513 = n4245 & n4466 ;
  assign n10514 = ( n4303 & n4466 ) | ( n4303 & n10513 ) | ( n4466 & n10513 ) ;
  assign n10515 = n4468 & n5192 ;
  assign n10516 = ( n4468 & n5179 ) | ( n4468 & n10515 ) | ( n5179 & n10515 ) ;
  assign n10517 = n10514 | n10516 ;
  assign n10518 = n4471 & n5117 ;
  assign n10519 = ( n4471 & ~n5037 ) | ( n4471 & n10518 ) | ( ~n5037 & n10518 ) ;
  assign n10520 = n10517 | n10519 ;
  assign n10521 = n4475 | n10519 ;
  assign n10522 = n10517 | n10521 ;
  assign n10523 = ( ~n5270 & n10520 ) | ( ~n5270 & n10522 ) | ( n10520 & n10522 ) ;
  assign n10524 = ~x17 & n10522 ;
  assign n10525 = ~x17 & n10520 ;
  assign n10526 = ( ~n5270 & n10524 ) | ( ~n5270 & n10525 ) | ( n10524 & n10525 ) ;
  assign n10527 = x17 | n10525 ;
  assign n10528 = x17 | n10524 ;
  assign n10529 = ( ~n5270 & n10527 ) | ( ~n5270 & n10528 ) | ( n10527 & n10528 ) ;
  assign n10530 = ( ~n10523 & n10526 ) | ( ~n10523 & n10529 ) | ( n10526 & n10529 ) ;
  assign n10531 = n10512 & n10530 ;
  assign n10532 = n10512 | n10530 ;
  assign n10533 = ~n10531 & n10532 ;
  assign n10534 = n9322 | n9324 ;
  assign n10535 = ( n9322 & n9326 ) | ( n9322 & n10534 ) | ( n9326 & n10534 ) ;
  assign n10536 = n10533 & n10535 ;
  assign n10537 = n10533 | n10535 ;
  assign n10538 = ~n10536 & n10537 ;
  assign n10539 = n5108 & n5237 ;
  assign n10540 = n5231 & n5997 ;
  assign n10541 = ( n5231 & n5979 ) | ( n5231 & n10540 ) | ( n5979 & n10540 ) ;
  assign n10542 = n10539 | n10541 ;
  assign n10543 = n5234 & n5857 ;
  assign n10544 = ( n5234 & ~n5899 ) | ( n5234 & n10543 ) | ( ~n5899 & n10543 ) ;
  assign n10545 = n10542 | n10544 ;
  assign n10546 = n5227 | n10545 ;
  assign n10547 = ( ~n6151 & n10545 ) | ( ~n6151 & n10546 ) | ( n10545 & n10546 ) ;
  assign n10548 = ~x14 & n10546 ;
  assign n10549 = ~x14 & n10545 ;
  assign n10550 = ( ~n6151 & n10548 ) | ( ~n6151 & n10549 ) | ( n10548 & n10549 ) ;
  assign n10551 = x14 | n10548 ;
  assign n10552 = x14 | n10549 ;
  assign n10553 = ( ~n6151 & n10551 ) | ( ~n6151 & n10552 ) | ( n10551 & n10552 ) ;
  assign n10554 = ( ~n10547 & n10550 ) | ( ~n10547 & n10553 ) | ( n10550 & n10553 ) ;
  assign n10555 = n10538 & n10554 ;
  assign n10556 = n10538 | n10554 ;
  assign n10557 = ~n10555 & n10556 ;
  assign n10558 = n9347 & n10557 ;
  assign n10559 = ( n9351 & n10557 ) | ( n9351 & n10558 ) | ( n10557 & n10558 ) ;
  assign n10560 = n9347 | n10557 ;
  assign n10561 = n9351 | n10560 ;
  assign n10562 = ~n10559 & n10561 ;
  assign n10563 = ~n6091 & n6125 ;
  assign n10564 = n6119 & n7036 ;
  assign n10565 = ( n6119 & n7023 ) | ( n6119 & n10564 ) | ( n7023 & n10564 ) ;
  assign n10566 = n10563 | n10565 ;
  assign n10567 = n6122 & n6950 ;
  assign n10568 = n10566 | n10567 ;
  assign n10569 = n6115 | n10568 ;
  assign n10570 = ( ~n7107 & n10568 ) | ( ~n7107 & n10569 ) | ( n10568 & n10569 ) ;
  assign n10571 = ~x11 & n10569 ;
  assign n10572 = ~x11 & n10568 ;
  assign n10573 = ( ~n7107 & n10571 ) | ( ~n7107 & n10572 ) | ( n10571 & n10572 ) ;
  assign n10574 = x11 | n10571 ;
  assign n10575 = x11 | n10572 ;
  assign n10576 = ( ~n7107 & n10574 ) | ( ~n7107 & n10575 ) | ( n10574 & n10575 ) ;
  assign n10577 = ( ~n10570 & n10573 ) | ( ~n10570 & n10576 ) | ( n10573 & n10576 ) ;
  assign n10578 = n10562 & n10577 ;
  assign n10579 = n10562 | n10577 ;
  assign n10580 = ~n10578 & n10579 ;
  assign n10581 = n9372 & n10580 ;
  assign n10582 = ( n9379 & n10580 ) | ( n9379 & n10581 ) | ( n10580 & n10581 ) ;
  assign n10583 = n10327 & ~n10582 ;
  assign n10584 = n6889 & n7074 ;
  assign n10585 = ( ~n6884 & n7074 ) | ( ~n6884 & n10584 ) | ( n7074 & n10584 ) ;
  assign n10586 = n7068 & n7907 ;
  assign n10587 = ( n7068 & n7902 ) | ( n7068 & n10586 ) | ( n7902 & n10586 ) ;
  assign n10588 = n7079 & n8079 ;
  assign n10589 = ( n7079 & ~n8070 ) | ( n7079 & n10588 ) | ( ~n8070 & n10588 ) ;
  assign n10590 = n10587 | n10589 ;
  assign n10591 = n10585 | n10590 ;
  assign n10592 = n7078 | n10591 ;
  assign n10593 = ( ~n8156 & n10591 ) | ( ~n8156 & n10592 ) | ( n10591 & n10592 ) ;
  assign n10594 = ~x8 & n10592 ;
  assign n10595 = ~x8 & n10591 ;
  assign n10596 = ( ~n8156 & n10594 ) | ( ~n8156 & n10595 ) | ( n10594 & n10595 ) ;
  assign n10597 = x8 | n10594 ;
  assign n10598 = x8 | n10595 ;
  assign n10599 = ( ~n8156 & n10597 ) | ( ~n8156 & n10598 ) | ( n10597 & n10598 ) ;
  assign n10600 = ( ~n10593 & n10596 ) | ( ~n10593 & n10599 ) | ( n10596 & n10599 ) ;
  assign n10601 = ~n9372 & n10580 ;
  assign n10602 = ~n9379 & n10601 ;
  assign n10603 = n10600 | n10602 ;
  assign n10604 = n10583 | n10603 ;
  assign n10605 = n10600 & n10602 ;
  assign n10606 = ( n10583 & n10600 ) | ( n10583 & n10605 ) | ( n10600 & n10605 ) ;
  assign n10607 = n10604 & ~n10606 ;
  assign n10608 = n9400 & n10607 ;
  assign n10609 = ( n9406 & n10607 ) | ( n9406 & n10608 ) | ( n10607 & n10608 ) ;
  assign n10610 = n10326 & ~n10609 ;
  assign n10611 = n10607 & ~n10609 ;
  assign n10612 = n10610 | n10611 ;
  assign n10613 = n8122 & ~n8982 ;
  assign n10614 = ( n8122 & n9051 ) | ( n8122 & n10613 ) | ( n9051 & n10613 ) ;
  assign n10615 = n8118 & n9022 ;
  assign n10616 = n10614 | n10615 ;
  assign n10617 = n8118 | n10614 ;
  assign n10618 = ( ~n9019 & n10616 ) | ( ~n9019 & n10617 ) | ( n10616 & n10617 ) ;
  assign n10619 = n8115 | n10618 ;
  assign n10620 = ( ~n8017 & n10618 ) | ( ~n8017 & n10619 ) | ( n10618 & n10619 ) ;
  assign n10621 = n8125 | n10620 ;
  assign n10622 = ( ~n10242 & n10620 ) | ( ~n10242 & n10621 ) | ( n10620 & n10621 ) ;
  assign n10623 = ~x5 & n10621 ;
  assign n10624 = ~x5 & n10620 ;
  assign n10625 = ( ~n10242 & n10623 ) | ( ~n10242 & n10624 ) | ( n10623 & n10624 ) ;
  assign n10626 = x5 | n10623 ;
  assign n10627 = x5 | n10624 ;
  assign n10628 = ( ~n10242 & n10626 ) | ( ~n10242 & n10627 ) | ( n10626 & n10627 ) ;
  assign n10629 = ( ~n10622 & n10625 ) | ( ~n10622 & n10628 ) | ( n10625 & n10628 ) ;
  assign n10630 = n10612 & n10629 ;
  assign n10631 = n10607 | n10629 ;
  assign n10632 = ( ~n10609 & n10629 ) | ( ~n10609 & n10631 ) | ( n10629 & n10631 ) ;
  assign n10633 = n10610 | n10632 ;
  assign n10634 = n9457 | n9460 ;
  assign n10635 = ( n9409 & n9457 ) | ( n9409 & n10634 ) | ( n9457 & n10634 ) ;
  assign n10636 = n10633 & n10635 ;
  assign n10637 = ~n10630 & n10636 ;
  assign n10638 = n10633 | n10635 ;
  assign n10639 = ( ~n10630 & n10635 ) | ( ~n10630 & n10638 ) | ( n10635 & n10638 ) ;
  assign n10640 = ~n10637 & n10639 ;
  assign n10641 = n9465 & n10640 ;
  assign n10642 = ( n9467 & n10640 ) | ( n9467 & n10641 ) | ( n10640 & n10641 ) ;
  assign n10643 = ( n9087 & n10640 ) | ( n9087 & n10641 ) | ( n10640 & n10641 ) ;
  assign n10644 = ( n10322 & n10642 ) | ( n10322 & n10643 ) | ( n10642 & n10643 ) ;
  assign n10645 = n9465 | n10640 ;
  assign n10646 = n9467 | n10645 ;
  assign n10647 = n9087 | n10645 ;
  assign n10648 = ( n10322 & n10646 ) | ( n10322 & n10647 ) | ( n10646 & n10647 ) ;
  assign n10649 = ~n10644 & n10648 ;
  assign n10650 = n10325 | n10649 ;
  assign n10651 = n10237 | n10313 ;
  assign n10652 = n10237 | n10320 ;
  assign n10653 = ( n10235 & n10651 ) | ( n10235 & n10652 ) | ( n10651 & n10652 ) ;
  assign n10654 = ~n10322 & n10653 ;
  assign n10655 = n10325 & n10654 ;
  assign n10656 = n10325 | n10654 ;
  assign n10657 = ~n10655 & n10656 ;
  assign n10658 = ( n10235 & n10312 ) | ( n10235 & n10319 ) | ( n10312 & n10319 ) ;
  assign n10659 = n10262 & ~n10311 ;
  assign n10660 = n10262 & ~n10318 ;
  assign n10661 = ( ~n10235 & n10659 ) | ( ~n10235 & n10660 ) | ( n10659 & n10660 ) ;
  assign n10662 = n10658 | n10661 ;
  assign n10663 = ( n10235 & n10310 ) | ( n10235 & n10317 ) | ( n10310 & n10317 ) ;
  assign n10664 = n10285 | n10316 ;
  assign n10665 = ~n10285 & n10309 ;
  assign n10666 = ( n10235 & n10664 ) | ( n10235 & ~n10665 ) | ( n10664 & ~n10665 ) ;
  assign n10667 = ~n10663 & n10666 ;
  assign n10668 = ~n10662 & n10667 ;
  assign n10669 = n10662 & ~n10667 ;
  assign n10670 = n10668 | n10669 ;
  assign n10671 = n9490 & ~n10308 ;
  assign n10672 = ( n10235 & ~n10308 ) | ( n10235 & n10671 ) | ( ~n10308 & n10671 ) ;
  assign n10673 = ~n9490 & n10308 ;
  assign n10674 = ~n10235 & n10673 ;
  assign n10675 = n10672 | n10674 ;
  assign n10676 = n9493 & ~n10233 ;
  assign n10677 = ~n10231 & n10676 ;
  assign n10678 = n10235 | n10677 ;
  assign n10679 = ~n10667 & n10678 ;
  assign n10680 = n10675 | n10679 ;
  assign n10681 = n10670 | n10680 ;
  assign n10682 = n10654 & ~n10662 ;
  assign n10683 = ~n10654 & n10662 ;
  assign n10684 = n10682 | n10683 ;
  assign n10685 = n10668 & ~n10684 ;
  assign n10686 = ( n10681 & n10684 ) | ( n10681 & ~n10685 ) | ( n10684 & ~n10685 ) ;
  assign n10687 = n10657 & n10682 ;
  assign n10688 = ( n10657 & ~n10686 ) | ( n10657 & n10687 ) | ( ~n10686 & n10687 ) ;
  assign n10689 = n10325 & n10649 ;
  assign n10690 = n10650 & ~n10689 ;
  assign n10691 = n10655 & n10690 ;
  assign n10692 = n10689 | n10691 ;
  assign n10693 = n10689 | n10690 ;
  assign n10694 = ( n10688 & n10692 ) | ( n10688 & n10693 ) | ( n10692 & n10693 ) ;
  assign n10695 = n10650 & ~n10694 ;
  assign n10696 = n1829 & n10649 ;
  assign n10697 = n1826 & n10654 ;
  assign n10698 = n1823 & n10325 ;
  assign n10699 = n10697 | n10698 ;
  assign n10700 = n10696 | n10699 ;
  assign n10701 = n10655 & ~n10690 ;
  assign n10702 = ( n10688 & ~n10690 ) | ( n10688 & n10701 ) | ( ~n10690 & n10701 ) ;
  assign n10703 = n1821 | n10696 ;
  assign n10704 = n10699 | n10703 ;
  assign n10705 = ( n10700 & n10702 ) | ( n10700 & n10704 ) | ( n10702 & n10704 ) ;
  assign n10706 = n10700 | n10704 ;
  assign n10707 = ( n10695 & n10705 ) | ( n10695 & n10706 ) | ( n10705 & n10706 ) ;
  assign n10708 = ~x29 & n10707 ;
  assign n10709 = x29 & n10704 ;
  assign n10710 = x29 & n10696 ;
  assign n10711 = ( x29 & n10699 ) | ( x29 & n10710 ) | ( n10699 & n10710 ) ;
  assign n10712 = ( n10702 & n10709 ) | ( n10702 & n10711 ) | ( n10709 & n10711 ) ;
  assign n10713 = n10709 | n10711 ;
  assign n10714 = ( n10695 & n10712 ) | ( n10695 & n10713 ) | ( n10712 & n10713 ) ;
  assign n10715 = x29 & ~n10714 ;
  assign n10716 = n10708 | n10715 ;
  assign n10717 = n1283 | n1340 ;
  assign n10718 = n619 | n10717 ;
  assign n10719 = n123 | n247 ;
  assign n10720 = n1521 | n10719 ;
  assign n10721 = n432 | n10720 ;
  assign n10722 = n2096 | n10721 ;
  assign n10723 = n10718 | n10722 ;
  assign n10724 = n2155 & ~n10723 ;
  assign n10725 = n401 | n638 ;
  assign n10726 = n273 | n758 ;
  assign n10727 = n10725 | n10726 ;
  assign n10728 = ( n4142 & ~n9136 ) | ( n4142 & n10727 ) | ( ~n9136 & n10727 ) ;
  assign n10729 = n438 | n9136 ;
  assign n10730 = n10728 | n10729 ;
  assign n10731 = n10724 & ~n10730 ;
  assign n10732 = n233 | n313 ;
  assign n10733 = n607 | n10732 ;
  assign n10734 = n6034 | n10733 ;
  assign n10735 = n1282 | n2116 ;
  assign n10736 = n178 | n418 ;
  assign n10737 = n141 | n10736 ;
  assign n10738 = n646 | n4184 ;
  assign n10739 = n10737 | n10738 ;
  assign n10740 = n771 | n2135 ;
  assign n10741 = n10739 | n10740 ;
  assign n10742 = n270 | n347 ;
  assign n10743 = n354 | n10742 ;
  assign n10744 = n2047 | n2053 ;
  assign n10745 = n171 | n246 ;
  assign n10746 = n10744 | n10745 ;
  assign n10747 = n10743 | n10746 ;
  assign n10748 = n10741 | n10747 ;
  assign n10749 = ( n10734 & n10735 ) | ( n10734 & ~n10748 ) | ( n10735 & ~n10748 ) ;
  assign n10750 = n202 | n667 ;
  assign n10751 = n3430 | n10750 ;
  assign n10752 = n405 | n654 ;
  assign n10753 = n886 | n10752 ;
  assign n10754 = n10751 | n10753 ;
  assign n10755 = n10748 | n10754 ;
  assign n10756 = n10749 | n10755 ;
  assign n10757 = n10731 & ~n10756 ;
  assign n10758 = n128 | n461 ;
  assign n10759 = n214 | n370 ;
  assign n10760 = n10758 | n10759 ;
  assign n10761 = n297 | n402 ;
  assign n10762 = n424 | n10761 ;
  assign n10763 = n10760 | n10762 ;
  assign n10764 = n390 | n10763 ;
  assign n10765 = n375 | n806 ;
  assign n10766 = n6853 | n10765 ;
  assign n10767 = n179 | n406 ;
  assign n10768 = n480 | n10767 ;
  assign n10769 = n10766 | n10768 ;
  assign n10770 = n133 | n223 ;
  assign n10771 = n118 | n277 ;
  assign n10772 = n10770 | n10771 ;
  assign n10773 = n555 | n820 ;
  assign n10774 = n39 | n10773 ;
  assign n10775 = n10772 | n10774 ;
  assign n10776 = n10769 | n10775 ;
  assign n10777 = n140 | n952 ;
  assign n10778 = n170 | n10777 ;
  assign n10779 = n10776 | n10778 ;
  assign n10780 = n10764 | n10779 ;
  assign n10781 = n10757 & ~n10780 ;
  assign n10782 = ~n10675 & n10678 ;
  assign n10783 = n10675 & ~n10678 ;
  assign n10784 = n10782 | n10783 ;
  assign n10785 = n646 | n3444 ;
  assign n10786 = n1620 | n10785 ;
  assign n10787 = n2255 | n7866 ;
  assign n10788 = n10786 | n10787 ;
  assign n10789 = n1296 | n10788 ;
  assign n10790 = n362 & ~n10789 ;
  assign n10791 = n305 | n886 ;
  assign n10792 = n1126 | n10791 ;
  assign n10793 = n375 | n10792 ;
  assign n10794 = n1499 | n7948 ;
  assign n10795 = n10793 | n10794 ;
  assign n10796 = n371 | n374 ;
  assign n10797 = n8038 | n10796 ;
  assign n10798 = n10795 | n10797 ;
  assign n10799 = n282 | n2135 ;
  assign n10800 = n152 | n228 ;
  assign n10801 = n277 | n10800 ;
  assign n10802 = n10799 | n10801 ;
  assign n10803 = n566 | n10802 ;
  assign n10804 = n457 | n1165 ;
  assign n10805 = n4328 | n10804 ;
  assign n10806 = n330 | n1039 ;
  assign n10807 = n198 | n434 ;
  assign n10808 = n10806 | n10807 ;
  assign n10809 = n10805 | n10808 ;
  assign n10810 = n10803 | n10809 ;
  assign n10811 = n10798 | n10810 ;
  assign n10812 = n177 | n764 ;
  assign n10813 = n183 | n643 ;
  assign n10814 = n568 | n10813 ;
  assign n10815 = n10812 | n10814 ;
  assign n10816 = n182 | n10815 ;
  assign n10817 = n1114 | n1723 ;
  assign n10818 = n2230 | n10817 ;
  assign n10819 = n10816 | n10818 ;
  assign n10820 = n10811 | n10819 ;
  assign n10821 = n10790 & ~n10820 ;
  assign n10822 = n214 | n406 ;
  assign n10823 = n4262 | n10822 ;
  assign n10824 = n424 | n10823 ;
  assign n10825 = n10821 & ~n10824 ;
  assign n10826 = n1062 | n1065 ;
  assign n10827 = ( n1062 & ~n10678 ) | ( n1062 & n10826 ) | ( ~n10678 & n10826 ) ;
  assign n10828 = n1057 & ~n10825 ;
  assign n10829 = ~n10675 & n10828 ;
  assign n10830 = ( ~n10825 & n10827 ) | ( ~n10825 & n10829 ) | ( n10827 & n10829 ) ;
  assign n10831 = n1065 & ~n10678 ;
  assign n10832 = ( ~n10825 & n10829 ) | ( ~n10825 & n10831 ) | ( n10829 & n10831 ) ;
  assign n10833 = ( n10784 & n10830 ) | ( n10784 & n10832 ) | ( n10830 & n10832 ) ;
  assign n10834 = ~n10781 & n10833 ;
  assign n10835 = ~n10667 & n10782 ;
  assign n10836 = n10667 & ~n10782 ;
  assign n10837 = n10835 | n10836 ;
  assign n10838 = n1062 & n10837 ;
  assign n10839 = n1057 & n10667 ;
  assign n10840 = n1060 & ~n10678 ;
  assign n10841 = n1065 & ~n10675 ;
  assign n10842 = n10840 | n10841 ;
  assign n10843 = n10839 | n10842 ;
  assign n10844 = n10838 | n10843 ;
  assign n10845 = n10781 & ~n10833 ;
  assign n10846 = n10834 | n10845 ;
  assign n10847 = n10844 & ~n10846 ;
  assign n10848 = n10834 | n10847 ;
  assign n10849 = n10670 & n10680 ;
  assign n10850 = n10681 & ~n10849 ;
  assign n10851 = n839 | n1016 ;
  assign n10852 = n168 | n938 ;
  assign n10853 = n480 | n10852 ;
  assign n10854 = n10851 | n10853 ;
  assign n10855 = n3412 | n10854 ;
  assign n10856 = n3295 | n3298 ;
  assign n10857 = n10855 | n10856 ;
  assign n10858 = n1521 | n5983 ;
  assign n10859 = n246 | n311 ;
  assign n10860 = n10858 | n10859 ;
  assign n10861 = n59 | n820 ;
  assign n10862 = n203 | n372 ;
  assign n10863 = n10861 | n10862 ;
  assign n10864 = n566 | n623 ;
  assign n10865 = n348 | n758 ;
  assign n10866 = n10864 | n10865 ;
  assign n10867 = n10863 | n10866 ;
  assign n10868 = n10860 | n10867 ;
  assign n10869 = n1675 | n2053 ;
  assign n10870 = n236 | n1785 ;
  assign n10871 = n10869 | n10870 ;
  assign n10872 = n71 | n171 ;
  assign n10873 = n10871 | n10872 ;
  assign n10874 = n10868 | n10873 ;
  assign n10875 = n10857 | n10874 ;
  assign n10876 = n497 | n10875 ;
  assign n10877 = n53 | n648 ;
  assign n10878 = n2117 | n10877 ;
  assign n10879 = n141 | n654 ;
  assign n10880 = n363 | n10879 ;
  assign n10881 = n10878 | n10880 ;
  assign n10882 = n155 | n448 ;
  assign n10883 = n443 | n10882 ;
  assign n10884 = n10881 | n10883 ;
  assign n10885 = n4008 | n4009 ;
  assign n10886 = n163 | n292 ;
  assign n10887 = n234 | n10886 ;
  assign n10888 = n533 | n10887 ;
  assign n10889 = n605 | n10888 ;
  assign n10890 = n10885 | n10889 ;
  assign n10891 = n10884 | n10890 ;
  assign n10892 = n402 | n434 ;
  assign n10893 = n254 | n10892 ;
  assign n10894 = n4314 | n10893 ;
  assign n10895 = n357 | n722 ;
  assign n10896 = n5946 | n10895 ;
  assign n10897 = n10894 | n10896 ;
  assign n10898 = n2696 | n2856 ;
  assign n10899 = n296 | n457 ;
  assign n10900 = n10898 | n10899 ;
  assign n10901 = n616 | n720 ;
  assign n10902 = n278 | n303 ;
  assign n10903 = n10901 | n10902 ;
  assign n10904 = n159 | n405 ;
  assign n10905 = n10903 | n10904 ;
  assign n10906 = n10900 | n10905 ;
  assign n10907 = n10897 | n10906 ;
  assign n10908 = n1002 | n5923 ;
  assign n10909 = n6891 | n10908 ;
  assign n10910 = n179 | n1172 ;
  assign n10911 = n340 | n388 ;
  assign n10912 = n10910 | n10911 ;
  assign n10913 = n10909 | n10912 ;
  assign n10914 = n237 | n489 ;
  assign n10915 = n515 | n10914 ;
  assign n10916 = n263 | n10915 ;
  assign n10917 = n245 | n10916 ;
  assign n10918 = n10913 | n10917 ;
  assign n10919 = n10907 | n10918 ;
  assign n10920 = n7954 | n10919 ;
  assign n10921 = ( ~n10876 & n10891 ) | ( ~n10876 & n10920 ) | ( n10891 & n10920 ) ;
  assign n10922 = n923 | n2188 ;
  assign n10923 = n344 | n418 ;
  assign n10924 = n297 | n10923 ;
  assign n10925 = n10922 | n10924 ;
  assign n10926 = n302 | n10925 ;
  assign n10927 = n10876 | n10926 ;
  assign n10928 = n10921 | n10927 ;
  assign n10929 = n1065 & n10667 ;
  assign n10930 = n1060 & ~n10675 ;
  assign n10931 = n10929 | n10930 ;
  assign n10932 = n1057 & ~n10662 ;
  assign n10933 = n1062 | n10932 ;
  assign n10934 = n10931 | n10933 ;
  assign n10935 = n10928 & n10934 ;
  assign n10936 = n10931 | n10932 ;
  assign n10937 = n10928 & n10936 ;
  assign n10938 = ( n10850 & n10935 ) | ( n10850 & n10937 ) | ( n10935 & n10937 ) ;
  assign n10939 = n10928 | n10934 ;
  assign n10940 = n10928 | n10936 ;
  assign n10941 = ( n10850 & n10939 ) | ( n10850 & n10940 ) | ( n10939 & n10940 ) ;
  assign n10942 = ~n10938 & n10941 ;
  assign n10943 = n10848 & ~n10942 ;
  assign n10944 = ~n10848 & n10942 ;
  assign n10945 = n10943 | n10944 ;
  assign n10946 = n10716 & n10945 ;
  assign n10947 = n10716 | n10945 ;
  assign n10948 = ~n10946 & n10947 ;
  assign n10949 = n10657 & ~n10688 ;
  assign n10950 = n1829 & n10325 ;
  assign n10951 = n1826 & ~n10662 ;
  assign n10952 = n1823 & n10654 ;
  assign n10953 = n10951 | n10952 ;
  assign n10954 = n10950 | n10953 ;
  assign n10955 = n1821 | n10954 ;
  assign n10956 = ~n10657 & n10682 ;
  assign n10957 = ( n10657 & n10686 ) | ( n10657 & ~n10956 ) | ( n10686 & ~n10956 ) ;
  assign n10958 = ( n10954 & n10955 ) | ( n10954 & ~n10957 ) | ( n10955 & ~n10957 ) ;
  assign n10959 = n10954 | n10955 ;
  assign n10960 = ( n10949 & n10958 ) | ( n10949 & n10959 ) | ( n10958 & n10959 ) ;
  assign n10961 = ~x29 & n10960 ;
  assign n10962 = x29 & n10954 ;
  assign n10963 = x29 & n1821 ;
  assign n10964 = ( x29 & n10954 ) | ( x29 & n10963 ) | ( n10954 & n10963 ) ;
  assign n10965 = ( ~n10957 & n10962 ) | ( ~n10957 & n10964 ) | ( n10962 & n10964 ) ;
  assign n10966 = n10962 | n10964 ;
  assign n10967 = ( n10949 & n10965 ) | ( n10949 & n10966 ) | ( n10965 & n10966 ) ;
  assign n10968 = x29 & ~n10967 ;
  assign n10969 = n10961 | n10968 ;
  assign n10970 = n10844 & ~n10847 ;
  assign n10971 = n10846 | n10847 ;
  assign n10972 = ~n10970 & n10971 ;
  assign n10973 = n10969 & ~n10972 ;
  assign n10974 = ~n10969 & n10972 ;
  assign n10975 = n10973 | n10974 ;
  assign n10976 = ~n10668 & n10684 ;
  assign n10977 = n10681 & n10976 ;
  assign n10978 = n10686 & ~n10977 ;
  assign n10979 = n1826 & n10667 ;
  assign n10980 = n1823 & ~n10662 ;
  assign n10981 = n10979 | n10980 ;
  assign n10982 = n1829 & n10654 ;
  assign n10983 = n1821 | n10982 ;
  assign n10984 = n10981 | n10983 ;
  assign n10985 = ~x29 & n10984 ;
  assign n10986 = n10981 | n10982 ;
  assign n10987 = ~x29 & n10986 ;
  assign n10988 = ( n10978 & n10985 ) | ( n10978 & n10987 ) | ( n10985 & n10987 ) ;
  assign n10989 = x29 & n10984 ;
  assign n10990 = x29 & ~n10989 ;
  assign n10991 = x29 & n10982 ;
  assign n10992 = ( x29 & n10981 ) | ( x29 & n10991 ) | ( n10981 & n10991 ) ;
  assign n10993 = x29 & ~n10992 ;
  assign n10994 = ( ~n10978 & n10990 ) | ( ~n10978 & n10993 ) | ( n10990 & n10993 ) ;
  assign n10995 = n10988 | n10994 ;
  assign n10996 = n1057 & ~n10675 ;
  assign n10997 = n10827 | n10996 ;
  assign n10998 = n10831 | n10996 ;
  assign n10999 = ( n10784 & n10997 ) | ( n10784 & n10998 ) | ( n10997 & n10998 ) ;
  assign n11000 = n10825 | n10999 ;
  assign n11001 = ~n10825 & n10999 ;
  assign n11002 = ( ~n10999 & n11000 ) | ( ~n10999 & n11001 ) | ( n11000 & n11001 ) ;
  assign n11003 = n10995 & ~n11002 ;
  assign n11004 = ~n10995 & n11002 ;
  assign n11005 = n11003 | n11004 ;
  assign n11006 = n2005 & ~n10678 ;
  assign n11007 = n1829 & ~n10662 ;
  assign n11008 = n1826 & ~n10675 ;
  assign n11009 = n1823 & n10667 ;
  assign n11010 = n11008 | n11009 ;
  assign n11011 = n11007 | n11010 ;
  assign n11012 = n1821 | n11007 ;
  assign n11013 = n11010 | n11012 ;
  assign n11014 = ( n10850 & n11011 ) | ( n10850 & n11013 ) | ( n11011 & n11013 ) ;
  assign n11015 = x29 & n11013 ;
  assign n11016 = x29 & n11011 ;
  assign n11017 = ( n10850 & n11015 ) | ( n10850 & n11016 ) | ( n11015 & n11016 ) ;
  assign n11018 = x29 & ~n11017 ;
  assign n11019 = ( n11014 & ~n11017 ) | ( n11014 & n11018 ) | ( ~n11017 & n11018 ) ;
  assign n11020 = n1829 & n10667 ;
  assign n11021 = n1826 & ~n10678 ;
  assign n11022 = n1823 & ~n10675 ;
  assign n11023 = n11021 | n11022 ;
  assign n11024 = n11020 | n11023 ;
  assign n11025 = n10837 | n11024 ;
  assign n11026 = n1821 | n11020 ;
  assign n11027 = n11023 | n11026 ;
  assign n11028 = n11025 & n11027 ;
  assign n11029 = ~x29 & n11027 ;
  assign n11030 = n11025 & n11029 ;
  assign n11031 = x29 | n11030 ;
  assign n11032 = ( ~n11028 & n11030 ) | ( ~n11028 & n11031 ) | ( n11030 & n11031 ) ;
  assign n11033 = n1821 & n10784 ;
  assign n11034 = n1823 & ~n10678 ;
  assign n11035 = n1829 & ~n10675 ;
  assign n11036 = n11034 | n11035 ;
  assign n11037 = x29 | n11036 ;
  assign n11038 = n11033 | n11037 ;
  assign n11039 = ~x29 & n11038 ;
  assign n11040 = x29 & ~n1820 ;
  assign n11041 = ( x29 & n10678 ) | ( x29 & n11040 ) | ( n10678 & n11040 ) ;
  assign n11042 = n11038 & n11041 ;
  assign n11043 = n11033 | n11036 ;
  assign n11044 = n11041 & ~n11043 ;
  assign n11045 = ( n11039 & n11042 ) | ( n11039 & n11044 ) | ( n11042 & n11044 ) ;
  assign n11046 = n11032 & n11045 ;
  assign n11047 = ( n11006 & n11019 ) | ( n11006 & n11046 ) | ( n11019 & n11046 ) ;
  assign n11048 = ~n11005 & n11047 ;
  assign n11049 = n11003 | n11048 ;
  assign n11050 = ~n10975 & n11049 ;
  assign n11051 = n10973 | n11050 ;
  assign n11052 = n10948 & n11051 ;
  assign n11053 = n10948 | n11051 ;
  assign n11054 = ~n11052 & n11053 ;
  assign n11055 = n8115 & ~n9022 ;
  assign n11056 = n8118 & ~n8982 ;
  assign n11057 = ( n8118 & n9051 ) | ( n8118 & n11056 ) | ( n9051 & n11056 ) ;
  assign n11058 = ( n8115 & ~n11055 ) | ( n8115 & n11057 ) | ( ~n11055 & n11057 ) ;
  assign n11059 = n8115 | n11057 ;
  assign n11060 = ( ~n9019 & n11058 ) | ( ~n9019 & n11059 ) | ( n11058 & n11059 ) ;
  assign n11061 = n8125 | n11060 ;
  assign n11062 = ( n9078 & n11060 ) | ( n9078 & n11061 ) | ( n11060 & n11061 ) ;
  assign n11063 = x5 & n11061 ;
  assign n11064 = x5 & n11060 ;
  assign n11065 = ( n9078 & n11063 ) | ( n9078 & n11064 ) | ( n11063 & n11064 ) ;
  assign n11066 = x5 & ~n11063 ;
  assign n11067 = x5 & ~n11064 ;
  assign n11068 = ( ~n9078 & n11066 ) | ( ~n9078 & n11067 ) | ( n11066 & n11067 ) ;
  assign n11069 = ( n11062 & ~n11065 ) | ( n11062 & n11068 ) | ( ~n11065 & n11068 ) ;
  assign n11070 = n10582 & n11069 ;
  assign n11071 = ( n10606 & n11069 ) | ( n10606 & n11070 ) | ( n11069 & n11070 ) ;
  assign n11072 = n10582 | n11069 ;
  assign n11073 = n10606 | n11072 ;
  assign n11074 = ~n11071 & n11073 ;
  assign n11151 = n10408 | n10427 ;
  assign n11152 = ( n10408 & n10412 ) | ( n10408 & n11151 ) | ( n10412 & n11151 ) ;
  assign n11075 = ( n1814 & n10399 ) | ( n1814 & n10402 ) | ( n10399 & n10402 ) ;
  assign n11076 = n340 | n447 ;
  assign n11077 = n5072 | n11076 ;
  assign n11078 = n1662 | n9150 ;
  assign n11079 = n11077 | n11078 ;
  assign n11080 = n950 | n11079 ;
  assign n11081 = n757 | n1364 ;
  assign n11082 = n67 | n209 ;
  assign n11083 = n341 | n11082 ;
  assign n11084 = n11081 | n11083 ;
  assign n11085 = n255 | n607 ;
  assign n11086 = n192 | n11085 ;
  assign n11087 = n725 | n841 ;
  assign n11088 = n310 | n344 ;
  assign n11089 = n11087 | n11088 ;
  assign n11090 = n11086 | n11089 ;
  assign n11091 = n11084 | n11090 ;
  assign n11092 = ( ~n758 & n11080 ) | ( ~n758 & n11091 ) | ( n11080 & n11091 ) ;
  assign n11093 = n11080 & n11091 ;
  assign n11094 = ( ~n5873 & n11092 ) | ( ~n5873 & n11093 ) | ( n11092 & n11093 ) ;
  assign n11095 = n5874 | n11094 ;
  assign n11096 = n1270 | n3987 ;
  assign n11097 = n457 | n720 ;
  assign n11098 = n270 | n11097 ;
  assign n11099 = n11096 | n11098 ;
  assign n11100 = n375 | n11099 ;
  assign n11101 = n6013 | n6014 ;
  assign n11102 = n496 | n11101 ;
  assign n11103 = n11100 | n11102 ;
  assign n11104 = n1607 | n1615 ;
  assign n11105 = n2053 | n11104 ;
  assign n11106 = n11103 | n11105 ;
  assign n11107 = ( ~n587 & n11095 ) | ( ~n587 & n11106 ) | ( n11095 & n11106 ) ;
  assign n11108 = n388 | n762 ;
  assign n11109 = n807 | n11108 ;
  assign n11110 = n104 | n349 ;
  assign n11111 = n413 | n11110 ;
  assign n11112 = n11109 | n11111 ;
  assign n11113 = x2 | n110 ;
  assign n11114 = n11112 | n11113 ;
  assign n11115 = n587 | n11114 ;
  assign n11116 = n11107 | n11115 ;
  assign n11117 = x2 & n110 ;
  assign n11118 = ( x2 & n11112 ) | ( x2 & n11117 ) | ( n11112 & n11117 ) ;
  assign n11119 = ( x2 & n587 ) | ( x2 & n11118 ) | ( n587 & n11118 ) ;
  assign n11120 = x2 | n11118 ;
  assign n11121 = ( n11107 & n11119 ) | ( n11107 & n11120 ) | ( n11119 & n11120 ) ;
  assign n11122 = n11116 & ~n11121 ;
  assign n11123 = n10402 & n11122 ;
  assign n11124 = n10391 & n11122 ;
  assign n11125 = ( n10395 & n11122 ) | ( n10395 & n11124 ) | ( n11122 & n11124 ) ;
  assign n11126 = ( n1814 & n11123 ) | ( n1814 & n11125 ) | ( n11123 & n11125 ) ;
  assign n11127 = n11075 & ~n11126 ;
  assign n11128 = n11121 | n11123 ;
  assign n11129 = n11116 & ~n11128 ;
  assign n11130 = n11121 | n11125 ;
  assign n11131 = n11116 & ~n11130 ;
  assign n11132 = ( ~n1814 & n11129 ) | ( ~n1814 & n11131 ) | ( n11129 & n11131 ) ;
  assign n11133 = n11127 | n11132 ;
  assign n11134 = n1057 & n2279 ;
  assign n11135 = ( n1057 & ~n2269 ) | ( n1057 & n11134 ) | ( ~n2269 & n11134 ) ;
  assign n11136 = n1060 & n1708 ;
  assign n11137 = n1065 & n1634 ;
  assign n11138 = ( n1065 & n1630 ) | ( n1065 & n11137 ) | ( n1630 & n11137 ) ;
  assign n11139 = n1062 | n11138 ;
  assign n11140 = n11136 | n11139 ;
  assign n11141 = n11135 | n11140 ;
  assign n11142 = n11136 | n11138 ;
  assign n11143 = n11135 | n11142 ;
  assign n11144 = ( ~n2343 & n11141 ) | ( ~n2343 & n11143 ) | ( n11141 & n11143 ) ;
  assign n11145 = n11132 & n11144 ;
  assign n11146 = ( n11127 & n11144 ) | ( n11127 & n11145 ) | ( n11144 & n11145 ) ;
  assign n11147 = n11133 & ~n11146 ;
  assign n11148 = ~n11132 & n11144 ;
  assign n11149 = ~n11127 & n11148 ;
  assign n11150 = n11147 | n11149 ;
  assign n11153 = n11150 & n11152 ;
  assign n11154 = n11152 & ~n11153 ;
  assign n11155 = n1826 & n2090 ;
  assign n11156 = ( n1826 & ~n2082 ) | ( n1826 & n11155 ) | ( ~n2082 & n11155 ) ;
  assign n11157 = n1829 & n2691 ;
  assign n11158 = ( n1829 & n2678 ) | ( n1829 & n11157 ) | ( n2678 & n11157 ) ;
  assign n11159 = n1823 & n2199 ;
  assign n11160 = ( n1823 & ~n2185 ) | ( n1823 & n11159 ) | ( ~n2185 & n11159 ) ;
  assign n11161 = n11158 | n11160 ;
  assign n11162 = n11156 | n11161 ;
  assign n11163 = n1821 | n11162 ;
  assign n11164 = ( n2985 & n11162 ) | ( n2985 & n11163 ) | ( n11162 & n11163 ) ;
  assign n11165 = x29 & n11163 ;
  assign n11166 = x29 & n11162 ;
  assign n11167 = ( n2985 & n11165 ) | ( n2985 & n11166 ) | ( n11165 & n11166 ) ;
  assign n11168 = x29 & ~n11165 ;
  assign n11169 = x29 & ~n11166 ;
  assign n11170 = ( ~n2985 & n11168 ) | ( ~n2985 & n11169 ) | ( n11168 & n11169 ) ;
  assign n11171 = ( n11164 & ~n11167 ) | ( n11164 & n11170 ) | ( ~n11167 & n11170 ) ;
  assign n11172 = n11150 & n11171 ;
  assign n11173 = ~n11152 & n11172 ;
  assign n11174 = ( n11154 & n11171 ) | ( n11154 & n11173 ) | ( n11171 & n11173 ) ;
  assign n11175 = n11150 | n11171 ;
  assign n11176 = ( ~n11152 & n11171 ) | ( ~n11152 & n11175 ) | ( n11171 & n11175 ) ;
  assign n11177 = n11154 | n11176 ;
  assign n11178 = ~n11174 & n11177 ;
  assign n11179 = n2308 & n2893 ;
  assign n11180 = ( n2308 & ~n2886 ) | ( n2308 & n11179 ) | ( ~n2886 & n11179 ) ;
  assign n11181 = n2312 & n2701 ;
  assign n11182 = ( n2312 & ~n2784 ) | ( n2312 & n11181 ) | ( ~n2784 & n11181 ) ;
  assign n11183 = n2315 & n3507 ;
  assign n11184 = ( n2315 & n3483 ) | ( n2315 & n11183 ) | ( n3483 & n11183 ) ;
  assign n11185 = n11182 | n11184 ;
  assign n11186 = n11180 | n11185 ;
  assign n11187 = n2306 | n11186 ;
  assign n11188 = ( n3603 & n11186 ) | ( n3603 & n11187 ) | ( n11186 & n11187 ) ;
  assign n11189 = x26 & n11187 ;
  assign n11190 = x26 & n11186 ;
  assign n11191 = ( n3603 & n11189 ) | ( n3603 & n11190 ) | ( n11189 & n11190 ) ;
  assign n11192 = x26 & ~n11189 ;
  assign n11193 = x26 & ~n11190 ;
  assign n11194 = ( ~n3603 & n11192 ) | ( ~n3603 & n11193 ) | ( n11192 & n11193 ) ;
  assign n11195 = ( n11188 & ~n11191 ) | ( n11188 & n11194 ) | ( ~n11191 & n11194 ) ;
  assign n11196 = n11178 & ~n11195 ;
  assign n11197 = n11178 | n11195 ;
  assign n11198 = ( ~n11178 & n11196 ) | ( ~n11178 & n11197 ) | ( n11196 & n11197 ) ;
  assign n11199 = n10432 | n10452 ;
  assign n11200 = ( n10432 & n10435 ) | ( n10432 & n11199 ) | ( n10435 & n11199 ) ;
  assign n11201 = n11198 & n11200 ;
  assign n11202 = n11198 | n11200 ;
  assign n11203 = ~n11201 & n11202 ;
  assign n11204 = n2932 & n4206 ;
  assign n11205 = n2925 & n3386 ;
  assign n11206 = n2928 & n3439 ;
  assign n11207 = ( n2928 & ~n3420 ) | ( n2928 & n11206 ) | ( ~n3420 & n11206 ) ;
  assign n11208 = n11205 | n11207 ;
  assign n11209 = n11204 | n11208 ;
  assign n11210 = n2936 | n11204 ;
  assign n11211 = n11208 | n11210 ;
  assign n11212 = ( ~n4220 & n11209 ) | ( ~n4220 & n11211 ) | ( n11209 & n11211 ) ;
  assign n11213 = ~x23 & n11211 ;
  assign n11214 = ~x23 & n11209 ;
  assign n11215 = ( ~n4220 & n11213 ) | ( ~n4220 & n11214 ) | ( n11213 & n11214 ) ;
  assign n11216 = x23 | n11214 ;
  assign n11217 = x23 | n11213 ;
  assign n11218 = ( ~n4220 & n11216 ) | ( ~n4220 & n11217 ) | ( n11216 & n11217 ) ;
  assign n11219 = ( ~n11212 & n11215 ) | ( ~n11212 & n11218 ) | ( n11215 & n11218 ) ;
  assign n11220 = n11203 & ~n11219 ;
  assign n11221 = n11203 | n11219 ;
  assign n11222 = ( ~n11203 & n11220 ) | ( ~n11203 & n11221 ) | ( n11220 & n11221 ) ;
  assign n11223 = n10460 | n10480 ;
  assign n11224 = ( n10460 & n10464 ) | ( n10460 & n11223 ) | ( n10464 & n11223 ) ;
  assign n11225 = n11222 & n11224 ;
  assign n11226 = n11222 | n11224 ;
  assign n11227 = ~n11225 & n11226 ;
  assign n11228 = n3544 & ~n4429 ;
  assign n11229 = n3541 & n4396 ;
  assign n11230 = n11228 | n11229 ;
  assign n11231 = n3547 & n4245 ;
  assign n11232 = ( n3547 & n4303 ) | ( n3547 & n11231 ) | ( n4303 & n11231 ) ;
  assign n11233 = n11230 | n11232 ;
  assign n11234 = n3537 | n11232 ;
  assign n11235 = n11230 | n11234 ;
  assign n11236 = ( n4455 & n11233 ) | ( n4455 & n11235 ) | ( n11233 & n11235 ) ;
  assign n11237 = x20 & n11235 ;
  assign n11238 = x20 & n11233 ;
  assign n11239 = ( n4455 & n11237 ) | ( n4455 & n11238 ) | ( n11237 & n11238 ) ;
  assign n11240 = x20 & ~n11238 ;
  assign n11241 = x20 & ~n11237 ;
  assign n11242 = ( ~n4455 & n11240 ) | ( ~n4455 & n11241 ) | ( n11240 & n11241 ) ;
  assign n11243 = ( n11236 & ~n11239 ) | ( n11236 & n11242 ) | ( ~n11239 & n11242 ) ;
  assign n11244 = n11227 & ~n11243 ;
  assign n11245 = n11227 | n11243 ;
  assign n11246 = ( ~n11227 & n11244 ) | ( ~n11227 & n11245 ) | ( n11244 & n11245 ) ;
  assign n11247 = n10486 | n10504 ;
  assign n11248 = ( n10486 & n10488 ) | ( n10486 & n11247 ) | ( n10488 & n11247 ) ;
  assign n11249 = n11246 & n11248 ;
  assign n11250 = n11246 | n11248 ;
  assign n11251 = ~n11249 & n11250 ;
  assign n11252 = n4468 & n5117 ;
  assign n11253 = ( n4468 & ~n5037 ) | ( n4468 & n11252 ) | ( ~n5037 & n11252 ) ;
  assign n11254 = n4471 & n5108 ;
  assign n11255 = n4466 & n5192 ;
  assign n11256 = ( n4466 & n5179 ) | ( n4466 & n11255 ) | ( n5179 & n11255 ) ;
  assign n11257 = n11254 | n11256 ;
  assign n11258 = n11253 | n11257 ;
  assign n11259 = n4475 | n11258 ;
  assign n11260 = ( ~n5220 & n11258 ) | ( ~n5220 & n11259 ) | ( n11258 & n11259 ) ;
  assign n11261 = ~x17 & n11259 ;
  assign n11262 = ~x17 & n11258 ;
  assign n11263 = ( ~n5220 & n11261 ) | ( ~n5220 & n11262 ) | ( n11261 & n11262 ) ;
  assign n11264 = x17 | n11261 ;
  assign n11265 = x17 | n11262 ;
  assign n11266 = ( ~n5220 & n11264 ) | ( ~n5220 & n11265 ) | ( n11264 & n11265 ) ;
  assign n11267 = ( ~n11260 & n11263 ) | ( ~n11260 & n11266 ) | ( n11263 & n11266 ) ;
  assign n11268 = n11251 & ~n11267 ;
  assign n11269 = n11251 | n11267 ;
  assign n11270 = ( ~n11251 & n11268 ) | ( ~n11251 & n11269 ) | ( n11268 & n11269 ) ;
  assign n11271 = n10510 | n10530 ;
  assign n11272 = ( n10510 & n10512 ) | ( n10510 & n11271 ) | ( n10512 & n11271 ) ;
  assign n11273 = n11270 & n11272 ;
  assign n11274 = n11270 | n11272 ;
  assign n11275 = ~n11273 & n11274 ;
  assign n11276 = n5231 & n5857 ;
  assign n11277 = ( n5231 & ~n5899 ) | ( n5231 & n11276 ) | ( ~n5899 & n11276 ) ;
  assign n11278 = n5234 & ~n6091 ;
  assign n11279 = n5237 & n5997 ;
  assign n11280 = ( n5237 & n5979 ) | ( n5237 & n11279 ) | ( n5979 & n11279 ) ;
  assign n11281 = n11278 | n11280 ;
  assign n11282 = n11277 | n11281 ;
  assign n11283 = n5227 | n11282 ;
  assign n11284 = ( n6108 & n11282 ) | ( n6108 & n11283 ) | ( n11282 & n11283 ) ;
  assign n11285 = x14 & n11283 ;
  assign n11286 = x14 & n11282 ;
  assign n11287 = ( n6108 & n11285 ) | ( n6108 & n11286 ) | ( n11285 & n11286 ) ;
  assign n11288 = x14 & ~n11285 ;
  assign n11289 = x14 & ~n11286 ;
  assign n11290 = ( ~n6108 & n11288 ) | ( ~n6108 & n11289 ) | ( n11288 & n11289 ) ;
  assign n11291 = ( n11284 & ~n11287 ) | ( n11284 & n11290 ) | ( ~n11287 & n11290 ) ;
  assign n11292 = n11275 & ~n11291 ;
  assign n11293 = n11275 | n11291 ;
  assign n11294 = ( ~n11275 & n11292 ) | ( ~n11275 & n11293 ) | ( n11292 & n11293 ) ;
  assign n11295 = n10536 | n10554 ;
  assign n11296 = ( n10536 & n10538 ) | ( n10536 & n11295 ) | ( n10538 & n11295 ) ;
  assign n11297 = n11294 & n11296 ;
  assign n11298 = n11294 | n11296 ;
  assign n11299 = ~n11297 & n11298 ;
  assign n11300 = n6119 & n6950 ;
  assign n11301 = n6125 & n7036 ;
  assign n11302 = ( n6125 & n7023 ) | ( n6125 & n11301 ) | ( n7023 & n11301 ) ;
  assign n11303 = n11300 | n11302 ;
  assign n11304 = n6122 & n6889 ;
  assign n11305 = ( n6122 & ~n6884 ) | ( n6122 & n11304 ) | ( ~n6884 & n11304 ) ;
  assign n11306 = n11303 | n11305 ;
  assign n11307 = n6115 | n11305 ;
  assign n11308 = n11303 | n11307 ;
  assign n11309 = ( ~n7061 & n11306 ) | ( ~n7061 & n11308 ) | ( n11306 & n11308 ) ;
  assign n11310 = ~x11 & n11308 ;
  assign n11311 = ~x11 & n11306 ;
  assign n11312 = ( ~n7061 & n11310 ) | ( ~n7061 & n11311 ) | ( n11310 & n11311 ) ;
  assign n11313 = x11 | n11311 ;
  assign n11314 = x11 | n11310 ;
  assign n11315 = ( ~n7061 & n11313 ) | ( ~n7061 & n11314 ) | ( n11313 & n11314 ) ;
  assign n11316 = ( ~n11309 & n11312 ) | ( ~n11309 & n11315 ) | ( n11312 & n11315 ) ;
  assign n11317 = n11299 & ~n11316 ;
  assign n11318 = n11299 | n11316 ;
  assign n11319 = ( ~n11299 & n11317 ) | ( ~n11299 & n11318 ) | ( n11317 & n11318 ) ;
  assign n11320 = n10559 | n10577 ;
  assign n11321 = ( n10559 & n10562 ) | ( n10559 & n11320 ) | ( n10562 & n11320 ) ;
  assign n11322 = n11319 & n11321 ;
  assign n11323 = n11319 | n11321 ;
  assign n11324 = ~n11322 & n11323 ;
  assign n11325 = n7074 & n7907 ;
  assign n11326 = ( n7074 & n7902 ) | ( n7074 & n11325 ) | ( n7902 & n11325 ) ;
  assign n11327 = n7068 & n8079 ;
  assign n11328 = ( n7068 & ~n8070 ) | ( n7068 & n11327 ) | ( ~n8070 & n11327 ) ;
  assign n11329 = n11326 | n11328 ;
  assign n11330 = n7079 & ~n8017 ;
  assign n11331 = n11329 | n11330 ;
  assign n11332 = n7078 | n11329 ;
  assign n11333 = n11330 | n11332 ;
  assign n11334 = ( n8104 & n11331 ) | ( n8104 & n11333 ) | ( n11331 & n11333 ) ;
  assign n11335 = x8 & n11333 ;
  assign n11336 = x8 & n11331 ;
  assign n11337 = ( n8104 & n11335 ) | ( n8104 & n11336 ) | ( n11335 & n11336 ) ;
  assign n11338 = x8 & ~n11336 ;
  assign n11339 = x8 & ~n11335 ;
  assign n11340 = ( ~n8104 & n11338 ) | ( ~n8104 & n11339 ) | ( n11338 & n11339 ) ;
  assign n11341 = ( n11334 & ~n11337 ) | ( n11334 & n11340 ) | ( ~n11337 & n11340 ) ;
  assign n11342 = n11324 & ~n11341 ;
  assign n11343 = n11324 | n11341 ;
  assign n11344 = ( ~n11324 & n11342 ) | ( ~n11324 & n11343 ) | ( n11342 & n11343 ) ;
  assign n11345 = n11074 & n11344 ;
  assign n11346 = n11074 | n11344 ;
  assign n11347 = ~n11345 & n11346 ;
  assign n11348 = n10609 | n10629 ;
  assign n11349 = n11347 & n11348 ;
  assign n11350 = n10609 & n11347 ;
  assign n11351 = ( n10612 & n11349 ) | ( n10612 & n11350 ) | ( n11349 & n11350 ) ;
  assign n11352 = n11347 | n11348 ;
  assign n11353 = n10609 | n11347 ;
  assign n11354 = ( n10612 & n11352 ) | ( n10612 & n11353 ) | ( n11352 & n11353 ) ;
  assign n11355 = ~n11351 & n11354 ;
  assign n11356 = n10637 | n10641 ;
  assign n11357 = n10637 | n10640 ;
  assign n11358 = ( n9467 & n11356 ) | ( n9467 & n11357 ) | ( n11356 & n11357 ) ;
  assign n11359 = ( n9087 & n11356 ) | ( n9087 & n11357 ) | ( n11356 & n11357 ) ;
  assign n11360 = ( n10322 & n11358 ) | ( n10322 & n11359 ) | ( n11358 & n11359 ) ;
  assign n11361 = n11355 & n11360 ;
  assign n11362 = n11355 | n11360 ;
  assign n11363 = ~n11361 & n11362 ;
  assign n11364 = n8115 & ~n8982 ;
  assign n11365 = ( n8115 & n9051 ) | ( n8115 & n11364 ) | ( n9051 & n11364 ) ;
  assign n11366 = n8125 | n11365 ;
  assign n11367 = n9442 & ~n11365 ;
  assign n11368 = n9074 & ~n11365 ;
  assign n11369 = ( ~n9440 & n11367 ) | ( ~n9440 & n11368 ) | ( n11367 & n11368 ) ;
  assign n11370 = n11366 & ~n11369 ;
  assign n11371 = n11365 & n11366 ;
  assign n11372 = ( ~n9442 & n11366 ) | ( ~n9442 & n11371 ) | ( n11366 & n11371 ) ;
  assign n11373 = ( ~n9072 & n11370 ) | ( ~n9072 & n11372 ) | ( n11370 & n11372 ) ;
  assign n11374 = ~x5 & n11370 ;
  assign n11375 = ~x5 & n11372 ;
  assign n11376 = ( ~n9072 & n11374 ) | ( ~n9072 & n11375 ) | ( n11374 & n11375 ) ;
  assign n11377 = x5 | n11374 ;
  assign n11378 = x5 | n11375 ;
  assign n11379 = ( ~n9072 & n11377 ) | ( ~n9072 & n11378 ) | ( n11377 & n11378 ) ;
  assign n11380 = ( ~n11373 & n11376 ) | ( ~n11373 & n11379 ) | ( n11376 & n11379 ) ;
  assign n11381 = n11322 | n11341 ;
  assign n11382 = ( n11322 & n11324 ) | ( n11322 & n11381 ) | ( n11324 & n11381 ) ;
  assign n11383 = n11380 & n11382 ;
  assign n11384 = n11380 | n11382 ;
  assign n11385 = ~n11383 & n11384 ;
  assign n11386 = ( n1814 & n11128 ) | ( n1814 & n11130 ) | ( n11128 & n11130 ) ;
  assign n11387 = x2 & n568 ;
  assign n11388 = n511 | n644 ;
  assign n11389 = n283 | n581 ;
  assign n11390 = n414 | n11389 ;
  assign n11391 = n11388 | n11390 ;
  assign n11392 = n4020 | n11391 ;
  assign n11393 = n4364 | n11392 ;
  assign n11394 = n6905 | n11393 ;
  assign n11395 = n2241 | n11394 ;
  assign n11396 = n834 | n960 ;
  assign n11397 = n168 | n777 ;
  assign n11398 = n11396 | n11397 ;
  assign n11399 = n278 | n758 ;
  assign n11400 = n2794 | n11399 ;
  assign n11401 = n11398 | n11400 ;
  assign n11402 = n149 & ~n11401 ;
  assign n11403 = n258 | n1172 ;
  assign n11404 = n481 | n11403 ;
  assign n11405 = n450 | n560 ;
  assign n11406 = n240 | n11405 ;
  assign n11407 = n11404 | n11406 ;
  assign n11408 = n2666 | n10379 ;
  assign n11409 = n11407 | n11408 ;
  assign n11410 = n192 | n1662 ;
  assign n11411 = n212 | n11410 ;
  assign n11412 = n887 | n11411 ;
  assign n11413 = n11409 | n11412 ;
  assign n11414 = n11402 & ~n11413 ;
  assign n11415 = ~n11395 & n11414 ;
  assign n11416 = ( x2 & n11387 ) | ( x2 & ~n11415 ) | ( n11387 & ~n11415 ) ;
  assign n11417 = x2 | n568 ;
  assign n11418 = n11415 & ~n11417 ;
  assign n11419 = n11416 | n11418 ;
  assign n11420 = n11121 & ~n11419 ;
  assign n11421 = ( n11125 & ~n11419 ) | ( n11125 & n11420 ) | ( ~n11419 & n11420 ) ;
  assign n11422 = ( n11123 & ~n11419 ) | ( n11123 & n11420 ) | ( ~n11419 & n11420 ) ;
  assign n11423 = ( n1814 & n11421 ) | ( n1814 & n11422 ) | ( n11421 & n11422 ) ;
  assign n11424 = n11386 & ~n11423 ;
  assign n11425 = n1065 & n2279 ;
  assign n11426 = ( n1065 & ~n2269 ) | ( n1065 & n11425 ) | ( ~n2269 & n11425 ) ;
  assign n11427 = n1060 & n1634 ;
  assign n11428 = ( n1060 & n1630 ) | ( n1060 & n11427 ) | ( n1630 & n11427 ) ;
  assign n11429 = n11426 | n11428 ;
  assign n11430 = n1062 | n11429 ;
  assign n11431 = n1057 & n2090 ;
  assign n11432 = ( n1057 & ~n2082 ) | ( n1057 & n11431 ) | ( ~n2082 & n11431 ) ;
  assign n11433 = n11430 | n11432 ;
  assign n11434 = n11429 | n11432 ;
  assign n11435 = ( n2568 & n11433 ) | ( n2568 & n11434 ) | ( n11433 & n11434 ) ;
  assign n11436 = n11121 | n11416 ;
  assign n11437 = ( n11416 & ~n11419 ) | ( n11416 & n11436 ) | ( ~n11419 & n11436 ) ;
  assign n11438 = n11418 | n11437 ;
  assign n11439 = n11125 | n11438 ;
  assign n11440 = n11123 | n11438 ;
  assign n11441 = ( n1814 & n11439 ) | ( n1814 & n11440 ) | ( n11439 & n11440 ) ;
  assign n11442 = n11435 & ~n11441 ;
  assign n11443 = ( n11424 & n11435 ) | ( n11424 & n11442 ) | ( n11435 & n11442 ) ;
  assign n11444 = ~n11435 & n11441 ;
  assign n11445 = ~n11424 & n11444 ;
  assign n11446 = n11443 | n11445 ;
  assign n11447 = n11146 | n11149 ;
  assign n11448 = n11147 | n11447 ;
  assign n11449 = ~n11446 & n11448 ;
  assign n11450 = n11146 & ~n11446 ;
  assign n11451 = ( n11152 & n11449 ) | ( n11152 & n11450 ) | ( n11449 & n11450 ) ;
  assign n11452 = n11446 & ~n11448 ;
  assign n11453 = ~n11146 & n11446 ;
  assign n11454 = ( ~n11152 & n11452 ) | ( ~n11152 & n11453 ) | ( n11452 & n11453 ) ;
  assign n11455 = n11451 | n11454 ;
  assign n11456 = n1829 & n2701 ;
  assign n11457 = ( n1829 & ~n2784 ) | ( n1829 & n11456 ) | ( ~n2784 & n11456 ) ;
  assign n11458 = n1823 & n2691 ;
  assign n11459 = ( n1823 & n2678 ) | ( n1823 & n11458 ) | ( n2678 & n11458 ) ;
  assign n11460 = n11457 | n11459 ;
  assign n11461 = n1826 & n2199 ;
  assign n11462 = ( n1826 & ~n2185 ) | ( n1826 & n11461 ) | ( ~n2185 & n11461 ) ;
  assign n11463 = n11460 | n11462 ;
  assign n11464 = n1821 | n11462 ;
  assign n11465 = n11460 | n11464 ;
  assign n11466 = ( n2960 & n11463 ) | ( n2960 & n11465 ) | ( n11463 & n11465 ) ;
  assign n11467 = x29 & n11465 ;
  assign n11468 = x29 & n11463 ;
  assign n11469 = ( n2960 & n11467 ) | ( n2960 & n11468 ) | ( n11467 & n11468 ) ;
  assign n11470 = x29 & ~n11468 ;
  assign n11471 = x29 & ~n11467 ;
  assign n11472 = ( ~n2960 & n11470 ) | ( ~n2960 & n11471 ) | ( n11470 & n11471 ) ;
  assign n11473 = ( n11466 & ~n11469 ) | ( n11466 & n11472 ) | ( ~n11469 & n11472 ) ;
  assign n11474 = ~n11455 & n11473 ;
  assign n11475 = n11455 & ~n11473 ;
  assign n11476 = n11474 | n11475 ;
  assign n11477 = n2312 & n2893 ;
  assign n11478 = ( n2312 & ~n2886 ) | ( n2312 & n11477 ) | ( ~n2886 & n11477 ) ;
  assign n11479 = n2308 & n3507 ;
  assign n11480 = ( n2308 & n3483 ) | ( n2308 & n11479 ) | ( n3483 & n11479 ) ;
  assign n11481 = n11478 | n11480 ;
  assign n11482 = n2315 & n3386 ;
  assign n11483 = n11481 | n11482 ;
  assign n11484 = n2306 | n11482 ;
  assign n11485 = n11481 | n11484 ;
  assign n11486 = ( ~n3568 & n11483 ) | ( ~n3568 & n11485 ) | ( n11483 & n11485 ) ;
  assign n11487 = ~x26 & n11485 ;
  assign n11488 = ~x26 & n11483 ;
  assign n11489 = ( ~n3568 & n11487 ) | ( ~n3568 & n11488 ) | ( n11487 & n11488 ) ;
  assign n11490 = x26 | n11488 ;
  assign n11491 = x26 | n11487 ;
  assign n11492 = ( ~n3568 & n11490 ) | ( ~n3568 & n11491 ) | ( n11490 & n11491 ) ;
  assign n11493 = ( ~n11486 & n11489 ) | ( ~n11486 & n11492 ) | ( n11489 & n11492 ) ;
  assign n11494 = ~n11476 & n11493 ;
  assign n11495 = n11476 | n11494 ;
  assign n11497 = n11174 | n11195 ;
  assign n11498 = ( n11174 & n11178 ) | ( n11174 & n11497 ) | ( n11178 & n11497 ) ;
  assign n11496 = n11476 & n11493 ;
  assign n11499 = n11496 & n11498 ;
  assign n11500 = ( ~n11495 & n11498 ) | ( ~n11495 & n11499 ) | ( n11498 & n11499 ) ;
  assign n11501 = n11496 | n11498 ;
  assign n11502 = n11495 & ~n11501 ;
  assign n11503 = n11500 | n11502 ;
  assign n11504 = n2928 & n4206 ;
  assign n11505 = n2932 & ~n4429 ;
  assign n11506 = n2925 & n3439 ;
  assign n11507 = ( n2925 & ~n3420 ) | ( n2925 & n11506 ) | ( ~n3420 & n11506 ) ;
  assign n11508 = n11505 | n11507 ;
  assign n11509 = n11504 | n11508 ;
  assign n11510 = n2936 | n11504 ;
  assign n11511 = n11508 | n11510 ;
  assign n11512 = ( ~n4527 & n11509 ) | ( ~n4527 & n11511 ) | ( n11509 & n11511 ) ;
  assign n11513 = ~x23 & n11511 ;
  assign n11514 = ~x23 & n11509 ;
  assign n11515 = ( ~n4527 & n11513 ) | ( ~n4527 & n11514 ) | ( n11513 & n11514 ) ;
  assign n11516 = x23 | n11514 ;
  assign n11517 = x23 | n11513 ;
  assign n11518 = ( ~n4527 & n11516 ) | ( ~n4527 & n11517 ) | ( n11516 & n11517 ) ;
  assign n11519 = ( ~n11512 & n11515 ) | ( ~n11512 & n11518 ) | ( n11515 & n11518 ) ;
  assign n11520 = ~n11503 & n11519 ;
  assign n11521 = n11503 | n11520 ;
  assign n11523 = n11201 | n11219 ;
  assign n11524 = ( n11201 & n11203 ) | ( n11201 & n11523 ) | ( n11203 & n11523 ) ;
  assign n11522 = n11503 & n11519 ;
  assign n11525 = n11522 & n11524 ;
  assign n11526 = ( ~n11521 & n11524 ) | ( ~n11521 & n11525 ) | ( n11524 & n11525 ) ;
  assign n11527 = n11522 | n11524 ;
  assign n11528 = n11521 & ~n11527 ;
  assign n11529 = n11526 | n11528 ;
  assign n11530 = n3544 & n4396 ;
  assign n11531 = n3541 & n4245 ;
  assign n11532 = ( n3541 & n4303 ) | ( n3541 & n11531 ) | ( n4303 & n11531 ) ;
  assign n11533 = n11530 | n11532 ;
  assign n11534 = n3547 & n5192 ;
  assign n11535 = ( n3547 & n5179 ) | ( n3547 & n11534 ) | ( n5179 & n11534 ) ;
  assign n11536 = n11533 | n11535 ;
  assign n11537 = n3537 | n11535 ;
  assign n11538 = n11533 | n11537 ;
  assign n11539 = ( n5306 & n11536 ) | ( n5306 & n11538 ) | ( n11536 & n11538 ) ;
  assign n11540 = x20 & n11538 ;
  assign n11541 = x20 & n11536 ;
  assign n11542 = ( n5306 & n11540 ) | ( n5306 & n11541 ) | ( n11540 & n11541 ) ;
  assign n11543 = x20 & ~n11541 ;
  assign n11544 = x20 & ~n11540 ;
  assign n11545 = ( ~n5306 & n11543 ) | ( ~n5306 & n11544 ) | ( n11543 & n11544 ) ;
  assign n11546 = ( n11539 & ~n11542 ) | ( n11539 & n11545 ) | ( ~n11542 & n11545 ) ;
  assign n11547 = n11529 | n11546 ;
  assign n11548 = n11529 & ~n11546 ;
  assign n11549 = ( ~n11529 & n11547 ) | ( ~n11529 & n11548 ) | ( n11547 & n11548 ) ;
  assign n11550 = n11225 | n11243 ;
  assign n11551 = ( n11225 & n11227 ) | ( n11225 & n11550 ) | ( n11227 & n11550 ) ;
  assign n11552 = ~n11549 & n11551 ;
  assign n11553 = n11549 & ~n11551 ;
  assign n11554 = n11552 | n11553 ;
  assign n11555 = n4466 & n5117 ;
  assign n11556 = ( n4466 & ~n5037 ) | ( n4466 & n11555 ) | ( ~n5037 & n11555 ) ;
  assign n11557 = n4468 & n5108 ;
  assign n11558 = n4471 & n5997 ;
  assign n11559 = ( n4471 & n5979 ) | ( n4471 & n11558 ) | ( n5979 & n11558 ) ;
  assign n11560 = n11557 | n11559 ;
  assign n11561 = n11556 | n11560 ;
  assign n11562 = n4475 | n11561 ;
  assign n11563 = ( n6181 & n11561 ) | ( n6181 & n11562 ) | ( n11561 & n11562 ) ;
  assign n11564 = x17 & n11562 ;
  assign n11565 = x17 & n11561 ;
  assign n11566 = ( n6181 & n11564 ) | ( n6181 & n11565 ) | ( n11564 & n11565 ) ;
  assign n11567 = x17 & ~n11564 ;
  assign n11568 = x17 & ~n11565 ;
  assign n11569 = ( ~n6181 & n11567 ) | ( ~n6181 & n11568 ) | ( n11567 & n11568 ) ;
  assign n11570 = ( n11563 & ~n11566 ) | ( n11563 & n11569 ) | ( ~n11566 & n11569 ) ;
  assign n11571 = n11554 | n11570 ;
  assign n11572 = n11554 & ~n11570 ;
  assign n11573 = ( ~n11554 & n11571 ) | ( ~n11554 & n11572 ) | ( n11571 & n11572 ) ;
  assign n11574 = n11249 | n11267 ;
  assign n11575 = ( n11249 & n11251 ) | ( n11249 & n11574 ) | ( n11251 & n11574 ) ;
  assign n11576 = ~n11573 & n11575 ;
  assign n11577 = n11573 & ~n11575 ;
  assign n11578 = n11576 | n11577 ;
  assign n11579 = n5237 & n5857 ;
  assign n11580 = ( n5237 & ~n5899 ) | ( n5237 & n11579 ) | ( ~n5899 & n11579 ) ;
  assign n11581 = n5231 & ~n6091 ;
  assign n11582 = n5234 & n7036 ;
  assign n11583 = ( n5234 & n7023 ) | ( n5234 & n11582 ) | ( n7023 & n11582 ) ;
  assign n11584 = n11581 | n11583 ;
  assign n11585 = n11580 | n11584 ;
  assign n11586 = n5227 | n11585 ;
  assign n11587 = ( n7136 & n11585 ) | ( n7136 & n11586 ) | ( n11585 & n11586 ) ;
  assign n11588 = x14 & n11586 ;
  assign n11589 = x14 & n11585 ;
  assign n11590 = ( n7136 & n11588 ) | ( n7136 & n11589 ) | ( n11588 & n11589 ) ;
  assign n11591 = x14 & ~n11588 ;
  assign n11592 = x14 & ~n11589 ;
  assign n11593 = ( ~n7136 & n11591 ) | ( ~n7136 & n11592 ) | ( n11591 & n11592 ) ;
  assign n11594 = ( n11587 & ~n11590 ) | ( n11587 & n11593 ) | ( ~n11590 & n11593 ) ;
  assign n11595 = n11578 | n11594 ;
  assign n11596 = n11578 & ~n11594 ;
  assign n11597 = ( ~n11578 & n11595 ) | ( ~n11578 & n11596 ) | ( n11595 & n11596 ) ;
  assign n11598 = n11273 | n11291 ;
  assign n11599 = ( n11273 & n11275 ) | ( n11273 & n11598 ) | ( n11275 & n11598 ) ;
  assign n11600 = ~n11597 & n11599 ;
  assign n11601 = n11597 & ~n11599 ;
  assign n11602 = n11600 | n11601 ;
  assign n11603 = n6125 & n6950 ;
  assign n11604 = n6119 & n6889 ;
  assign n11605 = ( n6119 & ~n6884 ) | ( n6119 & n11604 ) | ( ~n6884 & n11604 ) ;
  assign n11606 = n11603 | n11605 ;
  assign n11607 = n6122 & n7907 ;
  assign n11608 = ( n6122 & n7902 ) | ( n6122 & n11607 ) | ( n7902 & n11607 ) ;
  assign n11609 = n11606 | n11608 ;
  assign n11610 = n6115 | n11608 ;
  assign n11611 = n11606 | n11610 ;
  assign n11612 = ( ~n8193 & n11609 ) | ( ~n8193 & n11611 ) | ( n11609 & n11611 ) ;
  assign n11613 = ~x11 & n11611 ;
  assign n11614 = ~x11 & n11609 ;
  assign n11615 = ( ~n8193 & n11613 ) | ( ~n8193 & n11614 ) | ( n11613 & n11614 ) ;
  assign n11616 = x11 | n11614 ;
  assign n11617 = x11 | n11613 ;
  assign n11618 = ( ~n8193 & n11616 ) | ( ~n8193 & n11617 ) | ( n11616 & n11617 ) ;
  assign n11619 = ( ~n11612 & n11615 ) | ( ~n11612 & n11618 ) | ( n11615 & n11618 ) ;
  assign n11620 = n11602 | n11619 ;
  assign n11621 = n11602 & ~n11619 ;
  assign n11622 = ( ~n11602 & n11620 ) | ( ~n11602 & n11621 ) | ( n11620 & n11621 ) ;
  assign n11623 = n11297 | n11316 ;
  assign n11624 = ( n11297 & n11299 ) | ( n11297 & n11623 ) | ( n11299 & n11623 ) ;
  assign n11625 = ~n11622 & n11624 ;
  assign n11626 = n11622 & ~n11624 ;
  assign n11627 = n11625 | n11626 ;
  assign n11628 = n7074 & n8079 ;
  assign n11629 = ( n7074 & ~n8070 ) | ( n7074 & n11628 ) | ( ~n8070 & n11628 ) ;
  assign n11630 = n7068 | n11629 ;
  assign n11631 = ( ~n8017 & n11629 ) | ( ~n8017 & n11630 ) | ( n11629 & n11630 ) ;
  assign n11632 = n7079 & n9022 ;
  assign n11633 = ( n7079 & ~n9019 ) | ( n7079 & n11632 ) | ( ~n9019 & n11632 ) ;
  assign n11634 = n11631 | n11633 ;
  assign n11635 = n7078 | n11633 ;
  assign n11636 = n11631 | n11635 ;
  assign n11637 = ( ~n9416 & n11634 ) | ( ~n9416 & n11636 ) | ( n11634 & n11636 ) ;
  assign n11638 = ~x8 & n11636 ;
  assign n11639 = ~x8 & n11634 ;
  assign n11640 = ( ~n9416 & n11638 ) | ( ~n9416 & n11639 ) | ( n11638 & n11639 ) ;
  assign n11641 = x8 | n11639 ;
  assign n11642 = x8 | n11638 ;
  assign n11643 = ( ~n9416 & n11641 ) | ( ~n9416 & n11642 ) | ( n11641 & n11642 ) ;
  assign n11644 = ( ~n11637 & n11640 ) | ( ~n11637 & n11643 ) | ( n11640 & n11643 ) ;
  assign n11645 = n11627 | n11644 ;
  assign n11646 = n11627 & ~n11644 ;
  assign n11647 = ( ~n11627 & n11645 ) | ( ~n11627 & n11646 ) | ( n11645 & n11646 ) ;
  assign n11648 = n11385 & ~n11647 ;
  assign n11649 = n11385 | n11647 ;
  assign n11650 = ( ~n11385 & n11648 ) | ( ~n11385 & n11649 ) | ( n11648 & n11649 ) ;
  assign n11651 = n11071 | n11344 ;
  assign n11652 = ( n11071 & n11074 ) | ( n11071 & n11651 ) | ( n11074 & n11651 ) ;
  assign n11653 = ~n11650 & n11652 ;
  assign n11654 = n11650 & ~n11652 ;
  assign n11655 = n11653 | n11654 ;
  assign n11656 = n11351 & ~n11655 ;
  assign n11657 = ( n11355 & ~n11655 ) | ( n11355 & n11656 ) | ( ~n11655 & n11656 ) ;
  assign n11658 = ~n11655 & n11656 ;
  assign n11659 = ( n11360 & n11657 ) | ( n11360 & n11658 ) | ( n11657 & n11658 ) ;
  assign n11660 = ~n11351 & n11655 ;
  assign n11661 = ~n11355 & n11660 ;
  assign n11662 = ( ~n11360 & n11660 ) | ( ~n11360 & n11661 ) | ( n11660 & n11661 ) ;
  assign n11663 = n11659 | n11662 ;
  assign n11664 = n11363 & ~n11663 ;
  assign n11665 = ~n11363 & n11663 ;
  assign n11666 = n10649 & n11363 ;
  assign n11667 = n10649 | n11363 ;
  assign n11668 = ~n11666 & n11667 ;
  assign n11669 = n11666 | n11668 ;
  assign n11670 = ~n11665 & n11669 ;
  assign n11671 = ~n11665 & n11666 ;
  assign n11672 = ( n10694 & n11670 ) | ( n10694 & n11671 ) | ( n11670 & n11671 ) ;
  assign n11673 = n11664 | n11672 ;
  assign n11691 = n11625 | n11644 ;
  assign n11692 = ( n11625 & ~n11627 ) | ( n11625 & n11691 ) | ( ~n11627 & n11691 ) ;
  assign n11674 = n7079 & ~n8982 ;
  assign n11675 = ( n7079 & n9051 ) | ( n7079 & n11674 ) | ( n9051 & n11674 ) ;
  assign n11676 = n7068 & n9022 ;
  assign n11677 = n11675 | n11676 ;
  assign n11678 = n7068 | n11675 ;
  assign n11679 = ( ~n9019 & n11677 ) | ( ~n9019 & n11678 ) | ( n11677 & n11678 ) ;
  assign n11680 = n7074 | n11679 ;
  assign n11681 = ( ~n8017 & n11679 ) | ( ~n8017 & n11680 ) | ( n11679 & n11680 ) ;
  assign n11682 = n7078 | n11681 ;
  assign n11683 = ( ~n10242 & n11681 ) | ( ~n10242 & n11682 ) | ( n11681 & n11682 ) ;
  assign n11684 = ~x8 & n11682 ;
  assign n11685 = ~x8 & n11681 ;
  assign n11686 = ( ~n10242 & n11684 ) | ( ~n10242 & n11685 ) | ( n11684 & n11685 ) ;
  assign n11687 = x8 | n11684 ;
  assign n11688 = x8 | n11685 ;
  assign n11689 = ( ~n10242 & n11687 ) | ( ~n10242 & n11688 ) | ( n11687 & n11688 ) ;
  assign n11690 = ( ~n11683 & n11686 ) | ( ~n11683 & n11689 ) | ( n11686 & n11689 ) ;
  assign n11693 = n11690 & n11692 ;
  assign n11694 = n11692 & ~n11693 ;
  assign n11695 = n6125 & n6889 ;
  assign n11696 = ( n6125 & ~n6884 ) | ( n6125 & n11695 ) | ( ~n6884 & n11695 ) ;
  assign n11697 = n6119 & n7907 ;
  assign n11698 = ( n6119 & n7902 ) | ( n6119 & n11697 ) | ( n7902 & n11697 ) ;
  assign n11699 = n6122 & n8079 ;
  assign n11700 = ( n6122 & ~n8070 ) | ( n6122 & n11699 ) | ( ~n8070 & n11699 ) ;
  assign n11701 = n11698 | n11700 ;
  assign n11702 = n11696 | n11701 ;
  assign n11703 = n6115 | n11702 ;
  assign n11704 = n11702 & n11703 ;
  assign n11705 = ( ~n8156 & n11703 ) | ( ~n8156 & n11704 ) | ( n11703 & n11704 ) ;
  assign n11706 = ~x11 & n11704 ;
  assign n11707 = ~x11 & n11703 ;
  assign n11708 = ( ~n8156 & n11706 ) | ( ~n8156 & n11707 ) | ( n11706 & n11707 ) ;
  assign n11709 = x11 | n11706 ;
  assign n11710 = x11 | n11707 ;
  assign n11711 = ( ~n8156 & n11709 ) | ( ~n8156 & n11710 ) | ( n11709 & n11710 ) ;
  assign n11712 = ( ~n11705 & n11708 ) | ( ~n11705 & n11711 ) | ( n11708 & n11711 ) ;
  assign n11713 = n11600 | n11619 ;
  assign n11714 = ( n11600 & ~n11602 ) | ( n11600 & n11713 ) | ( ~n11602 & n11713 ) ;
  assign n11715 = n11712 & n11714 ;
  assign n11716 = n11712 | n11714 ;
  assign n11717 = ~n11715 & n11716 ;
  assign n11718 = n374 | n489 ;
  assign n11719 = n307 | n11718 ;
  assign n11720 = n3312 | n4180 ;
  assign n11721 = ( ~n9107 & n11719 ) | ( ~n9107 & n11720 ) | ( n11719 & n11720 ) ;
  assign n11722 = n11719 & n11720 ;
  assign n11723 = ( ~n9105 & n11721 ) | ( ~n9105 & n11722 ) | ( n11721 & n11722 ) ;
  assign n11724 = n9108 | n11723 ;
  assign n11725 = n126 | n280 ;
  assign n11726 = n500 | n11725 ;
  assign n11727 = n209 | n588 ;
  assign n11728 = n1678 | n11727 ;
  assign n11729 = n262 | n1039 ;
  assign n11730 = n226 | n11729 ;
  assign n11731 = n11728 | n11730 ;
  assign n11732 = n6878 | n11731 ;
  assign n11733 = n11726 | n11732 ;
  assign n11734 = n11724 | n11733 ;
  assign n11735 = n170 | n175 ;
  assign n11736 = n820 | n11735 ;
  assign n11737 = n9113 | n11736 ;
  assign n11738 = n263 | n303 ;
  assign n11739 = n333 | n11738 ;
  assign n11740 = n112 | n581 ;
  assign n11741 = n355 | n735 ;
  assign n11742 = n11740 | n11741 ;
  assign n11743 = n11739 | n11742 ;
  assign n11744 = n11737 | n11743 ;
  assign n11745 = n461 | n901 ;
  assign n11746 = n594 | n11745 ;
  assign n11747 = n39 | n312 ;
  assign n11748 = n229 | n289 ;
  assign n11749 = n11747 | n11748 ;
  assign n11750 = n11746 | n11749 ;
  assign n11751 = n967 | n1494 ;
  assign n11752 = n11750 | n11751 ;
  assign n11753 = n11744 | n11752 ;
  assign n11754 = n1171 | n1404 ;
  assign n11755 = n258 | n992 ;
  assign n11756 = n11754 | n11755 ;
  assign n11757 = n83 | n249 ;
  assign n11758 = n11756 | n11757 ;
  assign n11759 = n110 | n168 ;
  assign n11760 = n390 | n11759 ;
  assign n11761 = n383 | n491 ;
  assign n11762 = n277 | n431 ;
  assign n11763 = n11761 | n11762 ;
  assign n11764 = n11760 | n11763 ;
  assign n11765 = n6038 | n11764 ;
  assign n11766 = n11758 | n11765 ;
  assign n11767 = n11753 | n11766 ;
  assign n11768 = n11734 | n11767 ;
  assign n11769 = n1116 | n7011 ;
  assign n11770 = n114 | n208 ;
  assign n11771 = n99 | n11770 ;
  assign n11772 = n11769 | n11771 ;
  assign n11773 = n469 | n517 ;
  assign n11774 = n5091 | n11773 ;
  assign n11775 = n11772 | n11774 ;
  assign n11776 = n617 | n11775 ;
  assign n11777 = n987 | n6063 ;
  assign n11778 = n11776 | n11777 ;
  assign n11779 = n412 | n11778 ;
  assign n11780 = n178 | n458 ;
  assign n11781 = n160 | n190 ;
  assign n11782 = n11780 | n11781 ;
  assign n11783 = n513 | n762 ;
  assign n11784 = n568 | n11783 ;
  assign n11785 = n11782 | n11784 ;
  assign n11786 = x2 & n182 ;
  assign n11787 = ( x2 & n11785 ) | ( x2 & n11786 ) | ( n11785 & n11786 ) ;
  assign n11788 = ( x2 & n11779 ) | ( x2 & n11787 ) | ( n11779 & n11787 ) ;
  assign n11789 = x2 | n11787 ;
  assign n11790 = ( n11768 & n11788 ) | ( n11768 & n11789 ) | ( n11788 & n11789 ) ;
  assign n11791 = x2 | n182 ;
  assign n11792 = n11785 | n11791 ;
  assign n11793 = n11779 | n11792 ;
  assign n11794 = n11768 | n11793 ;
  assign n11795 = ~n11790 & n11794 ;
  assign n11796 = x5 | n11795 ;
  assign n11797 = x5 & n11795 ;
  assign n11798 = n11796 & ~n11797 ;
  assign n11799 = ~n11416 & n11419 ;
  assign n11800 = ( n11123 & n11437 ) | ( n11123 & ~n11799 ) | ( n11437 & ~n11799 ) ;
  assign n11801 = n11798 & n11800 ;
  assign n11802 = ( n11125 & n11437 ) | ( n11125 & ~n11799 ) | ( n11437 & ~n11799 ) ;
  assign n11803 = n11798 & n11802 ;
  assign n11804 = ( n1814 & n11801 ) | ( n1814 & n11803 ) | ( n11801 & n11803 ) ;
  assign n11805 = n11798 | n11800 ;
  assign n11806 = n11798 | n11802 ;
  assign n11807 = ( n1814 & n11805 ) | ( n1814 & n11806 ) | ( n11805 & n11806 ) ;
  assign n11808 = ~n11804 & n11807 ;
  assign n11809 = n1065 & n2090 ;
  assign n11810 = ( n1065 & ~n2082 ) | ( n1065 & n11809 ) | ( ~n2082 & n11809 ) ;
  assign n11811 = n1060 & n2279 ;
  assign n11812 = ( n1060 & ~n2269 ) | ( n1060 & n11811 ) | ( ~n2269 & n11811 ) ;
  assign n11813 = n1057 & n2199 ;
  assign n11814 = ( n1057 & ~n2185 ) | ( n1057 & n11813 ) | ( ~n2185 & n11813 ) ;
  assign n11815 = n11812 | n11814 ;
  assign n11816 = n11810 | n11815 ;
  assign n11817 = n1062 | n11816 ;
  assign n11818 = ( ~n2325 & n11816 ) | ( ~n2325 & n11817 ) | ( n11816 & n11817 ) ;
  assign n11819 = n11816 & n11817 ;
  assign n11820 = ( ~n2299 & n11818 ) | ( ~n2299 & n11819 ) | ( n11818 & n11819 ) ;
  assign n11821 = ~n11808 & n11820 ;
  assign n11822 = n11808 & ~n11820 ;
  assign n11823 = n11821 | n11822 ;
  assign n11824 = n11443 & n11823 ;
  assign n11825 = ( n11449 & n11823 ) | ( n11449 & n11824 ) | ( n11823 & n11824 ) ;
  assign n11826 = ( n11450 & n11823 ) | ( n11450 & n11824 ) | ( n11823 & n11824 ) ;
  assign n11827 = ( n11152 & n11825 ) | ( n11152 & n11826 ) | ( n11825 & n11826 ) ;
  assign n11828 = n11443 | n11823 ;
  assign n11829 = n11449 | n11828 ;
  assign n11830 = n11450 | n11828 ;
  assign n11831 = ( n11152 & n11829 ) | ( n11152 & n11830 ) | ( n11829 & n11830 ) ;
  assign n11832 = ~n11827 & n11831 ;
  assign n11833 = n1826 & n2691 ;
  assign n11834 = ( n1826 & n2678 ) | ( n1826 & n11833 ) | ( n2678 & n11833 ) ;
  assign n11835 = n1823 & n2701 ;
  assign n11836 = ( n1823 & ~n2784 ) | ( n1823 & n11835 ) | ( ~n2784 & n11835 ) ;
  assign n11837 = n11834 | n11836 ;
  assign n11838 = n1829 & n2893 ;
  assign n11839 = ( n1829 & ~n2886 ) | ( n1829 & n11838 ) | ( ~n2886 & n11838 ) ;
  assign n11840 = n11837 | n11839 ;
  assign n11841 = n1821 | n11840 ;
  assign n11842 = ( ~n2914 & n11840 ) | ( ~n2914 & n11841 ) | ( n11840 & n11841 ) ;
  assign n11843 = ~x29 & n11841 ;
  assign n11844 = ~x29 & n11840 ;
  assign n11845 = ( ~n2914 & n11843 ) | ( ~n2914 & n11844 ) | ( n11843 & n11844 ) ;
  assign n11846 = x29 | n11843 ;
  assign n11847 = x29 | n11844 ;
  assign n11848 = ( ~n2914 & n11846 ) | ( ~n2914 & n11847 ) | ( n11846 & n11847 ) ;
  assign n11849 = ( ~n11842 & n11845 ) | ( ~n11842 & n11848 ) | ( n11845 & n11848 ) ;
  assign n11850 = n11832 & n11849 ;
  assign n11851 = n11832 & ~n11850 ;
  assign n11852 = n2308 & n3386 ;
  assign n11853 = n2312 & n3507 ;
  assign n11854 = ( n2312 & n3483 ) | ( n2312 & n11853 ) | ( n3483 & n11853 ) ;
  assign n11855 = n2315 & n3439 ;
  assign n11856 = ( n2315 & ~n3420 ) | ( n2315 & n11855 ) | ( ~n3420 & n11855 ) ;
  assign n11857 = n11854 | n11856 ;
  assign n11858 = n11852 | n11857 ;
  assign n11859 = n2306 | n11858 ;
  assign n11860 = n11858 & n11859 ;
  assign n11861 = ( ~n3530 & n11859 ) | ( ~n3530 & n11860 ) | ( n11859 & n11860 ) ;
  assign n11862 = ~x26 & n11860 ;
  assign n11863 = ~x26 & n11859 ;
  assign n11864 = ( ~n3530 & n11862 ) | ( ~n3530 & n11863 ) | ( n11862 & n11863 ) ;
  assign n11865 = x26 | n11862 ;
  assign n11866 = x26 | n11863 ;
  assign n11867 = ( ~n3530 & n11865 ) | ( ~n3530 & n11866 ) | ( n11865 & n11866 ) ;
  assign n11868 = ( ~n11861 & n11864 ) | ( ~n11861 & n11867 ) | ( n11864 & n11867 ) ;
  assign n11869 = n11849 & n11868 ;
  assign n11870 = ~n11832 & n11869 ;
  assign n11871 = ( n11851 & n11868 ) | ( n11851 & n11870 ) | ( n11868 & n11870 ) ;
  assign n11872 = n11849 | n11868 ;
  assign n11873 = ( ~n11832 & n11868 ) | ( ~n11832 & n11872 ) | ( n11868 & n11872 ) ;
  assign n11874 = n11851 | n11873 ;
  assign n11875 = ~n11871 & n11874 ;
  assign n11876 = n11474 | n11493 ;
  assign n11877 = ( n11474 & ~n11476 ) | ( n11474 & n11876 ) | ( ~n11476 & n11876 ) ;
  assign n11878 = n11875 & n11877 ;
  assign n11879 = n11875 | n11877 ;
  assign n11880 = ~n11878 & n11879 ;
  assign n11881 = n2928 & ~n4429 ;
  assign n11882 = n2925 | n2928 ;
  assign n11883 = ( n2925 & ~n4429 ) | ( n2925 & n11882 ) | ( ~n4429 & n11882 ) ;
  assign n11884 = ( n4206 & n11881 ) | ( n4206 & n11883 ) | ( n11881 & n11883 ) ;
  assign n11885 = n2932 & n4396 ;
  assign n11886 = n11884 | n11885 ;
  assign n11887 = n2936 | n11885 ;
  assign n11888 = n11884 | n11887 ;
  assign n11889 = ( ~n4501 & n11886 ) | ( ~n4501 & n11888 ) | ( n11886 & n11888 ) ;
  assign n11890 = ~x23 & n11888 ;
  assign n11891 = ~x23 & n11886 ;
  assign n11892 = ( ~n4501 & n11890 ) | ( ~n4501 & n11891 ) | ( n11890 & n11891 ) ;
  assign n11893 = x23 | n11891 ;
  assign n11894 = x23 | n11890 ;
  assign n11895 = ( ~n4501 & n11893 ) | ( ~n4501 & n11894 ) | ( n11893 & n11894 ) ;
  assign n11896 = ( ~n11889 & n11892 ) | ( ~n11889 & n11895 ) | ( n11892 & n11895 ) ;
  assign n11897 = n11880 & n11896 ;
  assign n11898 = n11880 & ~n11897 ;
  assign n11900 = n11500 | n11519 ;
  assign n11901 = ( n11500 & ~n11503 ) | ( n11500 & n11900 ) | ( ~n11503 & n11900 ) ;
  assign n11899 = ~n11880 & n11896 ;
  assign n11902 = n11899 & n11901 ;
  assign n11903 = ( n11898 & n11901 ) | ( n11898 & n11902 ) | ( n11901 & n11902 ) ;
  assign n11904 = n11899 | n11901 ;
  assign n11905 = n11898 | n11904 ;
  assign n11906 = ~n11903 & n11905 ;
  assign n11907 = n3544 & n4245 ;
  assign n11908 = ( n3544 & n4303 ) | ( n3544 & n11907 ) | ( n4303 & n11907 ) ;
  assign n11909 = n3541 & n5192 ;
  assign n11910 = ( n3541 & n5179 ) | ( n3541 & n11909 ) | ( n5179 & n11909 ) ;
  assign n11911 = n11908 | n11910 ;
  assign n11912 = n3547 & n5117 ;
  assign n11913 = ( n3547 & ~n5037 ) | ( n3547 & n11912 ) | ( ~n5037 & n11912 ) ;
  assign n11915 = n3537 | n11913 ;
  assign n11916 = n11911 | n11915 ;
  assign n11914 = n11911 | n11913 ;
  assign n11917 = n11914 & n11916 ;
  assign n11918 = ( ~n5270 & n11916 ) | ( ~n5270 & n11917 ) | ( n11916 & n11917 ) ;
  assign n11919 = ~x20 & n11917 ;
  assign n11920 = ~x20 & n11916 ;
  assign n11921 = ( ~n5270 & n11919 ) | ( ~n5270 & n11920 ) | ( n11919 & n11920 ) ;
  assign n11922 = x20 | n11919 ;
  assign n11923 = x20 | n11920 ;
  assign n11924 = ( ~n5270 & n11922 ) | ( ~n5270 & n11923 ) | ( n11922 & n11923 ) ;
  assign n11925 = ( ~n11918 & n11921 ) | ( ~n11918 & n11924 ) | ( n11921 & n11924 ) ;
  assign n11926 = n11906 & n11925 ;
  assign n11927 = n11906 | n11925 ;
  assign n11928 = ~n11926 & n11927 ;
  assign n11929 = n11526 | n11546 ;
  assign n11930 = ( n11526 & ~n11529 ) | ( n11526 & n11929 ) | ( ~n11529 & n11929 ) ;
  assign n11931 = n11928 & n11930 ;
  assign n11932 = n11928 | n11930 ;
  assign n11933 = ~n11931 & n11932 ;
  assign n11934 = n4466 & n5108 ;
  assign n11935 = n4468 & n5997 ;
  assign n11936 = ( n4468 & n5979 ) | ( n4468 & n11935 ) | ( n5979 & n11935 ) ;
  assign n11937 = n11934 | n11936 ;
  assign n11938 = n4471 & n5857 ;
  assign n11939 = ( n4471 & ~n5899 ) | ( n4471 & n11938 ) | ( ~n5899 & n11938 ) ;
  assign n11940 = n11937 | n11939 ;
  assign n11941 = n4475 | n11940 ;
  assign n11942 = ( ~n6151 & n11940 ) | ( ~n6151 & n11941 ) | ( n11940 & n11941 ) ;
  assign n11943 = ~x17 & n11941 ;
  assign n11944 = ~x17 & n11940 ;
  assign n11945 = ( ~n6151 & n11943 ) | ( ~n6151 & n11944 ) | ( n11943 & n11944 ) ;
  assign n11946 = x17 | n11943 ;
  assign n11947 = x17 | n11944 ;
  assign n11948 = ( ~n6151 & n11946 ) | ( ~n6151 & n11947 ) | ( n11946 & n11947 ) ;
  assign n11949 = ( ~n11942 & n11945 ) | ( ~n11942 & n11948 ) | ( n11945 & n11948 ) ;
  assign n11950 = n11933 & n11949 ;
  assign n11951 = ~n11933 & n11949 ;
  assign n11952 = ( n11933 & ~n11950 ) | ( n11933 & n11951 ) | ( ~n11950 & n11951 ) ;
  assign n11953 = n11552 | n11570 ;
  assign n11954 = ( n11552 & ~n11554 ) | ( n11552 & n11953 ) | ( ~n11554 & n11953 ) ;
  assign n11955 = n11952 & n11954 ;
  assign n11956 = n11952 | n11954 ;
  assign n11957 = ~n11955 & n11956 ;
  assign n11958 = n5237 & ~n6091 ;
  assign n11959 = n5231 & n7036 ;
  assign n11960 = ( n5231 & n7023 ) | ( n5231 & n11959 ) | ( n7023 & n11959 ) ;
  assign n11961 = n11958 | n11960 ;
  assign n11962 = n5234 & n6950 ;
  assign n11963 = n11961 | n11962 ;
  assign n11964 = n5227 | n11963 ;
  assign n11965 = n11963 & n11964 ;
  assign n11966 = ( ~n7107 & n11964 ) | ( ~n7107 & n11965 ) | ( n11964 & n11965 ) ;
  assign n11967 = ~x14 & n11965 ;
  assign n11968 = ~x14 & n11964 ;
  assign n11969 = ( ~n7107 & n11967 ) | ( ~n7107 & n11968 ) | ( n11967 & n11968 ) ;
  assign n11970 = x14 | n11967 ;
  assign n11971 = x14 | n11968 ;
  assign n11972 = ( ~n7107 & n11970 ) | ( ~n7107 & n11971 ) | ( n11970 & n11971 ) ;
  assign n11973 = ( ~n11966 & n11969 ) | ( ~n11966 & n11972 ) | ( n11969 & n11972 ) ;
  assign n11974 = n11957 & n11973 ;
  assign n11975 = n11957 | n11973 ;
  assign n11976 = ~n11974 & n11975 ;
  assign n11977 = n11576 | n11594 ;
  assign n11978 = ( n11576 & ~n11578 ) | ( n11576 & n11977 ) | ( ~n11578 & n11977 ) ;
  assign n11979 = n11976 & n11978 ;
  assign n11980 = n11976 | n11978 ;
  assign n11981 = ~n11979 & n11980 ;
  assign n11982 = n11717 & n11981 ;
  assign n11983 = n11717 | n11981 ;
  assign n11984 = ~n11982 & n11983 ;
  assign n11985 = n11690 & n11984 ;
  assign n11986 = ~n11692 & n11985 ;
  assign n11987 = ( n11694 & n11984 ) | ( n11694 & n11986 ) | ( n11984 & n11986 ) ;
  assign n11988 = n11690 | n11984 ;
  assign n11989 = ( ~n11692 & n11984 ) | ( ~n11692 & n11988 ) | ( n11984 & n11988 ) ;
  assign n11990 = n11694 | n11989 ;
  assign n11991 = ~n11987 & n11990 ;
  assign n11992 = ~n11383 & n11647 ;
  assign n11993 = ( n11383 & n11385 ) | ( n11383 & ~n11992 ) | ( n11385 & ~n11992 ) ;
  assign n11994 = n11991 & n11993 ;
  assign n11995 = n11991 | n11993 ;
  assign n11996 = ~n11994 & n11995 ;
  assign n11997 = ~n11653 & n11655 ;
  assign n11998 = ( n11351 & n11653 ) | ( n11351 & ~n11997 ) | ( n11653 & ~n11997 ) ;
  assign n11999 = n11996 & n11998 ;
  assign n12000 = n11653 & n11996 ;
  assign n12001 = ( ~n11655 & n11996 ) | ( ~n11655 & n12000 ) | ( n11996 & n12000 ) ;
  assign n12002 = ( n11355 & n11999 ) | ( n11355 & n12001 ) | ( n11999 & n12001 ) ;
  assign n12003 = n11999 & n12001 ;
  assign n12004 = ( n11360 & n12002 ) | ( n11360 & n12003 ) | ( n12002 & n12003 ) ;
  assign n12005 = ~n11997 & n11998 ;
  assign n12006 = n11996 | n12005 ;
  assign n12007 = ( n11355 & ~n11997 ) | ( n11355 & n11998 ) | ( ~n11997 & n11998 ) ;
  assign n12008 = n11996 | n12007 ;
  assign n12009 = ( n11360 & n12006 ) | ( n11360 & n12008 ) | ( n12006 & n12008 ) ;
  assign n12010 = ~n12004 & n12009 ;
  assign n12011 = ~n11663 & n12010 ;
  assign n12012 = n11663 & ~n12010 ;
  assign n12013 = n11664 & ~n12012 ;
  assign n12014 = ~n12011 & n12013 ;
  assign n12015 = n12011 | n12012 ;
  assign n12016 = ( n11672 & n12014 ) | ( n11672 & ~n12015 ) | ( n12014 & ~n12015 ) ;
  assign n12017 = n11673 & ~n12016 ;
  assign n12019 = n2315 & n12010 ;
  assign n12020 = n2308 & ~n11663 ;
  assign n12021 = n12019 | n12020 ;
  assign n12018 = n2312 & n11363 ;
  assign n12023 = n2306 | n12018 ;
  assign n12024 = n12021 | n12023 ;
  assign n12022 = n12018 | n12021 ;
  assign n12025 = n12022 & n12024 ;
  assign n12026 = ( ~n11663 & n11664 ) | ( ~n11663 & n12010 ) | ( n11664 & n12010 ) ;
  assign n12027 = n12012 | n12026 ;
  assign n12028 = n11672 | n12027 ;
  assign n12029 = ( n12024 & n12025 ) | ( n12024 & ~n12028 ) | ( n12025 & ~n12028 ) ;
  assign n12030 = n12024 | n12025 ;
  assign n12031 = ( n12017 & n12029 ) | ( n12017 & n12030 ) | ( n12029 & n12030 ) ;
  assign n12032 = ~x26 & n12031 ;
  assign n12033 = x26 | n12031 ;
  assign n12034 = ( ~n12031 & n12032 ) | ( ~n12031 & n12033 ) | ( n12032 & n12033 ) ;
  assign n12035 = n11054 & n12034 ;
  assign n12036 = n10975 & ~n11049 ;
  assign n12037 = n11050 | n12036 ;
  assign n12038 = n10694 & n11668 ;
  assign n12039 = ~n11664 & n11672 ;
  assign n12040 = ( n11666 & n12038 ) | ( n11666 & ~n12039 ) | ( n12038 & ~n12039 ) ;
  assign n12041 = n2308 & n11363 ;
  assign n12042 = n2312 & n10649 ;
  assign n12043 = n12041 | n12042 ;
  assign n12044 = n2315 & ~n11663 ;
  assign n12045 = n2306 | n12044 ;
  assign n12046 = n12043 | n12045 ;
  assign n12047 = n12043 | n12044 ;
  assign n12048 = n11664 | n11665 ;
  assign n12049 = ~n12047 & n12048 ;
  assign n12050 = ( n11672 & ~n12047 ) | ( n11672 & n12049 ) | ( ~n12047 & n12049 ) ;
  assign n12051 = n12046 & ~n12050 ;
  assign n12052 = ( n12040 & n12046 ) | ( n12040 & n12051 ) | ( n12046 & n12051 ) ;
  assign n12053 = x26 & n12052 ;
  assign n12054 = x26 & ~n12052 ;
  assign n12055 = ( n12052 & ~n12053 ) | ( n12052 & n12054 ) | ( ~n12053 & n12054 ) ;
  assign n12056 = ~n12037 & n12055 ;
  assign n12057 = n11005 | n11048 ;
  assign n12058 = n10694 | n11668 ;
  assign n12059 = ~n12038 & n12058 ;
  assign n12060 = n2315 & n11363 ;
  assign n12061 = n2312 & n10325 ;
  assign n12062 = n2308 & n10649 ;
  assign n12063 = n12061 | n12062 ;
  assign n12064 = n12060 | n12063 ;
  assign n12065 = n2306 | n12064 ;
  assign n12066 = n12064 & n12065 ;
  assign n12067 = ( n12059 & n12065 ) | ( n12059 & n12066 ) | ( n12065 & n12066 ) ;
  assign n12068 = x26 & n12066 ;
  assign n12069 = x26 & n12065 ;
  assign n12070 = ( n12059 & n12068 ) | ( n12059 & n12069 ) | ( n12068 & n12069 ) ;
  assign n12071 = x26 & ~n12068 ;
  assign n12072 = x26 & ~n12069 ;
  assign n12073 = ( ~n12059 & n12071 ) | ( ~n12059 & n12072 ) | ( n12071 & n12072 ) ;
  assign n12074 = ( n12067 & ~n12070 ) | ( n12067 & n12073 ) | ( ~n12070 & n12073 ) ;
  assign n12075 = n11005 & n11047 ;
  assign n12076 = n12074 & n12075 ;
  assign n12077 = ( ~n12057 & n12074 ) | ( ~n12057 & n12076 ) | ( n12074 & n12076 ) ;
  assign n12078 = n2308 & n10325 ;
  assign n12079 = n2312 & n10654 ;
  assign n12080 = n2312 | n2315 ;
  assign n12081 = ( n2315 & n10654 ) | ( n2315 & n12080 ) | ( n10654 & n12080 ) ;
  assign n12082 = ( n10649 & n12079 ) | ( n10649 & n12081 ) | ( n12079 & n12081 ) ;
  assign n12083 = n12078 | n12082 ;
  assign n12084 = n2306 | n12083 ;
  assign n12085 = ( n10702 & n12083 ) | ( n10702 & n12084 ) | ( n12083 & n12084 ) ;
  assign n12086 = n12083 | n12084 ;
  assign n12087 = ( n10695 & n12085 ) | ( n10695 & n12086 ) | ( n12085 & n12086 ) ;
  assign n12088 = ~x26 & n12087 ;
  assign n12089 = x26 & n12083 ;
  assign n12090 = x26 & n2306 ;
  assign n12091 = ( x26 & n12083 ) | ( x26 & n12090 ) | ( n12083 & n12090 ) ;
  assign n12092 = ( n10702 & n12089 ) | ( n10702 & n12091 ) | ( n12089 & n12091 ) ;
  assign n12093 = n12089 | n12091 ;
  assign n12094 = ( n10695 & n12092 ) | ( n10695 & n12093 ) | ( n12092 & n12093 ) ;
  assign n12095 = x26 & ~n12094 ;
  assign n12096 = n12088 | n12095 ;
  assign n12097 = ~n11006 & n11030 ;
  assign n12098 = n11006 | n11028 ;
  assign n12099 = ( n11031 & n12097 ) | ( n11031 & ~n12098 ) | ( n12097 & ~n12098 ) ;
  assign n12100 = n11045 & n12099 ;
  assign n12101 = n11006 & ~n11030 ;
  assign n12102 = n11006 & n11028 ;
  assign n12103 = ( ~n11031 & n12101 ) | ( ~n11031 & n12102 ) | ( n12101 & n12102 ) ;
  assign n12104 = ( n11006 & ~n11045 ) | ( n11006 & n12103 ) | ( ~n11045 & n12103 ) ;
  assign n12105 = n12100 | n12104 ;
  assign n12106 = n11019 & n12105 ;
  assign n12107 = n11019 | n12105 ;
  assign n12108 = ~n12106 & n12107 ;
  assign n12109 = n12096 & n12108 ;
  assign n12110 = n12096 | n12108 ;
  assign n12111 = ~n12109 & n12110 ;
  assign n12112 = n2315 & n10325 ;
  assign n12113 = n2312 & ~n10662 ;
  assign n12114 = n2308 & n10654 ;
  assign n12115 = n12113 | n12114 ;
  assign n12116 = n12112 | n12115 ;
  assign n12117 = n2306 | n12116 ;
  assign n12118 = ( ~n10957 & n12116 ) | ( ~n10957 & n12117 ) | ( n12116 & n12117 ) ;
  assign n12119 = n12116 | n12117 ;
  assign n12120 = ( n10949 & n12118 ) | ( n10949 & n12119 ) | ( n12118 & n12119 ) ;
  assign n12121 = ~x26 & n12120 ;
  assign n12122 = x26 & n12116 ;
  assign n12123 = ( x26 & n12090 ) | ( x26 & n12116 ) | ( n12090 & n12116 ) ;
  assign n12124 = ( ~n10957 & n12122 ) | ( ~n10957 & n12123 ) | ( n12122 & n12123 ) ;
  assign n12125 = n12122 | n12123 ;
  assign n12126 = ( n10949 & n12124 ) | ( n10949 & n12125 ) | ( n12124 & n12125 ) ;
  assign n12127 = x26 & ~n12126 ;
  assign n12128 = n12121 | n12127 ;
  assign n12129 = n11032 | n11045 ;
  assign n12130 = ~n11046 & n12129 ;
  assign n12131 = n12128 & n12130 ;
  assign n12132 = n12128 | n12130 ;
  assign n12133 = ~n12131 & n12132 ;
  assign n12134 = n11038 | n11041 ;
  assign n12135 = ~n11041 & n11043 ;
  assign n12136 = ( n11039 & n12134 ) | ( n11039 & ~n12135 ) | ( n12134 & ~n12135 ) ;
  assign n12137 = ~n11045 & n12136 ;
  assign n12138 = n2315 & n10654 ;
  assign n12139 = n2312 & n10667 ;
  assign n12140 = n2308 & ~n10662 ;
  assign n12141 = n12139 | n12140 ;
  assign n12142 = n12138 | n12141 ;
  assign n12143 = n2306 | n12138 ;
  assign n12144 = n12141 | n12143 ;
  assign n12145 = ( n10978 & n12142 ) | ( n10978 & n12144 ) | ( n12142 & n12144 ) ;
  assign n12146 = x26 & n12144 ;
  assign n12147 = x26 & n12142 ;
  assign n12148 = ( n10978 & n12146 ) | ( n10978 & n12147 ) | ( n12146 & n12147 ) ;
  assign n12149 = x26 & ~n12147 ;
  assign n12150 = x26 & ~n12146 ;
  assign n12151 = ( ~n10978 & n12149 ) | ( ~n10978 & n12150 ) | ( n12149 & n12150 ) ;
  assign n12152 = ( n12145 & ~n12148 ) | ( n12145 & n12151 ) | ( ~n12148 & n12151 ) ;
  assign n12153 = n12137 & n12152 ;
  assign n12154 = n2306 & n10784 ;
  assign n12155 = n2315 & ~n10675 ;
  assign n12156 = n2308 & ~n10678 ;
  assign n12157 = n12155 | n12156 ;
  assign n12158 = x26 | n12157 ;
  assign n12159 = n12154 | n12158 ;
  assign n12160 = ~x26 & n12159 ;
  assign n12161 = x26 & ~n2302 ;
  assign n12162 = ( x26 & n10678 ) | ( x26 & n12161 ) | ( n10678 & n12161 ) ;
  assign n12163 = n12159 & n12162 ;
  assign n12164 = n12154 | n12157 ;
  assign n12165 = n12162 & ~n12164 ;
  assign n12166 = ( n12160 & n12163 ) | ( n12160 & n12165 ) | ( n12163 & n12165 ) ;
  assign n12167 = n2312 & ~n10678 ;
  assign n12168 = n2315 & n10667 ;
  assign n12169 = n2308 & ~n10675 ;
  assign n12170 = n12168 | n12169 ;
  assign n12171 = n12167 | n12170 ;
  assign n12172 = n10837 | n12171 ;
  assign n12173 = n2306 | n12167 ;
  assign n12174 = n12170 | n12173 ;
  assign n12175 = ~x26 & n12174 ;
  assign n12176 = n12172 & n12175 ;
  assign n12177 = x26 | n12176 ;
  assign n12178 = n1820 & ~n10678 ;
  assign n12179 = n12176 & n12178 ;
  assign n12180 = n12172 & n12174 ;
  assign n12181 = n12178 & ~n12180 ;
  assign n12182 = ( n12177 & n12179 ) | ( n12177 & n12181 ) | ( n12179 & n12181 ) ;
  assign n12183 = n12166 & n12182 ;
  assign n12184 = ( n12176 & n12177 ) | ( n12176 & ~n12180 ) | ( n12177 & ~n12180 ) ;
  assign n12185 = n12166 | n12178 ;
  assign n12186 = ( n12178 & n12184 ) | ( n12178 & n12185 ) | ( n12184 & n12185 ) ;
  assign n12187 = ~n12183 & n12186 ;
  assign n12188 = n2315 & ~n10662 ;
  assign n12189 = n2312 & ~n10675 ;
  assign n12190 = n2308 & n10667 ;
  assign n12191 = n12189 | n12190 ;
  assign n12192 = n12188 | n12191 ;
  assign n12193 = ( n2306 & n10850 ) | ( n2306 & n12192 ) | ( n10850 & n12192 ) ;
  assign n12194 = ( x26 & n2306 ) | ( x26 & ~n12192 ) | ( n2306 & ~n12192 ) ;
  assign n12195 = ( x26 & n10850 ) | ( x26 & n12194 ) | ( n10850 & n12194 ) ;
  assign n12196 = ~n12193 & n12195 ;
  assign n12197 = n12192 | n12195 ;
  assign n12198 = ( ~x26 & n12196 ) | ( ~x26 & n12197 ) | ( n12196 & n12197 ) ;
  assign n12199 = n12183 | n12198 ;
  assign n12200 = ( n12183 & n12187 ) | ( n12183 & n12199 ) | ( n12187 & n12199 ) ;
  assign n12201 = n12137 | n12152 ;
  assign n12202 = ~n12153 & n12201 ;
  assign n12203 = n12153 | n12202 ;
  assign n12204 = ( n12153 & n12200 ) | ( n12153 & n12203 ) | ( n12200 & n12203 ) ;
  assign n12205 = n12133 & n12204 ;
  assign n12206 = n12131 | n12205 ;
  assign n12207 = n12111 & n12206 ;
  assign n12208 = n12074 | n12075 ;
  assign n12209 = n12057 & ~n12208 ;
  assign n12210 = n12077 | n12209 ;
  assign n12211 = n12109 & ~n12210 ;
  assign n12212 = ( n12207 & ~n12210 ) | ( n12207 & n12211 ) | ( ~n12210 & n12211 ) ;
  assign n12213 = n12077 | n12212 ;
  assign n12214 = n12037 | n12056 ;
  assign n12215 = n12037 & n12055 ;
  assign n12216 = n12214 & ~n12215 ;
  assign n12217 = n12213 & ~n12216 ;
  assign n12218 = n12056 | n12217 ;
  assign n12219 = n11054 & ~n12035 ;
  assign n12220 = ~n11054 & n12034 ;
  assign n12221 = n12219 | n12220 ;
  assign n12222 = n12218 & n12221 ;
  assign n12223 = n12035 | n12222 ;
  assign n12224 = n1829 & n11363 ;
  assign n12225 = n1826 & n10325 ;
  assign n12226 = n1823 & n10649 ;
  assign n12227 = n12225 | n12226 ;
  assign n12228 = n12224 | n12227 ;
  assign n12229 = n1821 | n12228 ;
  assign n12230 = ( n12059 & n12228 ) | ( n12059 & n12229 ) | ( n12228 & n12229 ) ;
  assign n12231 = x29 & n12229 ;
  assign n12232 = x29 & n12228 ;
  assign n12233 = ( n12059 & n12231 ) | ( n12059 & n12232 ) | ( n12231 & n12232 ) ;
  assign n12234 = x29 & ~n12231 ;
  assign n12235 = x29 & ~n12232 ;
  assign n12236 = ( ~n12059 & n12234 ) | ( ~n12059 & n12235 ) | ( n12234 & n12235 ) ;
  assign n12237 = ( n12230 & ~n12233 ) | ( n12230 & n12236 ) | ( ~n12233 & n12236 ) ;
  assign n12238 = n1057 & n10654 ;
  assign n12239 = n1065 & ~n10662 ;
  assign n12240 = n1060 & n10667 ;
  assign n12241 = n12239 | n12240 ;
  assign n12242 = n12238 | n12241 ;
  assign n12243 = n1062 | n12238 ;
  assign n12244 = n12241 | n12243 ;
  assign n12245 = ( n10978 & n12242 ) | ( n10978 & n12244 ) | ( n12242 & n12244 ) ;
  assign n12246 = n272 | n608 ;
  assign n12247 = n470 | n12246 ;
  assign n12248 = n196 | n12247 ;
  assign n12249 = n1673 | n3393 ;
  assign n12250 = n2787 | n12249 ;
  assign n12251 = n12248 | n12250 ;
  assign n12252 = n324 | n5956 ;
  assign n12253 = n12251 | n12252 ;
  assign n12254 = n1733 | n12253 ;
  assign n12255 = n90 | n12254 ;
  assign n12256 = n3337 | n12255 ;
  assign n12257 = n205 | n288 ;
  assign n12258 = n341 | n489 ;
  assign n12259 = n12257 | n12258 ;
  assign n12260 = n607 | n12259 ;
  assign n12261 = n227 | n1583 ;
  assign n12262 = n317 | n382 ;
  assign n12263 = n12261 | n12262 ;
  assign n12264 = n399 | n648 ;
  assign n12265 = n237 | n720 ;
  assign n12266 = n12264 | n12265 ;
  assign n12267 = n12263 | n12266 ;
  assign n12268 = n168 | n450 ;
  assign n12269 = n766 | n12268 ;
  assign n12270 = n239 | n501 ;
  assign n12271 = n447 | n12270 ;
  assign n12272 = n12269 | n12271 ;
  assign n12273 = n12267 | n12272 ;
  assign n12274 = n184 | n590 ;
  assign n12275 = n839 | n12274 ;
  assign n12276 = n6848 & ~n12275 ;
  assign n12277 = n206 | n581 ;
  assign n12278 = n5946 | n12277 ;
  assign n12279 = n12276 & ~n12278 ;
  assign n12280 = n349 | n365 ;
  assign n12281 = n419 | n764 ;
  assign n12282 = n12280 | n12281 ;
  assign n12283 = n53 | n406 ;
  assign n12284 = n12282 | n12283 ;
  assign n12285 = n12279 & ~n12284 ;
  assign n12286 = ~n12273 & n12285 ;
  assign n12287 = n92 | n696 ;
  assign n12288 = n139 | n278 ;
  assign n12289 = n12287 | n12288 ;
  assign n12290 = n229 | n513 ;
  assign n12291 = n12289 | n12290 ;
  assign n12292 = n1013 | n12291 ;
  assign n12293 = n12286 & ~n12292 ;
  assign n12294 = ~n12260 & n12293 ;
  assign n12295 = ~n12256 & n12294 ;
  assign n12296 = n12244 & ~n12295 ;
  assign n12297 = n12238 & ~n12295 ;
  assign n12298 = ( n12241 & ~n12295 ) | ( n12241 & n12297 ) | ( ~n12295 & n12297 ) ;
  assign n12299 = ( n10978 & n12296 ) | ( n10978 & n12298 ) | ( n12296 & n12298 ) ;
  assign n12300 = n12245 & ~n12299 ;
  assign n12301 = n12244 | n12295 ;
  assign n12302 = n12242 | n12295 ;
  assign n12303 = ( n10978 & n12301 ) | ( n10978 & n12302 ) | ( n12301 & n12302 ) ;
  assign n12304 = ~n12300 & n12303 ;
  assign n12305 = n10938 | n10942 ;
  assign n12306 = ( n10848 & n10938 ) | ( n10848 & n12305 ) | ( n10938 & n12305 ) ;
  assign n12307 = n12304 & n12306 ;
  assign n12308 = n12304 | n12306 ;
  assign n12309 = ~n12307 & n12308 ;
  assign n12310 = n12237 & ~n12309 ;
  assign n12311 = n12237 & ~n12310 ;
  assign n12312 = n12309 | n12310 ;
  assign n12313 = ~n12311 & n12312 ;
  assign n12314 = n10946 | n10948 ;
  assign n12315 = ( n10946 & n11051 ) | ( n10946 & n12314 ) | ( n11051 & n12314 ) ;
  assign n12316 = ~n12313 & n12315 ;
  assign n12317 = n12313 & ~n12315 ;
  assign n12318 = n12316 | n12317 ;
  assign n12319 = n7068 & ~n8982 ;
  assign n12320 = ( n7068 & n9051 ) | ( n7068 & n12319 ) | ( n9051 & n12319 ) ;
  assign n12321 = n7074 & ~n9022 ;
  assign n12322 = ( n7074 & n12320 ) | ( n7074 & ~n12321 ) | ( n12320 & ~n12321 ) ;
  assign n12323 = n7074 | n12320 ;
  assign n12324 = ( ~n9019 & n12322 ) | ( ~n9019 & n12323 ) | ( n12322 & n12323 ) ;
  assign n12325 = n7078 | n12324 ;
  assign n12326 = ( n9078 & n12324 ) | ( n9078 & n12325 ) | ( n12324 & n12325 ) ;
  assign n12327 = x8 & n12325 ;
  assign n12328 = x8 & n12324 ;
  assign n12329 = ( n9078 & n12327 ) | ( n9078 & n12328 ) | ( n12327 & n12328 ) ;
  assign n12330 = x8 & ~n12327 ;
  assign n12331 = x8 & ~n12328 ;
  assign n12332 = ( ~n9078 & n12330 ) | ( ~n9078 & n12331 ) | ( n12330 & n12331 ) ;
  assign n12333 = ( n12326 & ~n12329 ) | ( n12326 & n12332 ) | ( ~n12329 & n12332 ) ;
  assign n12334 = n11715 | n11981 ;
  assign n12335 = ( n11715 & n11717 ) | ( n11715 & n12334 ) | ( n11717 & n12334 ) ;
  assign n12336 = n12333 & n12335 ;
  assign n12337 = n12333 | n12335 ;
  assign n12338 = ~n12336 & n12337 ;
  assign n12339 = n11897 | n11903 ;
  assign n12340 = n1060 & n2090 ;
  assign n12341 = ( n1060 & ~n2082 ) | ( n1060 & n12340 ) | ( ~n2082 & n12340 ) ;
  assign n12342 = n1057 & n2691 ;
  assign n12343 = ( n1057 & n2678 ) | ( n1057 & n12342 ) | ( n2678 & n12342 ) ;
  assign n12344 = n1065 & n2199 ;
  assign n12345 = ( n1065 & ~n2185 ) | ( n1065 & n12344 ) | ( ~n2185 & n12344 ) ;
  assign n12346 = n12343 | n12345 ;
  assign n12347 = n12341 | n12346 ;
  assign n12348 = n1062 | n12347 ;
  assign n12349 = ( n2985 & n12347 ) | ( n2985 & n12348 ) | ( n12347 & n12348 ) ;
  assign n12350 = n182 | n11785 ;
  assign n12351 = n11779 | n12350 ;
  assign n12352 = n11768 | n12351 ;
  assign n12353 = ( x2 & x5 ) | ( x2 & ~n12352 ) | ( x5 & ~n12352 ) ;
  assign n12354 = n176 | n412 ;
  assign n12355 = n720 | n12354 ;
  assign n12356 = n5042 | n12355 ;
  assign n12357 = n2706 | n12356 ;
  assign n12358 = n880 | n2846 ;
  assign n12359 = n179 | n318 ;
  assign n12360 = n222 | n12359 ;
  assign n12361 = n12358 | n12360 ;
  assign n12362 = n333 | n383 ;
  assign n12363 = n12361 | n12362 ;
  assign n12364 = n12357 | n12363 ;
  assign n12365 = n986 | n2256 ;
  assign n12366 = n695 | n3425 ;
  assign n12367 = n12365 | n12366 ;
  assign n12368 = n168 | n223 ;
  assign n12369 = n118 | n363 ;
  assign n12370 = n12368 | n12369 ;
  assign n12371 = n569 | n12370 ;
  assign n12372 = n12367 | n12371 ;
  assign n12373 = n1133 | n12372 ;
  assign n12374 = n12364 | n12373 ;
  assign n12375 = n1113 & ~n12374 ;
  assign n12376 = n170 | n355 ;
  assign n12377 = n1005 | n12376 ;
  assign n12378 = n1652 | n12377 ;
  assign n12379 = n1384 | n12378 ;
  assign n12380 = n510 | n1172 ;
  assign n12381 = n229 | n12380 ;
  assign n12382 = ( n202 & ~n2806 ) | ( n202 & n12381 ) | ( ~n2806 & n12381 ) ;
  assign n12383 = n624 | n2806 ;
  assign n12384 = n12382 | n12383 ;
  assign n12385 = n12379 | n12384 ;
  assign n12386 = n937 | n2129 ;
  assign n12387 = n255 | n581 ;
  assign n12388 = n442 | n12387 ;
  assign n12389 = n12386 | n12388 ;
  assign n12390 = n775 | n12389 ;
  assign n12391 = n321 | n340 ;
  assign n12392 = n134 | n226 ;
  assign n12393 = n12391 | n12392 ;
  assign n12394 = n281 | n468 ;
  assign n12395 = n348 | n12394 ;
  assign n12396 = n12393 | n12395 ;
  assign n12397 = n12390 | n12396 ;
  assign n12398 = n12385 | n12397 ;
  assign n12399 = n10341 | n12398 ;
  assign n12400 = n152 | n387 ;
  assign n12401 = n9118 | n12400 ;
  assign n12402 = n131 | n280 ;
  assign n12403 = n517 | n12402 ;
  assign n12404 = n12401 | n12403 ;
  assign n12405 = n154 | n354 ;
  assign n12406 = n12404 | n12405 ;
  assign n12407 = n12399 | n12406 ;
  assign n12408 = n12375 & ~n12407 ;
  assign n12409 = ~n12353 & n12408 ;
  assign n12410 = n12353 & ~n12408 ;
  assign n12411 = n12409 | n12410 ;
  assign n12412 = n12348 & n12411 ;
  assign n12413 = n12347 & n12411 ;
  assign n12414 = ( n2985 & n12412 ) | ( n2985 & n12413 ) | ( n12412 & n12413 ) ;
  assign n12415 = n12411 & ~n12413 ;
  assign n12416 = n12411 & ~n12412 ;
  assign n12417 = ( ~n2985 & n12415 ) | ( ~n2985 & n12416 ) | ( n12415 & n12416 ) ;
  assign n12418 = ( n12349 & ~n12414 ) | ( n12349 & n12417 ) | ( ~n12414 & n12417 ) ;
  assign n12419 = n11804 | n11820 ;
  assign n12420 = ( n11804 & n11808 ) | ( n11804 & n12419 ) | ( n11808 & n12419 ) ;
  assign n12421 = ~n12418 & n12420 ;
  assign n12422 = n12418 & ~n12420 ;
  assign n12423 = n12421 | n12422 ;
  assign n12424 = n1823 & n2893 ;
  assign n12425 = ( n1823 & ~n2886 ) | ( n1823 & n12424 ) | ( ~n2886 & n12424 ) ;
  assign n12426 = n1826 & n2701 ;
  assign n12427 = ( n1826 & ~n2784 ) | ( n1826 & n12426 ) | ( ~n2784 & n12426 ) ;
  assign n12428 = n1829 & n3507 ;
  assign n12429 = ( n1829 & n3483 ) | ( n1829 & n12428 ) | ( n3483 & n12428 ) ;
  assign n12430 = n12427 | n12429 ;
  assign n12431 = n12425 | n12430 ;
  assign n12432 = n1821 | n12431 ;
  assign n12433 = n12431 & n12432 ;
  assign n12434 = ( n3603 & n12432 ) | ( n3603 & n12433 ) | ( n12432 & n12433 ) ;
  assign n12435 = x29 & n12433 ;
  assign n12436 = x29 & n12432 ;
  assign n12437 = ( n3603 & n12435 ) | ( n3603 & n12436 ) | ( n12435 & n12436 ) ;
  assign n12438 = x29 & ~n12435 ;
  assign n12439 = x29 & ~n12436 ;
  assign n12440 = ( ~n3603 & n12438 ) | ( ~n3603 & n12439 ) | ( n12438 & n12439 ) ;
  assign n12441 = ( n12434 & ~n12437 ) | ( n12434 & n12440 ) | ( ~n12437 & n12440 ) ;
  assign n12442 = ~n12423 & n12441 ;
  assign n12443 = n12423 & ~n12441 ;
  assign n12444 = n12442 | n12443 ;
  assign n12445 = n11827 | n11849 ;
  assign n12446 = ( n11827 & n11832 ) | ( n11827 & n12445 ) | ( n11832 & n12445 ) ;
  assign n12447 = ~n12444 & n12446 ;
  assign n12448 = n12444 & ~n12446 ;
  assign n12449 = n12447 | n12448 ;
  assign n12450 = n2315 & n4206 ;
  assign n12451 = n2312 & n3386 ;
  assign n12452 = n2308 & n3439 ;
  assign n12453 = ( n2308 & ~n3420 ) | ( n2308 & n12452 ) | ( ~n3420 & n12452 ) ;
  assign n12454 = n12451 | n12453 ;
  assign n12455 = n12450 | n12454 ;
  assign n12456 = n2306 | n12450 ;
  assign n12457 = n12454 | n12456 ;
  assign n12458 = ( ~n4220 & n12455 ) | ( ~n4220 & n12457 ) | ( n12455 & n12457 ) ;
  assign n12459 = ~x26 & n12457 ;
  assign n12460 = ~x26 & n12455 ;
  assign n12461 = ( ~n4220 & n12459 ) | ( ~n4220 & n12460 ) | ( n12459 & n12460 ) ;
  assign n12462 = x26 | n12460 ;
  assign n12463 = x26 | n12459 ;
  assign n12464 = ( ~n4220 & n12462 ) | ( ~n4220 & n12463 ) | ( n12462 & n12463 ) ;
  assign n12465 = ( ~n12458 & n12461 ) | ( ~n12458 & n12464 ) | ( n12461 & n12464 ) ;
  assign n12466 = n12449 | n12465 ;
  assign n12467 = n12449 & ~n12465 ;
  assign n12468 = ( ~n12449 & n12466 ) | ( ~n12449 & n12467 ) | ( n12466 & n12467 ) ;
  assign n12469 = n11871 | n11877 ;
  assign n12470 = ( n11871 & n11875 ) | ( n11871 & n12469 ) | ( n11875 & n12469 ) ;
  assign n12471 = ~n12468 & n12470 ;
  assign n12472 = n12468 & ~n12470 ;
  assign n12473 = n12471 | n12472 ;
  assign n12474 = n2925 & ~n4429 ;
  assign n12475 = n2928 & n4396 ;
  assign n12476 = n12474 | n12475 ;
  assign n12477 = n2932 & n4245 ;
  assign n12478 = ( n2932 & n4303 ) | ( n2932 & n12477 ) | ( n4303 & n12477 ) ;
  assign n12479 = n12476 | n12478 ;
  assign n12480 = n2936 | n12478 ;
  assign n12481 = n12476 | n12480 ;
  assign n12482 = ( n4455 & n12479 ) | ( n4455 & n12481 ) | ( n12479 & n12481 ) ;
  assign n12483 = x23 & n12481 ;
  assign n12484 = x23 & n12479 ;
  assign n12485 = ( n4455 & n12483 ) | ( n4455 & n12484 ) | ( n12483 & n12484 ) ;
  assign n12486 = x23 & ~n12484 ;
  assign n12487 = x23 & ~n12483 ;
  assign n12488 = ( ~n4455 & n12486 ) | ( ~n4455 & n12487 ) | ( n12486 & n12487 ) ;
  assign n12489 = ( n12482 & ~n12485 ) | ( n12482 & n12488 ) | ( ~n12485 & n12488 ) ;
  assign n12490 = n12473 | n12489 ;
  assign n12491 = n12473 & ~n12489 ;
  assign n12492 = ( ~n12473 & n12490 ) | ( ~n12473 & n12491 ) | ( n12490 & n12491 ) ;
  assign n12493 = n12339 & ~n12492 ;
  assign n12494 = ~n12339 & n12492 ;
  assign n12495 = n12493 | n12494 ;
  assign n12496 = n3541 & n5117 ;
  assign n12497 = ( n3541 & ~n5037 ) | ( n3541 & n12496 ) | ( ~n5037 & n12496 ) ;
  assign n12498 = n3547 & n5108 ;
  assign n12499 = n3544 & n5192 ;
  assign n12500 = ( n3544 & n5179 ) | ( n3544 & n12499 ) | ( n5179 & n12499 ) ;
  assign n12501 = n12498 | n12500 ;
  assign n12502 = n12497 | n12501 ;
  assign n12503 = n3537 | n12502 ;
  assign n12504 = ( ~n5220 & n12502 ) | ( ~n5220 & n12503 ) | ( n12502 & n12503 ) ;
  assign n12505 = ~x20 & n12503 ;
  assign n12506 = ~x20 & n12502 ;
  assign n12507 = ( ~n5220 & n12505 ) | ( ~n5220 & n12506 ) | ( n12505 & n12506 ) ;
  assign n12508 = x20 | n12505 ;
  assign n12509 = x20 | n12506 ;
  assign n12510 = ( ~n5220 & n12508 ) | ( ~n5220 & n12509 ) | ( n12508 & n12509 ) ;
  assign n12511 = ( ~n12504 & n12507 ) | ( ~n12504 & n12510 ) | ( n12507 & n12510 ) ;
  assign n12512 = ~n12495 & n12511 ;
  assign n12513 = n12495 | n12512 ;
  assign n12515 = n11926 | n11930 ;
  assign n12516 = ( n11926 & n11928 ) | ( n11926 & n12515 ) | ( n11928 & n12515 ) ;
  assign n12514 = n12495 & n12511 ;
  assign n12517 = n12514 & n12516 ;
  assign n12518 = ( ~n12513 & n12516 ) | ( ~n12513 & n12517 ) | ( n12516 & n12517 ) ;
  assign n12519 = n12514 | n12516 ;
  assign n12520 = n12513 & ~n12519 ;
  assign n12521 = n12518 | n12520 ;
  assign n12522 = n4468 & n5857 ;
  assign n12523 = ( n4468 & ~n5899 ) | ( n4468 & n12522 ) | ( ~n5899 & n12522 ) ;
  assign n12524 = n4471 & ~n6091 ;
  assign n12525 = n4466 & n5997 ;
  assign n12526 = ( n4466 & n5979 ) | ( n4466 & n12525 ) | ( n5979 & n12525 ) ;
  assign n12527 = n12524 | n12526 ;
  assign n12528 = n12523 | n12527 ;
  assign n12529 = n4475 | n12528 ;
  assign n12530 = ( n6108 & n12528 ) | ( n6108 & n12529 ) | ( n12528 & n12529 ) ;
  assign n12531 = x17 & n12529 ;
  assign n12532 = x17 & n12528 ;
  assign n12533 = ( n6108 & n12531 ) | ( n6108 & n12532 ) | ( n12531 & n12532 ) ;
  assign n12534 = x17 & ~n12531 ;
  assign n12535 = x17 & ~n12532 ;
  assign n12536 = ( ~n6108 & n12534 ) | ( ~n6108 & n12535 ) | ( n12534 & n12535 ) ;
  assign n12537 = ( n12530 & ~n12533 ) | ( n12530 & n12536 ) | ( ~n12533 & n12536 ) ;
  assign n12538 = ~n12521 & n12537 ;
  assign n12539 = n12521 | n12538 ;
  assign n12541 = n11950 | n11954 ;
  assign n12542 = ( n11950 & n11952 ) | ( n11950 & n12541 ) | ( n11952 & n12541 ) ;
  assign n12540 = n12521 & n12537 ;
  assign n12543 = n12540 & n12542 ;
  assign n12544 = ( ~n12539 & n12542 ) | ( ~n12539 & n12543 ) | ( n12542 & n12543 ) ;
  assign n12545 = n12540 | n12542 ;
  assign n12546 = n12539 & ~n12545 ;
  assign n12547 = n12544 | n12546 ;
  assign n12548 = n5231 & n6950 ;
  assign n12549 = n5237 & n7036 ;
  assign n12550 = ( n5237 & n7023 ) | ( n5237 & n12549 ) | ( n7023 & n12549 ) ;
  assign n12551 = n12548 | n12550 ;
  assign n12552 = n5234 & n6889 ;
  assign n12553 = ( n5234 & ~n6884 ) | ( n5234 & n12552 ) | ( ~n6884 & n12552 ) ;
  assign n12554 = n12551 | n12553 ;
  assign n12555 = n5227 | n12553 ;
  assign n12556 = n12551 | n12555 ;
  assign n12557 = ( ~n7061 & n12554 ) | ( ~n7061 & n12556 ) | ( n12554 & n12556 ) ;
  assign n12558 = ~x14 & n12556 ;
  assign n12559 = ~x14 & n12554 ;
  assign n12560 = ( ~n7061 & n12558 ) | ( ~n7061 & n12559 ) | ( n12558 & n12559 ) ;
  assign n12561 = x14 | n12559 ;
  assign n12562 = x14 | n12558 ;
  assign n12563 = ( ~n7061 & n12561 ) | ( ~n7061 & n12562 ) | ( n12561 & n12562 ) ;
  assign n12564 = ( ~n12557 & n12560 ) | ( ~n12557 & n12563 ) | ( n12560 & n12563 ) ;
  assign n12565 = n12547 | n12564 ;
  assign n12566 = n12547 & ~n12564 ;
  assign n12567 = ( ~n12547 & n12565 ) | ( ~n12547 & n12566 ) | ( n12565 & n12566 ) ;
  assign n12568 = n11974 | n11976 ;
  assign n12569 = ( n11974 & n11978 ) | ( n11974 & n12568 ) | ( n11978 & n12568 ) ;
  assign n12570 = ~n12567 & n12569 ;
  assign n12571 = n12567 & ~n12569 ;
  assign n12572 = n12570 | n12571 ;
  assign n12573 = n6125 & n7907 ;
  assign n12574 = ( n6125 & n7902 ) | ( n6125 & n12573 ) | ( n7902 & n12573 ) ;
  assign n12575 = n6119 & n8079 ;
  assign n12576 = ( n6119 & ~n8070 ) | ( n6119 & n12575 ) | ( ~n8070 & n12575 ) ;
  assign n12577 = n12574 | n12576 ;
  assign n12578 = n6122 & ~n8017 ;
  assign n12579 = n12577 | n12578 ;
  assign n12580 = n6115 | n12577 ;
  assign n12581 = n12578 | n12580 ;
  assign n12582 = ( n8104 & n12579 ) | ( n8104 & n12581 ) | ( n12579 & n12581 ) ;
  assign n12583 = x11 & n12581 ;
  assign n12584 = x11 & n12579 ;
  assign n12585 = ( n8104 & n12583 ) | ( n8104 & n12584 ) | ( n12583 & n12584 ) ;
  assign n12586 = x11 & ~n12584 ;
  assign n12587 = x11 & ~n12583 ;
  assign n12588 = ( ~n8104 & n12586 ) | ( ~n8104 & n12587 ) | ( n12586 & n12587 ) ;
  assign n12589 = ( n12582 & ~n12585 ) | ( n12582 & n12588 ) | ( ~n12585 & n12588 ) ;
  assign n12590 = n12572 | n12589 ;
  assign n12591 = n12572 & ~n12589 ;
  assign n12592 = ( ~n12572 & n12590 ) | ( ~n12572 & n12591 ) | ( n12590 & n12591 ) ;
  assign n12593 = n12338 & ~n12592 ;
  assign n12594 = ~n12338 & n12592 ;
  assign n12595 = n12593 | n12594 ;
  assign n12596 = n11693 & ~n12595 ;
  assign n12597 = ( n11987 & ~n12595 ) | ( n11987 & n12596 ) | ( ~n12595 & n12596 ) ;
  assign n12598 = ~n11693 & n12595 ;
  assign n12599 = ~n11987 & n12598 ;
  assign n12600 = n12597 | n12599 ;
  assign n12601 = n11994 | n11996 ;
  assign n12602 = ~n12600 & n12601 ;
  assign n12603 = n11994 & ~n12600 ;
  assign n12604 = ( n11998 & n12602 ) | ( n11998 & n12603 ) | ( n12602 & n12603 ) ;
  assign n12605 = ( n12001 & ~n12600 ) | ( n12001 & n12603 ) | ( ~n12600 & n12603 ) ;
  assign n12606 = ( n11355 & n12604 ) | ( n11355 & n12605 ) | ( n12604 & n12605 ) ;
  assign n12607 = n12604 & n12605 ;
  assign n12608 = ( n11360 & n12606 ) | ( n11360 & n12607 ) | ( n12606 & n12607 ) ;
  assign n12609 = n11994 | n12001 ;
  assign n12610 = ( n11994 & n11998 ) | ( n11994 & n12601 ) | ( n11998 & n12601 ) ;
  assign n12611 = n12609 & n12610 ;
  assign n12612 = n12600 & ~n12611 ;
  assign n12613 = ( n11355 & n12609 ) | ( n11355 & n12610 ) | ( n12609 & n12610 ) ;
  assign n12614 = n12600 & ~n12613 ;
  assign n12615 = ( ~n11360 & n12612 ) | ( ~n11360 & n12614 ) | ( n12612 & n12614 ) ;
  assign n12616 = n12608 | n12615 ;
  assign n12617 = n12010 & ~n12616 ;
  assign n12618 = ~n12010 & n12616 ;
  assign n12619 = n12617 | n12618 ;
  assign n12620 = n12026 & ~n12619 ;
  assign n12621 = n12012 | n12619 ;
  assign n12622 = ( n11672 & n12620 ) | ( n11672 & ~n12621 ) | ( n12620 & ~n12621 ) ;
  assign n12623 = ~n12026 & n12619 ;
  assign n12624 = n12012 & n12619 ;
  assign n12625 = ( ~n11672 & n12623 ) | ( ~n11672 & n12624 ) | ( n12623 & n12624 ) ;
  assign n12626 = n12622 | n12625 ;
  assign n12628 = n2308 & n12010 ;
  assign n12629 = n2315 & ~n12616 ;
  assign n12630 = n12628 | n12629 ;
  assign n12627 = n2312 & ~n11663 ;
  assign n12632 = n2306 | n12627 ;
  assign n12633 = n12630 | n12632 ;
  assign n12631 = n12627 | n12630 ;
  assign n12634 = n12631 & n12633 ;
  assign n12635 = ( ~n12626 & n12633 ) | ( ~n12626 & n12634 ) | ( n12633 & n12634 ) ;
  assign n12636 = ~x26 & n12634 ;
  assign n12637 = ~x26 & n12633 ;
  assign n12638 = ( ~n12626 & n12636 ) | ( ~n12626 & n12637 ) | ( n12636 & n12637 ) ;
  assign n12639 = x26 | n12636 ;
  assign n12640 = x26 | n12637 ;
  assign n12641 = ( ~n12626 & n12639 ) | ( ~n12626 & n12640 ) | ( n12639 & n12640 ) ;
  assign n12642 = ( ~n12635 & n12638 ) | ( ~n12635 & n12641 ) | ( n12638 & n12641 ) ;
  assign n12643 = ~n12318 & n12642 ;
  assign n12644 = n12318 | n12643 ;
  assign n12645 = n12318 & n12642 ;
  assign n12646 = n12644 & ~n12645 ;
  assign n12647 = n12223 & ~n12646 ;
  assign n12648 = n12223 & ~n12647 ;
  assign n12649 = n12223 | n12646 ;
  assign n12650 = ~n12648 & n12649 ;
  assign n12651 = n7074 & ~n8982 ;
  assign n12652 = ( n7074 & n9051 ) | ( n7074 & n12651 ) | ( n9051 & n12651 ) ;
  assign n12653 = n7078 | n12652 ;
  assign n12654 = n9442 & ~n12652 ;
  assign n12655 = n9074 & ~n12652 ;
  assign n12656 = ( ~n9440 & n12654 ) | ( ~n9440 & n12655 ) | ( n12654 & n12655 ) ;
  assign n12657 = n12653 & ~n12656 ;
  assign n12658 = n12652 & n12653 ;
  assign n12659 = ( ~n9442 & n12653 ) | ( ~n9442 & n12658 ) | ( n12653 & n12658 ) ;
  assign n12660 = ( ~n9072 & n12657 ) | ( ~n9072 & n12659 ) | ( n12657 & n12659 ) ;
  assign n12661 = ~x8 & n12657 ;
  assign n12662 = ~x8 & n12659 ;
  assign n12663 = ( ~n9072 & n12661 ) | ( ~n9072 & n12662 ) | ( n12661 & n12662 ) ;
  assign n12664 = x8 | n12661 ;
  assign n12665 = x8 | n12662 ;
  assign n12666 = ( ~n9072 & n12664 ) | ( ~n9072 & n12665 ) | ( n12664 & n12665 ) ;
  assign n12667 = ( ~n12660 & n12663 ) | ( ~n12660 & n12666 ) | ( n12663 & n12666 ) ;
  assign n12668 = n12570 | n12589 ;
  assign n12669 = ( n12570 & ~n12572 ) | ( n12570 & n12668 ) | ( ~n12572 & n12668 ) ;
  assign n12670 = n12667 & n12669 ;
  assign n12671 = n12667 | n12669 ;
  assign n12672 = ~n12670 & n12671 ;
  assign n12749 = n12421 | n12441 ;
  assign n12750 = ( n12421 & ~n12423 ) | ( n12421 & n12749 ) | ( ~n12423 & n12749 ) ;
  assign n12673 = n12348 & ~n12411 ;
  assign n12674 = n12409 | n12673 ;
  assign n12675 = n12347 | n12409 ;
  assign n12676 = ( n12409 & ~n12411 ) | ( n12409 & n12675 ) | ( ~n12411 & n12675 ) ;
  assign n12677 = ( n2985 & n12674 ) | ( n2985 & n12676 ) | ( n12674 & n12676 ) ;
  assign n12678 = n702 | n966 ;
  assign n12679 = n676 | n3288 ;
  assign n12680 = n12678 | n12679 ;
  assign n12681 = n500 | n12680 ;
  assign n12682 = n228 | n1172 ;
  assign n12683 = n355 | n12682 ;
  assign n12684 = n2116 | n12683 ;
  assign n12685 = n12681 | n12684 ;
  assign n12686 = n756 | n12685 ;
  assign n12687 = n484 | n1030 ;
  assign n12688 = n262 | n12687 ;
  assign n12689 = n250 | n277 ;
  assign n12690 = n438 | n12689 ;
  assign n12691 = n6916 | n12690 ;
  assign n12692 = n12688 | n12691 ;
  assign n12693 = n1149 | n12274 ;
  assign n12694 = n561 | n3495 ;
  assign n12695 = n12693 | n12694 ;
  assign n12696 = n138 | n735 ;
  assign n12697 = n96 | n469 ;
  assign n12698 = n12696 | n12697 ;
  assign n12699 = n110 | n332 ;
  assign n12700 = n12698 | n12699 ;
  assign n12701 = n12695 | n12700 ;
  assign n12702 = n12692 | n12701 ;
  assign n12703 = n12363 | n12702 ;
  assign n12704 = n12686 | n12703 ;
  assign n12705 = n10876 | n12704 ;
  assign n12706 = n325 | n401 ;
  assign n12707 = n384 | n4249 ;
  assign n12708 = n661 | n2233 ;
  assign n12709 = ( n296 & ~n12707 ) | ( n296 & n12708 ) | ( ~n12707 & n12708 ) ;
  assign n12710 = n631 | n12707 ;
  assign n12711 = n12709 | n12710 ;
  assign n12712 = n344 | n444 ;
  assign n12713 = n447 | n12712 ;
  assign n12714 = n12711 | n12713 ;
  assign n12715 = n12706 | n12714 ;
  assign n12716 = n12705 | n12715 ;
  assign n12717 = n12408 | n12716 ;
  assign n12718 = n12408 & n12716 ;
  assign n12719 = n12409 & ~n12718 ;
  assign n12720 = n12717 & n12719 ;
  assign n12721 = n12717 & ~n12718 ;
  assign n12722 = ( n12673 & n12720 ) | ( n12673 & n12721 ) | ( n12720 & n12721 ) ;
  assign n12723 = n12676 & n12721 ;
  assign n12724 = ( n2985 & n12722 ) | ( n2985 & n12723 ) | ( n12722 & n12723 ) ;
  assign n12725 = n12677 & ~n12724 ;
  assign n12726 = n12718 | n12722 ;
  assign n12727 = n12717 & ~n12726 ;
  assign n12728 = n12718 | n12723 ;
  assign n12729 = n12717 & ~n12728 ;
  assign n12730 = ( ~n2985 & n12727 ) | ( ~n2985 & n12729 ) | ( n12727 & n12729 ) ;
  assign n12731 = n12725 | n12730 ;
  assign n12732 = n1065 & n2691 ;
  assign n12733 = ( n1065 & n2678 ) | ( n1065 & n12732 ) | ( n2678 & n12732 ) ;
  assign n12734 = n1060 & n2199 ;
  assign n12735 = ( n1060 & ~n2185 ) | ( n1060 & n12734 ) | ( ~n2185 & n12734 ) ;
  assign n12736 = n12733 | n12735 ;
  assign n12737 = n1062 | n12736 ;
  assign n12738 = n1057 & n2701 ;
  assign n12739 = ( n1057 & ~n2784 ) | ( n1057 & n12738 ) | ( ~n2784 & n12738 ) ;
  assign n12740 = n12737 | n12739 ;
  assign n12741 = n12736 | n12739 ;
  assign n12742 = ( n2960 & n12740 ) | ( n2960 & n12741 ) | ( n12740 & n12741 ) ;
  assign n12743 = n12730 & n12742 ;
  assign n12744 = ( n12725 & n12742 ) | ( n12725 & n12743 ) | ( n12742 & n12743 ) ;
  assign n12745 = n12731 & ~n12744 ;
  assign n12746 = ~n12730 & n12742 ;
  assign n12747 = ~n12725 & n12746 ;
  assign n12748 = n12745 | n12747 ;
  assign n12751 = n12748 & n12750 ;
  assign n12752 = n12750 & ~n12751 ;
  assign n12753 = n12748 & ~n12751 ;
  assign n12754 = n12752 | n12753 ;
  assign n12755 = n1826 & n2893 ;
  assign n12756 = ( n1826 & ~n2886 ) | ( n1826 & n12755 ) | ( ~n2886 & n12755 ) ;
  assign n12757 = n1823 & n3507 ;
  assign n12758 = ( n1823 & n3483 ) | ( n1823 & n12757 ) | ( n3483 & n12757 ) ;
  assign n12759 = n12756 | n12758 ;
  assign n12760 = n1829 & n3386 ;
  assign n12762 = n1821 | n12760 ;
  assign n12763 = n12759 | n12762 ;
  assign n12761 = n12759 | n12760 ;
  assign n12764 = n12761 & n12763 ;
  assign n12765 = ( ~n3568 & n12763 ) | ( ~n3568 & n12764 ) | ( n12763 & n12764 ) ;
  assign n12766 = ~x29 & n12764 ;
  assign n12767 = ~x29 & n12763 ;
  assign n12768 = ( ~n3568 & n12766 ) | ( ~n3568 & n12767 ) | ( n12766 & n12767 ) ;
  assign n12769 = x29 | n12766 ;
  assign n12770 = x29 | n12767 ;
  assign n12771 = ( ~n3568 & n12769 ) | ( ~n3568 & n12770 ) | ( n12769 & n12770 ) ;
  assign n12772 = ( ~n12765 & n12768 ) | ( ~n12765 & n12771 ) | ( n12768 & n12771 ) ;
  assign n12773 = n12754 & n12772 ;
  assign n12774 = n12754 | n12772 ;
  assign n12775 = ~n12773 & n12774 ;
  assign n12776 = n2308 & n4206 ;
  assign n12777 = n2315 & ~n4429 ;
  assign n12778 = n2312 & n3439 ;
  assign n12779 = ( n2312 & ~n3420 ) | ( n2312 & n12778 ) | ( ~n3420 & n12778 ) ;
  assign n12780 = n12777 | n12779 ;
  assign n12781 = n12776 | n12780 ;
  assign n12782 = n2306 | n12776 ;
  assign n12783 = n12780 | n12782 ;
  assign n12784 = ( ~n4527 & n12781 ) | ( ~n4527 & n12783 ) | ( n12781 & n12783 ) ;
  assign n12785 = ~x26 & n12783 ;
  assign n12786 = ~x26 & n12781 ;
  assign n12787 = ( ~n4527 & n12785 ) | ( ~n4527 & n12786 ) | ( n12785 & n12786 ) ;
  assign n12788 = x26 | n12786 ;
  assign n12789 = x26 | n12785 ;
  assign n12790 = ( ~n4527 & n12788 ) | ( ~n4527 & n12789 ) | ( n12788 & n12789 ) ;
  assign n12791 = ( ~n12784 & n12787 ) | ( ~n12784 & n12790 ) | ( n12787 & n12790 ) ;
  assign n12792 = n12775 & ~n12791 ;
  assign n12793 = n12775 | n12791 ;
  assign n12794 = ( ~n12775 & n12792 ) | ( ~n12775 & n12793 ) | ( n12792 & n12793 ) ;
  assign n12795 = n12447 | n12465 ;
  assign n12796 = ( n12447 & ~n12449 ) | ( n12447 & n12795 ) | ( ~n12449 & n12795 ) ;
  assign n12797 = n12794 & n12796 ;
  assign n12798 = n12794 | n12796 ;
  assign n12799 = ~n12797 & n12798 ;
  assign n12800 = n2925 & n4396 ;
  assign n12801 = n2928 & n4245 ;
  assign n12802 = ( n2928 & n4303 ) | ( n2928 & n12801 ) | ( n4303 & n12801 ) ;
  assign n12803 = n12800 | n12802 ;
  assign n12804 = n2932 & n5192 ;
  assign n12805 = ( n2932 & n5179 ) | ( n2932 & n12804 ) | ( n5179 & n12804 ) ;
  assign n12806 = n12803 | n12805 ;
  assign n12807 = n2936 | n12805 ;
  assign n12808 = n12803 | n12807 ;
  assign n12809 = ( n5306 & n12806 ) | ( n5306 & n12808 ) | ( n12806 & n12808 ) ;
  assign n12810 = x23 & n12808 ;
  assign n12811 = x23 & n12806 ;
  assign n12812 = ( n5306 & n12810 ) | ( n5306 & n12811 ) | ( n12810 & n12811 ) ;
  assign n12813 = x23 & ~n12811 ;
  assign n12814 = x23 & ~n12810 ;
  assign n12815 = ( ~n5306 & n12813 ) | ( ~n5306 & n12814 ) | ( n12813 & n12814 ) ;
  assign n12816 = ( n12809 & ~n12812 ) | ( n12809 & n12815 ) | ( ~n12812 & n12815 ) ;
  assign n12817 = n12799 & ~n12816 ;
  assign n12818 = n12799 | n12816 ;
  assign n12819 = ( ~n12799 & n12817 ) | ( ~n12799 & n12818 ) | ( n12817 & n12818 ) ;
  assign n12820 = n12471 | n12489 ;
  assign n12821 = ( n12471 & ~n12473 ) | ( n12471 & n12820 ) | ( ~n12473 & n12820 ) ;
  assign n12822 = n12819 & n12821 ;
  assign n12823 = n12819 | n12821 ;
  assign n12824 = ~n12822 & n12823 ;
  assign n12825 = n3544 & n5117 ;
  assign n12826 = ( n3544 & ~n5037 ) | ( n3544 & n12825 ) | ( ~n5037 & n12825 ) ;
  assign n12827 = n3541 & n5108 ;
  assign n12828 = n3547 & n5997 ;
  assign n12829 = ( n3547 & n5979 ) | ( n3547 & n12828 ) | ( n5979 & n12828 ) ;
  assign n12830 = n12827 | n12829 ;
  assign n12831 = n12826 | n12830 ;
  assign n12832 = n3537 | n12831 ;
  assign n12833 = ( n6181 & n12831 ) | ( n6181 & n12832 ) | ( n12831 & n12832 ) ;
  assign n12834 = x20 & n12832 ;
  assign n12835 = x20 & n12831 ;
  assign n12836 = ( n6181 & n12834 ) | ( n6181 & n12835 ) | ( n12834 & n12835 ) ;
  assign n12837 = x20 & ~n12834 ;
  assign n12838 = x20 & ~n12835 ;
  assign n12839 = ( ~n6181 & n12837 ) | ( ~n6181 & n12838 ) | ( n12837 & n12838 ) ;
  assign n12840 = ( n12833 & ~n12836 ) | ( n12833 & n12839 ) | ( ~n12836 & n12839 ) ;
  assign n12841 = n12824 & ~n12840 ;
  assign n12842 = n12824 | n12840 ;
  assign n12843 = ( ~n12824 & n12841 ) | ( ~n12824 & n12842 ) | ( n12841 & n12842 ) ;
  assign n12844 = n12493 | n12511 ;
  assign n12845 = ( n12493 & ~n12495 ) | ( n12493 & n12844 ) | ( ~n12495 & n12844 ) ;
  assign n12846 = n12843 & n12845 ;
  assign n12847 = n12843 | n12845 ;
  assign n12848 = ~n12846 & n12847 ;
  assign n12849 = n4466 & n5857 ;
  assign n12850 = ( n4466 & ~n5899 ) | ( n4466 & n12849 ) | ( ~n5899 & n12849 ) ;
  assign n12851 = n4468 & ~n6091 ;
  assign n12852 = n4471 & n7036 ;
  assign n12853 = ( n4471 & n7023 ) | ( n4471 & n12852 ) | ( n7023 & n12852 ) ;
  assign n12854 = n12851 | n12853 ;
  assign n12855 = n12850 | n12854 ;
  assign n12856 = n4475 | n12855 ;
  assign n12857 = ( n7136 & n12855 ) | ( n7136 & n12856 ) | ( n12855 & n12856 ) ;
  assign n12858 = x17 & n12856 ;
  assign n12859 = x17 & n12855 ;
  assign n12860 = ( n7136 & n12858 ) | ( n7136 & n12859 ) | ( n12858 & n12859 ) ;
  assign n12861 = x17 & ~n12858 ;
  assign n12862 = x17 & ~n12859 ;
  assign n12863 = ( ~n7136 & n12861 ) | ( ~n7136 & n12862 ) | ( n12861 & n12862 ) ;
  assign n12864 = ( n12857 & ~n12860 ) | ( n12857 & n12863 ) | ( ~n12860 & n12863 ) ;
  assign n12865 = n12848 & ~n12864 ;
  assign n12866 = n12848 | n12864 ;
  assign n12867 = ( ~n12848 & n12865 ) | ( ~n12848 & n12866 ) | ( n12865 & n12866 ) ;
  assign n12868 = n12518 | n12537 ;
  assign n12869 = ( n12518 & ~n12521 ) | ( n12518 & n12868 ) | ( ~n12521 & n12868 ) ;
  assign n12870 = n12867 & n12869 ;
  assign n12871 = n12867 | n12869 ;
  assign n12872 = ~n12870 & n12871 ;
  assign n12873 = n5237 & n6950 ;
  assign n12874 = n5231 & n6889 ;
  assign n12875 = ( n5231 & ~n6884 ) | ( n5231 & n12874 ) | ( ~n6884 & n12874 ) ;
  assign n12876 = n12873 | n12875 ;
  assign n12877 = n5234 & n7907 ;
  assign n12878 = ( n5234 & n7902 ) | ( n5234 & n12877 ) | ( n7902 & n12877 ) ;
  assign n12879 = n12876 | n12878 ;
  assign n12880 = n5227 | n12878 ;
  assign n12881 = n12876 | n12880 ;
  assign n12882 = ( ~n8193 & n12879 ) | ( ~n8193 & n12881 ) | ( n12879 & n12881 ) ;
  assign n12883 = ~x14 & n12881 ;
  assign n12884 = ~x14 & n12879 ;
  assign n12885 = ( ~n8193 & n12883 ) | ( ~n8193 & n12884 ) | ( n12883 & n12884 ) ;
  assign n12886 = x14 | n12884 ;
  assign n12887 = x14 | n12883 ;
  assign n12888 = ( ~n8193 & n12886 ) | ( ~n8193 & n12887 ) | ( n12886 & n12887 ) ;
  assign n12889 = ( ~n12882 & n12885 ) | ( ~n12882 & n12888 ) | ( n12885 & n12888 ) ;
  assign n12890 = n12872 & n12889 ;
  assign n12891 = n12872 & ~n12890 ;
  assign n12893 = n12544 | n12564 ;
  assign n12894 = ( n12544 & ~n12547 ) | ( n12544 & n12893 ) | ( ~n12547 & n12893 ) ;
  assign n12892 = ~n12872 & n12889 ;
  assign n12895 = n12892 & n12894 ;
  assign n12896 = ( n12891 & n12894 ) | ( n12891 & n12895 ) | ( n12894 & n12895 ) ;
  assign n12897 = n12892 | n12894 ;
  assign n12898 = n12891 | n12897 ;
  assign n12899 = ~n12896 & n12898 ;
  assign n12900 = n6125 & n8079 ;
  assign n12901 = ( n6125 & ~n8070 ) | ( n6125 & n12900 ) | ( ~n8070 & n12900 ) ;
  assign n12902 = n6119 | n12901 ;
  assign n12903 = ( ~n8017 & n12901 ) | ( ~n8017 & n12902 ) | ( n12901 & n12902 ) ;
  assign n12904 = n6122 & n9022 ;
  assign n12905 = ( n6122 & ~n9019 ) | ( n6122 & n12904 ) | ( ~n9019 & n12904 ) ;
  assign n12906 = n12903 | n12905 ;
  assign n12907 = n6115 | n12905 ;
  assign n12908 = n12903 | n12907 ;
  assign n12909 = ( ~n9416 & n12906 ) | ( ~n9416 & n12908 ) | ( n12906 & n12908 ) ;
  assign n12910 = ~x11 & n12908 ;
  assign n12911 = ~x11 & n12906 ;
  assign n12912 = ( ~n9416 & n12910 ) | ( ~n9416 & n12911 ) | ( n12910 & n12911 ) ;
  assign n12913 = x11 | n12911 ;
  assign n12914 = x11 | n12910 ;
  assign n12915 = ( ~n9416 & n12913 ) | ( ~n9416 & n12914 ) | ( n12913 & n12914 ) ;
  assign n12916 = ( ~n12909 & n12912 ) | ( ~n12909 & n12915 ) | ( n12912 & n12915 ) ;
  assign n12917 = n12899 & ~n12916 ;
  assign n12918 = n12899 | n12916 ;
  assign n12919 = ( ~n12899 & n12917 ) | ( ~n12899 & n12918 ) | ( n12917 & n12918 ) ;
  assign n12920 = n12672 & ~n12919 ;
  assign n12921 = n12672 | n12919 ;
  assign n12922 = ( ~n12672 & n12920 ) | ( ~n12672 & n12921 ) | ( n12920 & n12921 ) ;
  assign n12923 = ~n12336 & n12592 ;
  assign n12924 = ( n12336 & n12338 ) | ( n12336 & ~n12923 ) | ( n12338 & ~n12923 ) ;
  assign n12925 = n12922 & n12924 ;
  assign n12926 = n12922 | n12924 ;
  assign n12927 = ~n12925 & n12926 ;
  assign n12928 = n12597 | n12606 ;
  assign n12929 = n12927 & n12928 ;
  assign n12930 = n12597 | n12607 ;
  assign n12931 = n12927 & n12930 ;
  assign n12932 = ( n11360 & n12929 ) | ( n11360 & n12931 ) | ( n12929 & n12931 ) ;
  assign n12933 = n12927 | n12928 ;
  assign n12934 = n12927 | n12930 ;
  assign n12935 = ( n11360 & n12933 ) | ( n11360 & n12934 ) | ( n12933 & n12934 ) ;
  assign n12936 = ~n12932 & n12935 ;
  assign n12937 = n6122 & ~n8982 ;
  assign n12938 = ( n6122 & n9051 ) | ( n6122 & n12937 ) | ( n9051 & n12937 ) ;
  assign n12939 = n6119 & n9022 ;
  assign n12940 = n12938 | n12939 ;
  assign n12941 = n6119 | n12938 ;
  assign n12942 = ( ~n9019 & n12940 ) | ( ~n9019 & n12941 ) | ( n12940 & n12941 ) ;
  assign n12943 = n6125 | n12942 ;
  assign n12944 = ( ~n8017 & n12942 ) | ( ~n8017 & n12943 ) | ( n12942 & n12943 ) ;
  assign n12945 = n6115 | n12944 ;
  assign n12946 = ( ~n10242 & n12944 ) | ( ~n10242 & n12945 ) | ( n12944 & n12945 ) ;
  assign n12947 = ~x11 & n12945 ;
  assign n12948 = ~x11 & n12944 ;
  assign n12949 = ( ~n10242 & n12947 ) | ( ~n10242 & n12948 ) | ( n12947 & n12948 ) ;
  assign n12950 = x11 | n12947 ;
  assign n12951 = x11 | n12948 ;
  assign n12952 = ( ~n10242 & n12950 ) | ( ~n10242 & n12951 ) | ( n12950 & n12951 ) ;
  assign n12953 = ( ~n12946 & n12949 ) | ( ~n12946 & n12952 ) | ( n12949 & n12952 ) ;
  assign n12954 = n12896 | n12916 ;
  assign n12955 = ( n12896 & n12899 ) | ( n12896 & n12954 ) | ( n12899 & n12954 ) ;
  assign n12956 = n12953 & n12955 ;
  assign n12957 = n12953 | n12955 ;
  assign n12958 = ~n12956 & n12957 ;
  assign n12959 = n233 | n517 ;
  assign n12960 = n296 | n476 ;
  assign n12961 = n2156 | n12960 ;
  assign n12962 = n12959 | n12961 ;
  assign n12963 = n182 | n610 ;
  assign n12964 = n12962 | n12963 ;
  assign n12965 = n10884 | n12964 ;
  assign n12966 = n1028 | n12965 ;
  assign n12967 = n234 | n9130 ;
  assign n12968 = n7013 | n10893 ;
  assign n12969 = n1287 | n12968 ;
  assign n12970 = n12967 | n12969 ;
  assign n12971 = n85 | n202 ;
  assign n12972 = n163 | n590 ;
  assign n12973 = n12971 | n12972 ;
  assign n12974 = n222 | n383 ;
  assign n12975 = n134 | n12974 ;
  assign n12976 = n12973 | n12975 ;
  assign n12977 = n324 | n758 ;
  assign n12978 = n3376 | n12977 ;
  assign n12979 = n12976 | n12978 ;
  assign n12980 = n888 | n1607 ;
  assign n12981 = n1016 | n2053 ;
  assign n12982 = n12980 | n12981 ;
  assign n12983 = n295 | n312 ;
  assign n12984 = n12982 | n12983 ;
  assign n12985 = n12979 | n12984 ;
  assign n12986 = n12970 | n12985 ;
  assign n12987 = n12966 | n12986 ;
  assign n12988 = n210 | n3465 ;
  assign n12989 = n382 | n4184 ;
  assign n12990 = n12988 | n12989 ;
  assign n12991 = n237 | n600 ;
  assign n12992 = n689 | n12991 ;
  assign n12993 = n460 | n643 ;
  assign n12994 = n313 | n355 ;
  assign n12995 = n12993 | n12994 ;
  assign n12996 = n12992 | n12995 ;
  assign n12997 = n12990 | n12996 ;
  assign n12998 = n3445 | n3986 ;
  assign n12999 = n5092 | n12998 ;
  assign n13000 = n12997 | n12999 ;
  assign n13001 = n12987 | n13000 ;
  assign n13002 = n1005 | n1349 ;
  assign n13003 = n566 | n13002 ;
  assign n13004 = n370 | n375 ;
  assign n13005 = n282 | n13004 ;
  assign n13006 = n1081 | n13005 ;
  assign n13007 = n13003 | n13006 ;
  assign n13008 = n12681 | n13007 ;
  assign n13009 = n80 | n7880 ;
  assign n13010 = n228 | n411 ;
  assign n13011 = n13009 | n13010 ;
  assign n13012 = n309 | n895 ;
  assign n13013 = n110 | n13012 ;
  assign n13014 = n384 | n735 ;
  assign n13015 = n9140 | n13014 ;
  assign n13016 = n13013 | n13015 ;
  assign n13017 = n13011 | n13016 ;
  assign n13018 = n551 | n1723 ;
  assign n13019 = n5183 | n13018 ;
  assign n13020 = n259 | n3495 ;
  assign n13021 = n13019 | n13020 ;
  assign n13022 = n13017 | n13021 ;
  assign n13023 = n13008 | n13022 ;
  assign n13024 = n117 | n806 ;
  assign n13025 = ( n801 & ~n4245 ) | ( n801 & n13024 ) | ( ~n4245 & n13024 ) ;
  assign n13026 = n212 | n4245 ;
  assign n13027 = n13025 | n13026 ;
  assign n13028 = n1171 | n13027 ;
  assign n13029 = n13023 | n13028 ;
  assign n13030 = n162 | n720 ;
  assign n13031 = n133 | n262 ;
  assign n13032 = n13030 | n13031 ;
  assign n13033 = n310 | n354 ;
  assign n13034 = n13032 | n13033 ;
  assign n13035 = n13029 | n13034 ;
  assign n13036 = n13001 | n13035 ;
  assign n13037 = n12408 & ~n13036 ;
  assign n13038 = ( x8 & n12408 ) | ( x8 & ~n13036 ) | ( n12408 & ~n13036 ) ;
  assign n13039 = ~n13037 & n13038 ;
  assign n13040 = ~n12408 & n13036 ;
  assign n13041 = n13037 | n13040 ;
  assign n13042 = ~x8 & n13041 ;
  assign n13043 = n13039 | n13042 ;
  assign n13044 = n12726 & n13043 ;
  assign n13045 = n12728 & n13043 ;
  assign n13046 = ( n2985 & n13044 ) | ( n2985 & n13045 ) | ( n13044 & n13045 ) ;
  assign n13047 = n12726 | n13043 ;
  assign n13048 = n12728 | n13043 ;
  assign n13049 = ( n2985 & n13047 ) | ( n2985 & n13048 ) | ( n13047 & n13048 ) ;
  assign n13050 = ~n13046 & n13049 ;
  assign n13051 = n1060 & n2691 ;
  assign n13052 = ( n1060 & n2678 ) | ( n1060 & n13051 ) | ( n2678 & n13051 ) ;
  assign n13053 = n1065 & n2701 ;
  assign n13054 = ( n1065 & ~n2784 ) | ( n1065 & n13053 ) | ( ~n2784 & n13053 ) ;
  assign n13055 = n13052 | n13054 ;
  assign n13056 = n1057 & n2893 ;
  assign n13057 = ( n1057 & ~n2886 ) | ( n1057 & n13056 ) | ( ~n2886 & n13056 ) ;
  assign n13058 = n13055 | n13057 ;
  assign n13059 = n1062 | n13058 ;
  assign n13060 = ( ~n2914 & n13058 ) | ( ~n2914 & n13059 ) | ( n13058 & n13059 ) ;
  assign n13061 = ~n13050 & n13060 ;
  assign n13062 = n13050 & ~n13060 ;
  assign n13063 = n13061 | n13062 ;
  assign n13064 = n1823 & n3386 ;
  assign n13065 = n1826 & n3507 ;
  assign n13066 = ( n1826 & n3483 ) | ( n1826 & n13065 ) | ( n3483 & n13065 ) ;
  assign n13067 = n1829 & n3439 ;
  assign n13068 = ( n1829 & ~n3420 ) | ( n1829 & n13067 ) | ( ~n3420 & n13067 ) ;
  assign n13069 = n13066 | n13068 ;
  assign n13070 = n13064 | n13069 ;
  assign n13071 = n1821 | n13070 ;
  assign n13072 = ( ~n3530 & n13070 ) | ( ~n3530 & n13071 ) | ( n13070 & n13071 ) ;
  assign n13073 = ~x29 & n13071 ;
  assign n13074 = ~x29 & n13070 ;
  assign n13075 = ( ~n3530 & n13073 ) | ( ~n3530 & n13074 ) | ( n13073 & n13074 ) ;
  assign n13076 = x29 | n13073 ;
  assign n13077 = x29 | n13074 ;
  assign n13078 = ( ~n3530 & n13076 ) | ( ~n3530 & n13077 ) | ( n13076 & n13077 ) ;
  assign n13079 = ( ~n13072 & n13075 ) | ( ~n13072 & n13078 ) | ( n13075 & n13078 ) ;
  assign n13080 = n13063 & n13079 ;
  assign n13081 = n13063 & ~n13080 ;
  assign n13082 = ~n13063 & n13079 ;
  assign n13083 = n13081 | n13082 ;
  assign n13084 = n12744 | n12751 ;
  assign n13085 = n13083 & n13084 ;
  assign n13086 = n13083 | n13084 ;
  assign n13087 = ~n13085 & n13086 ;
  assign n13088 = n2308 & ~n4429 ;
  assign n13089 = n2308 | n2312 ;
  assign n13090 = ( n2312 & ~n4429 ) | ( n2312 & n13089 ) | ( ~n4429 & n13089 ) ;
  assign n13091 = ( n4206 & n13088 ) | ( n4206 & n13090 ) | ( n13088 & n13090 ) ;
  assign n13092 = n2315 & n4396 ;
  assign n13094 = n2306 | n13092 ;
  assign n13095 = n13091 | n13094 ;
  assign n13093 = n13091 | n13092 ;
  assign n13096 = n13093 & n13095 ;
  assign n13097 = ( ~n4501 & n13095 ) | ( ~n4501 & n13096 ) | ( n13095 & n13096 ) ;
  assign n13098 = ~x26 & n13096 ;
  assign n13099 = ~x26 & n13095 ;
  assign n13100 = ( ~n4501 & n13098 ) | ( ~n4501 & n13099 ) | ( n13098 & n13099 ) ;
  assign n13101 = x26 | n13098 ;
  assign n13102 = x26 | n13099 ;
  assign n13103 = ( ~n4501 & n13101 ) | ( ~n4501 & n13102 ) | ( n13101 & n13102 ) ;
  assign n13104 = ( ~n13097 & n13100 ) | ( ~n13097 & n13103 ) | ( n13100 & n13103 ) ;
  assign n13105 = n13087 & n13104 ;
  assign n13106 = n13087 | n13104 ;
  assign n13107 = ~n13105 & n13106 ;
  assign n13108 = n12773 | n12791 ;
  assign n13109 = ( n12773 & n12775 ) | ( n12773 & n13108 ) | ( n12775 & n13108 ) ;
  assign n13110 = n13107 & n13109 ;
  assign n13111 = n13107 | n13109 ;
  assign n13112 = ~n13110 & n13111 ;
  assign n13113 = n2925 & n4245 ;
  assign n13114 = ( n2925 & n4303 ) | ( n2925 & n13113 ) | ( n4303 & n13113 ) ;
  assign n13115 = n2928 & n5192 ;
  assign n13116 = ( n2928 & n5179 ) | ( n2928 & n13115 ) | ( n5179 & n13115 ) ;
  assign n13117 = n13114 | n13116 ;
  assign n13118 = n2932 & n5117 ;
  assign n13119 = ( n2932 & ~n5037 ) | ( n2932 & n13118 ) | ( ~n5037 & n13118 ) ;
  assign n13120 = n13117 | n13119 ;
  assign n13121 = n2936 | n13119 ;
  assign n13122 = n13117 | n13121 ;
  assign n13123 = ( ~n5270 & n13120 ) | ( ~n5270 & n13122 ) | ( n13120 & n13122 ) ;
  assign n13124 = ~x23 & n13122 ;
  assign n13125 = ~x23 & n13120 ;
  assign n13126 = ( ~n5270 & n13124 ) | ( ~n5270 & n13125 ) | ( n13124 & n13125 ) ;
  assign n13127 = x23 | n13125 ;
  assign n13128 = x23 | n13124 ;
  assign n13129 = ( ~n5270 & n13127 ) | ( ~n5270 & n13128 ) | ( n13127 & n13128 ) ;
  assign n13130 = ( ~n13123 & n13126 ) | ( ~n13123 & n13129 ) | ( n13126 & n13129 ) ;
  assign n13131 = n13112 & n13130 ;
  assign n13132 = ~n13112 & n13130 ;
  assign n13133 = ( n13112 & ~n13131 ) | ( n13112 & n13132 ) | ( ~n13131 & n13132 ) ;
  assign n13134 = n12797 | n12816 ;
  assign n13135 = ( n12797 & n12799 ) | ( n12797 & n13134 ) | ( n12799 & n13134 ) ;
  assign n13136 = n13133 & n13135 ;
  assign n13137 = n13133 | n13135 ;
  assign n13138 = ~n13136 & n13137 ;
  assign n13139 = n3544 & n5108 ;
  assign n13140 = n3541 & n5997 ;
  assign n13141 = ( n3541 & n5979 ) | ( n3541 & n13140 ) | ( n5979 & n13140 ) ;
  assign n13142 = n13139 | n13141 ;
  assign n13143 = n3547 & n5857 ;
  assign n13144 = ( n3547 & ~n5899 ) | ( n3547 & n13143 ) | ( ~n5899 & n13143 ) ;
  assign n13145 = n13142 | n13144 ;
  assign n13146 = n3537 | n13145 ;
  assign n13147 = n13145 & n13146 ;
  assign n13148 = ( ~n6151 & n13146 ) | ( ~n6151 & n13147 ) | ( n13146 & n13147 ) ;
  assign n13149 = ~x20 & n13147 ;
  assign n13150 = ~x20 & n13146 ;
  assign n13151 = ( ~n6151 & n13149 ) | ( ~n6151 & n13150 ) | ( n13149 & n13150 ) ;
  assign n13152 = x20 | n13149 ;
  assign n13153 = x20 | n13150 ;
  assign n13154 = ( ~n6151 & n13152 ) | ( ~n6151 & n13153 ) | ( n13152 & n13153 ) ;
  assign n13155 = ( ~n13148 & n13151 ) | ( ~n13148 & n13154 ) | ( n13151 & n13154 ) ;
  assign n13156 = n13138 & n13155 ;
  assign n13157 = n13138 | n13155 ;
  assign n13158 = ~n13156 & n13157 ;
  assign n13159 = n12822 | n12840 ;
  assign n13160 = ( n12822 & n12824 ) | ( n12822 & n13159 ) | ( n12824 & n13159 ) ;
  assign n13161 = n13158 & n13160 ;
  assign n13162 = n13158 | n13160 ;
  assign n13163 = ~n13161 & n13162 ;
  assign n13164 = n4466 & ~n6091 ;
  assign n13165 = n4468 & n7036 ;
  assign n13166 = ( n4468 & n7023 ) | ( n4468 & n13165 ) | ( n7023 & n13165 ) ;
  assign n13167 = n13164 | n13166 ;
  assign n13168 = n4471 & n6950 ;
  assign n13169 = n13167 | n13168 ;
  assign n13170 = n4475 | n13169 ;
  assign n13171 = ( ~n7107 & n13169 ) | ( ~n7107 & n13170 ) | ( n13169 & n13170 ) ;
  assign n13172 = ~x17 & n13170 ;
  assign n13173 = ~x17 & n13169 ;
  assign n13174 = ( ~n7107 & n13172 ) | ( ~n7107 & n13173 ) | ( n13172 & n13173 ) ;
  assign n13175 = x17 | n13172 ;
  assign n13176 = x17 | n13173 ;
  assign n13177 = ( ~n7107 & n13175 ) | ( ~n7107 & n13176 ) | ( n13175 & n13176 ) ;
  assign n13178 = ( ~n13171 & n13174 ) | ( ~n13171 & n13177 ) | ( n13174 & n13177 ) ;
  assign n13179 = n13163 & n13178 ;
  assign n13180 = ~n13163 & n13178 ;
  assign n13181 = ( n13163 & ~n13179 ) | ( n13163 & n13180 ) | ( ~n13179 & n13180 ) ;
  assign n13182 = n12846 | n12864 ;
  assign n13183 = ( n12846 & n12848 ) | ( n12846 & n13182 ) | ( n12848 & n13182 ) ;
  assign n13184 = n13181 & n13183 ;
  assign n13185 = n13181 | n13183 ;
  assign n13186 = ~n13184 & n13185 ;
  assign n13187 = n5237 & n6889 ;
  assign n13188 = ( n5237 & ~n6884 ) | ( n5237 & n13187 ) | ( ~n6884 & n13187 ) ;
  assign n13189 = n5231 & n7907 ;
  assign n13190 = ( n5231 & n7902 ) | ( n5231 & n13189 ) | ( n7902 & n13189 ) ;
  assign n13191 = n5234 & n8079 ;
  assign n13192 = ( n5234 & ~n8070 ) | ( n5234 & n13191 ) | ( ~n8070 & n13191 ) ;
  assign n13193 = n13190 | n13192 ;
  assign n13194 = n13188 | n13193 ;
  assign n13195 = n5227 | n13194 ;
  assign n13196 = n13194 & n13195 ;
  assign n13197 = ( ~n8156 & n13195 ) | ( ~n8156 & n13196 ) | ( n13195 & n13196 ) ;
  assign n13198 = ~x14 & n13196 ;
  assign n13199 = ~x14 & n13195 ;
  assign n13200 = ( ~n8156 & n13198 ) | ( ~n8156 & n13199 ) | ( n13198 & n13199 ) ;
  assign n13201 = x14 | n13198 ;
  assign n13202 = x14 | n13199 ;
  assign n13203 = ( ~n8156 & n13201 ) | ( ~n8156 & n13202 ) | ( n13201 & n13202 ) ;
  assign n13204 = ( ~n13197 & n13200 ) | ( ~n13197 & n13203 ) | ( n13200 & n13203 ) ;
  assign n13205 = n13186 & n13204 ;
  assign n13206 = n13186 & ~n13205 ;
  assign n13207 = ~n13186 & n13204 ;
  assign n13208 = n13206 | n13207 ;
  assign n13209 = n12870 | n12889 ;
  assign n13210 = ( n12870 & n12872 ) | ( n12870 & n13209 ) | ( n12872 & n13209 ) ;
  assign n13211 = n13208 & n13210 ;
  assign n13212 = n13208 & ~n13211 ;
  assign n13213 = ~n13208 & n13210 ;
  assign n13214 = n13212 | n13213 ;
  assign n13215 = ~n12958 & n13214 ;
  assign n13216 = n12958 & ~n13214 ;
  assign n13217 = n13215 | n13216 ;
  assign n13218 = n12670 | n12919 ;
  assign n13219 = ( n12670 & n12672 ) | ( n12670 & n13218 ) | ( n12672 & n13218 ) ;
  assign n13220 = n13217 & n13219 ;
  assign n13221 = n13217 | n13219 ;
  assign n13222 = ~n13220 & n13221 ;
  assign n13223 = n12922 & n13222 ;
  assign n13224 = n12924 & n13223 ;
  assign n13225 = ( n12927 & n13222 ) | ( n12927 & n13224 ) | ( n13222 & n13224 ) ;
  assign n13226 = ( n12928 & n13224 ) | ( n12928 & n13225 ) | ( n13224 & n13225 ) ;
  assign n13227 = ( n12930 & n13224 ) | ( n12930 & n13225 ) | ( n13224 & n13225 ) ;
  assign n13228 = ( n11360 & n13226 ) | ( n11360 & n13227 ) | ( n13226 & n13227 ) ;
  assign n13229 = n12925 | n12927 ;
  assign n13230 = ( n12925 & n12930 ) | ( n12925 & n13229 ) | ( n12930 & n13229 ) ;
  assign n13231 = n13222 | n13230 ;
  assign n13232 = ( n12925 & n12928 ) | ( n12925 & n13229 ) | ( n12928 & n13229 ) ;
  assign n13233 = n13222 | n13232 ;
  assign n13234 = ( n11360 & n13231 ) | ( n11360 & n13233 ) | ( n13231 & n13233 ) ;
  assign n13235 = ~n13228 & n13234 ;
  assign n13236 = n12936 & n13235 ;
  assign n13237 = n12936 | n13235 ;
  assign n13238 = ~n13236 & n13237 ;
  assign n13239 = n13236 | n13238 ;
  assign n13240 = ~n12617 & n12619 ;
  assign n13241 = ~n12616 & n12936 ;
  assign n13242 = n12616 & ~n12936 ;
  assign n13243 = n13241 | n13242 ;
  assign n13244 = n13240 | n13243 ;
  assign n13245 = n12617 & ~n13243 ;
  assign n13246 = ( n12026 & ~n13244 ) | ( n12026 & n13245 ) | ( ~n13244 & n13245 ) ;
  assign n13247 = ( n12012 & n13244 ) | ( n12012 & ~n13245 ) | ( n13244 & ~n13245 ) ;
  assign n13248 = ( n11672 & n13246 ) | ( n11672 & ~n13247 ) | ( n13246 & ~n13247 ) ;
  assign n13249 = n13236 | n13241 ;
  assign n13250 = ( n13236 & n13238 ) | ( n13236 & n13249 ) | ( n13238 & n13249 ) ;
  assign n13251 = ( n13239 & n13248 ) | ( n13239 & n13250 ) | ( n13248 & n13250 ) ;
  assign n13252 = n6119 & ~n8982 ;
  assign n13253 = ( n6119 & n9051 ) | ( n6119 & n13252 ) | ( n9051 & n13252 ) ;
  assign n13254 = n6125 & ~n9022 ;
  assign n13255 = ( n6125 & n13253 ) | ( n6125 & ~n13254 ) | ( n13253 & ~n13254 ) ;
  assign n13256 = n6125 | n13253 ;
  assign n13257 = ( ~n9019 & n13255 ) | ( ~n9019 & n13256 ) | ( n13255 & n13256 ) ;
  assign n13258 = n6115 | n13257 ;
  assign n13259 = ( n9078 & n13257 ) | ( n9078 & n13258 ) | ( n13257 & n13258 ) ;
  assign n13260 = x11 & n13258 ;
  assign n13261 = x11 & n13257 ;
  assign n13262 = ( n9078 & n13260 ) | ( n9078 & n13261 ) | ( n13260 & n13261 ) ;
  assign n13263 = x11 & ~n13260 ;
  assign n13264 = x11 & ~n13261 ;
  assign n13265 = ( ~n9078 & n13263 ) | ( ~n9078 & n13264 ) | ( n13263 & n13264 ) ;
  assign n13266 = ( n13259 & ~n13262 ) | ( n13259 & n13265 ) | ( ~n13262 & n13265 ) ;
  assign n13267 = n13204 & n13266 ;
  assign n13268 = n13186 & n13267 ;
  assign n13269 = ( n13210 & n13266 ) | ( n13210 & n13268 ) | ( n13266 & n13268 ) ;
  assign n13270 = n13266 & n13268 ;
  assign n13271 = ( n13208 & n13269 ) | ( n13208 & n13270 ) | ( n13269 & n13270 ) ;
  assign n13272 = n13204 | n13266 ;
  assign n13273 = ( n13186 & n13266 ) | ( n13186 & n13272 ) | ( n13266 & n13272 ) ;
  assign n13274 = n13210 | n13273 ;
  assign n13275 = ( n13208 & n13273 ) | ( n13208 & n13274 ) | ( n13273 & n13274 ) ;
  assign n13276 = ~n13271 & n13275 ;
  assign n13277 = n13156 | n13161 ;
  assign n13278 = n1065 & n2893 ;
  assign n13279 = ( n1065 & ~n2886 ) | ( n1065 & n13278 ) | ( ~n2886 & n13278 ) ;
  assign n13280 = n1060 & n2701 ;
  assign n13281 = ( n1060 & ~n2784 ) | ( n1060 & n13280 ) | ( ~n2784 & n13280 ) ;
  assign n13282 = n1057 & n3507 ;
  assign n13283 = ( n1057 & n3483 ) | ( n1057 & n13282 ) | ( n3483 & n13282 ) ;
  assign n13284 = n13281 | n13283 ;
  assign n13285 = n13279 | n13284 ;
  assign n13286 = n1062 | n13285 ;
  assign n13287 = ( n3603 & n13285 ) | ( n3603 & n13286 ) | ( n13285 & n13286 ) ;
  assign n13288 = n270 | n321 ;
  assign n13289 = n498 | n682 ;
  assign n13290 = n261 | n749 ;
  assign n13291 = n13289 | n13290 ;
  assign n13292 = n370 | n694 ;
  assign n13293 = n273 | n13292 ;
  assign n13294 = n152 | n503 ;
  assign n13295 = n325 | n13294 ;
  assign n13296 = n13293 | n13295 ;
  assign n13297 = n13291 | n13296 ;
  assign n13298 = n13288 | n13297 ;
  assign n13299 = n3469 | n3471 ;
  assign n13300 = n139 | n959 ;
  assign n13301 = n487 | n13300 ;
  assign n13302 = n606 | n923 ;
  assign n13303 = n13301 | n13302 ;
  assign n13304 = n461 | n477 ;
  assign n13305 = n197 | n13304 ;
  assign n13306 = n13303 | n13305 ;
  assign n13307 = n13299 | n13306 ;
  assign n13308 = n13298 | n13307 ;
  assign n13309 = n6028 | n13308 ;
  assign n13310 = n67 | n560 ;
  assign n13311 = n9151 | n13310 ;
  assign n13312 = n793 | n13311 ;
  assign n13313 = n1398 | n6827 ;
  assign n13314 = n1035 | n13313 ;
  assign n13315 = n13312 | n13314 ;
  assign n13316 = n313 | n696 ;
  assign n13317 = n967 | n13316 ;
  assign n13318 = n141 | n13317 ;
  assign n13319 = n302 | n374 ;
  assign n13320 = n13318 | n13319 ;
  assign n13321 = n13315 | n13320 ;
  assign n13322 = n228 | n249 ;
  assign n13323 = n929 | n13322 ;
  assign n13324 = n118 | n395 ;
  assign n13325 = n184 | n13324 ;
  assign n13326 = n13323 | n13325 ;
  assign n13327 = n333 | n13326 ;
  assign n13328 = n2623 | n2753 ;
  assign n13329 = n660 | n4028 ;
  assign n13330 = n13328 | n13329 ;
  assign n13331 = n13327 | n13330 ;
  assign n13332 = n53 | n288 ;
  assign n13333 = n12387 | n13332 ;
  assign n13334 = n94 | n720 ;
  assign n13335 = n13333 | n13334 ;
  assign n13336 = n239 | n320 ;
  assign n13337 = n182 | n306 ;
  assign n13338 = n13336 | n13337 ;
  assign n13339 = n13335 | n13338 ;
  assign n13340 = n13331 | n13339 ;
  assign n13341 = n13321 | n13340 ;
  assign n13342 = n13309 | n13341 ;
  assign n13343 = n457 | n638 ;
  assign n13344 = n280 | n624 ;
  assign n13345 = n13343 | n13344 ;
  assign n13346 = n13342 | n13345 ;
  assign n13347 = n13038 | n13346 ;
  assign n13348 = n13038 & n13346 ;
  assign n13349 = n13347 & ~n13348 ;
  assign n13350 = n13286 & n13349 ;
  assign n13351 = n13285 & n13349 ;
  assign n13352 = ( n3603 & n13350 ) | ( n3603 & n13351 ) | ( n13350 & n13351 ) ;
  assign n13353 = n13349 & ~n13351 ;
  assign n13354 = n13349 & ~n13350 ;
  assign n13355 = ( ~n3603 & n13353 ) | ( ~n3603 & n13354 ) | ( n13353 & n13354 ) ;
  assign n13356 = ( n13287 & ~n13352 ) | ( n13287 & n13355 ) | ( ~n13352 & n13355 ) ;
  assign n13357 = n13046 | n13060 ;
  assign n13358 = ( n13046 & n13050 ) | ( n13046 & n13357 ) | ( n13050 & n13357 ) ;
  assign n13359 = n13356 & n13358 ;
  assign n13360 = n13356 | n13358 ;
  assign n13361 = ~n13359 & n13360 ;
  assign n13362 = n1829 & n4206 ;
  assign n13363 = n1826 & n3386 ;
  assign n13364 = n1823 & n3439 ;
  assign n13365 = ( n1823 & ~n3420 ) | ( n1823 & n13364 ) | ( ~n3420 & n13364 ) ;
  assign n13366 = n13363 | n13365 ;
  assign n13367 = n13362 | n13366 ;
  assign n13368 = n1821 | n13362 ;
  assign n13369 = n13366 | n13368 ;
  assign n13370 = ( ~n4220 & n13367 ) | ( ~n4220 & n13369 ) | ( n13367 & n13369 ) ;
  assign n13371 = ~x29 & n13369 ;
  assign n13372 = ~x29 & n13367 ;
  assign n13373 = ( ~n4220 & n13371 ) | ( ~n4220 & n13372 ) | ( n13371 & n13372 ) ;
  assign n13374 = x29 | n13372 ;
  assign n13375 = x29 | n13371 ;
  assign n13376 = ( ~n4220 & n13374 ) | ( ~n4220 & n13375 ) | ( n13374 & n13375 ) ;
  assign n13377 = ( ~n13370 & n13373 ) | ( ~n13370 & n13376 ) | ( n13373 & n13376 ) ;
  assign n13378 = n13361 & n13377 ;
  assign n13379 = n13361 | n13377 ;
  assign n13380 = ~n13378 & n13379 ;
  assign n13381 = n13080 & n13380 ;
  assign n13382 = ( n13085 & n13380 ) | ( n13085 & n13381 ) | ( n13380 & n13381 ) ;
  assign n13383 = n13080 | n13380 ;
  assign n13384 = n13085 | n13383 ;
  assign n13385 = ~n13382 & n13384 ;
  assign n13386 = n2312 & ~n4429 ;
  assign n13387 = n2308 & n4396 ;
  assign n13388 = n13386 | n13387 ;
  assign n13389 = n2315 & n4245 ;
  assign n13390 = ( n2315 & n4303 ) | ( n2315 & n13389 ) | ( n4303 & n13389 ) ;
  assign n13391 = n13388 | n13390 ;
  assign n13392 = n2306 | n13390 ;
  assign n13393 = n13388 | n13392 ;
  assign n13394 = ( n4455 & n13391 ) | ( n4455 & n13393 ) | ( n13391 & n13393 ) ;
  assign n13395 = x26 & n13393 ;
  assign n13396 = x26 & n13391 ;
  assign n13397 = ( n4455 & n13395 ) | ( n4455 & n13396 ) | ( n13395 & n13396 ) ;
  assign n13398 = x26 & ~n13396 ;
  assign n13399 = x26 & ~n13395 ;
  assign n13400 = ( ~n4455 & n13398 ) | ( ~n4455 & n13399 ) | ( n13398 & n13399 ) ;
  assign n13401 = ( n13394 & ~n13397 ) | ( n13394 & n13400 ) | ( ~n13397 & n13400 ) ;
  assign n13402 = n13385 & ~n13401 ;
  assign n13403 = n13385 | n13401 ;
  assign n13404 = ( ~n13385 & n13402 ) | ( ~n13385 & n13403 ) | ( n13402 & n13403 ) ;
  assign n13405 = n13105 | n13110 ;
  assign n13406 = n13404 & n13405 ;
  assign n13407 = n13404 | n13405 ;
  assign n13408 = ~n13406 & n13407 ;
  assign n13409 = n2928 & n5117 ;
  assign n13410 = ( n2928 & ~n5037 ) | ( n2928 & n13409 ) | ( ~n5037 & n13409 ) ;
  assign n13411 = n2932 & n5108 ;
  assign n13412 = n2925 & n5192 ;
  assign n13413 = ( n2925 & n5179 ) | ( n2925 & n13412 ) | ( n5179 & n13412 ) ;
  assign n13414 = n13411 | n13413 ;
  assign n13415 = n13410 | n13414 ;
  assign n13416 = n2936 | n13415 ;
  assign n13417 = ( ~n5220 & n13415 ) | ( ~n5220 & n13416 ) | ( n13415 & n13416 ) ;
  assign n13418 = ~x23 & n13416 ;
  assign n13419 = ~x23 & n13415 ;
  assign n13420 = ( ~n5220 & n13418 ) | ( ~n5220 & n13419 ) | ( n13418 & n13419 ) ;
  assign n13421 = x23 | n13418 ;
  assign n13422 = x23 | n13419 ;
  assign n13423 = ( ~n5220 & n13421 ) | ( ~n5220 & n13422 ) | ( n13421 & n13422 ) ;
  assign n13424 = ( ~n13417 & n13420 ) | ( ~n13417 & n13423 ) | ( n13420 & n13423 ) ;
  assign n13425 = n13408 & ~n13424 ;
  assign n13426 = n13408 | n13424 ;
  assign n13427 = ( ~n13408 & n13425 ) | ( ~n13408 & n13426 ) | ( n13425 & n13426 ) ;
  assign n13428 = n13131 | n13133 ;
  assign n13429 = ( n13131 & n13135 ) | ( n13131 & n13428 ) | ( n13135 & n13428 ) ;
  assign n13430 = n13427 & n13429 ;
  assign n13431 = n13427 | n13429 ;
  assign n13432 = ~n13430 & n13431 ;
  assign n13433 = n3541 & n5857 ;
  assign n13434 = ( n3541 & ~n5899 ) | ( n3541 & n13433 ) | ( ~n5899 & n13433 ) ;
  assign n13435 = n3547 & ~n6091 ;
  assign n13436 = n3544 & n5997 ;
  assign n13437 = ( n3544 & n5979 ) | ( n3544 & n13436 ) | ( n5979 & n13436 ) ;
  assign n13438 = n13435 | n13437 ;
  assign n13439 = n13434 | n13438 ;
  assign n13440 = n3537 | n13439 ;
  assign n13441 = ( n6108 & n13439 ) | ( n6108 & n13440 ) | ( n13439 & n13440 ) ;
  assign n13442 = x20 & n13440 ;
  assign n13443 = x20 & n13439 ;
  assign n13444 = ( n6108 & n13442 ) | ( n6108 & n13443 ) | ( n13442 & n13443 ) ;
  assign n13445 = x20 & ~n13442 ;
  assign n13446 = x20 & ~n13443 ;
  assign n13447 = ( ~n6108 & n13445 ) | ( ~n6108 & n13446 ) | ( n13445 & n13446 ) ;
  assign n13448 = ( n13441 & ~n13444 ) | ( n13441 & n13447 ) | ( ~n13444 & n13447 ) ;
  assign n13449 = n13432 & ~n13448 ;
  assign n13450 = n13432 | n13448 ;
  assign n13451 = ( ~n13432 & n13449 ) | ( ~n13432 & n13450 ) | ( n13449 & n13450 ) ;
  assign n13452 = n13277 & n13451 ;
  assign n13453 = n13277 | n13451 ;
  assign n13454 = ~n13452 & n13453 ;
  assign n13455 = n4468 & n6950 ;
  assign n13456 = n4466 & n7036 ;
  assign n13457 = ( n4466 & n7023 ) | ( n4466 & n13456 ) | ( n7023 & n13456 ) ;
  assign n13458 = n13455 | n13457 ;
  assign n13459 = n4471 & n6889 ;
  assign n13460 = ( n4471 & ~n6884 ) | ( n4471 & n13459 ) | ( ~n6884 & n13459 ) ;
  assign n13461 = n13458 | n13460 ;
  assign n13462 = n4475 | n13460 ;
  assign n13463 = n13458 | n13462 ;
  assign n13464 = ( ~n7061 & n13461 ) | ( ~n7061 & n13463 ) | ( n13461 & n13463 ) ;
  assign n13465 = ~x17 & n13463 ;
  assign n13466 = ~x17 & n13461 ;
  assign n13467 = ( ~n7061 & n13465 ) | ( ~n7061 & n13466 ) | ( n13465 & n13466 ) ;
  assign n13468 = x17 | n13466 ;
  assign n13469 = x17 | n13465 ;
  assign n13470 = ( ~n7061 & n13468 ) | ( ~n7061 & n13469 ) | ( n13468 & n13469 ) ;
  assign n13471 = ( ~n13464 & n13467 ) | ( ~n13464 & n13470 ) | ( n13467 & n13470 ) ;
  assign n13472 = n13454 & ~n13471 ;
  assign n13473 = n13454 | n13471 ;
  assign n13474 = ( ~n13454 & n13472 ) | ( ~n13454 & n13473 ) | ( n13472 & n13473 ) ;
  assign n13475 = n13179 | n13181 ;
  assign n13476 = ( n13179 & n13183 ) | ( n13179 & n13475 ) | ( n13183 & n13475 ) ;
  assign n13477 = n13474 & n13476 ;
  assign n13478 = n13474 | n13476 ;
  assign n13479 = ~n13477 & n13478 ;
  assign n13480 = n5237 & n7907 ;
  assign n13481 = ( n5237 & n7902 ) | ( n5237 & n13480 ) | ( n7902 & n13480 ) ;
  assign n13482 = n5231 & n8079 ;
  assign n13483 = ( n5231 & ~n8070 ) | ( n5231 & n13482 ) | ( ~n8070 & n13482 ) ;
  assign n13484 = n13481 | n13483 ;
  assign n13485 = n5234 & ~n8017 ;
  assign n13486 = n13484 | n13485 ;
  assign n13487 = n5227 | n13484 ;
  assign n13488 = n13485 | n13487 ;
  assign n13489 = ( n8104 & n13486 ) | ( n8104 & n13488 ) | ( n13486 & n13488 ) ;
  assign n13490 = x14 & n13488 ;
  assign n13491 = x14 & n13486 ;
  assign n13492 = ( n8104 & n13490 ) | ( n8104 & n13491 ) | ( n13490 & n13491 ) ;
  assign n13493 = x14 & ~n13491 ;
  assign n13494 = x14 & ~n13490 ;
  assign n13495 = ( ~n8104 & n13493 ) | ( ~n8104 & n13494 ) | ( n13493 & n13494 ) ;
  assign n13496 = ( n13489 & ~n13492 ) | ( n13489 & n13495 ) | ( ~n13492 & n13495 ) ;
  assign n13497 = n13479 & ~n13496 ;
  assign n13498 = n13479 | n13496 ;
  assign n13499 = ( ~n13479 & n13497 ) | ( ~n13479 & n13498 ) | ( n13497 & n13498 ) ;
  assign n13500 = n13276 & n13499 ;
  assign n13501 = n13276 | n13499 ;
  assign n13502 = ~n13500 & n13501 ;
  assign n13503 = n12956 | n13214 ;
  assign n13504 = ( n12956 & n12958 ) | ( n12956 & n13503 ) | ( n12958 & n13503 ) ;
  assign n13505 = n13502 & n13504 ;
  assign n13506 = n13502 | n13504 ;
  assign n13507 = ~n13505 & n13506 ;
  assign n13508 = n13220 | n13222 ;
  assign n13509 = n13220 | n13223 ;
  assign n13510 = ( n12924 & n13220 ) | ( n12924 & n13509 ) | ( n13220 & n13509 ) ;
  assign n13511 = ( n12927 & n13508 ) | ( n12927 & n13510 ) | ( n13508 & n13510 ) ;
  assign n13512 = n13507 & n13511 ;
  assign n13513 = n13507 & n13510 ;
  assign n13514 = ( n12928 & n13512 ) | ( n12928 & n13513 ) | ( n13512 & n13513 ) ;
  assign n13515 = ( n12930 & n13512 ) | ( n12930 & n13513 ) | ( n13512 & n13513 ) ;
  assign n13516 = ( n11360 & n13514 ) | ( n11360 & n13515 ) | ( n13514 & n13515 ) ;
  assign n13517 = ( n12930 & n13510 ) | ( n12930 & n13511 ) | ( n13510 & n13511 ) ;
  assign n13518 = n13507 | n13517 ;
  assign n13519 = ( n12928 & n13510 ) | ( n12928 & n13511 ) | ( n13510 & n13511 ) ;
  assign n13520 = n13507 | n13519 ;
  assign n13521 = ( n11360 & n13518 ) | ( n11360 & n13520 ) | ( n13518 & n13520 ) ;
  assign n13522 = ~n13516 & n13521 ;
  assign n13523 = n13235 & n13522 ;
  assign n13524 = n13235 | n13522 ;
  assign n13525 = n13239 & n13524 ;
  assign n13526 = ~n13523 & n13525 ;
  assign n13527 = n13250 & n13524 ;
  assign n13528 = ~n13523 & n13527 ;
  assign n13529 = ( n13248 & n13526 ) | ( n13248 & n13528 ) | ( n13526 & n13528 ) ;
  assign n13530 = n13251 & ~n13529 ;
  assign n13531 = n2932 & n13522 ;
  assign n13532 = n2925 & n12936 ;
  assign n13533 = n2928 & n13235 ;
  assign n13534 = n13532 | n13533 ;
  assign n13535 = n13531 | n13534 ;
  assign n13536 = ~n13523 & n13524 ;
  assign n13537 = ~n13527 & n13536 ;
  assign n13538 = n2936 & n13537 ;
  assign n13539 = ~n13525 & n13536 ;
  assign n13540 = n2936 & n13539 ;
  assign n13541 = ( ~n13248 & n13538 ) | ( ~n13248 & n13540 ) | ( n13538 & n13540 ) ;
  assign n13542 = n13535 | n13541 ;
  assign n13543 = n2936 | n13535 ;
  assign n13544 = ( n13530 & n13542 ) | ( n13530 & n13543 ) | ( n13542 & n13543 ) ;
  assign n13545 = x23 | n13544 ;
  assign n13546 = ~x23 & n13544 ;
  assign n13547 = ( ~n13544 & n13545 ) | ( ~n13544 & n13546 ) | ( n13545 & n13546 ) ;
  assign n13548 = ~n12649 & n13547 ;
  assign n13549 = ( n12648 & n13547 ) | ( n12648 & n13548 ) | ( n13547 & n13548 ) ;
  assign n13550 = n12650 | n13549 ;
  assign n13551 = n12649 & n13547 ;
  assign n13552 = ~n12648 & n13551 ;
  assign n13553 = n13550 & ~n13552 ;
  assign n13554 = ~n12218 & n12221 ;
  assign n13555 = n12218 & ~n12221 ;
  assign n13556 = n13554 | n13555 ;
  assign n13557 = n13238 & n13241 ;
  assign n13558 = ( n13238 & n13248 ) | ( n13238 & n13557 ) | ( n13248 & n13557 ) ;
  assign n13559 = n13238 | n13241 ;
  assign n13560 = n13248 | n13559 ;
  assign n13561 = ~n13558 & n13560 ;
  assign n13562 = n2932 & n13235 ;
  assign n13563 = n2925 & ~n12616 ;
  assign n13564 = n2928 & n12936 ;
  assign n13565 = n13563 | n13564 ;
  assign n13566 = n13562 | n13565 ;
  assign n13567 = n2936 | n13562 ;
  assign n13568 = n13565 | n13567 ;
  assign n13569 = ( n13561 & n13566 ) | ( n13561 & n13568 ) | ( n13566 & n13568 ) ;
  assign n13570 = x23 & n13568 ;
  assign n13571 = x23 & n13566 ;
  assign n13572 = ( n13561 & n13570 ) | ( n13561 & n13571 ) | ( n13570 & n13571 ) ;
  assign n13573 = x23 & ~n13571 ;
  assign n13574 = x23 & ~n13570 ;
  assign n13575 = ( ~n13561 & n13573 ) | ( ~n13561 & n13574 ) | ( n13573 & n13574 ) ;
  assign n13576 = ( n13569 & ~n13572 ) | ( n13569 & n13575 ) | ( ~n13572 & n13575 ) ;
  assign n13577 = n13556 & n13576 ;
  assign n13578 = n12213 & ~n12217 ;
  assign n13579 = n12216 | n12217 ;
  assign n13580 = ~n13578 & n13579 ;
  assign n13581 = n2932 & n12936 ;
  assign n13582 = n2925 & n12010 ;
  assign n13583 = n2928 & ~n12616 ;
  assign n13584 = n13582 | n13583 ;
  assign n13585 = n13581 | n13584 ;
  assign n13586 = ( n12012 & ~n12617 ) | ( n12012 & n13240 ) | ( ~n12617 & n13240 ) ;
  assign n13587 = n13243 & n13586 ;
  assign n13588 = ( n12026 & n12617 ) | ( n12026 & ~n13240 ) | ( n12617 & ~n13240 ) ;
  assign n13589 = n13243 & ~n13588 ;
  assign n13590 = ( ~n11672 & n13587 ) | ( ~n11672 & n13589 ) | ( n13587 & n13589 ) ;
  assign n13591 = n13248 | n13590 ;
  assign n13592 = n2936 | n13581 ;
  assign n13593 = n13584 | n13592 ;
  assign n13594 = ( n13585 & ~n13591 ) | ( n13585 & n13593 ) | ( ~n13591 & n13593 ) ;
  assign n13595 = ~x23 & n13593 ;
  assign n13596 = ~x23 & n13585 ;
  assign n13597 = ( ~n13591 & n13595 ) | ( ~n13591 & n13596 ) | ( n13595 & n13596 ) ;
  assign n13598 = x23 | n13596 ;
  assign n13599 = x23 | n13595 ;
  assign n13600 = ( ~n13591 & n13598 ) | ( ~n13591 & n13599 ) | ( n13598 & n13599 ) ;
  assign n13601 = ( ~n13594 & n13597 ) | ( ~n13594 & n13600 ) | ( n13597 & n13600 ) ;
  assign n13602 = ~n13580 & n13601 ;
  assign n13603 = n13580 | n13602 ;
  assign n13604 = n13580 & n13601 ;
  assign n13605 = n13603 & ~n13604 ;
  assign n13606 = n12109 | n12207 ;
  assign n13607 = ~n12212 & n13606 ;
  assign n13608 = n12210 | n12212 ;
  assign n13609 = ~n13607 & n13608 ;
  assign n13610 = n2932 & ~n12616 ;
  assign n13611 = n2925 & ~n11663 ;
  assign n13612 = n2928 & n12010 ;
  assign n13613 = n13611 | n13612 ;
  assign n13614 = n13610 | n13613 ;
  assign n13615 = n2936 | n13610 ;
  assign n13616 = n13613 | n13615 ;
  assign n13617 = ( ~n12626 & n13614 ) | ( ~n12626 & n13616 ) | ( n13614 & n13616 ) ;
  assign n13618 = ~x23 & n13616 ;
  assign n13619 = ~x23 & n13614 ;
  assign n13620 = ( ~n12626 & n13618 ) | ( ~n12626 & n13619 ) | ( n13618 & n13619 ) ;
  assign n13621 = x23 | n13619 ;
  assign n13622 = x23 | n13618 ;
  assign n13623 = ( ~n12626 & n13621 ) | ( ~n12626 & n13622 ) | ( n13621 & n13622 ) ;
  assign n13624 = ( ~n13617 & n13620 ) | ( ~n13617 & n13623 ) | ( n13620 & n13623 ) ;
  assign n13625 = n13609 & n13624 ;
  assign n13626 = n12111 | n12206 ;
  assign n13627 = ~n12207 & n13626 ;
  assign n13629 = n2925 & n11363 ;
  assign n13630 = n2928 & ~n11663 ;
  assign n13631 = n13629 | n13630 ;
  assign n13628 = n2932 & n12010 ;
  assign n13633 = n2936 | n13628 ;
  assign n13634 = n13631 | n13633 ;
  assign n13632 = n13628 | n13631 ;
  assign n13635 = n13632 & n13634 ;
  assign n13636 = ( ~n12028 & n13634 ) | ( ~n12028 & n13635 ) | ( n13634 & n13635 ) ;
  assign n13637 = n13634 | n13635 ;
  assign n13638 = ( n12017 & n13636 ) | ( n12017 & n13637 ) | ( n13636 & n13637 ) ;
  assign n13639 = ~x23 & n13638 ;
  assign n13640 = x23 | n13638 ;
  assign n13641 = ( ~n13638 & n13639 ) | ( ~n13638 & n13640 ) | ( n13639 & n13640 ) ;
  assign n13642 = n13627 & n13641 ;
  assign n13643 = n12133 | n12204 ;
  assign n13644 = ~n12205 & n13643 ;
  assign n13645 = n2925 & n10649 ;
  assign n13646 = n2928 & n11363 ;
  assign n13647 = n13645 | n13646 ;
  assign n13648 = n2932 & ~n11663 ;
  assign n13649 = n2936 | n13648 ;
  assign n13650 = n13647 | n13649 ;
  assign n13651 = n13647 | n13648 ;
  assign n13652 = n12048 & ~n13651 ;
  assign n13653 = ( n11672 & ~n13651 ) | ( n11672 & n13652 ) | ( ~n13651 & n13652 ) ;
  assign n13654 = n13650 & ~n13653 ;
  assign n13655 = ( n12040 & n13650 ) | ( n12040 & n13654 ) | ( n13650 & n13654 ) ;
  assign n13656 = x23 & n13655 ;
  assign n13657 = x23 & ~n13655 ;
  assign n13658 = ( n13655 & ~n13656 ) | ( n13655 & n13657 ) | ( ~n13656 & n13657 ) ;
  assign n13659 = n13644 & n13658 ;
  assign n13660 = n13644 & ~n13659 ;
  assign n13661 = ~n13644 & n13658 ;
  assign n13662 = n13660 | n13661 ;
  assign n13663 = n12200 & n12202 ;
  assign n13664 = n12200 | n12202 ;
  assign n13665 = ~n13663 & n13664 ;
  assign n13666 = n2932 & n11363 ;
  assign n13667 = n2925 & n10325 ;
  assign n13668 = n2928 & n10649 ;
  assign n13669 = n13667 | n13668 ;
  assign n13670 = n13666 | n13669 ;
  assign n13671 = n2936 | n13670 ;
  assign n13672 = ( n12059 & n13670 ) | ( n12059 & n13671 ) | ( n13670 & n13671 ) ;
  assign n13673 = x23 & n13671 ;
  assign n13674 = x23 & n13670 ;
  assign n13675 = ( n12059 & n13673 ) | ( n12059 & n13674 ) | ( n13673 & n13674 ) ;
  assign n13676 = x23 & ~n13673 ;
  assign n13677 = x23 & ~n13674 ;
  assign n13678 = ( ~n12059 & n13676 ) | ( ~n12059 & n13677 ) | ( n13676 & n13677 ) ;
  assign n13679 = ( n13672 & ~n13675 ) | ( n13672 & n13678 ) | ( ~n13675 & n13678 ) ;
  assign n13680 = n13665 & n13679 ;
  assign n13681 = n12187 & n12198 ;
  assign n13682 = n12187 & ~n13681 ;
  assign n13683 = n2932 & n10649 ;
  assign n13684 = n2925 & n10654 ;
  assign n13685 = n2928 & n10325 ;
  assign n13686 = n13684 | n13685 ;
  assign n13687 = n13683 | n13686 ;
  assign n13688 = n2936 | n13683 ;
  assign n13689 = n13686 | n13688 ;
  assign n13690 = ( n10702 & n13687 ) | ( n10702 & n13689 ) | ( n13687 & n13689 ) ;
  assign n13691 = n13687 | n13689 ;
  assign n13692 = ( n10695 & n13690 ) | ( n10695 & n13691 ) | ( n13690 & n13691 ) ;
  assign n13693 = x23 & n13692 ;
  assign n13694 = x23 & ~n13692 ;
  assign n13695 = ( n13692 & ~n13693 ) | ( n13692 & n13694 ) | ( ~n13693 & n13694 ) ;
  assign n13696 = ~n12187 & n12198 ;
  assign n13697 = n13695 & n13696 ;
  assign n13698 = ( n13682 & n13695 ) | ( n13682 & n13697 ) | ( n13695 & n13697 ) ;
  assign n13699 = n13695 | n13696 ;
  assign n13700 = n13682 | n13699 ;
  assign n13701 = ~n13698 & n13700 ;
  assign n13702 = n2932 & n10325 ;
  assign n13703 = n2925 & ~n10662 ;
  assign n13704 = n2928 & n10654 ;
  assign n13705 = n13703 | n13704 ;
  assign n13706 = n13702 | n13705 ;
  assign n13707 = n2936 | n13706 ;
  assign n13708 = ( ~n10957 & n13706 ) | ( ~n10957 & n13707 ) | ( n13706 & n13707 ) ;
  assign n13709 = n13706 | n13707 ;
  assign n13710 = ( n10949 & n13708 ) | ( n10949 & n13709 ) | ( n13708 & n13709 ) ;
  assign n13711 = ~x23 & n13710 ;
  assign n13712 = x23 & n13706 ;
  assign n13713 = x23 & n2936 ;
  assign n13714 = ( x23 & n13706 ) | ( x23 & n13713 ) | ( n13706 & n13713 ) ;
  assign n13715 = ( ~n10957 & n13712 ) | ( ~n10957 & n13714 ) | ( n13712 & n13714 ) ;
  assign n13716 = n13712 | n13714 ;
  assign n13717 = ( n10949 & n13715 ) | ( n10949 & n13716 ) | ( n13715 & n13716 ) ;
  assign n13718 = x23 & ~n13717 ;
  assign n13719 = n13711 | n13718 ;
  assign n13720 = n12166 & n12184 ;
  assign n13721 = n12166 | n12184 ;
  assign n13722 = ~n13720 & n13721 ;
  assign n13723 = n13719 & n13722 ;
  assign n13724 = n13719 | n13722 ;
  assign n13725 = ~n13723 & n13724 ;
  assign n13726 = n12159 | n12162 ;
  assign n13727 = ~n12162 & n12164 ;
  assign n13728 = ( n12160 & n13726 ) | ( n12160 & ~n13727 ) | ( n13726 & ~n13727 ) ;
  assign n13729 = ~n12166 & n13728 ;
  assign n13730 = n2932 & n10654 ;
  assign n13731 = n2925 & n10667 ;
  assign n13732 = n2928 & ~n10662 ;
  assign n13733 = n13731 | n13732 ;
  assign n13734 = n13730 | n13733 ;
  assign n13735 = n2936 | n13730 ;
  assign n13736 = n13733 | n13735 ;
  assign n13737 = ( n10978 & n13734 ) | ( n10978 & n13736 ) | ( n13734 & n13736 ) ;
  assign n13738 = x23 & n13736 ;
  assign n13739 = x23 & n13734 ;
  assign n13740 = ( n10978 & n13738 ) | ( n10978 & n13739 ) | ( n13738 & n13739 ) ;
  assign n13741 = x23 & ~n13739 ;
  assign n13742 = x23 & ~n13738 ;
  assign n13743 = ( ~n10978 & n13741 ) | ( ~n10978 & n13742 ) | ( n13741 & n13742 ) ;
  assign n13744 = ( n13737 & ~n13740 ) | ( n13737 & n13743 ) | ( ~n13740 & n13743 ) ;
  assign n13745 = n13729 & n13744 ;
  assign n13746 = n2936 & n10784 ;
  assign n13747 = n2928 & ~n10678 ;
  assign n13748 = n2932 & ~n10675 ;
  assign n13749 = n13747 | n13748 ;
  assign n13750 = x23 | n13749 ;
  assign n13751 = n13746 | n13750 ;
  assign n13752 = ~x23 & n13751 ;
  assign n13753 = x23 & ~n2920 ;
  assign n13754 = ( x23 & n10678 ) | ( x23 & n13753 ) | ( n10678 & n13753 ) ;
  assign n13755 = n13751 & n13754 ;
  assign n13756 = n13746 | n13749 ;
  assign n13757 = n13754 & ~n13756 ;
  assign n13758 = ( n13752 & n13755 ) | ( n13752 & n13757 ) | ( n13755 & n13757 ) ;
  assign n13759 = n2932 & n10667 ;
  assign n13760 = n2925 & ~n10678 ;
  assign n13761 = n2928 & ~n10675 ;
  assign n13762 = n13760 | n13761 ;
  assign n13763 = n13759 | n13762 ;
  assign n13764 = n10837 | n13763 ;
  assign n13765 = n2936 | n13759 ;
  assign n13766 = n13762 | n13765 ;
  assign n13767 = ~x23 & n13766 ;
  assign n13768 = n13764 & n13767 ;
  assign n13769 = x23 | n13768 ;
  assign n13770 = n2302 & ~n10678 ;
  assign n13771 = n13768 & n13770 ;
  assign n13772 = n13764 & n13766 ;
  assign n13773 = n13770 & ~n13772 ;
  assign n13774 = ( n13769 & n13771 ) | ( n13769 & n13773 ) | ( n13771 & n13773 ) ;
  assign n13775 = n13758 & n13774 ;
  assign n13776 = ( n13768 & n13769 ) | ( n13768 & ~n13772 ) | ( n13769 & ~n13772 ) ;
  assign n13777 = n13758 | n13770 ;
  assign n13778 = ( n13770 & n13776 ) | ( n13770 & n13777 ) | ( n13776 & n13777 ) ;
  assign n13779 = ~n13775 & n13778 ;
  assign n13780 = n2932 & ~n10662 ;
  assign n13781 = n2925 & ~n10675 ;
  assign n13782 = n2928 & n10667 ;
  assign n13783 = n13781 | n13782 ;
  assign n13784 = n13780 | n13783 ;
  assign n13785 = ( n2936 & n10850 ) | ( n2936 & n13784 ) | ( n10850 & n13784 ) ;
  assign n13786 = ( x23 & n2936 ) | ( x23 & ~n13784 ) | ( n2936 & ~n13784 ) ;
  assign n13787 = ( x23 & n10850 ) | ( x23 & n13786 ) | ( n10850 & n13786 ) ;
  assign n13788 = ~n13785 & n13787 ;
  assign n13789 = n13784 | n13787 ;
  assign n13790 = ( ~x23 & n13788 ) | ( ~x23 & n13789 ) | ( n13788 & n13789 ) ;
  assign n13791 = n13775 | n13790 ;
  assign n13792 = ( n13775 & n13779 ) | ( n13775 & n13791 ) | ( n13779 & n13791 ) ;
  assign n13793 = n13729 | n13744 ;
  assign n13794 = ~n13745 & n13793 ;
  assign n13795 = n13745 | n13794 ;
  assign n13796 = ( n13745 & n13792 ) | ( n13745 & n13795 ) | ( n13792 & n13795 ) ;
  assign n13797 = n13725 & n13796 ;
  assign n13798 = n13723 | n13797 ;
  assign n13799 = n13701 & n13798 ;
  assign n13800 = n13698 | n13799 ;
  assign n13801 = ~n13665 & n13679 ;
  assign n13802 = ( n13665 & ~n13680 ) | ( n13665 & n13801 ) | ( ~n13680 & n13801 ) ;
  assign n13803 = n13680 | n13802 ;
  assign n13804 = ( n13680 & n13800 ) | ( n13680 & n13803 ) | ( n13800 & n13803 ) ;
  assign n13805 = n13662 & n13804 ;
  assign n13806 = n13659 | n13805 ;
  assign n13807 = n13627 | n13641 ;
  assign n13808 = ~n13642 & n13807 ;
  assign n13809 = n13642 | n13808 ;
  assign n13810 = ( n13642 & n13806 ) | ( n13642 & n13809 ) | ( n13806 & n13809 ) ;
  assign n13811 = n13625 & n13810 ;
  assign n13812 = ~n13609 & n13624 ;
  assign n13813 = n13810 | n13812 ;
  assign n13814 = n13609 | n13812 ;
  assign n13815 = ~n13812 & n13814 ;
  assign n13816 = ( n13811 & n13813 ) | ( n13811 & ~n13815 ) | ( n13813 & ~n13815 ) ;
  assign n13817 = n13602 | n13816 ;
  assign n13818 = ( n13602 & ~n13605 ) | ( n13602 & n13817 ) | ( ~n13605 & n13817 ) ;
  assign n13819 = n13556 | n13576 ;
  assign n13820 = ~n13577 & n13819 ;
  assign n13821 = n13577 | n13820 ;
  assign n13822 = ( n13577 & n13818 ) | ( n13577 & n13821 ) | ( n13818 & n13821 ) ;
  assign n13823 = ~n13553 & n13822 ;
  assign n13824 = n13553 & ~n13822 ;
  assign n13825 = n13823 | n13824 ;
  assign n13826 = n297 | n566 ;
  assign n13827 = n1483 | n13826 ;
  assign n13828 = ( ~n4024 & n12355 ) | ( ~n4024 & n13827 ) | ( n12355 & n13827 ) ;
  assign n13829 = n12355 & n13827 ;
  assign n13830 = ( ~n4023 & n13828 ) | ( ~n4023 & n13829 ) | ( n13828 & n13829 ) ;
  assign n13831 = n4025 | n13830 ;
  assign n13832 = n162 | n590 ;
  assign n13833 = n96 | n600 ;
  assign n13834 = n13832 | n13833 ;
  assign n13835 = n333 | n13834 ;
  assign n13836 = n332 | n417 ;
  assign n13837 = n5056 | n13836 ;
  assign n13838 = n442 | n502 ;
  assign n13839 = n317 | n2696 ;
  assign n13840 = n13838 | n13839 ;
  assign n13841 = n167 | n399 ;
  assign n13842 = n13840 | n13841 ;
  assign n13843 = n13837 | n13842 ;
  assign n13844 = n13835 | n13843 ;
  assign n13845 = n13831 | n13844 ;
  assign n13846 = n645 | n3414 ;
  assign n13847 = n6992 | n11076 ;
  assign n13848 = n13846 | n13847 ;
  assign n13849 = n179 | n503 ;
  assign n13850 = n222 | n458 ;
  assign n13851 = n13849 | n13850 ;
  assign n13852 = n444 | n13851 ;
  assign n13853 = n13848 | n13852 ;
  assign n13854 = n2214 | n4342 ;
  assign n13855 = n59 | n239 ;
  assign n13856 = n405 | n487 ;
  assign n13857 = n13855 | n13856 ;
  assign n13858 = n649 | n13857 ;
  assign n13859 = n13854 | n13858 ;
  assign n13860 = n13853 | n13859 ;
  assign n13861 = n349 | n820 ;
  assign n13862 = n518 | n13861 ;
  assign n13863 = n3313 | n5092 ;
  assign n13864 = n13862 | n13863 ;
  assign n13865 = n443 | n9128 ;
  assign n13866 = n202 | n288 ;
  assign n13867 = n170 | n320 ;
  assign n13868 = n13866 | n13867 ;
  assign n13869 = n13865 | n13868 ;
  assign n13870 = n13864 | n13869 ;
  assign n13871 = n660 | n13870 ;
  assign n13872 = n796 | n10772 ;
  assign n13873 = n13871 | n13872 ;
  assign n13874 = n13860 | n13873 ;
  assign n13875 = n13845 | n13874 ;
  assign n13876 = n1251 | n1631 ;
  assign n13877 = n952 | n13876 ;
  assign n13878 = n13321 | n13877 ;
  assign n13879 = n83 | n654 ;
  assign n13880 = n189 | n356 ;
  assign n13881 = n13879 | n13880 ;
  assign n13882 = n39 | n432 ;
  assign n13883 = n151 | n13882 ;
  assign n13884 = n13881 | n13883 ;
  assign n13885 = n12405 | n13884 ;
  assign n13886 = n13878 | n13885 ;
  assign n13887 = n13875 | n13886 ;
  assign n13888 = n13346 | n13887 ;
  assign n13889 = ( ~x11 & n13346 ) | ( ~x11 & n13887 ) | ( n13346 & n13887 ) ;
  assign n13890 = n13888 & ~n13889 ;
  assign n13891 = n13346 & n13887 ;
  assign n13892 = n13888 & ~n13891 ;
  assign n13893 = x11 | n13892 ;
  assign n13894 = ~n13890 & n13893 ;
  assign n13895 = n1057 & n3439 ;
  assign n13896 = ( n1057 & ~n3420 ) | ( n1057 & n13895 ) | ( ~n3420 & n13895 ) ;
  assign n13897 = n1065 & n3386 ;
  assign n13898 = n1060 & n3507 ;
  assign n13899 = ( n1060 & n3483 ) | ( n1060 & n13898 ) | ( n3483 & n13898 ) ;
  assign n13900 = n1062 | n13899 ;
  assign n13901 = n13897 | n13900 ;
  assign n13902 = n13896 | n13901 ;
  assign n13903 = ~n13894 & n13902 ;
  assign n13904 = n13896 | n13899 ;
  assign n13905 = n13897 | n13904 ;
  assign n13906 = ~n13894 & n13905 ;
  assign n13907 = ( ~n3530 & n13903 ) | ( ~n3530 & n13906 ) | ( n13903 & n13906 ) ;
  assign n13908 = n13894 & ~n13902 ;
  assign n13909 = n13894 & ~n13905 ;
  assign n13910 = ( n3530 & n13908 ) | ( n3530 & n13909 ) | ( n13908 & n13909 ) ;
  assign n13911 = n13907 | n13910 ;
  assign n13912 = n203 | n501 ;
  assign n13913 = n282 | n13912 ;
  assign n13914 = n85 | n451 ;
  assign n13915 = n542 | n13914 ;
  assign n13916 = n13913 | n13915 ;
  assign n13917 = n192 | n225 ;
  assign n13918 = n13916 | n13917 ;
  assign n13919 = n10342 | n11390 ;
  assign n13920 = n5139 | n13919 ;
  assign n13921 = n1160 | n3455 ;
  assign n13922 = n13920 | n13921 ;
  assign n13923 = n13918 | n13922 ;
  assign n13924 = n3481 | n13923 ;
  assign n13925 = n235 | n2044 ;
  assign n13926 = n271 | n13925 ;
  assign n13927 = n2042 | n13926 ;
  assign n13928 = n13924 | n13927 ;
  assign n13929 = n5026 | n13928 ;
  assign n13930 = n236 | n261 ;
  assign n13931 = n133 | n320 ;
  assign n13932 = n13930 | n13931 ;
  assign n13933 = n469 | n527 ;
  assign n13934 = n184 | n13933 ;
  assign n13935 = n13932 | n13934 ;
  assign n13936 = n13929 | n13935 ;
  assign n13937 = ~n13346 & n13936 ;
  assign n13938 = ~n13285 & n13347 ;
  assign n13939 = ( n13347 & ~n13349 ) | ( n13347 & n13938 ) | ( ~n13349 & n13938 ) ;
  assign n13940 = n13346 & ~n13936 ;
  assign n13941 = n13937 | n13940 ;
  assign n13942 = n13939 | n13941 ;
  assign n13943 = ~n13937 & n13942 ;
  assign n13944 = n13347 | n13937 ;
  assign n13945 = n13940 | n13944 ;
  assign n13946 = ( ~n13350 & n13941 ) | ( ~n13350 & n13945 ) | ( n13941 & n13945 ) ;
  assign n13947 = ~n13937 & n13946 ;
  assign n13948 = ( ~n3603 & n13943 ) | ( ~n3603 & n13947 ) | ( n13943 & n13947 ) ;
  assign n13949 = n13911 | n13948 ;
  assign n13950 = n13911 & n13948 ;
  assign n13951 = n13949 & ~n13950 ;
  assign n13952 = n13347 & ~n13350 ;
  assign n13953 = ( ~n3603 & n13939 ) | ( ~n3603 & n13952 ) | ( n13939 & n13952 ) ;
  assign n13954 = ( ~n3603 & n13942 ) | ( ~n3603 & n13946 ) | ( n13942 & n13946 ) ;
  assign n13955 = ~n13953 & n13954 ;
  assign n13956 = ~n13940 & n13947 ;
  assign n13957 = ~n13940 & n13943 ;
  assign n13958 = ( ~n3603 & n13956 ) | ( ~n3603 & n13957 ) | ( n13956 & n13957 ) ;
  assign n13959 = n13955 | n13958 ;
  assign n13960 = n1057 & n3386 ;
  assign n13961 = n1060 & n2893 ;
  assign n13962 = ( n1060 & ~n2886 ) | ( n1060 & n13961 ) | ( ~n2886 & n13961 ) ;
  assign n13963 = n1065 & n3507 ;
  assign n13964 = ( n1065 & n3483 ) | ( n1065 & n13963 ) | ( n3483 & n13963 ) ;
  assign n13965 = n1062 | n13964 ;
  assign n13966 = n13962 | n13965 ;
  assign n13967 = n13960 | n13966 ;
  assign n13968 = n13962 | n13964 ;
  assign n13969 = n13960 | n13968 ;
  assign n13970 = ( ~n3568 & n13967 ) | ( ~n3568 & n13969 ) | ( n13967 & n13969 ) ;
  assign n13971 = n13959 & n13970 ;
  assign n13972 = n13951 & n13971 ;
  assign n13973 = n13959 & ~n13971 ;
  assign n13974 = n1823 & n4206 ;
  assign n13975 = n1829 & ~n4429 ;
  assign n13976 = n1826 & n3439 ;
  assign n13977 = ( n1826 & ~n3420 ) | ( n1826 & n13976 ) | ( ~n3420 & n13976 ) ;
  assign n13978 = n13975 | n13977 ;
  assign n13979 = n13974 | n13978 ;
  assign n13980 = n1821 | n13974 ;
  assign n13981 = n13978 | n13980 ;
  assign n13982 = ( ~n4527 & n13979 ) | ( ~n4527 & n13981 ) | ( n13979 & n13981 ) ;
  assign n13983 = ~x29 & n13981 ;
  assign n13984 = ~x29 & n13979 ;
  assign n13985 = ( ~n4527 & n13983 ) | ( ~n4527 & n13984 ) | ( n13983 & n13984 ) ;
  assign n13986 = x29 | n13984 ;
  assign n13987 = x29 | n13983 ;
  assign n13988 = ( ~n4527 & n13986 ) | ( ~n4527 & n13987 ) | ( n13986 & n13987 ) ;
  assign n13989 = ( ~n13982 & n13985 ) | ( ~n13982 & n13988 ) | ( n13985 & n13988 ) ;
  assign n13990 = ~n13959 & n13970 ;
  assign n13991 = n13989 & n13990 ;
  assign n13992 = ( n13973 & n13989 ) | ( n13973 & n13991 ) | ( n13989 & n13991 ) ;
  assign n13993 = ( n13951 & n13972 ) | ( n13951 & n13992 ) | ( n13972 & n13992 ) ;
  assign n13994 = n13951 | n13971 ;
  assign n13995 = n13992 | n13994 ;
  assign n13996 = ~n13993 & n13995 ;
  assign n13997 = n1823 & ~n4429 ;
  assign n13998 = n1823 | n1826 ;
  assign n13999 = ( n1826 & ~n4429 ) | ( n1826 & n13998 ) | ( ~n4429 & n13998 ) ;
  assign n14000 = ( n4206 & n13997 ) | ( n4206 & n13999 ) | ( n13997 & n13999 ) ;
  assign n14001 = n1829 & n4396 ;
  assign n14002 = n14000 | n14001 ;
  assign n14003 = n1821 | n14001 ;
  assign n14004 = n14000 | n14003 ;
  assign n14005 = ( ~n4501 & n14002 ) | ( ~n4501 & n14004 ) | ( n14002 & n14004 ) ;
  assign n14006 = ~x29 & n14004 ;
  assign n14007 = ~x29 & n14002 ;
  assign n14008 = ( ~n4501 & n14006 ) | ( ~n4501 & n14007 ) | ( n14006 & n14007 ) ;
  assign n14009 = x29 | n14007 ;
  assign n14010 = x29 | n14006 ;
  assign n14011 = ( ~n4501 & n14009 ) | ( ~n4501 & n14010 ) | ( n14009 & n14010 ) ;
  assign n14012 = ( ~n14005 & n14008 ) | ( ~n14005 & n14011 ) | ( n14008 & n14011 ) ;
  assign n14013 = n13996 & n14012 ;
  assign n14014 = n13996 & ~n14013 ;
  assign n14015 = n2312 & n4245 ;
  assign n14016 = ( n2312 & n4303 ) | ( n2312 & n14015 ) | ( n4303 & n14015 ) ;
  assign n14017 = n2308 & n5192 ;
  assign n14018 = ( n2308 & n5179 ) | ( n2308 & n14017 ) | ( n5179 & n14017 ) ;
  assign n14019 = n14016 | n14018 ;
  assign n14020 = n2315 & n5117 ;
  assign n14021 = ( n2315 & ~n5037 ) | ( n2315 & n14020 ) | ( ~n5037 & n14020 ) ;
  assign n14023 = n2306 | n14021 ;
  assign n14024 = n14019 | n14023 ;
  assign n14022 = n14019 | n14021 ;
  assign n14025 = n14022 & n14024 ;
  assign n14026 = ( ~n5270 & n14024 ) | ( ~n5270 & n14025 ) | ( n14024 & n14025 ) ;
  assign n14027 = ~x26 & n14025 ;
  assign n14028 = ~x26 & n14024 ;
  assign n14029 = ( ~n5270 & n14027 ) | ( ~n5270 & n14028 ) | ( n14027 & n14028 ) ;
  assign n14030 = x26 | n14027 ;
  assign n14031 = x26 | n14028 ;
  assign n14032 = ( ~n5270 & n14030 ) | ( ~n5270 & n14031 ) | ( n14030 & n14031 ) ;
  assign n14033 = ( ~n14026 & n14029 ) | ( ~n14026 & n14032 ) | ( n14029 & n14032 ) ;
  assign n14034 = n14012 & n14033 ;
  assign n14035 = ~n13996 & n14034 ;
  assign n14036 = ( n14014 & n14033 ) | ( n14014 & n14035 ) | ( n14033 & n14035 ) ;
  assign n14037 = n14012 | n14033 ;
  assign n14038 = ( ~n13996 & n14033 ) | ( ~n13996 & n14037 ) | ( n14033 & n14037 ) ;
  assign n14039 = n14014 | n14038 ;
  assign n14040 = ~n14036 & n14039 ;
  assign n14041 = n13989 | n13990 ;
  assign n14042 = n13973 | n14041 ;
  assign n14043 = ~n13992 & n14042 ;
  assign n14044 = n13359 | n13377 ;
  assign n14045 = ( n13359 & n13361 ) | ( n13359 & n14044 ) | ( n13361 & n14044 ) ;
  assign n14046 = n14043 & n14045 ;
  assign n14047 = n14043 | n14045 ;
  assign n14048 = ~n14046 & n14047 ;
  assign n14049 = n2312 & n4396 ;
  assign n14050 = n2308 & n4245 ;
  assign n14051 = ( n2308 & n4303 ) | ( n2308 & n14050 ) | ( n4303 & n14050 ) ;
  assign n14052 = n14049 | n14051 ;
  assign n14053 = n2315 & n5192 ;
  assign n14054 = ( n2315 & n5179 ) | ( n2315 & n14053 ) | ( n5179 & n14053 ) ;
  assign n14055 = n14052 | n14054 ;
  assign n14056 = n2306 | n14054 ;
  assign n14057 = n14052 | n14056 ;
  assign n14058 = ( n5306 & n14055 ) | ( n5306 & n14057 ) | ( n14055 & n14057 ) ;
  assign n14059 = x26 & n14057 ;
  assign n14060 = x26 & n14055 ;
  assign n14061 = ( n5306 & n14059 ) | ( n5306 & n14060 ) | ( n14059 & n14060 ) ;
  assign n14062 = x26 & ~n14060 ;
  assign n14063 = x26 & ~n14059 ;
  assign n14064 = ( ~n5306 & n14062 ) | ( ~n5306 & n14063 ) | ( n14062 & n14063 ) ;
  assign n14065 = ( n14058 & ~n14061 ) | ( n14058 & n14064 ) | ( ~n14061 & n14064 ) ;
  assign n14066 = n14046 | n14065 ;
  assign n14067 = ( n14046 & n14048 ) | ( n14046 & n14066 ) | ( n14048 & n14066 ) ;
  assign n14068 = n14040 & n14067 ;
  assign n14069 = n14040 | n14067 ;
  assign n14070 = ~n14068 & n14069 ;
  assign n14071 = n2925 & n5108 ;
  assign n14072 = n2928 & n5997 ;
  assign n14073 = ( n2928 & n5979 ) | ( n2928 & n14072 ) | ( n5979 & n14072 ) ;
  assign n14074 = n14071 | n14073 ;
  assign n14075 = n2932 & n5857 ;
  assign n14076 = ( n2932 & ~n5899 ) | ( n2932 & n14075 ) | ( ~n5899 & n14075 ) ;
  assign n14077 = n14074 | n14076 ;
  assign n14078 = n2936 | n14077 ;
  assign n14079 = ( ~n6151 & n14077 ) | ( ~n6151 & n14078 ) | ( n14077 & n14078 ) ;
  assign n14080 = ~x23 & n14078 ;
  assign n14081 = ~x23 & n14077 ;
  assign n14082 = ( ~n6151 & n14080 ) | ( ~n6151 & n14081 ) | ( n14080 & n14081 ) ;
  assign n14083 = x23 | n14080 ;
  assign n14084 = x23 | n14081 ;
  assign n14085 = ( ~n6151 & n14083 ) | ( ~n6151 & n14084 ) | ( n14083 & n14084 ) ;
  assign n14086 = ( ~n14079 & n14082 ) | ( ~n14079 & n14085 ) | ( n14082 & n14085 ) ;
  assign n14087 = n14070 & n14086 ;
  assign n14088 = ~n14070 & n14086 ;
  assign n14089 = ( n14070 & ~n14087 ) | ( n14070 & n14088 ) | ( ~n14087 & n14088 ) ;
  assign n14090 = n14048 & ~n14065 ;
  assign n14091 = n14048 | n14065 ;
  assign n14092 = ( ~n14048 & n14090 ) | ( ~n14048 & n14091 ) | ( n14090 & n14091 ) ;
  assign n14093 = n13382 | n13401 ;
  assign n14094 = ( n13382 & n13385 ) | ( n13382 & n14093 ) | ( n13385 & n14093 ) ;
  assign n14095 = n14092 & n14094 ;
  assign n14096 = n14092 | n14094 ;
  assign n14097 = ~n14095 & n14096 ;
  assign n14098 = n2925 & n5117 ;
  assign n14099 = ( n2925 & ~n5037 ) | ( n2925 & n14098 ) | ( ~n5037 & n14098 ) ;
  assign n14100 = n2928 & n5108 ;
  assign n14101 = n2932 & n5997 ;
  assign n14102 = ( n2932 & n5979 ) | ( n2932 & n14101 ) | ( n5979 & n14101 ) ;
  assign n14103 = n14100 | n14102 ;
  assign n14104 = n14099 | n14103 ;
  assign n14105 = n2936 | n14104 ;
  assign n14106 = ( n6181 & n14104 ) | ( n6181 & n14105 ) | ( n14104 & n14105 ) ;
  assign n14107 = x23 & n14105 ;
  assign n14108 = x23 & n14104 ;
  assign n14109 = ( n6181 & n14107 ) | ( n6181 & n14108 ) | ( n14107 & n14108 ) ;
  assign n14110 = x23 & ~n14107 ;
  assign n14111 = x23 & ~n14108 ;
  assign n14112 = ( ~n6181 & n14110 ) | ( ~n6181 & n14111 ) | ( n14110 & n14111 ) ;
  assign n14113 = ( n14106 & ~n14109 ) | ( n14106 & n14112 ) | ( ~n14109 & n14112 ) ;
  assign n14114 = n14095 | n14113 ;
  assign n14115 = ( n14095 & n14097 ) | ( n14095 & n14114 ) | ( n14097 & n14114 ) ;
  assign n14116 = n14089 & n14115 ;
  assign n14117 = n14089 | n14115 ;
  assign n14118 = ~n14116 & n14117 ;
  assign n14119 = n3544 & ~n6091 ;
  assign n14120 = n3541 & n7036 ;
  assign n14121 = ( n3541 & n7023 ) | ( n3541 & n14120 ) | ( n7023 & n14120 ) ;
  assign n14122 = n14119 | n14121 ;
  assign n14123 = n3547 & n6950 ;
  assign n14124 = n14122 | n14123 ;
  assign n14125 = n3537 | n14124 ;
  assign n14126 = n14124 & n14125 ;
  assign n14127 = ( ~n7107 & n14125 ) | ( ~n7107 & n14126 ) | ( n14125 & n14126 ) ;
  assign n14128 = ~x20 & n14126 ;
  assign n14129 = ~x20 & n14125 ;
  assign n14130 = ( ~n7107 & n14128 ) | ( ~n7107 & n14129 ) | ( n14128 & n14129 ) ;
  assign n14131 = x20 | n14128 ;
  assign n14132 = x20 | n14129 ;
  assign n14133 = ( ~n7107 & n14131 ) | ( ~n7107 & n14132 ) | ( n14131 & n14132 ) ;
  assign n14134 = ( ~n14127 & n14130 ) | ( ~n14127 & n14133 ) | ( n14130 & n14133 ) ;
  assign n14135 = n14118 & n14134 ;
  assign n14136 = n14118 | n14134 ;
  assign n14137 = ~n14135 & n14136 ;
  assign n14138 = n14097 & ~n14113 ;
  assign n14139 = n14097 | n14113 ;
  assign n14140 = ( ~n14097 & n14138 ) | ( ~n14097 & n14139 ) | ( n14138 & n14139 ) ;
  assign n14141 = n13406 | n13424 ;
  assign n14142 = ( n13406 & n13408 ) | ( n13406 & n14141 ) | ( n13408 & n14141 ) ;
  assign n14143 = n14140 & n14142 ;
  assign n14144 = n14140 | n14142 ;
  assign n14145 = ~n14143 & n14144 ;
  assign n14146 = n3544 & n5857 ;
  assign n14147 = ( n3544 & ~n5899 ) | ( n3544 & n14146 ) | ( ~n5899 & n14146 ) ;
  assign n14148 = n3541 & ~n6091 ;
  assign n14149 = n3547 & n7036 ;
  assign n14150 = ( n3547 & n7023 ) | ( n3547 & n14149 ) | ( n7023 & n14149 ) ;
  assign n14151 = n14148 | n14150 ;
  assign n14152 = n14147 | n14151 ;
  assign n14153 = n3537 | n14152 ;
  assign n14154 = ( n7136 & n14152 ) | ( n7136 & n14153 ) | ( n14152 & n14153 ) ;
  assign n14155 = x20 & n14153 ;
  assign n14156 = x20 & n14152 ;
  assign n14157 = ( n7136 & n14155 ) | ( n7136 & n14156 ) | ( n14155 & n14156 ) ;
  assign n14158 = x20 & ~n14155 ;
  assign n14159 = x20 & ~n14156 ;
  assign n14160 = ( ~n7136 & n14158 ) | ( ~n7136 & n14159 ) | ( n14158 & n14159 ) ;
  assign n14161 = ( n14154 & ~n14157 ) | ( n14154 & n14160 ) | ( ~n14157 & n14160 ) ;
  assign n14162 = n14143 | n14161 ;
  assign n14163 = ( n14143 & n14145 ) | ( n14143 & n14162 ) | ( n14145 & n14162 ) ;
  assign n14164 = n14137 & n14163 ;
  assign n14165 = n14137 | n14163 ;
  assign n14166 = ~n14164 & n14165 ;
  assign n14167 = n4466 & n6889 ;
  assign n14168 = ( n4466 & ~n6884 ) | ( n4466 & n14167 ) | ( ~n6884 & n14167 ) ;
  assign n14169 = n4468 & n7907 ;
  assign n14170 = ( n4468 & n7902 ) | ( n4468 & n14169 ) | ( n7902 & n14169 ) ;
  assign n14171 = n4471 & n8079 ;
  assign n14172 = ( n4471 & ~n8070 ) | ( n4471 & n14171 ) | ( ~n8070 & n14171 ) ;
  assign n14173 = n14170 | n14172 ;
  assign n14174 = n14168 | n14173 ;
  assign n14175 = n4475 | n14174 ;
  assign n14176 = ( ~n8156 & n14174 ) | ( ~n8156 & n14175 ) | ( n14174 & n14175 ) ;
  assign n14177 = ~x17 & n14175 ;
  assign n14178 = ~x17 & n14174 ;
  assign n14179 = ( ~n8156 & n14177 ) | ( ~n8156 & n14178 ) | ( n14177 & n14178 ) ;
  assign n14180 = x17 | n14177 ;
  assign n14181 = x17 | n14178 ;
  assign n14182 = ( ~n8156 & n14180 ) | ( ~n8156 & n14181 ) | ( n14180 & n14181 ) ;
  assign n14183 = ( ~n14176 & n14179 ) | ( ~n14176 & n14182 ) | ( n14179 & n14182 ) ;
  assign n14184 = n14166 & n14183 ;
  assign n14185 = n14166 & ~n14184 ;
  assign n14186 = n14145 & ~n14161 ;
  assign n14187 = n14145 | n14161 ;
  assign n14188 = ( ~n14145 & n14186 ) | ( ~n14145 & n14187 ) | ( n14186 & n14187 ) ;
  assign n14189 = n13430 | n13448 ;
  assign n14190 = ( n13430 & n13432 ) | ( n13430 & n14189 ) | ( n13432 & n14189 ) ;
  assign n14191 = n14188 & n14190 ;
  assign n14192 = n14188 | n14190 ;
  assign n14193 = ~n14191 & n14192 ;
  assign n14194 = n4466 & n6950 ;
  assign n14195 = n4468 & n6889 ;
  assign n14196 = ( n4468 & ~n6884 ) | ( n4468 & n14195 ) | ( ~n6884 & n14195 ) ;
  assign n14197 = n14194 | n14196 ;
  assign n14198 = n4471 & n7907 ;
  assign n14199 = ( n4471 & n7902 ) | ( n4471 & n14198 ) | ( n7902 & n14198 ) ;
  assign n14200 = n14197 | n14199 ;
  assign n14201 = n4475 | n14199 ;
  assign n14202 = n14197 | n14201 ;
  assign n14203 = ( ~n8193 & n14200 ) | ( ~n8193 & n14202 ) | ( n14200 & n14202 ) ;
  assign n14204 = ~x17 & n14202 ;
  assign n14205 = ~x17 & n14200 ;
  assign n14206 = ( ~n8193 & n14204 ) | ( ~n8193 & n14205 ) | ( n14204 & n14205 ) ;
  assign n14207 = x17 | n14205 ;
  assign n14208 = x17 | n14204 ;
  assign n14209 = ( ~n8193 & n14207 ) | ( ~n8193 & n14208 ) | ( n14207 & n14208 ) ;
  assign n14210 = ( ~n14203 & n14206 ) | ( ~n14203 & n14209 ) | ( n14206 & n14209 ) ;
  assign n14211 = n14191 | n14210 ;
  assign n14212 = ( n14191 & n14193 ) | ( n14191 & n14211 ) | ( n14193 & n14211 ) ;
  assign n14213 = ~n14166 & n14183 ;
  assign n14214 = n14212 & n14213 ;
  assign n14215 = ( n14185 & n14212 ) | ( n14185 & n14214 ) | ( n14212 & n14214 ) ;
  assign n14216 = n14212 | n14213 ;
  assign n14217 = n14185 | n14216 ;
  assign n14218 = ~n14215 & n14217 ;
  assign n14236 = n14193 & ~n14210 ;
  assign n14237 = n14193 | n14210 ;
  assign n14238 = ( ~n14193 & n14236 ) | ( ~n14193 & n14237 ) | ( n14236 & n14237 ) ;
  assign n14239 = n13452 | n13471 ;
  assign n14240 = ( n13452 & n13454 ) | ( n13452 & n14239 ) | ( n13454 & n14239 ) ;
  assign n14241 = n14238 & n14240 ;
  assign n14242 = n14238 | n14240 ;
  assign n14243 = ~n14241 & n14242 ;
  assign n14244 = n5237 & n8079 ;
  assign n14245 = ( n5237 & ~n8070 ) | ( n5237 & n14244 ) | ( ~n8070 & n14244 ) ;
  assign n14246 = n5231 | n14245 ;
  assign n14247 = ( ~n8017 & n14245 ) | ( ~n8017 & n14246 ) | ( n14245 & n14246 ) ;
  assign n14248 = n5234 & n9022 ;
  assign n14249 = ( n5234 & ~n9019 ) | ( n5234 & n14248 ) | ( ~n9019 & n14248 ) ;
  assign n14250 = n14247 | n14249 ;
  assign n14251 = n5227 | n14249 ;
  assign n14252 = n14247 | n14251 ;
  assign n14253 = ( ~n9416 & n14250 ) | ( ~n9416 & n14252 ) | ( n14250 & n14252 ) ;
  assign n14254 = ~x14 & n14252 ;
  assign n14255 = ~x14 & n14250 ;
  assign n14256 = ( ~n9416 & n14254 ) | ( ~n9416 & n14255 ) | ( n14254 & n14255 ) ;
  assign n14257 = x14 | n14255 ;
  assign n14258 = x14 | n14254 ;
  assign n14259 = ( ~n9416 & n14257 ) | ( ~n9416 & n14258 ) | ( n14257 & n14258 ) ;
  assign n14260 = ( ~n14253 & n14256 ) | ( ~n14253 & n14259 ) | ( n14256 & n14259 ) ;
  assign n14261 = n14241 | n14260 ;
  assign n14262 = ( n14241 & n14243 ) | ( n14241 & n14261 ) | ( n14243 & n14261 ) ;
  assign n14219 = n5234 & ~n8982 ;
  assign n14220 = ( n5234 & n9051 ) | ( n5234 & n14219 ) | ( n9051 & n14219 ) ;
  assign n14221 = n5231 & n9022 ;
  assign n14222 = n14220 | n14221 ;
  assign n14223 = n5231 | n14220 ;
  assign n14224 = ( ~n9019 & n14222 ) | ( ~n9019 & n14223 ) | ( n14222 & n14223 ) ;
  assign n14225 = n5237 | n14224 ;
  assign n14226 = ( ~n8017 & n14224 ) | ( ~n8017 & n14225 ) | ( n14224 & n14225 ) ;
  assign n14227 = n5227 | n14226 ;
  assign n14228 = ( ~n10242 & n14226 ) | ( ~n10242 & n14227 ) | ( n14226 & n14227 ) ;
  assign n14229 = ~x14 & n14227 ;
  assign n14230 = ~x14 & n14226 ;
  assign n14231 = ( ~n10242 & n14229 ) | ( ~n10242 & n14230 ) | ( n14229 & n14230 ) ;
  assign n14232 = x14 | n14229 ;
  assign n14233 = x14 | n14230 ;
  assign n14234 = ( ~n10242 & n14232 ) | ( ~n10242 & n14233 ) | ( n14232 & n14233 ) ;
  assign n14235 = ( ~n14228 & n14231 ) | ( ~n14228 & n14234 ) | ( n14231 & n14234 ) ;
  assign n14263 = n14235 & n14262 ;
  assign n14264 = n14262 & ~n14263 ;
  assign n14265 = n14218 & n14235 ;
  assign n14266 = ~n14262 & n14265 ;
  assign n14267 = ( n14218 & n14264 ) | ( n14218 & n14266 ) | ( n14264 & n14266 ) ;
  assign n14268 = n14218 | n14235 ;
  assign n14269 = ( n14218 & ~n14262 ) | ( n14218 & n14268 ) | ( ~n14262 & n14268 ) ;
  assign n14270 = n14264 | n14269 ;
  assign n14271 = ~n14267 & n14270 ;
  assign n14272 = n6125 & ~n8982 ;
  assign n14273 = ( n6125 & n9051 ) | ( n6125 & n14272 ) | ( n9051 & n14272 ) ;
  assign n14274 = n6115 | n14273 ;
  assign n14275 = n9442 & ~n14273 ;
  assign n14276 = n9074 & ~n14273 ;
  assign n14277 = ( ~n9440 & n14275 ) | ( ~n9440 & n14276 ) | ( n14275 & n14276 ) ;
  assign n14278 = n14274 & ~n14277 ;
  assign n14279 = n14273 & n14274 ;
  assign n14280 = ( ~n9442 & n14274 ) | ( ~n9442 & n14279 ) | ( n14274 & n14279 ) ;
  assign n14281 = ( ~n9072 & n14278 ) | ( ~n9072 & n14280 ) | ( n14278 & n14280 ) ;
  assign n14282 = ~x11 & n14278 ;
  assign n14283 = ~x11 & n14280 ;
  assign n14284 = ( ~n9072 & n14282 ) | ( ~n9072 & n14283 ) | ( n14282 & n14283 ) ;
  assign n14285 = x11 | n14282 ;
  assign n14286 = x11 | n14283 ;
  assign n14287 = ( ~n9072 & n14285 ) | ( ~n9072 & n14286 ) | ( n14285 & n14286 ) ;
  assign n14288 = ( ~n14281 & n14284 ) | ( ~n14281 & n14287 ) | ( n14284 & n14287 ) ;
  assign n14289 = n13477 | n13496 ;
  assign n14290 = ( n13477 & n13479 ) | ( n13477 & n14289 ) | ( n13479 & n14289 ) ;
  assign n14291 = n14288 & n14290 ;
  assign n14292 = n14288 | n14290 ;
  assign n14293 = ~n14291 & n14292 ;
  assign n14294 = n14243 & ~n14260 ;
  assign n14295 = n14243 | n14260 ;
  assign n14296 = ( ~n14243 & n14294 ) | ( ~n14243 & n14295 ) | ( n14294 & n14295 ) ;
  assign n14297 = n14291 | n14296 ;
  assign n14298 = ( n14291 & n14293 ) | ( n14291 & n14297 ) | ( n14293 & n14297 ) ;
  assign n14299 = n14271 & n14298 ;
  assign n14300 = n14271 | n14298 ;
  assign n14301 = ~n14299 & n14300 ;
  assign n14302 = n14293 & ~n14296 ;
  assign n14303 = n14293 | n14296 ;
  assign n14304 = ( ~n14293 & n14302 ) | ( ~n14293 & n14303 ) | ( n14302 & n14303 ) ;
  assign n14305 = n13271 | n13499 ;
  assign n14306 = ( n13271 & n13276 ) | ( n13271 & n14305 ) | ( n13276 & n14305 ) ;
  assign n14307 = n14304 & n14306 ;
  assign n14308 = n14304 | n14306 ;
  assign n14309 = ~n14307 & n14308 ;
  assign n14310 = n13505 | n13507 ;
  assign n14311 = n14309 & n14310 ;
  assign n14312 = n14307 | n14311 ;
  assign n14313 = n14301 & n14312 ;
  assign n14314 = n13505 & n14309 ;
  assign n14315 = n14307 | n14314 ;
  assign n14316 = n14301 & n14315 ;
  assign n14317 = ( n13511 & n14313 ) | ( n13511 & n14316 ) | ( n14313 & n14316 ) ;
  assign n14318 = ( n13510 & n14313 ) | ( n13510 & n14316 ) | ( n14313 & n14316 ) ;
  assign n14319 = ( n12928 & n14317 ) | ( n12928 & n14318 ) | ( n14317 & n14318 ) ;
  assign n14320 = ( n12930 & n14317 ) | ( n12930 & n14318 ) | ( n14317 & n14318 ) ;
  assign n14321 = ( n11360 & n14319 ) | ( n11360 & n14320 ) | ( n14319 & n14320 ) ;
  assign n14322 = ( n13511 & n14312 ) | ( n13511 & n14315 ) | ( n14312 & n14315 ) ;
  assign n14323 = ( n13510 & n14312 ) | ( n13510 & n14315 ) | ( n14312 & n14315 ) ;
  assign n14324 = ( n12930 & n14322 ) | ( n12930 & n14323 ) | ( n14322 & n14323 ) ;
  assign n14325 = n14301 | n14324 ;
  assign n14326 = ( n12928 & n14322 ) | ( n12928 & n14323 ) | ( n14322 & n14323 ) ;
  assign n14327 = n14301 | n14326 ;
  assign n14328 = ( n11360 & n14325 ) | ( n11360 & n14327 ) | ( n14325 & n14327 ) ;
  assign n14329 = ~n14321 & n14328 ;
  assign n14330 = n5231 & ~n8982 ;
  assign n14331 = ( n5231 & n9051 ) | ( n5231 & n14330 ) | ( n9051 & n14330 ) ;
  assign n14332 = n5237 & ~n9022 ;
  assign n14333 = ( n5237 & n14331 ) | ( n5237 & ~n14332 ) | ( n14331 & ~n14332 ) ;
  assign n14334 = n5237 | n14331 ;
  assign n14335 = ( ~n9019 & n14333 ) | ( ~n9019 & n14334 ) | ( n14333 & n14334 ) ;
  assign n14336 = n5227 | n14335 ;
  assign n14337 = ( n9078 & n14335 ) | ( n9078 & n14336 ) | ( n14335 & n14336 ) ;
  assign n14338 = x14 & n14336 ;
  assign n14339 = x14 & n14335 ;
  assign n14340 = ( n9078 & n14338 ) | ( n9078 & n14339 ) | ( n14338 & n14339 ) ;
  assign n14341 = x14 & ~n14338 ;
  assign n14342 = x14 & ~n14339 ;
  assign n14343 = ( ~n9078 & n14341 ) | ( ~n9078 & n14342 ) | ( n14341 & n14342 ) ;
  assign n14344 = ( n14337 & ~n14340 ) | ( n14337 & n14343 ) | ( ~n14340 & n14343 ) ;
  assign n14345 = n14183 & n14344 ;
  assign n14346 = n14166 & n14345 ;
  assign n14347 = ( n14215 & n14344 ) | ( n14215 & n14346 ) | ( n14344 & n14346 ) ;
  assign n14348 = n14183 | n14344 ;
  assign n14349 = ( n14166 & n14344 ) | ( n14166 & n14348 ) | ( n14344 & n14348 ) ;
  assign n14350 = n14215 | n14349 ;
  assign n14351 = ~n14347 & n14350 ;
  assign n14352 = n1057 & n4206 ;
  assign n14353 = n1060 & n3386 ;
  assign n14354 = n1065 & n3439 ;
  assign n14355 = ( n1065 & ~n3420 ) | ( n1065 & n14354 ) | ( ~n3420 & n14354 ) ;
  assign n14356 = n14353 | n14355 ;
  assign n14357 = n14352 | n14356 ;
  assign n14358 = n1062 | n14352 ;
  assign n14359 = n14356 | n14358 ;
  assign n14360 = ( ~n4220 & n14357 ) | ( ~n4220 & n14359 ) | ( n14357 & n14359 ) ;
  assign n14361 = n310 | n574 ;
  assign n14362 = n151 | n14361 ;
  assign n14363 = n542 | n901 ;
  assign n14364 = n1723 | n14363 ;
  assign n14365 = n11388 | n14364 ;
  assign n14366 = n14362 | n14365 ;
  assign n14367 = n13306 | n14366 ;
  assign n14368 = n1002 | n1608 ;
  assign n14369 = n14367 | n14368 ;
  assign n14370 = n573 | n5133 ;
  assign n14371 = n1079 | n14370 ;
  assign n14372 = n53 | n257 ;
  assign n14373 = n189 | n249 ;
  assign n14374 = n14372 | n14373 ;
  assign n14375 = n14371 | n14374 ;
  assign n14376 = n321 | n465 ;
  assign n14377 = n183 | n255 ;
  assign n14378 = n14376 | n14377 ;
  assign n14379 = n223 | n14378 ;
  assign n14380 = n349 | n14379 ;
  assign n14381 = n14375 | n14380 ;
  assign n14382 = n14369 | n14381 ;
  assign n14383 = n114 | n431 ;
  assign n14384 = n577 | n14383 ;
  assign n14385 = n4247 | n14384 ;
  assign n14386 = n635 | n14385 ;
  assign n14387 = n168 | n497 ;
  assign n14388 = n1581 | n14387 ;
  assign n14389 = n7029 | n14388 ;
  assign n14390 = n14386 | n14389 ;
  assign n14391 = n152 | n239 ;
  assign n14392 = n155 | n14391 ;
  assign n14393 = n460 | n1014 ;
  assign n14394 = n14392 | n14393 ;
  assign n14395 = n608 | n14394 ;
  assign n14396 = n383 | n388 ;
  assign n14397 = n208 | n372 ;
  assign n14398 = n14396 | n14397 ;
  assign n14399 = n448 | n14398 ;
  assign n14400 = n14395 | n14399 ;
  assign n14401 = n14390 | n14400 ;
  assign n14402 = n14382 | n14401 ;
  assign n14403 = n879 | n2163 ;
  assign n14404 = n9158 | n14403 ;
  assign n14405 = n11100 | n14404 ;
  assign n14406 = n181 | n182 ;
  assign n14407 = n539 | n561 ;
  assign n14408 = n405 | n14407 ;
  assign n14409 = ( n304 & ~n14406 ) | ( n304 & n14408 ) | ( ~n14406 & n14408 ) ;
  assign n14410 = n110 | n229 ;
  assign n14411 = n14406 | n14410 ;
  assign n14412 = n14409 | n14411 ;
  assign n14413 = n14405 | n14412 ;
  assign n14414 = n728 | n1031 ;
  assign n14415 = n654 | n967 ;
  assign n14416 = n14414 | n14415 ;
  assign n14417 = n313 | n1039 ;
  assign n14418 = n14416 | n14417 ;
  assign n14419 = n39 | n666 ;
  assign n14420 = n281 | n675 ;
  assign n14421 = n14419 | n14420 ;
  assign n14422 = n14418 | n14421 ;
  assign n14423 = n14413 | n14422 ;
  assign n14424 = n710 | n1479 ;
  assign n14425 = n306 | n456 ;
  assign n14426 = n689 | n14425 ;
  assign n14427 = n14424 | n14426 ;
  assign n14428 = n196 | n263 ;
  assign n14429 = n676 | n14428 ;
  assign n14430 = n14427 | n14429 ;
  assign n14431 = n14423 | n14430 ;
  assign n14432 = n14402 | n14431 ;
  assign n14433 = n13889 & ~n14432 ;
  assign n14434 = ~n13889 & n14432 ;
  assign n14435 = n14433 | n14434 ;
  assign n14436 = n14359 & n14435 ;
  assign n14437 = n14357 & n14435 ;
  assign n14438 = ( ~n4220 & n14436 ) | ( ~n4220 & n14437 ) | ( n14436 & n14437 ) ;
  assign n14439 = n14435 & ~n14437 ;
  assign n14440 = n14435 & ~n14436 ;
  assign n14441 = ( n4220 & n14439 ) | ( n4220 & n14440 ) | ( n14439 & n14440 ) ;
  assign n14442 = ( n14360 & ~n14438 ) | ( n14360 & n14441 ) | ( ~n14438 & n14441 ) ;
  assign n14443 = ~n13907 & n13948 ;
  assign n14444 = ( ~n13907 & n13911 ) | ( ~n13907 & n14443 ) | ( n13911 & n14443 ) ;
  assign n14445 = n14442 | n14444 ;
  assign n14446 = n14442 & n14444 ;
  assign n14447 = n14445 & ~n14446 ;
  assign n14448 = n1826 & ~n4429 ;
  assign n14449 = n1823 & n4396 ;
  assign n14450 = n14448 | n14449 ;
  assign n14451 = n1829 & n4245 ;
  assign n14452 = ( n1829 & n4303 ) | ( n1829 & n14451 ) | ( n4303 & n14451 ) ;
  assign n14454 = n1821 | n14452 ;
  assign n14455 = n14450 | n14454 ;
  assign n14453 = n14450 | n14452 ;
  assign n14456 = n14453 & n14455 ;
  assign n14457 = ( n4455 & n14455 ) | ( n4455 & n14456 ) | ( n14455 & n14456 ) ;
  assign n14458 = x29 & n14456 ;
  assign n14459 = x29 & n14455 ;
  assign n14460 = ( n4455 & n14458 ) | ( n4455 & n14459 ) | ( n14458 & n14459 ) ;
  assign n14461 = x29 & ~n14458 ;
  assign n14462 = x29 & ~n14459 ;
  assign n14463 = ( ~n4455 & n14461 ) | ( ~n4455 & n14462 ) | ( n14461 & n14462 ) ;
  assign n14464 = ( n14457 & ~n14460 ) | ( n14457 & n14463 ) | ( ~n14460 & n14463 ) ;
  assign n14465 = n14447 & n14464 ;
  assign n14466 = n14447 | n14464 ;
  assign n14467 = ~n14465 & n14466 ;
  assign n14468 = n13993 | n14012 ;
  assign n14469 = ( n13993 & n13996 ) | ( n13993 & n14468 ) | ( n13996 & n14468 ) ;
  assign n14470 = n14467 & n14469 ;
  assign n14471 = n14467 | n14469 ;
  assign n14472 = ~n14470 & n14471 ;
  assign n14473 = n2308 & n5117 ;
  assign n14474 = ( n2308 & ~n5037 ) | ( n2308 & n14473 ) | ( ~n5037 & n14473 ) ;
  assign n14475 = n2315 & n5108 ;
  assign n14476 = n2312 & n5192 ;
  assign n14477 = ( n2312 & n5179 ) | ( n2312 & n14476 ) | ( n5179 & n14476 ) ;
  assign n14478 = n14475 | n14477 ;
  assign n14479 = n14474 | n14478 ;
  assign n14480 = n2306 | n14479 ;
  assign n14481 = ( ~n5220 & n14479 ) | ( ~n5220 & n14480 ) | ( n14479 & n14480 ) ;
  assign n14482 = ~x26 & n14480 ;
  assign n14483 = ~x26 & n14479 ;
  assign n14484 = ( ~n5220 & n14482 ) | ( ~n5220 & n14483 ) | ( n14482 & n14483 ) ;
  assign n14485 = x26 | n14482 ;
  assign n14486 = x26 | n14483 ;
  assign n14487 = ( ~n5220 & n14485 ) | ( ~n5220 & n14486 ) | ( n14485 & n14486 ) ;
  assign n14488 = ( ~n14481 & n14484 ) | ( ~n14481 & n14487 ) | ( n14484 & n14487 ) ;
  assign n14489 = n14472 & ~n14488 ;
  assign n14490 = n14472 | n14488 ;
  assign n14491 = ( ~n14472 & n14489 ) | ( ~n14472 & n14490 ) | ( n14489 & n14490 ) ;
  assign n14492 = n14036 | n14067 ;
  assign n14493 = ( n14036 & n14040 ) | ( n14036 & n14492 ) | ( n14040 & n14492 ) ;
  assign n14494 = n14491 & n14493 ;
  assign n14495 = n14491 | n14493 ;
  assign n14496 = ~n14494 & n14495 ;
  assign n14497 = n2928 & n5857 ;
  assign n14498 = ( n2928 & ~n5899 ) | ( n2928 & n14497 ) | ( ~n5899 & n14497 ) ;
  assign n14499 = n2932 & ~n6091 ;
  assign n14500 = n2925 & n5997 ;
  assign n14501 = ( n2925 & n5979 ) | ( n2925 & n14500 ) | ( n5979 & n14500 ) ;
  assign n14502 = n14499 | n14501 ;
  assign n14503 = n14498 | n14502 ;
  assign n14504 = n2936 | n14503 ;
  assign n14505 = ( n6108 & n14503 ) | ( n6108 & n14504 ) | ( n14503 & n14504 ) ;
  assign n14506 = x23 & n14504 ;
  assign n14507 = x23 & n14503 ;
  assign n14508 = ( n6108 & n14506 ) | ( n6108 & n14507 ) | ( n14506 & n14507 ) ;
  assign n14509 = x23 & ~n14506 ;
  assign n14510 = x23 & ~n14507 ;
  assign n14511 = ( ~n6108 & n14509 ) | ( ~n6108 & n14510 ) | ( n14509 & n14510 ) ;
  assign n14512 = ( n14505 & ~n14508 ) | ( n14505 & n14511 ) | ( ~n14508 & n14511 ) ;
  assign n14513 = n14496 & ~n14512 ;
  assign n14514 = n14496 | n14512 ;
  assign n14515 = ( ~n14496 & n14513 ) | ( ~n14496 & n14514 ) | ( n14513 & n14514 ) ;
  assign n14516 = n14087 | n14115 ;
  assign n14517 = ( n14087 & n14089 ) | ( n14087 & n14516 ) | ( n14089 & n14516 ) ;
  assign n14518 = n14515 & n14517 ;
  assign n14519 = n14515 | n14517 ;
  assign n14520 = ~n14518 & n14519 ;
  assign n14521 = n3541 & n6950 ;
  assign n14522 = n3544 & n7036 ;
  assign n14523 = ( n3544 & n7023 ) | ( n3544 & n14522 ) | ( n7023 & n14522 ) ;
  assign n14524 = n14521 | n14523 ;
  assign n14525 = n3547 & n6889 ;
  assign n14526 = ( n3547 & ~n6884 ) | ( n3547 & n14525 ) | ( ~n6884 & n14525 ) ;
  assign n14527 = n14524 | n14526 ;
  assign n14528 = n3537 | n14526 ;
  assign n14529 = n14524 | n14528 ;
  assign n14530 = ( ~n7061 & n14527 ) | ( ~n7061 & n14529 ) | ( n14527 & n14529 ) ;
  assign n14531 = ~x20 & n14529 ;
  assign n14532 = ~x20 & n14527 ;
  assign n14533 = ( ~n7061 & n14531 ) | ( ~n7061 & n14532 ) | ( n14531 & n14532 ) ;
  assign n14534 = x20 | n14532 ;
  assign n14535 = x20 | n14531 ;
  assign n14536 = ( ~n7061 & n14534 ) | ( ~n7061 & n14535 ) | ( n14534 & n14535 ) ;
  assign n14537 = ( ~n14530 & n14533 ) | ( ~n14530 & n14536 ) | ( n14533 & n14536 ) ;
  assign n14538 = n14520 & ~n14537 ;
  assign n14539 = n14520 | n14537 ;
  assign n14540 = ( ~n14520 & n14538 ) | ( ~n14520 & n14539 ) | ( n14538 & n14539 ) ;
  assign n14541 = n14135 | n14163 ;
  assign n14542 = ( n14135 & n14137 ) | ( n14135 & n14541 ) | ( n14137 & n14541 ) ;
  assign n14543 = n14540 & n14542 ;
  assign n14544 = n14540 | n14542 ;
  assign n14545 = ~n14543 & n14544 ;
  assign n14546 = n4466 & n7907 ;
  assign n14547 = ( n4466 & n7902 ) | ( n4466 & n14546 ) | ( n7902 & n14546 ) ;
  assign n14548 = n4468 & n8079 ;
  assign n14549 = ( n4468 & ~n8070 ) | ( n4468 & n14548 ) | ( ~n8070 & n14548 ) ;
  assign n14550 = n14547 | n14549 ;
  assign n14551 = n4471 & ~n8017 ;
  assign n14552 = n14550 | n14551 ;
  assign n14553 = n4475 | n14550 ;
  assign n14554 = n14551 | n14553 ;
  assign n14555 = ( n8104 & n14552 ) | ( n8104 & n14554 ) | ( n14552 & n14554 ) ;
  assign n14556 = x17 & n14554 ;
  assign n14557 = x17 & n14552 ;
  assign n14558 = ( n8104 & n14556 ) | ( n8104 & n14557 ) | ( n14556 & n14557 ) ;
  assign n14559 = x17 & ~n14557 ;
  assign n14560 = x17 & ~n14556 ;
  assign n14561 = ( ~n8104 & n14559 ) | ( ~n8104 & n14560 ) | ( n14559 & n14560 ) ;
  assign n14562 = ( n14555 & ~n14558 ) | ( n14555 & n14561 ) | ( ~n14558 & n14561 ) ;
  assign n14563 = n14545 & ~n14562 ;
  assign n14564 = n14545 | n14562 ;
  assign n14565 = ( ~n14545 & n14563 ) | ( ~n14545 & n14564 ) | ( n14563 & n14564 ) ;
  assign n14566 = n14351 & n14565 ;
  assign n14567 = n14351 | n14565 ;
  assign n14568 = ~n14566 & n14567 ;
  assign n14569 = n14263 & n14568 ;
  assign n14570 = ( n14267 & n14568 ) | ( n14267 & n14569 ) | ( n14568 & n14569 ) ;
  assign n14571 = n14263 | n14568 ;
  assign n14572 = n14267 | n14571 ;
  assign n14573 = ~n14570 & n14572 ;
  assign n14574 = n14299 | n14313 ;
  assign n14575 = n14573 & n14574 ;
  assign n14576 = n14299 | n14316 ;
  assign n14577 = n14573 & n14576 ;
  assign n14578 = ( n13511 & n14575 ) | ( n13511 & n14577 ) | ( n14575 & n14577 ) ;
  assign n14579 = n14299 & n14573 ;
  assign n14580 = ( n14318 & n14573 ) | ( n14318 & n14579 ) | ( n14573 & n14579 ) ;
  assign n14581 = ( n12928 & n14578 ) | ( n12928 & n14580 ) | ( n14578 & n14580 ) ;
  assign n14582 = ( n12930 & n14578 ) | ( n12930 & n14580 ) | ( n14578 & n14580 ) ;
  assign n14583 = ( n11360 & n14581 ) | ( n11360 & n14582 ) | ( n14581 & n14582 ) ;
  assign n14584 = n14299 | n14318 ;
  assign n14585 = ( n13511 & n14574 ) | ( n13511 & n14576 ) | ( n14574 & n14576 ) ;
  assign n14586 = ( n12930 & n14584 ) | ( n12930 & n14585 ) | ( n14584 & n14585 ) ;
  assign n14587 = n14573 | n14586 ;
  assign n14588 = ( n12928 & n14584 ) | ( n12928 & n14585 ) | ( n14584 & n14585 ) ;
  assign n14589 = n14573 | n14588 ;
  assign n14590 = ( n11360 & n14587 ) | ( n11360 & n14589 ) | ( n14587 & n14589 ) ;
  assign n14591 = ~n14583 & n14590 ;
  assign n14592 = n14329 & n14591 ;
  assign n14593 = n14329 | n14591 ;
  assign n14594 = ~n14592 & n14593 ;
  assign n14595 = ( n13511 & n14311 ) | ( n13511 & n14314 ) | ( n14311 & n14314 ) ;
  assign n14596 = ( n13510 & n14311 ) | ( n13510 & n14314 ) | ( n14311 & n14314 ) ;
  assign n14597 = ( n12928 & n14595 ) | ( n12928 & n14596 ) | ( n14595 & n14596 ) ;
  assign n14598 = ( n12930 & n14595 ) | ( n12930 & n14596 ) | ( n14595 & n14596 ) ;
  assign n14599 = ( n11360 & n14597 ) | ( n11360 & n14598 ) | ( n14597 & n14598 ) ;
  assign n14600 = ( n13505 & n13511 ) | ( n13505 & n14310 ) | ( n13511 & n14310 ) ;
  assign n14601 = ( n13505 & n13510 ) | ( n13505 & n14310 ) | ( n13510 & n14310 ) ;
  assign n14602 = ( n12930 & n14600 ) | ( n12930 & n14601 ) | ( n14600 & n14601 ) ;
  assign n14603 = n14309 | n14602 ;
  assign n14604 = ( n12928 & n14600 ) | ( n12928 & n14601 ) | ( n14600 & n14601 ) ;
  assign n14605 = n14309 | n14604 ;
  assign n14606 = ( n11360 & n14603 ) | ( n11360 & n14605 ) | ( n14603 & n14605 ) ;
  assign n14607 = ~n14599 & n14606 ;
  assign n14608 = n14329 & n14607 ;
  assign n14609 = n14594 & n14608 ;
  assign n14610 = n14329 | n14607 ;
  assign n14611 = ~n14608 & n14610 ;
  assign n14612 = n13522 & n14607 ;
  assign n14613 = n13522 | n14607 ;
  assign n14614 = ~n14612 & n14613 ;
  assign n14615 = n13523 | n14612 ;
  assign n14616 = ( n14612 & n14614 ) | ( n14612 & n14615 ) | ( n14614 & n14615 ) ;
  assign n14617 = n14611 & n14616 ;
  assign n14618 = n14612 | n14614 ;
  assign n14619 = n14611 & n14618 ;
  assign n14620 = ( n13527 & n14617 ) | ( n13527 & n14619 ) | ( n14617 & n14619 ) ;
  assign n14621 = ( n14594 & n14609 ) | ( n14594 & n14620 ) | ( n14609 & n14620 ) ;
  assign n14622 = ( n13525 & n14617 ) | ( n13525 & n14619 ) | ( n14617 & n14619 ) ;
  assign n14623 = ( n14594 & n14609 ) | ( n14594 & n14622 ) | ( n14609 & n14622 ) ;
  assign n14624 = ( n13248 & n14621 ) | ( n13248 & n14623 ) | ( n14621 & n14623 ) ;
  assign n14625 = n14594 | n14608 ;
  assign n14626 = n14620 | n14625 ;
  assign n14627 = n14622 | n14625 ;
  assign n14628 = ( n13248 & n14626 ) | ( n13248 & n14627 ) | ( n14626 & n14627 ) ;
  assign n14629 = ~n14624 & n14628 ;
  assign n14631 = n3544 & n14607 ;
  assign n14632 = n3541 & n14329 ;
  assign n14633 = n14631 | n14632 ;
  assign n14630 = n3547 & n14591 ;
  assign n14635 = n3537 | n14630 ;
  assign n14636 = n14633 | n14635 ;
  assign n14634 = n14630 | n14633 ;
  assign n14637 = n14634 & n14636 ;
  assign n14638 = ( n14629 & n14636 ) | ( n14629 & n14637 ) | ( n14636 & n14637 ) ;
  assign n14639 = x20 & n14637 ;
  assign n14640 = x20 & n14636 ;
  assign n14641 = ( n14629 & n14639 ) | ( n14629 & n14640 ) | ( n14639 & n14640 ) ;
  assign n14642 = x20 & ~n14639 ;
  assign n14643 = x20 & ~n14640 ;
  assign n14644 = ( ~n14629 & n14642 ) | ( ~n14629 & n14643 ) | ( n14642 & n14643 ) ;
  assign n14645 = ( n14638 & ~n14641 ) | ( n14638 & n14644 ) | ( ~n14641 & n14644 ) ;
  assign n14646 = ~n13825 & n14645 ;
  assign n14647 = n13818 & n13820 ;
  assign n14648 = n13818 | n13820 ;
  assign n14649 = ~n14647 & n14648 ;
  assign n14650 = ( n13248 & n14620 ) | ( n13248 & n14622 ) | ( n14620 & n14622 ) ;
  assign n14651 = ( n13527 & n14616 ) | ( n13527 & n14618 ) | ( n14616 & n14618 ) ;
  assign n14652 = n14611 | n14651 ;
  assign n14653 = ( n13525 & n14616 ) | ( n13525 & n14618 ) | ( n14616 & n14618 ) ;
  assign n14654 = n14611 | n14653 ;
  assign n14655 = ( n13248 & n14652 ) | ( n13248 & n14654 ) | ( n14652 & n14654 ) ;
  assign n14656 = ~n14650 & n14655 ;
  assign n14658 = n3544 & n13522 ;
  assign n14659 = n3541 & n14607 ;
  assign n14660 = n14658 | n14659 ;
  assign n14657 = n3547 & n14329 ;
  assign n14662 = n3537 | n14657 ;
  assign n14663 = n14660 | n14662 ;
  assign n14661 = n14657 | n14660 ;
  assign n14664 = n14661 & n14663 ;
  assign n14665 = ( n14656 & n14663 ) | ( n14656 & n14664 ) | ( n14663 & n14664 ) ;
  assign n14666 = x20 & n14664 ;
  assign n14667 = x20 & n14663 ;
  assign n14668 = ( n14656 & n14666 ) | ( n14656 & n14667 ) | ( n14666 & n14667 ) ;
  assign n14669 = x20 & ~n14666 ;
  assign n14670 = x20 & ~n14667 ;
  assign n14671 = ( ~n14656 & n14669 ) | ( ~n14656 & n14670 ) | ( n14669 & n14670 ) ;
  assign n14672 = ( n14665 & ~n14668 ) | ( n14665 & n14671 ) | ( ~n14668 & n14671 ) ;
  assign n14673 = n14649 & n14672 ;
  assign n14674 = n14649 & ~n14673 ;
  assign n14675 = ~n14649 & n14672 ;
  assign n14676 = n14674 | n14675 ;
  assign n14677 = ~n13605 & n13816 ;
  assign n14678 = n13605 & ~n13816 ;
  assign n14679 = n14677 | n14678 ;
  assign n14680 = n13523 | n13525 ;
  assign n14681 = n13523 | n13527 ;
  assign n14682 = ( n13248 & n14680 ) | ( n13248 & n14681 ) | ( n14680 & n14681 ) ;
  assign n14683 = n13523 & n14614 ;
  assign n14684 = ( n13525 & n14614 ) | ( n13525 & n14683 ) | ( n14614 & n14683 ) ;
  assign n14685 = ( n13527 & n14614 ) | ( n13527 & n14683 ) | ( n14614 & n14683 ) ;
  assign n14686 = ( n13248 & n14684 ) | ( n13248 & n14685 ) | ( n14684 & n14685 ) ;
  assign n14687 = n14682 & ~n14686 ;
  assign n14688 = n3544 & n13235 ;
  assign n14689 = n3541 & n13522 ;
  assign n14690 = n14688 | n14689 ;
  assign n14691 = n3547 & n14607 ;
  assign n14692 = n3537 | n14691 ;
  assign n14693 = n14690 | n14692 ;
  assign n14694 = n14690 | n14691 ;
  assign n14695 = n14613 & ~n14616 ;
  assign n14696 = ~n13527 & n14695 ;
  assign n14697 = n14694 | n14696 ;
  assign n14698 = ~n13525 & n14695 ;
  assign n14699 = n14694 | n14698 ;
  assign n14700 = ( ~n13248 & n14697 ) | ( ~n13248 & n14699 ) | ( n14697 & n14699 ) ;
  assign n14701 = n14693 & n14700 ;
  assign n14702 = ( n14687 & n14693 ) | ( n14687 & n14701 ) | ( n14693 & n14701 ) ;
  assign n14703 = ~x20 & n14702 ;
  assign n14704 = x20 | n14702 ;
  assign n14705 = ( ~n14702 & n14703 ) | ( ~n14702 & n14704 ) | ( n14703 & n14704 ) ;
  assign n14706 = ~n14679 & n14705 ;
  assign n14707 = n14679 | n14706 ;
  assign n14708 = n14679 & n14705 ;
  assign n14709 = n14707 & ~n14708 ;
  assign n14710 = ( n13810 & n13811 ) | ( n13810 & ~n13814 ) | ( n13811 & ~n13814 ) ;
  assign n14711 = n13625 | n13810 ;
  assign n14712 = n13814 & ~n14711 ;
  assign n14713 = n14710 | n14712 ;
  assign n14714 = n3544 & n12936 ;
  assign n14715 = n3541 & n13235 ;
  assign n14716 = n14714 | n14715 ;
  assign n14717 = n3547 & n13522 ;
  assign n14718 = n3537 | n14717 ;
  assign n14719 = n14716 | n14718 ;
  assign n14720 = n14716 | n14717 ;
  assign n14721 = n13537 | n14720 ;
  assign n14722 = n13539 | n14720 ;
  assign n14723 = ( ~n13248 & n14721 ) | ( ~n13248 & n14722 ) | ( n14721 & n14722 ) ;
  assign n14724 = n14719 & n14723 ;
  assign n14725 = ( n13530 & n14719 ) | ( n13530 & n14724 ) | ( n14719 & n14724 ) ;
  assign n14726 = ~x20 & n14725 ;
  assign n14727 = x20 | n14725 ;
  assign n14728 = ( ~n14725 & n14726 ) | ( ~n14725 & n14727 ) | ( n14726 & n14727 ) ;
  assign n14729 = ~n14713 & n14728 ;
  assign n14730 = n14713 | n14729 ;
  assign n14731 = n14713 & n14728 ;
  assign n14732 = n14730 & ~n14731 ;
  assign n14733 = n13806 & n13808 ;
  assign n14734 = n13806 | n13808 ;
  assign n14735 = ~n14733 & n14734 ;
  assign n14736 = n3547 & n13235 ;
  assign n14737 = n3544 & ~n12616 ;
  assign n14738 = n3541 & n12936 ;
  assign n14739 = n14737 | n14738 ;
  assign n14740 = n14736 | n14739 ;
  assign n14741 = n3537 | n14736 ;
  assign n14742 = n14739 | n14741 ;
  assign n14743 = ( n13561 & n14740 ) | ( n13561 & n14742 ) | ( n14740 & n14742 ) ;
  assign n14744 = x20 & n14742 ;
  assign n14745 = x20 & n14740 ;
  assign n14746 = ( n13561 & n14744 ) | ( n13561 & n14745 ) | ( n14744 & n14745 ) ;
  assign n14747 = x20 & ~n14745 ;
  assign n14748 = x20 & ~n14744 ;
  assign n14749 = ( ~n13561 & n14747 ) | ( ~n13561 & n14748 ) | ( n14747 & n14748 ) ;
  assign n14750 = ( n14743 & ~n14746 ) | ( n14743 & n14749 ) | ( ~n14746 & n14749 ) ;
  assign n14751 = n14735 & n14750 ;
  assign n14752 = ~n14735 & n14750 ;
  assign n14753 = ( n14735 & ~n14751 ) | ( n14735 & n14752 ) | ( ~n14751 & n14752 ) ;
  assign n14754 = ~n13662 & n13804 ;
  assign n14755 = n13662 & ~n13804 ;
  assign n14756 = n14754 | n14755 ;
  assign n14757 = n3547 & n12936 ;
  assign n14758 = n3544 & n12010 ;
  assign n14759 = n3541 & ~n12616 ;
  assign n14760 = n14758 | n14759 ;
  assign n14761 = n14757 | n14760 ;
  assign n14762 = n3537 | n14757 ;
  assign n14763 = n14760 | n14762 ;
  assign n14764 = ( ~n13591 & n14761 ) | ( ~n13591 & n14763 ) | ( n14761 & n14763 ) ;
  assign n14765 = ~x20 & n14763 ;
  assign n14766 = ~x20 & n14761 ;
  assign n14767 = ( ~n13591 & n14765 ) | ( ~n13591 & n14766 ) | ( n14765 & n14766 ) ;
  assign n14768 = x20 | n14766 ;
  assign n14769 = x20 | n14765 ;
  assign n14770 = ( ~n13591 & n14768 ) | ( ~n13591 & n14769 ) | ( n14768 & n14769 ) ;
  assign n14771 = ( ~n14764 & n14767 ) | ( ~n14764 & n14770 ) | ( n14767 & n14770 ) ;
  assign n14772 = n14756 & n14771 ;
  assign n14773 = n13800 & n13802 ;
  assign n14774 = n13800 | n13802 ;
  assign n14775 = ~n14773 & n14774 ;
  assign n14777 = n3544 & ~n11663 ;
  assign n14778 = n3541 & n12010 ;
  assign n14779 = n14777 | n14778 ;
  assign n14776 = n3547 & ~n12616 ;
  assign n14781 = n3537 | n14776 ;
  assign n14782 = n14779 | n14781 ;
  assign n14780 = n14776 | n14779 ;
  assign n14783 = n14780 & n14782 ;
  assign n14784 = ( ~n12626 & n14782 ) | ( ~n12626 & n14783 ) | ( n14782 & n14783 ) ;
  assign n14785 = ~x20 & n14783 ;
  assign n14786 = ~x20 & n14782 ;
  assign n14787 = ( ~n12626 & n14785 ) | ( ~n12626 & n14786 ) | ( n14785 & n14786 ) ;
  assign n14788 = x20 | n14785 ;
  assign n14789 = x20 | n14786 ;
  assign n14790 = ( ~n12626 & n14788 ) | ( ~n12626 & n14789 ) | ( n14788 & n14789 ) ;
  assign n14791 = ( ~n14784 & n14787 ) | ( ~n14784 & n14790 ) | ( n14787 & n14790 ) ;
  assign n14792 = n14775 & n14791 ;
  assign n14793 = n13701 | n13798 ;
  assign n14794 = ~n13799 & n14793 ;
  assign n14796 = n3544 & n11363 ;
  assign n14797 = n3541 & ~n11663 ;
  assign n14798 = n14796 | n14797 ;
  assign n14795 = n3547 & n12010 ;
  assign n14800 = n3537 | n14795 ;
  assign n14801 = n14798 | n14800 ;
  assign n14799 = n14795 | n14798 ;
  assign n14802 = n14799 & n14801 ;
  assign n14803 = ( ~n12028 & n14801 ) | ( ~n12028 & n14802 ) | ( n14801 & n14802 ) ;
  assign n14804 = n14801 | n14802 ;
  assign n14805 = ( n12017 & n14803 ) | ( n12017 & n14804 ) | ( n14803 & n14804 ) ;
  assign n14806 = ~x20 & n14805 ;
  assign n14807 = x20 | n14805 ;
  assign n14808 = ( ~n14805 & n14806 ) | ( ~n14805 & n14807 ) | ( n14806 & n14807 ) ;
  assign n14809 = n14794 & n14808 ;
  assign n14810 = n14794 & ~n14809 ;
  assign n14811 = ~n14794 & n14808 ;
  assign n14812 = n14810 | n14811 ;
  assign n14813 = n13725 | n13796 ;
  assign n14814 = ~n13797 & n14813 ;
  assign n14815 = n3544 & n10649 ;
  assign n14816 = n3541 & n11363 ;
  assign n14817 = n14815 | n14816 ;
  assign n14818 = n3547 & ~n11663 ;
  assign n14819 = n3537 | n14818 ;
  assign n14820 = n14817 | n14819 ;
  assign n14821 = n14817 | n14818 ;
  assign n14822 = n12048 & ~n14821 ;
  assign n14823 = ( n11672 & ~n14821 ) | ( n11672 & n14822 ) | ( ~n14821 & n14822 ) ;
  assign n14824 = n14820 & ~n14823 ;
  assign n14825 = ( n12040 & n14820 ) | ( n12040 & n14824 ) | ( n14820 & n14824 ) ;
  assign n14826 = x20 & n14825 ;
  assign n14827 = x20 & ~n14825 ;
  assign n14828 = ( n14825 & ~n14826 ) | ( n14825 & n14827 ) | ( ~n14826 & n14827 ) ;
  assign n14829 = n14814 & n14828 ;
  assign n14830 = n14814 & ~n14829 ;
  assign n14831 = ~n14814 & n14828 ;
  assign n14832 = n14830 | n14831 ;
  assign n14833 = n13792 & n13794 ;
  assign n14834 = n13792 | n13794 ;
  assign n14835 = ~n14833 & n14834 ;
  assign n14836 = n3547 & n11363 ;
  assign n14837 = n3544 & n10325 ;
  assign n14838 = n3541 & n10649 ;
  assign n14839 = n14837 | n14838 ;
  assign n14840 = n14836 | n14839 ;
  assign n14841 = n3537 | n14840 ;
  assign n14842 = ( n12059 & n14840 ) | ( n12059 & n14841 ) | ( n14840 & n14841 ) ;
  assign n14843 = x20 & n14841 ;
  assign n14844 = x20 & n14840 ;
  assign n14845 = ( n12059 & n14843 ) | ( n12059 & n14844 ) | ( n14843 & n14844 ) ;
  assign n14846 = x20 & ~n14843 ;
  assign n14847 = x20 & ~n14844 ;
  assign n14848 = ( ~n12059 & n14846 ) | ( ~n12059 & n14847 ) | ( n14846 & n14847 ) ;
  assign n14849 = ( n14842 & ~n14845 ) | ( n14842 & n14848 ) | ( ~n14845 & n14848 ) ;
  assign n14850 = n14835 & n14849 ;
  assign n14851 = n13779 & n13790 ;
  assign n14852 = n13779 & ~n14851 ;
  assign n14853 = n3547 & n10649 ;
  assign n14854 = n3544 & n10654 ;
  assign n14855 = n3541 & n10325 ;
  assign n14856 = n14854 | n14855 ;
  assign n14857 = n14853 | n14856 ;
  assign n14858 = n3537 | n14853 ;
  assign n14859 = n14856 | n14858 ;
  assign n14860 = ( n10702 & n14857 ) | ( n10702 & n14859 ) | ( n14857 & n14859 ) ;
  assign n14861 = n14857 | n14859 ;
  assign n14862 = ( n10695 & n14860 ) | ( n10695 & n14861 ) | ( n14860 & n14861 ) ;
  assign n14863 = x20 & n14862 ;
  assign n14864 = x20 & ~n14862 ;
  assign n14865 = ( n14862 & ~n14863 ) | ( n14862 & n14864 ) | ( ~n14863 & n14864 ) ;
  assign n14866 = ~n13779 & n13790 ;
  assign n14867 = n14865 & n14866 ;
  assign n14868 = ( n14852 & n14865 ) | ( n14852 & n14867 ) | ( n14865 & n14867 ) ;
  assign n14869 = n14865 | n14866 ;
  assign n14870 = n14852 | n14869 ;
  assign n14871 = ~n14868 & n14870 ;
  assign n14872 = n3547 & n10325 ;
  assign n14873 = n3544 & ~n10662 ;
  assign n14874 = n3541 & n10654 ;
  assign n14875 = n14873 | n14874 ;
  assign n14876 = n14872 | n14875 ;
  assign n14877 = n3537 | n14876 ;
  assign n14878 = ( ~n10957 & n14876 ) | ( ~n10957 & n14877 ) | ( n14876 & n14877 ) ;
  assign n14879 = n14876 | n14877 ;
  assign n14880 = ( n10949 & n14878 ) | ( n10949 & n14879 ) | ( n14878 & n14879 ) ;
  assign n14881 = ~x20 & n14880 ;
  assign n14882 = x20 & n14876 ;
  assign n14883 = x20 & n3537 ;
  assign n14884 = ( x20 & n14876 ) | ( x20 & n14883 ) | ( n14876 & n14883 ) ;
  assign n14885 = ( ~n10957 & n14882 ) | ( ~n10957 & n14884 ) | ( n14882 & n14884 ) ;
  assign n14886 = n14882 | n14884 ;
  assign n14887 = ( n10949 & n14885 ) | ( n10949 & n14886 ) | ( n14885 & n14886 ) ;
  assign n14888 = x20 & ~n14887 ;
  assign n14889 = n14881 | n14888 ;
  assign n14890 = n13758 & n13776 ;
  assign n14891 = n13758 | n13776 ;
  assign n14892 = ~n14890 & n14891 ;
  assign n14893 = n14889 & n14892 ;
  assign n14894 = n14889 | n14892 ;
  assign n14895 = ~n14893 & n14894 ;
  assign n14896 = n13751 | n13754 ;
  assign n14897 = ~n13754 & n13756 ;
  assign n14898 = ( n13752 & n14896 ) | ( n13752 & ~n14897 ) | ( n14896 & ~n14897 ) ;
  assign n14899 = ~n13758 & n14898 ;
  assign n14900 = n3547 & n10654 ;
  assign n14901 = n3544 & n10667 ;
  assign n14902 = n3541 & ~n10662 ;
  assign n14903 = n14901 | n14902 ;
  assign n14904 = n14900 | n14903 ;
  assign n14905 = n3537 | n14900 ;
  assign n14906 = n14903 | n14905 ;
  assign n14907 = ( n10978 & n14904 ) | ( n10978 & n14906 ) | ( n14904 & n14906 ) ;
  assign n14908 = x20 & n14906 ;
  assign n14909 = x20 & n14904 ;
  assign n14910 = ( n10978 & n14908 ) | ( n10978 & n14909 ) | ( n14908 & n14909 ) ;
  assign n14911 = x20 & ~n14909 ;
  assign n14912 = x20 & ~n14908 ;
  assign n14913 = ( ~n10978 & n14911 ) | ( ~n10978 & n14912 ) | ( n14911 & n14912 ) ;
  assign n14914 = ( n14907 & ~n14910 ) | ( n14907 & n14913 ) | ( ~n14910 & n14913 ) ;
  assign n14915 = n14899 & n14914 ;
  assign n14916 = n3537 & n10784 ;
  assign n14917 = n3541 & ~n10678 ;
  assign n14918 = n3547 & ~n10675 ;
  assign n14919 = n14917 | n14918 ;
  assign n14920 = x20 | n14919 ;
  assign n14921 = n14916 | n14920 ;
  assign n14922 = ~x20 & n14921 ;
  assign n14923 = x20 & ~n3536 ;
  assign n14924 = ( x20 & n10678 ) | ( x20 & n14923 ) | ( n10678 & n14923 ) ;
  assign n14925 = n14921 & n14924 ;
  assign n14926 = n14916 | n14919 ;
  assign n14927 = n14924 & ~n14926 ;
  assign n14928 = ( n14922 & n14925 ) | ( n14922 & n14927 ) | ( n14925 & n14927 ) ;
  assign n14929 = n3547 & n10667 ;
  assign n14930 = n3544 & ~n10678 ;
  assign n14931 = n3541 & ~n10675 ;
  assign n14932 = n14930 | n14931 ;
  assign n14933 = n14929 | n14932 ;
  assign n14934 = n10837 | n14933 ;
  assign n14935 = n3537 | n14929 ;
  assign n14936 = n14932 | n14935 ;
  assign n14937 = ~x20 & n14936 ;
  assign n14938 = n14934 & n14937 ;
  assign n14939 = x20 | n14938 ;
  assign n14940 = n2920 & ~n10678 ;
  assign n14941 = n14938 & n14940 ;
  assign n14942 = n14934 & n14936 ;
  assign n14943 = n14940 & ~n14942 ;
  assign n14944 = ( n14939 & n14941 ) | ( n14939 & n14943 ) | ( n14941 & n14943 ) ;
  assign n14945 = n14928 & n14944 ;
  assign n14946 = ( n14938 & n14939 ) | ( n14938 & ~n14942 ) | ( n14939 & ~n14942 ) ;
  assign n14947 = n14928 | n14940 ;
  assign n14948 = ( n14940 & n14946 ) | ( n14940 & n14947 ) | ( n14946 & n14947 ) ;
  assign n14949 = ~n14945 & n14948 ;
  assign n14950 = n3547 & ~n10662 ;
  assign n14951 = n3544 & ~n10675 ;
  assign n14952 = n3541 & n10667 ;
  assign n14953 = n14951 | n14952 ;
  assign n14954 = n14950 | n14953 ;
  assign n14955 = ( n3537 & n10850 ) | ( n3537 & n14954 ) | ( n10850 & n14954 ) ;
  assign n14956 = ( x20 & n3537 ) | ( x20 & ~n14954 ) | ( n3537 & ~n14954 ) ;
  assign n14957 = ( x20 & n10850 ) | ( x20 & n14956 ) | ( n10850 & n14956 ) ;
  assign n14958 = ~n14955 & n14957 ;
  assign n14959 = n14954 | n14957 ;
  assign n14960 = ( ~x20 & n14958 ) | ( ~x20 & n14959 ) | ( n14958 & n14959 ) ;
  assign n14961 = n14945 | n14960 ;
  assign n14962 = ( n14945 & n14949 ) | ( n14945 & n14961 ) | ( n14949 & n14961 ) ;
  assign n14963 = n14899 | n14914 ;
  assign n14964 = ~n14915 & n14963 ;
  assign n14965 = n14915 | n14964 ;
  assign n14966 = ( n14915 & n14962 ) | ( n14915 & n14965 ) | ( n14962 & n14965 ) ;
  assign n14967 = n14895 & n14966 ;
  assign n14968 = n14893 | n14967 ;
  assign n14969 = n14871 & n14968 ;
  assign n14970 = n14868 | n14969 ;
  assign n14971 = ~n14835 & n14849 ;
  assign n14972 = ( n14835 & ~n14850 ) | ( n14835 & n14971 ) | ( ~n14850 & n14971 ) ;
  assign n14973 = n14850 | n14972 ;
  assign n14974 = ( n14850 & n14970 ) | ( n14850 & n14973 ) | ( n14970 & n14973 ) ;
  assign n14975 = n14832 & n14974 ;
  assign n14976 = n14829 | n14975 ;
  assign n14977 = n14812 & n14976 ;
  assign n14978 = n14809 | n14977 ;
  assign n14979 = n14775 | n14791 ;
  assign n14980 = ~n14792 & n14979 ;
  assign n14981 = n14792 | n14980 ;
  assign n14982 = ( n14792 & n14978 ) | ( n14792 & n14981 ) | ( n14978 & n14981 ) ;
  assign n14983 = n14756 | n14771 ;
  assign n14984 = ~n14772 & n14983 ;
  assign n14985 = n14772 | n14984 ;
  assign n14986 = ( n14772 & n14982 ) | ( n14772 & n14985 ) | ( n14982 & n14985 ) ;
  assign n14987 = n14753 & n14986 ;
  assign n14988 = n14751 | n14987 ;
  assign n14989 = n14729 | n14988 ;
  assign n14990 = ( n14729 & ~n14732 ) | ( n14729 & n14989 ) | ( ~n14732 & n14989 ) ;
  assign n14991 = n14706 | n14990 ;
  assign n14992 = ( n14706 & ~n14709 ) | ( n14706 & n14991 ) | ( ~n14709 & n14991 ) ;
  assign n14993 = n14676 & n14992 ;
  assign n14994 = n14673 | n14993 ;
  assign n14995 = n13825 | n14646 ;
  assign n14996 = n13825 & n14645 ;
  assign n14997 = n14995 & ~n14996 ;
  assign n14998 = n14994 & ~n14997 ;
  assign n14999 = n14646 | n14998 ;
  assign n15000 = n1829 & ~n11663 ;
  assign n15001 = n1826 & n10649 ;
  assign n15002 = n1823 & n11363 ;
  assign n15003 = n15001 | n15002 ;
  assign n15004 = n15000 | n15003 ;
  assign n15005 = n1821 & ~n12048 ;
  assign n15006 = ~n11672 & n15005 ;
  assign n15007 = n15004 | n15006 ;
  assign n15008 = n1821 | n15004 ;
  assign n15009 = ( n12040 & n15007 ) | ( n12040 & n15008 ) | ( n15007 & n15008 ) ;
  assign n15010 = x29 | n15009 ;
  assign n15011 = ~x29 & n15009 ;
  assign n15012 = ( ~n15009 & n15010 ) | ( ~n15009 & n15011 ) | ( n15010 & n15011 ) ;
  assign n15013 = n1057 & n10325 ;
  assign n15014 = n1065 & n10654 ;
  assign n15015 = n1060 & ~n10662 ;
  assign n15016 = n15014 | n15015 ;
  assign n15017 = n15013 | n15016 ;
  assign n15018 = n1062 | n15016 ;
  assign n15019 = n15013 | n15018 ;
  assign n15020 = ( ~n10957 & n15017 ) | ( ~n10957 & n15019 ) | ( n15017 & n15019 ) ;
  assign n15021 = n15017 | n15019 ;
  assign n15022 = ( n10949 & n15020 ) | ( n10949 & n15021 ) | ( n15020 & n15021 ) ;
  assign n15023 = n711 | n4179 ;
  assign n15024 = n573 | n2789 ;
  assign n15025 = n2033 & ~n15024 ;
  assign n15026 = n748 | n3502 ;
  assign n15027 = n489 | n15026 ;
  assign n15028 = n15025 & ~n15027 ;
  assign n15029 = n83 | n369 ;
  assign n15030 = n401 | n15029 ;
  assign n15031 = n178 | n1039 ;
  assign n15032 = n887 | n15031 ;
  assign n15033 = n15030 | n15032 ;
  assign n15034 = n468 | n3986 ;
  assign n15035 = n15033 | n15034 ;
  assign n15036 = n4293 | n15035 ;
  assign n15037 = n15028 & ~n15036 ;
  assign n15038 = ~n15023 & n15037 ;
  assign n15039 = n1349 | n1460 ;
  assign n15040 = n314 | n966 ;
  assign n15041 = n15039 | n15040 ;
  assign n15042 = n306 | n441 ;
  assign n15043 = n349 | n15042 ;
  assign n15044 = n560 | n15043 ;
  assign n15045 = n15041 | n15044 ;
  assign n15046 = n15038 & ~n15045 ;
  assign n15047 = n96 | n581 ;
  assign n15048 = n2720 | n15047 ;
  assign n15049 = n1384 | n3296 ;
  assign n15050 = n15048 | n15049 ;
  assign n15051 = n189 | n477 ;
  assign n15052 = n484 | n15051 ;
  assign n15053 = n15050 | n15052 ;
  assign n15054 = n341 | n383 ;
  assign n15055 = n196 | n435 ;
  assign n15056 = n15054 | n15055 ;
  assign n15057 = n347 | n15056 ;
  assign n15058 = n15053 | n15057 ;
  assign n15059 = n229 | n365 ;
  assign n15060 = n2714 | n15059 ;
  assign n15061 = n407 | n15060 ;
  assign n15062 = n5913 | n11760 ;
  assign n15063 = n849 | n1124 ;
  assign n15064 = n796 | n15063 ;
  assign n15065 = n15062 | n15064 ;
  assign n15066 = n140 | n177 ;
  assign n15067 = n193 | n527 ;
  assign n15068 = n15066 | n15067 ;
  assign n15069 = n7876 | n15068 ;
  assign n15070 = n15065 | n15069 ;
  assign n15071 = ( n15058 & n15061 ) | ( n15058 & ~n15070 ) | ( n15061 & ~n15070 ) ;
  assign n15072 = n2053 | n15070 ;
  assign n15073 = n15071 | n15072 ;
  assign n15074 = n1304 | n15073 ;
  assign n15075 = n15046 & ~n15074 ;
  assign n15076 = n114 | n202 ;
  assign n15077 = n387 | n841 ;
  assign n15078 = n15076 | n15077 ;
  assign n15079 = n310 | n469 ;
  assign n15080 = n1114 | n15079 ;
  assign n15081 = n15078 | n15080 ;
  assign n15082 = n15075 & ~n15081 ;
  assign n15083 = n15017 & ~n15082 ;
  assign n15084 = n15013 & ~n15082 ;
  assign n15085 = ( n15018 & ~n15082 ) | ( n15018 & n15084 ) | ( ~n15082 & n15084 ) ;
  assign n15086 = ( ~n10957 & n15083 ) | ( ~n10957 & n15085 ) | ( n15083 & n15085 ) ;
  assign n15087 = n15083 | n15085 ;
  assign n15088 = ( n10949 & n15086 ) | ( n10949 & n15087 ) | ( n15086 & n15087 ) ;
  assign n15089 = n15022 & ~n15088 ;
  assign n15090 = n15022 | n15082 ;
  assign n15091 = ~n15089 & n15090 ;
  assign n15092 = ~n12304 & n12306 ;
  assign n15093 = n12299 | n15092 ;
  assign n15094 = n15091 & n15093 ;
  assign n15095 = n15091 | n15093 ;
  assign n15096 = ~n15094 & n15095 ;
  assign n15097 = n15012 & ~n15096 ;
  assign n15098 = n15012 & ~n15097 ;
  assign n15099 = n15096 | n15097 ;
  assign n15100 = ~n15098 & n15099 ;
  assign n15101 = ~n12310 & n12313 ;
  assign n15102 = ( n12310 & n12315 ) | ( n12310 & ~n15101 ) | ( n12315 & ~n15101 ) ;
  assign n15103 = ~n15100 & n15102 ;
  assign n15104 = n15100 & ~n15102 ;
  assign n15105 = n15103 | n15104 ;
  assign n15106 = n2315 & n12936 ;
  assign n15107 = n2312 & n12010 ;
  assign n15108 = n2308 & ~n12616 ;
  assign n15109 = n15107 | n15108 ;
  assign n15110 = n15106 | n15109 ;
  assign n15111 = n2306 | n15106 ;
  assign n15112 = n15109 | n15111 ;
  assign n15113 = ( ~n13591 & n15110 ) | ( ~n13591 & n15112 ) | ( n15110 & n15112 ) ;
  assign n15114 = ~x26 & n15112 ;
  assign n15115 = ~x26 & n15110 ;
  assign n15116 = ( ~n13591 & n15114 ) | ( ~n13591 & n15115 ) | ( n15114 & n15115 ) ;
  assign n15117 = x26 | n15115 ;
  assign n15118 = x26 | n15114 ;
  assign n15119 = ( ~n13591 & n15117 ) | ( ~n13591 & n15118 ) | ( n15117 & n15118 ) ;
  assign n15120 = ( ~n15113 & n15116 ) | ( ~n15113 & n15119 ) | ( n15116 & n15119 ) ;
  assign n15121 = ~n15105 & n15120 ;
  assign n15122 = n15105 | n15121 ;
  assign n15123 = n15105 & n15120 ;
  assign n15124 = n15122 & ~n15123 ;
  assign n15125 = ~n12643 & n12646 ;
  assign n15126 = ( n12223 & n12643 ) | ( n12223 & ~n15125 ) | ( n12643 & ~n15125 ) ;
  assign n15127 = n15124 | n15126 ;
  assign n15128 = n15124 & n15126 ;
  assign n15129 = n15127 & ~n15128 ;
  assign n15130 = n2932 & n14607 ;
  assign n15131 = n2925 & n13235 ;
  assign n15132 = n2928 & n13522 ;
  assign n15133 = n15131 | n15132 ;
  assign n15134 = n15130 | n15133 ;
  assign n15135 = n2936 & n14696 ;
  assign n15136 = n2936 & n14698 ;
  assign n15137 = ( ~n13248 & n15135 ) | ( ~n13248 & n15136 ) | ( n15135 & n15136 ) ;
  assign n15138 = n15134 | n15137 ;
  assign n15139 = n2936 | n15134 ;
  assign n15140 = ( n14687 & n15138 ) | ( n14687 & n15139 ) | ( n15138 & n15139 ) ;
  assign n15141 = x23 | n15140 ;
  assign n15142 = ~x23 & n15140 ;
  assign n15143 = ( ~n15140 & n15141 ) | ( ~n15140 & n15142 ) | ( n15141 & n15142 ) ;
  assign n15144 = ~n15129 & n15143 ;
  assign n15145 = n15129 & ~n15143 ;
  assign n15146 = n15144 | n15145 ;
  assign n15147 = n13549 | n13822 ;
  assign n15148 = ( n13549 & ~n13553 ) | ( n13549 & n15147 ) | ( ~n13553 & n15147 ) ;
  assign n15149 = ~n15146 & n15148 ;
  assign n15150 = n15146 & ~n15148 ;
  assign n15151 = n15149 | n15150 ;
  assign n15152 = n5237 & ~n8982 ;
  assign n15153 = ( n5237 & n9051 ) | ( n5237 & n15152 ) | ( n9051 & n15152 ) ;
  assign n15154 = n5227 | n15153 ;
  assign n15155 = n9442 & ~n15153 ;
  assign n15156 = n9074 & ~n15153 ;
  assign n15157 = ( ~n9440 & n15155 ) | ( ~n9440 & n15156 ) | ( n15155 & n15156 ) ;
  assign n15158 = n15154 & ~n15157 ;
  assign n15159 = n15153 & n15154 ;
  assign n15160 = ( ~n9442 & n15154 ) | ( ~n9442 & n15159 ) | ( n15154 & n15159 ) ;
  assign n15161 = ( ~n9072 & n15158 ) | ( ~n9072 & n15160 ) | ( n15158 & n15160 ) ;
  assign n15162 = ~x14 & n15158 ;
  assign n15163 = ~x14 & n15160 ;
  assign n15164 = ( ~n9072 & n15162 ) | ( ~n9072 & n15163 ) | ( n15162 & n15163 ) ;
  assign n15165 = x14 | n15162 ;
  assign n15166 = x14 | n15163 ;
  assign n15167 = ( ~n9072 & n15165 ) | ( ~n9072 & n15166 ) | ( n15165 & n15166 ) ;
  assign n15168 = ( ~n15161 & n15164 ) | ( ~n15161 & n15167 ) | ( n15164 & n15167 ) ;
  assign n15169 = n14543 | n14562 ;
  assign n15170 = ( n14543 & n14545 ) | ( n14543 & n15169 ) | ( n14545 & n15169 ) ;
  assign n15171 = n15168 & n15170 ;
  assign n15172 = n15168 | n15170 ;
  assign n15173 = ~n15171 & n15172 ;
  assign n15174 = n1065 & n4206 ;
  assign n15175 = n1057 & ~n4429 ;
  assign n15176 = n1060 & n3439 ;
  assign n15177 = ( n1060 & ~n3420 ) | ( n1060 & n15176 ) | ( ~n3420 & n15176 ) ;
  assign n15178 = n15175 | n15177 ;
  assign n15179 = n15174 | n15178 ;
  assign n15180 = n1062 | n15174 ;
  assign n15181 = n15178 | n15180 ;
  assign n15182 = ( ~n4527 & n15179 ) | ( ~n4527 & n15181 ) | ( n15179 & n15181 ) ;
  assign n15183 = n192 | n476 ;
  assign n15184 = n325 | n623 ;
  assign n15185 = n15183 | n15184 ;
  assign n15186 = n126 | n15185 ;
  assign n15187 = n433 | n3983 ;
  assign n15188 = n644 | n15187 ;
  assign n15189 = n99 | n901 ;
  assign n15190 = n303 | n500 ;
  assign n15191 = n15189 | n15190 ;
  assign n15192 = n2066 | n15191 ;
  assign n15193 = n15188 | n15192 ;
  assign n15194 = n3312 | n15193 ;
  assign n15195 = n461 | n600 ;
  assign n15196 = n694 | n15195 ;
  assign n15197 = n806 | n1583 ;
  assign n15198 = n15196 | n15197 ;
  assign n15199 = n331 | n667 ;
  assign n15200 = n198 | n511 ;
  assign n15201 = n15199 | n15200 ;
  assign n15202 = n10379 | n15201 ;
  assign n15203 = n15198 | n15202 ;
  assign n15204 = n153 | n663 ;
  assign n15205 = n1250 | n15204 ;
  assign n15206 = n138 | n938 ;
  assign n15207 = n15205 | n15206 ;
  assign n15208 = n15203 | n15207 ;
  assign n15209 = n15194 | n15208 ;
  assign n15210 = n85 | n387 ;
  assign n15211 = n418 | n725 ;
  assign n15212 = n15210 | n15211 ;
  assign n15213 = n309 | n349 ;
  assign n15214 = n15212 | n15213 ;
  assign n15215 = n15209 | n15214 ;
  assign n15216 = n540 | n854 ;
  assign n15217 = n12248 | n15216 ;
  assign n15218 = n2856 | n4249 ;
  assign n15219 = n320 | n839 ;
  assign n15220 = n15218 | n15219 ;
  assign n15221 = n15217 | n15220 ;
  assign n15222 = n295 | n762 ;
  assign n15223 = ( ~n405 & n9150 ) | ( ~n405 & n15222 ) | ( n9150 & n15222 ) ;
  assign n15224 = n9150 & n15222 ;
  assign n15225 = ( ~n2118 & n15223 ) | ( ~n2118 & n15224 ) | ( n15223 & n15224 ) ;
  assign n15226 = n2119 | n15225 ;
  assign n15227 = ( ~n15214 & n15221 ) | ( ~n15214 & n15226 ) | ( n15221 & n15226 ) ;
  assign n15228 = n15221 & n15226 ;
  assign n15229 = ( ~n15209 & n15227 ) | ( ~n15209 & n15228 ) | ( n15227 & n15228 ) ;
  assign n15230 = n15215 | n15229 ;
  assign n15231 = n249 | n5891 ;
  assign n15232 = n413 | n448 ;
  assign n15233 = n6979 | n15232 ;
  assign n15234 = n161 | n821 ;
  assign n15235 = n110 | n1136 ;
  assign n15236 = n15234 | n15235 ;
  assign n15237 = n15233 | n15236 ;
  assign n15238 = n15231 | n15237 ;
  assign n15239 = n1465 | n2147 ;
  assign n15240 = n1124 | n11076 ;
  assign n15241 = n15239 | n15240 ;
  assign n15242 = n1663 | n15241 ;
  assign n15243 = n189 | n402 ;
  assign n15244 = n575 | n15243 ;
  assign n15245 = n356 | n399 ;
  assign n15246 = n141 | n15245 ;
  assign n15247 = n15244 | n15246 ;
  assign n15248 = n283 | n15247 ;
  assign n15249 = n15242 | n15248 ;
  assign n15250 = n15238 | n15249 ;
  assign n15251 = n2167 | n15250 ;
  assign n15252 = n53 | n317 ;
  assign n15253 = n4016 | n15252 ;
  assign n15254 = n170 | n205 ;
  assign n15255 = n560 | n15254 ;
  assign n15256 = n15253 | n15255 ;
  assign n15257 = n517 | n2051 ;
  assign n15258 = n1607 | n15257 ;
  assign n15259 = n15256 | n15258 ;
  assign n15260 = n314 | n648 ;
  assign n15261 = n416 | n15260 ;
  assign n15262 = n15259 | n15261 ;
  assign n15263 = n15251 | n15262 ;
  assign n15264 = n15230 | n15263 ;
  assign n15265 = n15186 | n15264 ;
  assign n15266 = n14432 & ~n15265 ;
  assign n15267 = ~n14432 & n15265 ;
  assign n15268 = n15266 | n15267 ;
  assign n15269 = n15181 & ~n15268 ;
  assign n15270 = n15179 & ~n15268 ;
  assign n15271 = ( ~n4527 & n15269 ) | ( ~n4527 & n15270 ) | ( n15269 & n15270 ) ;
  assign n15272 = n15182 & ~n15271 ;
  assign n15273 = n14359 & ~n14435 ;
  assign n15274 = n14433 | n15273 ;
  assign n15275 = n14357 & ~n14435 ;
  assign n15276 = n14433 | n15275 ;
  assign n15277 = ( ~n4220 & n15274 ) | ( ~n4220 & n15276 ) | ( n15274 & n15276 ) ;
  assign n15278 = n15267 | n15270 ;
  assign n15279 = n15266 | n15278 ;
  assign n15280 = n15267 | n15269 ;
  assign n15281 = n15266 | n15280 ;
  assign n15282 = ( ~n4527 & n15279 ) | ( ~n4527 & n15281 ) | ( n15279 & n15281 ) ;
  assign n15283 = n15277 & ~n15282 ;
  assign n15284 = ( n15272 & n15277 ) | ( n15272 & n15283 ) | ( n15277 & n15283 ) ;
  assign n15285 = ~n15277 & n15282 ;
  assign n15286 = ~n15272 & n15285 ;
  assign n15287 = n15284 | n15286 ;
  assign n15288 = n14445 & ~n14464 ;
  assign n15289 = ( n14445 & ~n14447 ) | ( n14445 & n15288 ) | ( ~n14447 & n15288 ) ;
  assign n15290 = n15287 | n15289 ;
  assign n15291 = n15287 & n15289 ;
  assign n15292 = n15290 & ~n15291 ;
  assign n15293 = n1826 & n4396 ;
  assign n15294 = n1823 & n4245 ;
  assign n15295 = ( n1823 & n4303 ) | ( n1823 & n15294 ) | ( n4303 & n15294 ) ;
  assign n15296 = n15293 | n15295 ;
  assign n15297 = n1829 & n5192 ;
  assign n15298 = ( n1829 & n5179 ) | ( n1829 & n15297 ) | ( n5179 & n15297 ) ;
  assign n15300 = n1821 | n15298 ;
  assign n15301 = n15296 | n15300 ;
  assign n15299 = n15296 | n15298 ;
  assign n15302 = n15299 & n15301 ;
  assign n15303 = ( n5306 & n15301 ) | ( n5306 & n15302 ) | ( n15301 & n15302 ) ;
  assign n15304 = x29 & n15302 ;
  assign n15305 = x29 & n15301 ;
  assign n15306 = ( n5306 & n15304 ) | ( n5306 & n15305 ) | ( n15304 & n15305 ) ;
  assign n15307 = x29 & ~n15304 ;
  assign n15308 = x29 & ~n15305 ;
  assign n15309 = ( ~n5306 & n15307 ) | ( ~n5306 & n15308 ) | ( n15307 & n15308 ) ;
  assign n15310 = ( n15303 & ~n15306 ) | ( n15303 & n15309 ) | ( ~n15306 & n15309 ) ;
  assign n15311 = n15292 & n15310 ;
  assign n15312 = n15292 | n15310 ;
  assign n15313 = ~n15311 & n15312 ;
  assign n15314 = n2312 & n5117 ;
  assign n15315 = ( n2312 & ~n5037 ) | ( n2312 & n15314 ) | ( ~n5037 & n15314 ) ;
  assign n15316 = n2308 & n5108 ;
  assign n15317 = n2315 & n5997 ;
  assign n15318 = ( n2315 & n5979 ) | ( n2315 & n15317 ) | ( n5979 & n15317 ) ;
  assign n15319 = n15316 | n15318 ;
  assign n15320 = n15315 | n15319 ;
  assign n15321 = n2306 | n15320 ;
  assign n15322 = ( n6181 & n15320 ) | ( n6181 & n15321 ) | ( n15320 & n15321 ) ;
  assign n15323 = x26 & n15321 ;
  assign n15324 = x26 & n15320 ;
  assign n15325 = ( n6181 & n15323 ) | ( n6181 & n15324 ) | ( n15323 & n15324 ) ;
  assign n15326 = x26 & ~n15323 ;
  assign n15327 = x26 & ~n15324 ;
  assign n15328 = ( ~n6181 & n15326 ) | ( ~n6181 & n15327 ) | ( n15326 & n15327 ) ;
  assign n15329 = ( n15322 & ~n15325 ) | ( n15322 & n15328 ) | ( ~n15325 & n15328 ) ;
  assign n15330 = n15313 & n15329 ;
  assign n15331 = n15313 & ~n15330 ;
  assign n15333 = n14470 | n14488 ;
  assign n15334 = ( n14470 & n14472 ) | ( n14470 & n15333 ) | ( n14472 & n15333 ) ;
  assign n15332 = ~n15313 & n15329 ;
  assign n15335 = n15332 & n15334 ;
  assign n15336 = ( n15331 & n15334 ) | ( n15331 & n15335 ) | ( n15334 & n15335 ) ;
  assign n15337 = n15332 | n15334 ;
  assign n15338 = n15331 | n15337 ;
  assign n15339 = ~n15336 & n15338 ;
  assign n15340 = n2925 & n5857 ;
  assign n15341 = ( n2925 & ~n5899 ) | ( n2925 & n15340 ) | ( ~n5899 & n15340 ) ;
  assign n15342 = n2928 & ~n6091 ;
  assign n15343 = n2932 & n7036 ;
  assign n15344 = ( n2932 & n7023 ) | ( n2932 & n15343 ) | ( n7023 & n15343 ) ;
  assign n15345 = n15342 | n15344 ;
  assign n15346 = n15341 | n15345 ;
  assign n15347 = n2936 | n15346 ;
  assign n15348 = ( n7136 & n15346 ) | ( n7136 & n15347 ) | ( n15346 & n15347 ) ;
  assign n15349 = x23 & n15347 ;
  assign n15350 = x23 & n15346 ;
  assign n15351 = ( n7136 & n15349 ) | ( n7136 & n15350 ) | ( n15349 & n15350 ) ;
  assign n15352 = x23 & ~n15349 ;
  assign n15353 = x23 & ~n15350 ;
  assign n15354 = ( ~n7136 & n15352 ) | ( ~n7136 & n15353 ) | ( n15352 & n15353 ) ;
  assign n15355 = ( n15348 & ~n15351 ) | ( n15348 & n15354 ) | ( ~n15351 & n15354 ) ;
  assign n15356 = n15339 & ~n15355 ;
  assign n15357 = n15339 | n15355 ;
  assign n15358 = ( ~n15339 & n15356 ) | ( ~n15339 & n15357 ) | ( n15356 & n15357 ) ;
  assign n15359 = n14494 | n14512 ;
  assign n15360 = ( n14494 & n14496 ) | ( n14494 & n15359 ) | ( n14496 & n15359 ) ;
  assign n15361 = n15358 & n15360 ;
  assign n15362 = n15358 | n15360 ;
  assign n15363 = ~n15361 & n15362 ;
  assign n15364 = n3544 & n6950 ;
  assign n15365 = n3541 & n6889 ;
  assign n15366 = ( n3541 & ~n6884 ) | ( n3541 & n15365 ) | ( ~n6884 & n15365 ) ;
  assign n15367 = n15364 | n15366 ;
  assign n15368 = n3547 & n7907 ;
  assign n15369 = ( n3547 & n7902 ) | ( n3547 & n15368 ) | ( n7902 & n15368 ) ;
  assign n15370 = n15367 | n15369 ;
  assign n15371 = n3537 | n15369 ;
  assign n15372 = n15367 | n15371 ;
  assign n15373 = ( ~n8193 & n15370 ) | ( ~n8193 & n15372 ) | ( n15370 & n15372 ) ;
  assign n15374 = ~x20 & n15372 ;
  assign n15375 = ~x20 & n15370 ;
  assign n15376 = ( ~n8193 & n15374 ) | ( ~n8193 & n15375 ) | ( n15374 & n15375 ) ;
  assign n15377 = x20 | n15375 ;
  assign n15378 = x20 | n15374 ;
  assign n15379 = ( ~n8193 & n15377 ) | ( ~n8193 & n15378 ) | ( n15377 & n15378 ) ;
  assign n15380 = ( ~n15373 & n15376 ) | ( ~n15373 & n15379 ) | ( n15376 & n15379 ) ;
  assign n15381 = n15363 & ~n15380 ;
  assign n15382 = n15363 | n15380 ;
  assign n15383 = ( ~n15363 & n15381 ) | ( ~n15363 & n15382 ) | ( n15381 & n15382 ) ;
  assign n15384 = n14518 | n14537 ;
  assign n15385 = ( n14518 & n14520 ) | ( n14518 & n15384 ) | ( n14520 & n15384 ) ;
  assign n15386 = n15383 & n15385 ;
  assign n15387 = n15383 | n15385 ;
  assign n15388 = ~n15386 & n15387 ;
  assign n15389 = n4466 & n8079 ;
  assign n15390 = ( n4466 & ~n8070 ) | ( n4466 & n15389 ) | ( ~n8070 & n15389 ) ;
  assign n15391 = n4468 | n15390 ;
  assign n15392 = ( ~n8017 & n15390 ) | ( ~n8017 & n15391 ) | ( n15390 & n15391 ) ;
  assign n15393 = n4471 & n9022 ;
  assign n15394 = ( n4471 & ~n9019 ) | ( n4471 & n15393 ) | ( ~n9019 & n15393 ) ;
  assign n15395 = n15392 | n15394 ;
  assign n15396 = n4475 | n15394 ;
  assign n15397 = n15392 | n15396 ;
  assign n15398 = ( ~n9416 & n15395 ) | ( ~n9416 & n15397 ) | ( n15395 & n15397 ) ;
  assign n15399 = ~x17 & n15397 ;
  assign n15400 = ~x17 & n15395 ;
  assign n15401 = ( ~n9416 & n15399 ) | ( ~n9416 & n15400 ) | ( n15399 & n15400 ) ;
  assign n15402 = x17 | n15400 ;
  assign n15403 = x17 | n15399 ;
  assign n15404 = ( ~n9416 & n15402 ) | ( ~n9416 & n15403 ) | ( n15402 & n15403 ) ;
  assign n15405 = ( ~n15398 & n15401 ) | ( ~n15398 & n15404 ) | ( n15401 & n15404 ) ;
  assign n15406 = n15388 & ~n15405 ;
  assign n15407 = n15388 | n15405 ;
  assign n15408 = ( ~n15388 & n15406 ) | ( ~n15388 & n15407 ) | ( n15406 & n15407 ) ;
  assign n15409 = n15173 & ~n15408 ;
  assign n15410 = n15173 | n15408 ;
  assign n15411 = ( ~n15173 & n15409 ) | ( ~n15173 & n15410 ) | ( n15409 & n15410 ) ;
  assign n15412 = n14347 | n14565 ;
  assign n15413 = ( n14347 & n14351 ) | ( n14347 & n15412 ) | ( n14351 & n15412 ) ;
  assign n15414 = n15411 & n15413 ;
  assign n15415 = n15411 | n15413 ;
  assign n15416 = ~n15414 & n15415 ;
  assign n15417 = n14570 & n15416 ;
  assign n15418 = ( n14578 & n15416 ) | ( n14578 & n15417 ) | ( n15416 & n15417 ) ;
  assign n15419 = n14570 | n14579 ;
  assign n15420 = n15416 & n15419 ;
  assign n15421 = n14570 | n14573 ;
  assign n15422 = n15416 & n15421 ;
  assign n15423 = ( n14318 & n15420 ) | ( n14318 & n15422 ) | ( n15420 & n15422 ) ;
  assign n15424 = ( n12928 & n15418 ) | ( n12928 & n15423 ) | ( n15418 & n15423 ) ;
  assign n15425 = ( n12930 & n15418 ) | ( n12930 & n15423 ) | ( n15418 & n15423 ) ;
  assign n15426 = ( n11360 & n15424 ) | ( n11360 & n15425 ) | ( n15424 & n15425 ) ;
  assign n15427 = n14570 | n14578 ;
  assign n15428 = ( n14318 & n15419 ) | ( n14318 & n15421 ) | ( n15419 & n15421 ) ;
  assign n15429 = ( n12930 & n15427 ) | ( n12930 & n15428 ) | ( n15427 & n15428 ) ;
  assign n15430 = n15416 | n15429 ;
  assign n15431 = ( n12928 & n15427 ) | ( n12928 & n15428 ) | ( n15427 & n15428 ) ;
  assign n15432 = n15416 | n15431 ;
  assign n15433 = ( n11360 & n15430 ) | ( n11360 & n15432 ) | ( n15430 & n15432 ) ;
  assign n15434 = ~n15426 & n15433 ;
  assign n15435 = n14591 & n15434 ;
  assign n15436 = n14591 | n15434 ;
  assign n15437 = n14592 & n15436 ;
  assign n15438 = ( n14594 & n15436 ) | ( n14594 & n15437 ) | ( n15436 & n15437 ) ;
  assign n15439 = ~n15435 & n15438 ;
  assign n15440 = n14592 | n14608 ;
  assign n15441 = ( n14592 & n14594 ) | ( n14592 & n15440 ) | ( n14594 & n15440 ) ;
  assign n15442 = ~n15435 & n15436 ;
  assign n15443 = n15441 & n15442 ;
  assign n15444 = ( n14620 & n15439 ) | ( n14620 & n15443 ) | ( n15439 & n15443 ) ;
  assign n15445 = ( n14622 & n15439 ) | ( n14622 & n15443 ) | ( n15439 & n15443 ) ;
  assign n15446 = ( n13248 & n15444 ) | ( n13248 & n15445 ) | ( n15444 & n15445 ) ;
  assign n15447 = n14592 | n14594 ;
  assign n15448 = ( n14620 & n15441 ) | ( n14620 & n15447 ) | ( n15441 & n15447 ) ;
  assign n15449 = ( n14622 & n15441 ) | ( n14622 & n15447 ) | ( n15441 & n15447 ) ;
  assign n15450 = ( n13248 & n15448 ) | ( n13248 & n15449 ) | ( n15448 & n15449 ) ;
  assign n15451 = ~n15446 & n15450 ;
  assign n15452 = n15442 & ~n15446 ;
  assign n15453 = n15451 | n15452 ;
  assign n15455 = n3544 & n14329 ;
  assign n15456 = n3541 & n14591 ;
  assign n15457 = n15455 | n15456 ;
  assign n15454 = n3547 & n15434 ;
  assign n15459 = n3537 | n15454 ;
  assign n15460 = n15457 | n15459 ;
  assign n15458 = n15454 | n15457 ;
  assign n15461 = n15458 & n15460 ;
  assign n15462 = ( n15453 & n15460 ) | ( n15453 & n15461 ) | ( n15460 & n15461 ) ;
  assign n15463 = x20 & n15461 ;
  assign n15464 = x20 & n15460 ;
  assign n15465 = ( n15453 & n15463 ) | ( n15453 & n15464 ) | ( n15463 & n15464 ) ;
  assign n15466 = x20 & ~n15463 ;
  assign n15467 = x20 & ~n15464 ;
  assign n15468 = ( ~n15453 & n15466 ) | ( ~n15453 & n15467 ) | ( n15466 & n15467 ) ;
  assign n15469 = ( n15462 & ~n15465 ) | ( n15462 & n15468 ) | ( ~n15465 & n15468 ) ;
  assign n15470 = ~n15151 & n15469 ;
  assign n15471 = n15151 | n15470 ;
  assign n15472 = n15151 & n15469 ;
  assign n15473 = n15471 & ~n15472 ;
  assign n15474 = n14999 & ~n15473 ;
  assign n15475 = n14999 & ~n15474 ;
  assign n15476 = n14999 | n15473 ;
  assign n15477 = ~n15475 & n15476 ;
  assign n15478 = n1065 & ~n4429 ;
  assign n15479 = n1060 | n1065 ;
  assign n15480 = ( n1060 & ~n4429 ) | ( n1060 & n15479 ) | ( ~n4429 & n15479 ) ;
  assign n15481 = ( n4206 & n15478 ) | ( n4206 & n15480 ) | ( n15478 & n15480 ) ;
  assign n15482 = n1057 & n4396 ;
  assign n15483 = n15481 | n15482 ;
  assign n15484 = n1062 | n15482 ;
  assign n15485 = n15481 | n15484 ;
  assign n15486 = ( ~n4501 & n15483 ) | ( ~n4501 & n15485 ) | ( n15483 & n15485 ) ;
  assign n15487 = n2024 | n4144 ;
  assign n15488 = n4000 | n15487 ;
  assign n15489 = n2768 | n4266 ;
  assign n15490 = n15488 | n15489 ;
  assign n15491 = n9117 | n15490 ;
  assign n15492 = n9147 | n15491 ;
  assign n15493 = n11734 | n15492 ;
  assign n15494 = n114 | n667 ;
  assign n15495 = n162 | n344 ;
  assign n15496 = n15494 | n15495 ;
  assign n15497 = n254 | n15496 ;
  assign n15498 = n1736 | n4311 ;
  assign n15499 = n2696 | n9151 ;
  assign n15500 = n179 | n15499 ;
  assign n15501 = n15498 | n15500 ;
  assign n15502 = n318 | n820 ;
  assign n15503 = n247 | n330 ;
  assign n15504 = n15502 | n15503 ;
  assign n15505 = n143 & ~n15504 ;
  assign n15506 = ~n15501 & n15505 ;
  assign n15507 = n721 | n12384 ;
  assign n15508 = n15506 & ~n15507 ;
  assign n15509 = n869 | n4197 ;
  assign n15510 = n15508 & ~n15509 ;
  assign n15511 = ~n15497 & n15510 ;
  assign n15512 = ~n15493 & n15511 ;
  assign n15513 = ~n14432 & n15512 ;
  assign n15514 = ( x14 & ~n14432 ) | ( x14 & n15512 ) | ( ~n14432 & n15512 ) ;
  assign n15515 = ~n15513 & n15514 ;
  assign n15516 = n14432 & ~n15512 ;
  assign n15517 = n15513 | n15516 ;
  assign n15518 = ~x14 & n15517 ;
  assign n15519 = n15515 | n15518 ;
  assign n15520 = n15278 & n15519 ;
  assign n15521 = n15280 & n15519 ;
  assign n15522 = ( ~n4527 & n15520 ) | ( ~n4527 & n15521 ) | ( n15520 & n15521 ) ;
  assign n15523 = n15278 | n15519 ;
  assign n15524 = n15280 | n15519 ;
  assign n15525 = ( ~n4527 & n15523 ) | ( ~n4527 & n15524 ) | ( n15523 & n15524 ) ;
  assign n15526 = ~n15522 & n15525 ;
  assign n15527 = n15486 & n15526 ;
  assign n15528 = n15526 & ~n15527 ;
  assign n15529 = ( n15486 & ~n15527 ) | ( n15486 & n15528 ) | ( ~n15527 & n15528 ) ;
  assign n15530 = n1826 & n4245 ;
  assign n15531 = ( n1826 & n4303 ) | ( n1826 & n15530 ) | ( n4303 & n15530 ) ;
  assign n15532 = n1823 & n5192 ;
  assign n15533 = ( n1823 & n5179 ) | ( n1823 & n15532 ) | ( n5179 & n15532 ) ;
  assign n15534 = n15531 | n15533 ;
  assign n15535 = n1829 & n5117 ;
  assign n15536 = ( n1829 & ~n5037 ) | ( n1829 & n15535 ) | ( ~n5037 & n15535 ) ;
  assign n15537 = n15534 | n15536 ;
  assign n15538 = n1821 | n15536 ;
  assign n15539 = n15534 | n15538 ;
  assign n15540 = ( ~n5270 & n15537 ) | ( ~n5270 & n15539 ) | ( n15537 & n15539 ) ;
  assign n15541 = ~x29 & n15539 ;
  assign n15542 = ~x29 & n15537 ;
  assign n15543 = ( ~n5270 & n15541 ) | ( ~n5270 & n15542 ) | ( n15541 & n15542 ) ;
  assign n15544 = x29 | n15542 ;
  assign n15545 = x29 | n15541 ;
  assign n15546 = ( ~n5270 & n15544 ) | ( ~n5270 & n15545 ) | ( n15544 & n15545 ) ;
  assign n15547 = ( ~n15540 & n15543 ) | ( ~n15540 & n15546 ) | ( n15543 & n15546 ) ;
  assign n15548 = ~n15527 & n15547 ;
  assign n15549 = n15486 & n15547 ;
  assign n15550 = ( n15528 & n15548 ) | ( n15528 & n15549 ) | ( n15548 & n15549 ) ;
  assign n15551 = n15529 & ~n15550 ;
  assign n15552 = n15527 & n15547 ;
  assign n15553 = ~n15486 & n15547 ;
  assign n15554 = ( ~n15528 & n15552 ) | ( ~n15528 & n15553 ) | ( n15552 & n15553 ) ;
  assign n15555 = n15551 | n15554 ;
  assign n15556 = ~n15284 & n15287 ;
  assign n15557 = ( ~n15284 & n15289 ) | ( ~n15284 & n15556 ) | ( n15289 & n15556 ) ;
  assign n15558 = n15555 & ~n15557 ;
  assign n15559 = n1060 & ~n4429 ;
  assign n15560 = n1065 & n4396 ;
  assign n15561 = n15559 | n15560 ;
  assign n15562 = n1057 & n4245 ;
  assign n15563 = ( n1057 & n4303 ) | ( n1057 & n15562 ) | ( n4303 & n15562 ) ;
  assign n15564 = n15561 | n15563 ;
  assign n15565 = n1062 | n15563 ;
  assign n15566 = n15561 | n15565 ;
  assign n15567 = ( n4455 & n15564 ) | ( n4455 & n15566 ) | ( n15564 & n15566 ) ;
  assign n15568 = n443 | n1232 ;
  assign n15569 = n5921 | n15568 ;
  assign n15570 = n1747 | n15569 ;
  assign n15571 = n204 | n15570 ;
  assign n15572 = n718 | n8971 ;
  assign n15573 = n11719 | n15572 ;
  assign n15574 = n2027 | n15573 ;
  assign n15575 = n54 | n1002 ;
  assign n15576 = n451 | n460 ;
  assign n15577 = n15575 | n15576 ;
  assign n15578 = n384 | n511 ;
  assign n15579 = n134 | n255 ;
  assign n15580 = n15578 | n15579 ;
  assign n15581 = n497 | n801 ;
  assign n15582 = n15580 | n15581 ;
  assign n15583 = n15577 | n15582 ;
  assign n15584 = n15574 | n15583 ;
  assign n15585 = n15571 | n15584 ;
  assign n15586 = n14412 | n15585 ;
  assign n15587 = n13862 | n14384 ;
  assign n15588 = n13288 | n15587 ;
  assign n15589 = n1770 | n2211 ;
  assign n15590 = n15588 | n15589 ;
  assign n15591 = n1685 | n15590 ;
  assign n15592 = n94 | n331 ;
  assign n15593 = n363 | n15592 ;
  assign n15594 = n504 | n784 ;
  assign n15595 = n264 | n1404 ;
  assign n15596 = n15594 | n15595 ;
  assign n15597 = n289 | n648 ;
  assign n15598 = n15596 | n15597 ;
  assign n15599 = n15593 | n15598 ;
  assign n15600 = n15591 | n15599 ;
  assign n15601 = n15586 | n15600 ;
  assign n15602 = n283 | n632 ;
  assign n15603 = n891 | n15602 ;
  assign n15604 = n890 | n15603 ;
  assign n15605 = n588 | n1460 ;
  assign n15606 = n510 | n15605 ;
  assign n15607 = n594 | n15606 ;
  assign n15608 = n15604 | n15607 ;
  assign n15609 = n183 | n402 ;
  assign n15610 = n607 | n694 ;
  assign n15611 = n15609 | n15610 ;
  assign n15612 = n413 | n517 ;
  assign n15613 = n245 | n15612 ;
  assign n15614 = n15611 | n15613 ;
  assign n15615 = n15608 | n15614 ;
  assign n15616 = n15601 | n15615 ;
  assign n15617 = n15514 | n15616 ;
  assign n15618 = n15514 & n15616 ;
  assign n15619 = n15617 & ~n15618 ;
  assign n15620 = n15566 & n15619 ;
  assign n15621 = n15564 & n15619 ;
  assign n15622 = ( n4455 & n15620 ) | ( n4455 & n15621 ) | ( n15620 & n15621 ) ;
  assign n15623 = n15619 & ~n15621 ;
  assign n15624 = n15619 & ~n15620 ;
  assign n15625 = ( ~n4455 & n15623 ) | ( ~n4455 & n15624 ) | ( n15623 & n15624 ) ;
  assign n15626 = ( n15567 & ~n15622 ) | ( n15567 & n15625 ) | ( ~n15622 & n15625 ) ;
  assign n15627 = n15486 | n15522 ;
  assign n15628 = ( n15522 & n15526 ) | ( n15522 & n15627 ) | ( n15526 & n15627 ) ;
  assign n15629 = n15626 & n15628 ;
  assign n15630 = n15626 | n15628 ;
  assign n15631 = ~n15629 & n15630 ;
  assign n15632 = n1823 & n5117 ;
  assign n15633 = ( n1823 & ~n5037 ) | ( n1823 & n15632 ) | ( ~n5037 & n15632 ) ;
  assign n15634 = n1829 & n5108 ;
  assign n15635 = n1826 & n5192 ;
  assign n15636 = ( n1826 & n5179 ) | ( n1826 & n15635 ) | ( n5179 & n15635 ) ;
  assign n15637 = n15634 | n15636 ;
  assign n15638 = n15633 | n15637 ;
  assign n15639 = n1821 | n15638 ;
  assign n15640 = n15638 & n15639 ;
  assign n15641 = ( ~n5220 & n15639 ) | ( ~n5220 & n15640 ) | ( n15639 & n15640 ) ;
  assign n15642 = ~x29 & n15640 ;
  assign n15643 = ~x29 & n15639 ;
  assign n15644 = ( ~n5220 & n15642 ) | ( ~n5220 & n15643 ) | ( n15642 & n15643 ) ;
  assign n15645 = x29 | n15642 ;
  assign n15646 = x29 | n15643 ;
  assign n15647 = ( ~n5220 & n15645 ) | ( ~n5220 & n15646 ) | ( n15645 & n15646 ) ;
  assign n15648 = ( ~n15641 & n15644 ) | ( ~n15641 & n15647 ) | ( n15644 & n15647 ) ;
  assign n15649 = n15631 & n15648 ;
  assign n15650 = n15631 | n15648 ;
  assign n15651 = ~n15649 & n15650 ;
  assign n15652 = n15550 & n15651 ;
  assign n15653 = ( n15558 & n15651 ) | ( n15558 & n15652 ) | ( n15651 & n15652 ) ;
  assign n15654 = n15550 | n15651 ;
  assign n15655 = n15558 | n15654 ;
  assign n15656 = ~n15653 & n15655 ;
  assign n15657 = n2308 & n5857 ;
  assign n15658 = ( n2308 & ~n5899 ) | ( n2308 & n15657 ) | ( ~n5899 & n15657 ) ;
  assign n15659 = n2315 & ~n6091 ;
  assign n15660 = n2312 & n5997 ;
  assign n15661 = ( n2312 & n5979 ) | ( n2312 & n15660 ) | ( n5979 & n15660 ) ;
  assign n15662 = n15659 | n15661 ;
  assign n15663 = n15658 | n15662 ;
  assign n15664 = n2306 | n15663 ;
  assign n15665 = ( n6108 & n15663 ) | ( n6108 & n15664 ) | ( n15663 & n15664 ) ;
  assign n15666 = x26 & n15664 ;
  assign n15667 = x26 & n15663 ;
  assign n15668 = ( n6108 & n15666 ) | ( n6108 & n15667 ) | ( n15666 & n15667 ) ;
  assign n15669 = x26 & ~n15666 ;
  assign n15670 = x26 & ~n15667 ;
  assign n15671 = ( ~n6108 & n15669 ) | ( ~n6108 & n15670 ) | ( n15669 & n15670 ) ;
  assign n15672 = ( n15665 & ~n15668 ) | ( n15665 & n15671 ) | ( ~n15668 & n15671 ) ;
  assign n15673 = n15656 & ~n15672 ;
  assign n15674 = n15656 | n15672 ;
  assign n15675 = ( ~n15656 & n15673 ) | ( ~n15656 & n15674 ) | ( n15673 & n15674 ) ;
  assign n15676 = ~n15555 & n15557 ;
  assign n15677 = n15558 | n15676 ;
  assign n15678 = n2312 & n5108 ;
  assign n15679 = n2308 & n5997 ;
  assign n15680 = ( n2308 & n5979 ) | ( n2308 & n15679 ) | ( n5979 & n15679 ) ;
  assign n15681 = n15678 | n15680 ;
  assign n15682 = n2315 & n5857 ;
  assign n15683 = ( n2315 & ~n5899 ) | ( n2315 & n15682 ) | ( ~n5899 & n15682 ) ;
  assign n15684 = n15681 | n15683 ;
  assign n15685 = n2306 | n15684 ;
  assign n15686 = n15684 & n15685 ;
  assign n15687 = ( ~n6151 & n15685 ) | ( ~n6151 & n15686 ) | ( n15685 & n15686 ) ;
  assign n15688 = ~x26 & n15686 ;
  assign n15689 = ~x26 & n15685 ;
  assign n15690 = ( ~n6151 & n15688 ) | ( ~n6151 & n15689 ) | ( n15688 & n15689 ) ;
  assign n15691 = x26 | n15688 ;
  assign n15692 = x26 | n15689 ;
  assign n15693 = ( ~n6151 & n15691 ) | ( ~n6151 & n15692 ) | ( n15691 & n15692 ) ;
  assign n15694 = ( ~n15687 & n15690 ) | ( ~n15687 & n15693 ) | ( n15690 & n15693 ) ;
  assign n15695 = ~n15677 & n15694 ;
  assign n15696 = n15677 & ~n15694 ;
  assign n15697 = n15695 | n15696 ;
  assign n15698 = n15311 | n15329 ;
  assign n15699 = ( n15311 & n15313 ) | ( n15311 & n15698 ) | ( n15313 & n15698 ) ;
  assign n15700 = ~n15697 & n15699 ;
  assign n15701 = n15695 | n15700 ;
  assign n15702 = n15675 & n15701 ;
  assign n15703 = n15675 | n15701 ;
  assign n15704 = ~n15702 & n15703 ;
  assign n15705 = n2928 & n6950 ;
  assign n15706 = n2925 & n7036 ;
  assign n15707 = ( n2925 & n7023 ) | ( n2925 & n15706 ) | ( n7023 & n15706 ) ;
  assign n15708 = n15705 | n15707 ;
  assign n15709 = n2932 & n6889 ;
  assign n15710 = ( n2932 & ~n6884 ) | ( n2932 & n15709 ) | ( ~n6884 & n15709 ) ;
  assign n15711 = n15708 | n15710 ;
  assign n15712 = n2936 | n15710 ;
  assign n15713 = n15708 | n15712 ;
  assign n15714 = ( ~n7061 & n15711 ) | ( ~n7061 & n15713 ) | ( n15711 & n15713 ) ;
  assign n15715 = ~x23 & n15713 ;
  assign n15716 = ~x23 & n15711 ;
  assign n15717 = ( ~n7061 & n15715 ) | ( ~n7061 & n15716 ) | ( n15715 & n15716 ) ;
  assign n15718 = x23 | n15716 ;
  assign n15719 = x23 | n15715 ;
  assign n15720 = ( ~n7061 & n15718 ) | ( ~n7061 & n15719 ) | ( n15718 & n15719 ) ;
  assign n15721 = ( ~n15714 & n15717 ) | ( ~n15714 & n15720 ) | ( n15717 & n15720 ) ;
  assign n15722 = n15704 & ~n15721 ;
  assign n15723 = n15704 | n15721 ;
  assign n15724 = ( ~n15704 & n15722 ) | ( ~n15704 & n15723 ) | ( n15722 & n15723 ) ;
  assign n15725 = n15697 & ~n15699 ;
  assign n15726 = n15700 | n15725 ;
  assign n15727 = n2925 & ~n6091 ;
  assign n15728 = n2928 & n7036 ;
  assign n15729 = ( n2928 & n7023 ) | ( n2928 & n15728 ) | ( n7023 & n15728 ) ;
  assign n15730 = n15727 | n15729 ;
  assign n15731 = n2932 & n6950 ;
  assign n15732 = n15730 | n15731 ;
  assign n15733 = n2936 | n15732 ;
  assign n15734 = ( ~n7107 & n15732 ) | ( ~n7107 & n15733 ) | ( n15732 & n15733 ) ;
  assign n15735 = ~x23 & n15733 ;
  assign n15736 = ~x23 & n15732 ;
  assign n15737 = ( ~n7107 & n15735 ) | ( ~n7107 & n15736 ) | ( n15735 & n15736 ) ;
  assign n15738 = x23 | n15735 ;
  assign n15739 = x23 | n15736 ;
  assign n15740 = ( ~n7107 & n15738 ) | ( ~n7107 & n15739 ) | ( n15738 & n15739 ) ;
  assign n15741 = ( ~n15734 & n15737 ) | ( ~n15734 & n15740 ) | ( n15737 & n15740 ) ;
  assign n15742 = n15726 & n15741 ;
  assign n15743 = n15336 | n15355 ;
  assign n15744 = ( n15336 & n15339 ) | ( n15336 & n15743 ) | ( n15339 & n15743 ) ;
  assign n15745 = n15742 & n15744 ;
  assign n15746 = ~n15726 & n15741 ;
  assign n15747 = n15744 | n15746 ;
  assign n15748 = n15726 | n15746 ;
  assign n15749 = ~n15746 & n15748 ;
  assign n15750 = ( n15745 & n15747 ) | ( n15745 & ~n15749 ) | ( n15747 & ~n15749 ) ;
  assign n15751 = n15724 & n15750 ;
  assign n15752 = n15724 | n15750 ;
  assign n15753 = ~n15751 & n15752 ;
  assign n15754 = n3544 & n7907 ;
  assign n15755 = ( n3544 & n7902 ) | ( n3544 & n15754 ) | ( n7902 & n15754 ) ;
  assign n15756 = n3541 & n8079 ;
  assign n15757 = ( n3541 & ~n8070 ) | ( n3541 & n15756 ) | ( ~n8070 & n15756 ) ;
  assign n15758 = n15755 | n15757 ;
  assign n15759 = n3547 & ~n8017 ;
  assign n15760 = n15758 | n15759 ;
  assign n15761 = n3537 | n15758 ;
  assign n15762 = n15759 | n15761 ;
  assign n15763 = ( n8104 & n15760 ) | ( n8104 & n15762 ) | ( n15760 & n15762 ) ;
  assign n15764 = x20 & n15762 ;
  assign n15765 = x20 & n15760 ;
  assign n15766 = ( n8104 & n15764 ) | ( n8104 & n15765 ) | ( n15764 & n15765 ) ;
  assign n15767 = x20 & ~n15765 ;
  assign n15768 = x20 & ~n15764 ;
  assign n15769 = ( ~n8104 & n15767 ) | ( ~n8104 & n15768 ) | ( n15767 & n15768 ) ;
  assign n15770 = ( n15763 & ~n15766 ) | ( n15763 & n15769 ) | ( ~n15766 & n15769 ) ;
  assign n15771 = n15753 & n15770 ;
  assign n15772 = n15753 & ~n15771 ;
  assign n15774 = ( n15744 & n15745 ) | ( n15744 & ~n15748 ) | ( n15745 & ~n15748 ) ;
  assign n15775 = n15742 | n15744 ;
  assign n15776 = n15748 & ~n15775 ;
  assign n15777 = n15774 | n15776 ;
  assign n15778 = n3544 & n6889 ;
  assign n15779 = ( n3544 & ~n6884 ) | ( n3544 & n15778 ) | ( ~n6884 & n15778 ) ;
  assign n15780 = n3541 & n7907 ;
  assign n15781 = ( n3541 & n7902 ) | ( n3541 & n15780 ) | ( n7902 & n15780 ) ;
  assign n15782 = n3547 & n8079 ;
  assign n15783 = ( n3547 & ~n8070 ) | ( n3547 & n15782 ) | ( ~n8070 & n15782 ) ;
  assign n15784 = n15781 | n15783 ;
  assign n15785 = n15779 | n15784 ;
  assign n15786 = n3537 | n15785 ;
  assign n15787 = n15785 & n15786 ;
  assign n15788 = ( ~n8156 & n15786 ) | ( ~n8156 & n15787 ) | ( n15786 & n15787 ) ;
  assign n15789 = ~x20 & n15787 ;
  assign n15790 = ~x20 & n15786 ;
  assign n15791 = ( ~n8156 & n15789 ) | ( ~n8156 & n15790 ) | ( n15789 & n15790 ) ;
  assign n15792 = x20 | n15789 ;
  assign n15793 = x20 | n15790 ;
  assign n15794 = ( ~n8156 & n15792 ) | ( ~n8156 & n15793 ) | ( n15792 & n15793 ) ;
  assign n15795 = ( ~n15788 & n15791 ) | ( ~n15788 & n15794 ) | ( n15791 & n15794 ) ;
  assign n15796 = ~n15777 & n15795 ;
  assign n15797 = n15777 & ~n15795 ;
  assign n15798 = n15796 | n15797 ;
  assign n15799 = n15361 | n15380 ;
  assign n15800 = ( n15361 & n15363 ) | ( n15361 & n15799 ) | ( n15363 & n15799 ) ;
  assign n15801 = n15796 | n15800 ;
  assign n15802 = ( n15796 & ~n15798 ) | ( n15796 & n15801 ) | ( ~n15798 & n15801 ) ;
  assign n15773 = ~n15753 & n15770 ;
  assign n15803 = n15773 & n15802 ;
  assign n15804 = ( n15772 & n15802 ) | ( n15772 & n15803 ) | ( n15802 & n15803 ) ;
  assign n15805 = n15773 | n15802 ;
  assign n15806 = n15772 | n15805 ;
  assign n15807 = ~n15804 & n15806 ;
  assign n15808 = n4468 & ~n8982 ;
  assign n15809 = ( n4468 & n9051 ) | ( n4468 & n15808 ) | ( n9051 & n15808 ) ;
  assign n15810 = n4466 & ~n9022 ;
  assign n15811 = ( n4466 & n15809 ) | ( n4466 & ~n15810 ) | ( n15809 & ~n15810 ) ;
  assign n15812 = n4466 | n15809 ;
  assign n15813 = ( ~n9019 & n15811 ) | ( ~n9019 & n15812 ) | ( n15811 & n15812 ) ;
  assign n15814 = n4475 | n15813 ;
  assign n15815 = ( n9078 & n15813 ) | ( n9078 & n15814 ) | ( n15813 & n15814 ) ;
  assign n15816 = x17 & n15814 ;
  assign n15817 = x17 & n15813 ;
  assign n15818 = ( n9078 & n15816 ) | ( n9078 & n15817 ) | ( n15816 & n15817 ) ;
  assign n15819 = x17 & ~n15816 ;
  assign n15820 = x17 & ~n15817 ;
  assign n15821 = ( ~n9078 & n15819 ) | ( ~n9078 & n15820 ) | ( n15819 & n15820 ) ;
  assign n15822 = ( n15815 & ~n15818 ) | ( n15815 & n15821 ) | ( ~n15818 & n15821 ) ;
  assign n15823 = n15807 & ~n15822 ;
  assign n15824 = n15807 | n15822 ;
  assign n15825 = ( ~n15807 & n15823 ) | ( ~n15807 & n15824 ) | ( n15823 & n15824 ) ;
  assign n15826 = n4471 & ~n8982 ;
  assign n15827 = ( n4471 & n9051 ) | ( n4471 & n15826 ) | ( n9051 & n15826 ) ;
  assign n15828 = n4468 & n9022 ;
  assign n15829 = n15827 | n15828 ;
  assign n15830 = n4468 | n15827 ;
  assign n15831 = ( ~n9019 & n15829 ) | ( ~n9019 & n15830 ) | ( n15829 & n15830 ) ;
  assign n15832 = n4466 | n15831 ;
  assign n15833 = ( ~n8017 & n15831 ) | ( ~n8017 & n15832 ) | ( n15831 & n15832 ) ;
  assign n15834 = n4475 | n15833 ;
  assign n15835 = ( ~n10242 & n15833 ) | ( ~n10242 & n15834 ) | ( n15833 & n15834 ) ;
  assign n15836 = ~x17 & n15834 ;
  assign n15837 = ~x17 & n15833 ;
  assign n15838 = ( ~n10242 & n15836 ) | ( ~n10242 & n15837 ) | ( n15836 & n15837 ) ;
  assign n15839 = x17 | n15836 ;
  assign n15840 = x17 | n15837 ;
  assign n15841 = ( ~n10242 & n15839 ) | ( ~n10242 & n15840 ) | ( n15839 & n15840 ) ;
  assign n15842 = ( ~n15835 & n15838 ) | ( ~n15835 & n15841 ) | ( n15838 & n15841 ) ;
  assign n15843 = n15386 | n15405 ;
  assign n15844 = ( n15386 & n15388 ) | ( n15386 & n15843 ) | ( n15388 & n15843 ) ;
  assign n15845 = n15842 & n15844 ;
  assign n15846 = n15842 | n15844 ;
  assign n15847 = ~n15845 & n15846 ;
  assign n15848 = ~n15798 & n15800 ;
  assign n15849 = n15798 & ~n15800 ;
  assign n15850 = n15848 | n15849 ;
  assign n15851 = ~n15845 & n15850 ;
  assign n15852 = ( n15845 & n15847 ) | ( n15845 & ~n15851 ) | ( n15847 & ~n15851 ) ;
  assign n15853 = n15825 & n15852 ;
  assign n15854 = n15825 | n15852 ;
  assign n15855 = ~n15853 & n15854 ;
  assign n15856 = n15847 & ~n15850 ;
  assign n15857 = ~n15847 & n15850 ;
  assign n15858 = n15856 | n15857 ;
  assign n15859 = n15171 | n15408 ;
  assign n15860 = ( n15171 & n15173 ) | ( n15171 & n15859 ) | ( n15173 & n15859 ) ;
  assign n15861 = ~n15858 & n15860 ;
  assign n15862 = n15858 & ~n15860 ;
  assign n15863 = n15861 | n15862 ;
  assign n15864 = n15414 | n15417 ;
  assign n15865 = ~n15863 & n15864 ;
  assign n15866 = n15861 | n15865 ;
  assign n15867 = n15414 | n15416 ;
  assign n15868 = ~n15863 & n15867 ;
  assign n15869 = n15861 | n15868 ;
  assign n15870 = ( n14578 & n15866 ) | ( n14578 & n15869 ) | ( n15866 & n15869 ) ;
  assign n15871 = n15414 | n15420 ;
  assign n15872 = ~n15863 & n15871 ;
  assign n15873 = n15861 | n15872 ;
  assign n15874 = n15414 | n15422 ;
  assign n15875 = ~n15863 & n15874 ;
  assign n15876 = n15861 | n15875 ;
  assign n15877 = ( n14318 & n15873 ) | ( n14318 & n15876 ) | ( n15873 & n15876 ) ;
  assign n15878 = ( n12930 & n15870 ) | ( n12930 & n15877 ) | ( n15870 & n15877 ) ;
  assign n15879 = n15855 & n15878 ;
  assign n15880 = ( n12928 & n15870 ) | ( n12928 & n15877 ) | ( n15870 & n15877 ) ;
  assign n15881 = n15855 & n15880 ;
  assign n15882 = ( n11360 & n15879 ) | ( n11360 & n15881 ) | ( n15879 & n15881 ) ;
  assign n15883 = n15855 | n15878 ;
  assign n15884 = n15855 | n15880 ;
  assign n15885 = ( n11360 & n15883 ) | ( n11360 & n15884 ) | ( n15883 & n15884 ) ;
  assign n15886 = ~n15882 & n15885 ;
  assign n15887 = n4466 & ~n8982 ;
  assign n15888 = ( n4466 & n9051 ) | ( n4466 & n15887 ) | ( n9051 & n15887 ) ;
  assign n15889 = n4475 | n15888 ;
  assign n15890 = n9442 & ~n15888 ;
  assign n15891 = n9074 & ~n15888 ;
  assign n15892 = ( ~n9440 & n15890 ) | ( ~n9440 & n15891 ) | ( n15890 & n15891 ) ;
  assign n15893 = n15889 & ~n15892 ;
  assign n15894 = n15888 & n15889 ;
  assign n15895 = ( ~n9442 & n15889 ) | ( ~n9442 & n15894 ) | ( n15889 & n15894 ) ;
  assign n15896 = ( ~n9072 & n15893 ) | ( ~n9072 & n15895 ) | ( n15893 & n15895 ) ;
  assign n15897 = ~x17 & n15893 ;
  assign n15898 = ~x17 & n15895 ;
  assign n15899 = ( ~n9072 & n15897 ) | ( ~n9072 & n15898 ) | ( n15897 & n15898 ) ;
  assign n15900 = x17 | n15897 ;
  assign n15901 = x17 | n15898 ;
  assign n15902 = ( ~n9072 & n15900 ) | ( ~n9072 & n15901 ) | ( n15900 & n15901 ) ;
  assign n15903 = ( ~n15896 & n15899 ) | ( ~n15896 & n15902 ) | ( n15899 & n15902 ) ;
  assign n15904 = n15751 | n15770 ;
  assign n15905 = ( n15751 & n15753 ) | ( n15751 & n15904 ) | ( n15753 & n15904 ) ;
  assign n15906 = n15903 & n15905 ;
  assign n15907 = n15903 | n15905 ;
  assign n15908 = ~n15906 & n15907 ;
  assign n15909 = n15617 & ~n15620 ;
  assign n15910 = n15617 & ~n15621 ;
  assign n15911 = ( ~n4455 & n15909 ) | ( ~n4455 & n15910 ) | ( n15909 & n15910 ) ;
  assign n15912 = n296 | n839 ;
  assign n15913 = n291 | n631 ;
  assign n15914 = n15912 | n15913 ;
  assign n15915 = n2875 | n3987 ;
  assign n15916 = n1673 | n4410 ;
  assign n15917 = n15915 | n15916 ;
  assign n15918 = n15914 | n15917 ;
  assign n15919 = n497 | n2135 ;
  assign n15920 = n6065 | n15919 ;
  assign n15921 = n15918 | n15920 ;
  assign n15922 = n1701 | n15921 ;
  assign n15923 = n8067 | n15922 ;
  assign n15924 = n711 | n1016 ;
  assign n15925 = n268 | n15924 ;
  assign n15926 = n6868 & ~n15925 ;
  assign n15927 = ~n15923 & n15926 ;
  assign n15928 = n171 | n214 ;
  assign n15929 = n15243 | n15928 ;
  assign n15930 = n356 | n895 ;
  assign n15931 = n15929 | n15930 ;
  assign n15932 = n15927 & ~n15931 ;
  assign n15933 = n15616 | n15932 ;
  assign n15934 = n15616 & n15932 ;
  assign n15935 = n15617 | n15934 ;
  assign n15936 = n15933 & ~n15935 ;
  assign n15937 = n15933 & ~n15934 ;
  assign n15938 = ( n15620 & n15936 ) | ( n15620 & n15937 ) | ( n15936 & n15937 ) ;
  assign n15939 = ( n15621 & n15936 ) | ( n15621 & n15937 ) | ( n15936 & n15937 ) ;
  assign n15940 = ( n4455 & n15938 ) | ( n4455 & n15939 ) | ( n15938 & n15939 ) ;
  assign n15941 = n15911 | n15940 ;
  assign n15942 = n1060 & n4396 ;
  assign n15943 = n1065 & n4245 ;
  assign n15944 = ( n1065 & n4303 ) | ( n1065 & n15943 ) | ( n4303 & n15943 ) ;
  assign n15945 = n15942 | n15944 ;
  assign n15946 = n1062 | n15945 ;
  assign n15947 = n1057 & n5192 ;
  assign n15948 = ( n1057 & n5179 ) | ( n1057 & n15947 ) | ( n5179 & n15947 ) ;
  assign n15949 = n15946 | n15948 ;
  assign n15950 = n15945 | n15948 ;
  assign n15951 = ( n5306 & n15949 ) | ( n5306 & n15950 ) | ( n15949 & n15950 ) ;
  assign n15952 = n15934 | n15939 ;
  assign n15953 = n15933 & ~n15952 ;
  assign n15954 = n15934 | n15938 ;
  assign n15955 = n15933 & ~n15954 ;
  assign n15956 = ( ~n4455 & n15953 ) | ( ~n4455 & n15955 ) | ( n15953 & n15955 ) ;
  assign n15957 = n15951 & n15956 ;
  assign n15958 = ( ~n15941 & n15951 ) | ( ~n15941 & n15957 ) | ( n15951 & n15957 ) ;
  assign n15959 = n15951 | n15956 ;
  assign n15960 = n15941 & ~n15959 ;
  assign n15961 = n15958 | n15960 ;
  assign n15962 = n1826 & n5117 ;
  assign n15963 = ( n1826 & ~n5037 ) | ( n1826 & n15962 ) | ( ~n5037 & n15962 ) ;
  assign n15964 = n1823 & n5108 ;
  assign n15965 = n1829 & n5997 ;
  assign n15966 = ( n1829 & n5979 ) | ( n1829 & n15965 ) | ( n5979 & n15965 ) ;
  assign n15967 = n15964 | n15966 ;
  assign n15968 = n15963 | n15967 ;
  assign n15969 = n1821 | n15968 ;
  assign n15970 = ( n6181 & n15968 ) | ( n6181 & n15969 ) | ( n15968 & n15969 ) ;
  assign n15971 = x29 & n15969 ;
  assign n15972 = x29 & n15968 ;
  assign n15973 = ( n6181 & n15971 ) | ( n6181 & n15972 ) | ( n15971 & n15972 ) ;
  assign n15974 = x29 & ~n15971 ;
  assign n15975 = x29 & ~n15972 ;
  assign n15976 = ( ~n6181 & n15974 ) | ( ~n6181 & n15975 ) | ( n15974 & n15975 ) ;
  assign n15977 = ( n15970 & ~n15973 ) | ( n15970 & n15976 ) | ( ~n15973 & n15976 ) ;
  assign n15978 = ~n15961 & n15977 ;
  assign n15979 = n15961 | n15978 ;
  assign n15981 = n15629 | n15648 ;
  assign n15982 = ( n15629 & n15631 ) | ( n15629 & n15981 ) | ( n15631 & n15981 ) ;
  assign n15980 = n15961 & n15977 ;
  assign n15983 = n15980 & n15982 ;
  assign n15984 = ( ~n15979 & n15982 ) | ( ~n15979 & n15983 ) | ( n15982 & n15983 ) ;
  assign n15985 = n15980 | n15982 ;
  assign n15986 = n15979 & ~n15985 ;
  assign n15987 = n15984 | n15986 ;
  assign n15988 = n2312 & n5857 ;
  assign n15989 = ( n2312 & ~n5899 ) | ( n2312 & n15988 ) | ( ~n5899 & n15988 ) ;
  assign n15990 = n2308 & ~n6091 ;
  assign n15991 = n2315 & n7036 ;
  assign n15992 = ( n2315 & n7023 ) | ( n2315 & n15991 ) | ( n7023 & n15991 ) ;
  assign n15993 = n15990 | n15992 ;
  assign n15994 = n15989 | n15993 ;
  assign n15995 = n2306 | n15994 ;
  assign n15996 = ( n7136 & n15994 ) | ( n7136 & n15995 ) | ( n15994 & n15995 ) ;
  assign n15997 = x26 & n15995 ;
  assign n15998 = x26 & n15994 ;
  assign n15999 = ( n7136 & n15997 ) | ( n7136 & n15998 ) | ( n15997 & n15998 ) ;
  assign n16000 = x26 & ~n15997 ;
  assign n16001 = x26 & ~n15998 ;
  assign n16002 = ( ~n7136 & n16000 ) | ( ~n7136 & n16001 ) | ( n16000 & n16001 ) ;
  assign n16003 = ( n15996 & ~n15999 ) | ( n15996 & n16002 ) | ( ~n15999 & n16002 ) ;
  assign n16004 = n15987 | n16003 ;
  assign n16005 = n15987 & ~n16003 ;
  assign n16006 = ( ~n15987 & n16004 ) | ( ~n15987 & n16005 ) | ( n16004 & n16005 ) ;
  assign n16007 = n15653 | n15672 ;
  assign n16008 = ( n15653 & n15656 ) | ( n15653 & n16007 ) | ( n15656 & n16007 ) ;
  assign n16009 = ~n16006 & n16008 ;
  assign n16010 = n16006 & ~n16008 ;
  assign n16011 = n16009 | n16010 ;
  assign n16012 = n2925 & n6950 ;
  assign n16013 = n2928 & n6889 ;
  assign n16014 = ( n2928 & ~n6884 ) | ( n2928 & n16013 ) | ( ~n6884 & n16013 ) ;
  assign n16015 = n16012 | n16014 ;
  assign n16016 = n2932 & n7907 ;
  assign n16017 = ( n2932 & n7902 ) | ( n2932 & n16016 ) | ( n7902 & n16016 ) ;
  assign n16018 = n16015 | n16017 ;
  assign n16019 = n2936 | n16017 ;
  assign n16020 = n16015 | n16019 ;
  assign n16021 = ( ~n8193 & n16018 ) | ( ~n8193 & n16020 ) | ( n16018 & n16020 ) ;
  assign n16022 = ~x23 & n16020 ;
  assign n16023 = ~x23 & n16018 ;
  assign n16024 = ( ~n8193 & n16022 ) | ( ~n8193 & n16023 ) | ( n16022 & n16023 ) ;
  assign n16025 = x23 | n16023 ;
  assign n16026 = x23 | n16022 ;
  assign n16027 = ( ~n8193 & n16025 ) | ( ~n8193 & n16026 ) | ( n16025 & n16026 ) ;
  assign n16028 = ( ~n16021 & n16024 ) | ( ~n16021 & n16027 ) | ( n16024 & n16027 ) ;
  assign n16029 = n16011 | n16028 ;
  assign n16030 = n16011 & ~n16028 ;
  assign n16031 = ( ~n16011 & n16029 ) | ( ~n16011 & n16030 ) | ( n16029 & n16030 ) ;
  assign n16032 = n15702 | n15721 ;
  assign n16033 = ( n15702 & n15704 ) | ( n15702 & n16032 ) | ( n15704 & n16032 ) ;
  assign n16034 = ~n16031 & n16033 ;
  assign n16035 = n16031 & ~n16033 ;
  assign n16036 = n16034 | n16035 ;
  assign n16037 = n3544 & n8079 ;
  assign n16038 = ( n3544 & ~n8070 ) | ( n3544 & n16037 ) | ( ~n8070 & n16037 ) ;
  assign n16039 = n3541 | n16038 ;
  assign n16040 = ( ~n8017 & n16038 ) | ( ~n8017 & n16039 ) | ( n16038 & n16039 ) ;
  assign n16041 = n3547 & n9022 ;
  assign n16042 = ( n3547 & ~n9019 ) | ( n3547 & n16041 ) | ( ~n9019 & n16041 ) ;
  assign n16043 = n16040 | n16042 ;
  assign n16044 = n3537 | n16042 ;
  assign n16045 = n16040 | n16044 ;
  assign n16046 = ( ~n9416 & n16043 ) | ( ~n9416 & n16045 ) | ( n16043 & n16045 ) ;
  assign n16047 = ~x20 & n16045 ;
  assign n16048 = ~x20 & n16043 ;
  assign n16049 = ( ~n9416 & n16047 ) | ( ~n9416 & n16048 ) | ( n16047 & n16048 ) ;
  assign n16050 = x20 | n16048 ;
  assign n16051 = x20 | n16047 ;
  assign n16052 = ( ~n9416 & n16050 ) | ( ~n9416 & n16051 ) | ( n16050 & n16051 ) ;
  assign n16053 = ( ~n16046 & n16049 ) | ( ~n16046 & n16052 ) | ( n16049 & n16052 ) ;
  assign n16054 = n16036 | n16053 ;
  assign n16055 = n16036 & ~n16053 ;
  assign n16056 = ( ~n16036 & n16054 ) | ( ~n16036 & n16055 ) | ( n16054 & n16055 ) ;
  assign n16057 = n15908 & ~n16056 ;
  assign n16058 = n15908 | n16056 ;
  assign n16059 = ( ~n15908 & n16057 ) | ( ~n15908 & n16058 ) | ( n16057 & n16058 ) ;
  assign n16060 = n15804 | n15822 ;
  assign n16061 = ( n15804 & n15807 ) | ( n15804 & n16060 ) | ( n15807 & n16060 ) ;
  assign n16062 = ~n16059 & n16061 ;
  assign n16063 = n16059 & ~n16061 ;
  assign n16064 = n16062 | n16063 ;
  assign n16065 = n15853 & ~n16064 ;
  assign n16066 = ( n15882 & ~n16064 ) | ( n15882 & n16065 ) | ( ~n16064 & n16065 ) ;
  assign n16067 = ~n15853 & n16064 ;
  assign n16068 = ~n15882 & n16067 ;
  assign n16069 = n16066 | n16068 ;
  assign n16070 = n15886 & ~n16069 ;
  assign n16071 = ~n15886 & n16069 ;
  assign n16072 = n16070 | n16071 ;
  assign n16073 = ( n14578 & n15865 ) | ( n14578 & n15868 ) | ( n15865 & n15868 ) ;
  assign n16074 = ( n14318 & n15872 ) | ( n14318 & n15875 ) | ( n15872 & n15875 ) ;
  assign n16075 = ( n12928 & n16073 ) | ( n12928 & n16074 ) | ( n16073 & n16074 ) ;
  assign n16076 = ( n12930 & n16073 ) | ( n12930 & n16074 ) | ( n16073 & n16074 ) ;
  assign n16077 = ( n11360 & n16075 ) | ( n11360 & n16076 ) | ( n16075 & n16076 ) ;
  assign n16078 = ( n14578 & n15864 ) | ( n14578 & n15867 ) | ( n15864 & n15867 ) ;
  assign n16079 = ( n14318 & n15871 ) | ( n14318 & n15874 ) | ( n15871 & n15874 ) ;
  assign n16080 = ( n12930 & n16078 ) | ( n12930 & n16079 ) | ( n16078 & n16079 ) ;
  assign n16081 = n15863 & ~n16080 ;
  assign n16082 = ( n12928 & n16078 ) | ( n12928 & n16079 ) | ( n16078 & n16079 ) ;
  assign n16083 = n15863 & ~n16082 ;
  assign n16084 = ( ~n11360 & n16081 ) | ( ~n11360 & n16083 ) | ( n16081 & n16083 ) ;
  assign n16085 = n16077 | n16084 ;
  assign n16086 = n15886 & ~n16085 ;
  assign n16087 = n15434 & ~n16085 ;
  assign n16088 = ~n15434 & n16085 ;
  assign n16089 = n16087 | n16088 ;
  assign n16090 = ~n16087 & n16089 ;
  assign n16091 = ~n15886 & n16085 ;
  assign n16092 = n16086 | n16091 ;
  assign n16093 = ~n16086 & n16092 ;
  assign n16094 = ( ~n16086 & n16090 ) | ( ~n16086 & n16093 ) | ( n16090 & n16093 ) ;
  assign n16095 = n16072 | n16094 ;
  assign n16096 = n16086 | n16087 ;
  assign n16097 = ( n16086 & ~n16092 ) | ( n16086 & n16096 ) | ( ~n16092 & n16096 ) ;
  assign n16098 = ~n16072 & n16097 ;
  assign n16099 = ( n15435 & ~n16095 ) | ( n15435 & n16098 ) | ( ~n16095 & n16098 ) ;
  assign n16100 = n16095 & ~n16098 ;
  assign n16101 = ( n15446 & n16099 ) | ( n15446 & ~n16100 ) | ( n16099 & ~n16100 ) ;
  assign n16102 = n16094 & ~n16097 ;
  assign n16103 = n16072 & n16102 ;
  assign n16104 = ( n15435 & ~n16094 ) | ( n15435 & n16097 ) | ( ~n16094 & n16097 ) ;
  assign n16105 = n16072 & ~n16104 ;
  assign n16106 = ( ~n15446 & n16103 ) | ( ~n15446 & n16105 ) | ( n16103 & n16105 ) ;
  assign n16107 = n16101 | n16106 ;
  assign n16108 = n4471 & ~n16069 ;
  assign n16109 = n4466 & ~n16085 ;
  assign n16110 = n4468 & n15886 ;
  assign n16111 = n16109 | n16110 ;
  assign n16112 = n16108 | n16111 ;
  assign n16113 = n4475 | n16112 ;
  assign n16114 = ( ~n16107 & n16112 ) | ( ~n16107 & n16113 ) | ( n16112 & n16113 ) ;
  assign n16115 = ~x17 & n16113 ;
  assign n16116 = ~x17 & n16112 ;
  assign n16117 = ( ~n16107 & n16115 ) | ( ~n16107 & n16116 ) | ( n16115 & n16116 ) ;
  assign n16118 = x17 | n16115 ;
  assign n16119 = x17 | n16116 ;
  assign n16120 = ( ~n16107 & n16118 ) | ( ~n16107 & n16119 ) | ( n16118 & n16119 ) ;
  assign n16121 = ( ~n16114 & n16117 ) | ( ~n16114 & n16120 ) | ( n16117 & n16120 ) ;
  assign n16122 = ~n15476 & n16121 ;
  assign n16123 = ( n15475 & n16121 ) | ( n15475 & n16122 ) | ( n16121 & n16122 ) ;
  assign n16124 = n15477 | n16123 ;
  assign n16125 = n15476 & n16121 ;
  assign n16126 = ~n15475 & n16125 ;
  assign n16127 = n16124 & ~n16126 ;
  assign n16128 = n14994 & ~n14998 ;
  assign n16129 = n14997 | n14998 ;
  assign n16130 = ~n16128 & n16129 ;
  assign n16131 = n16090 | n16092 ;
  assign n16132 = n16087 & ~n16092 ;
  assign n16133 = ( n15435 & ~n16131 ) | ( n15435 & n16132 ) | ( ~n16131 & n16132 ) ;
  assign n16134 = n16131 & ~n16132 ;
  assign n16135 = ( n15446 & n16133 ) | ( n15446 & ~n16134 ) | ( n16133 & ~n16134 ) ;
  assign n16136 = ( n15434 & n15435 ) | ( n15434 & ~n16085 ) | ( n15435 & ~n16085 ) ;
  assign n16137 = n16092 & ~n16136 ;
  assign n16138 = n16088 & n16092 ;
  assign n16139 = ( ~n15446 & n16137 ) | ( ~n15446 & n16138 ) | ( n16137 & n16138 ) ;
  assign n16140 = n16135 | n16139 ;
  assign n16141 = n4471 & n15886 ;
  assign n16142 = n4466 & n15434 ;
  assign n16143 = n4468 & ~n16085 ;
  assign n16144 = n16142 | n16143 ;
  assign n16145 = n16141 | n16144 ;
  assign n16146 = n4475 | n16141 ;
  assign n16147 = n16144 | n16146 ;
  assign n16148 = ( ~n16140 & n16145 ) | ( ~n16140 & n16147 ) | ( n16145 & n16147 ) ;
  assign n16149 = ~x17 & n16147 ;
  assign n16150 = ~x17 & n16145 ;
  assign n16151 = ( ~n16140 & n16149 ) | ( ~n16140 & n16150 ) | ( n16149 & n16150 ) ;
  assign n16152 = x17 | n16150 ;
  assign n16153 = x17 | n16149 ;
  assign n16154 = ( ~n16140 & n16152 ) | ( ~n16140 & n16153 ) | ( n16152 & n16153 ) ;
  assign n16155 = ( ~n16148 & n16151 ) | ( ~n16148 & n16154 ) | ( n16151 & n16154 ) ;
  assign n16156 = ~n16130 & n16155 ;
  assign n16157 = n16130 | n16156 ;
  assign n16158 = n16130 & n16155 ;
  assign n16159 = n16157 & ~n16158 ;
  assign n16160 = n14992 & ~n14993 ;
  assign n16161 = n14676 & ~n14993 ;
  assign n16162 = n16160 | n16161 ;
  assign n16163 = n15435 & ~n16089 ;
  assign n16164 = ( n15446 & ~n16089 ) | ( n15446 & n16163 ) | ( ~n16089 & n16163 ) ;
  assign n16165 = ~n15435 & n16089 ;
  assign n16166 = ~n15446 & n16165 ;
  assign n16167 = n16164 | n16166 ;
  assign n16168 = n4471 & ~n16085 ;
  assign n16169 = n4466 & n14591 ;
  assign n16170 = n4468 & n15434 ;
  assign n16171 = n16169 | n16170 ;
  assign n16172 = n16168 | n16171 ;
  assign n16173 = n4475 | n16168 ;
  assign n16174 = n16171 | n16173 ;
  assign n16175 = ( ~n16167 & n16172 ) | ( ~n16167 & n16174 ) | ( n16172 & n16174 ) ;
  assign n16176 = ~x17 & n16174 ;
  assign n16177 = ~x17 & n16172 ;
  assign n16178 = ( ~n16167 & n16176 ) | ( ~n16167 & n16177 ) | ( n16176 & n16177 ) ;
  assign n16179 = x17 | n16177 ;
  assign n16180 = x17 | n16176 ;
  assign n16181 = ( ~n16167 & n16179 ) | ( ~n16167 & n16180 ) | ( n16179 & n16180 ) ;
  assign n16182 = ( ~n16175 & n16178 ) | ( ~n16175 & n16181 ) | ( n16178 & n16181 ) ;
  assign n16183 = n16162 & n16182 ;
  assign n16184 = n16162 & ~n16183 ;
  assign n16185 = ~n16162 & n16182 ;
  assign n16186 = n16184 | n16185 ;
  assign n16187 = n14709 & n14990 ;
  assign n16188 = n14709 | n14990 ;
  assign n16189 = ~n16187 & n16188 ;
  assign n16190 = n4471 & n15434 ;
  assign n16191 = n4466 & n14329 ;
  assign n16192 = n4468 & n14591 ;
  assign n16193 = n16191 | n16192 ;
  assign n16194 = n16190 | n16193 ;
  assign n16195 = n4475 | n16190 ;
  assign n16196 = n16193 | n16195 ;
  assign n16197 = ( n15453 & n16194 ) | ( n15453 & n16196 ) | ( n16194 & n16196 ) ;
  assign n16198 = x17 & n16196 ;
  assign n16199 = x17 & n16194 ;
  assign n16200 = ( n15453 & n16198 ) | ( n15453 & n16199 ) | ( n16198 & n16199 ) ;
  assign n16201 = x17 & ~n16199 ;
  assign n16202 = x17 & ~n16198 ;
  assign n16203 = ( ~n15453 & n16201 ) | ( ~n15453 & n16202 ) | ( n16201 & n16202 ) ;
  assign n16204 = ( n16197 & ~n16200 ) | ( n16197 & n16203 ) | ( ~n16200 & n16203 ) ;
  assign n16205 = ~n16189 & n16204 ;
  assign n16206 = n16189 & ~n16204 ;
  assign n16207 = n16205 | n16206 ;
  assign n16208 = ~n14732 & n14988 ;
  assign n16209 = n14732 | n16208 ;
  assign n16212 = n4471 & n14591 ;
  assign n16213 = n4466 & n14607 ;
  assign n16214 = n4468 & n14329 ;
  assign n16215 = n16213 | n16214 ;
  assign n16216 = n16212 | n16215 ;
  assign n16217 = n4475 | n16212 ;
  assign n16218 = n16215 | n16217 ;
  assign n16219 = ( n14629 & n16216 ) | ( n14629 & n16218 ) | ( n16216 & n16218 ) ;
  assign n16220 = x17 & n16218 ;
  assign n16221 = x17 & n16216 ;
  assign n16222 = ( n14629 & n16220 ) | ( n14629 & n16221 ) | ( n16220 & n16221 ) ;
  assign n16223 = x17 & ~n16221 ;
  assign n16224 = x17 & ~n16220 ;
  assign n16225 = ( ~n14629 & n16223 ) | ( ~n14629 & n16224 ) | ( n16223 & n16224 ) ;
  assign n16226 = ( n16219 & ~n16222 ) | ( n16219 & n16225 ) | ( ~n16222 & n16225 ) ;
  assign n16210 = n14732 & n14988 ;
  assign n16227 = n16210 & n16226 ;
  assign n16228 = ( ~n16209 & n16226 ) | ( ~n16209 & n16227 ) | ( n16226 & n16227 ) ;
  assign n16211 = n16209 & ~n16210 ;
  assign n16229 = n16211 | n16228 ;
  assign n16230 = ~n16210 & n16226 ;
  assign n16231 = n16209 & n16230 ;
  assign n16232 = n16229 & ~n16231 ;
  assign n16233 = n14753 | n14986 ;
  assign n16234 = ~n14987 & n16233 ;
  assign n16236 = n4466 & n13522 ;
  assign n16237 = n4468 & n14607 ;
  assign n16238 = n16236 | n16237 ;
  assign n16235 = n4471 & n14329 ;
  assign n16240 = n4475 | n16235 ;
  assign n16241 = n16238 | n16240 ;
  assign n16239 = n16235 | n16238 ;
  assign n16242 = n16239 & n16241 ;
  assign n16243 = ( n14656 & n16241 ) | ( n14656 & n16242 ) | ( n16241 & n16242 ) ;
  assign n16244 = x17 & n16242 ;
  assign n16245 = x17 & n16241 ;
  assign n16246 = ( n14656 & n16244 ) | ( n14656 & n16245 ) | ( n16244 & n16245 ) ;
  assign n16247 = x17 & ~n16244 ;
  assign n16248 = x17 & ~n16245 ;
  assign n16249 = ( ~n14656 & n16247 ) | ( ~n14656 & n16248 ) | ( n16247 & n16248 ) ;
  assign n16250 = ( n16243 & ~n16246 ) | ( n16243 & n16249 ) | ( ~n16246 & n16249 ) ;
  assign n16251 = n16234 & n16250 ;
  assign n16252 = n14982 & n14984 ;
  assign n16253 = n14982 | n14984 ;
  assign n16254 = ~n16252 & n16253 ;
  assign n16255 = n4466 & n13235 ;
  assign n16256 = n4468 & n13522 ;
  assign n16257 = n16255 | n16256 ;
  assign n16258 = n4471 & n14607 ;
  assign n16259 = n4475 | n16258 ;
  assign n16260 = n16257 | n16259 ;
  assign n16261 = n16257 | n16258 ;
  assign n16262 = n14696 | n16261 ;
  assign n16263 = n14698 | n16261 ;
  assign n16264 = ( ~n13248 & n16262 ) | ( ~n13248 & n16263 ) | ( n16262 & n16263 ) ;
  assign n16265 = n16260 & n16264 ;
  assign n16266 = ( n14687 & n16260 ) | ( n14687 & n16265 ) | ( n16260 & n16265 ) ;
  assign n16267 = ~x17 & n16266 ;
  assign n16268 = x17 | n16266 ;
  assign n16269 = ( ~n16266 & n16267 ) | ( ~n16266 & n16268 ) | ( n16267 & n16268 ) ;
  assign n16270 = n16254 & n16269 ;
  assign n16271 = n16254 & ~n16270 ;
  assign n16272 = ~n16254 & n16269 ;
  assign n16273 = n16271 | n16272 ;
  assign n16274 = n14978 & n14980 ;
  assign n16275 = n14978 | n14980 ;
  assign n16276 = ~n16274 & n16275 ;
  assign n16277 = n4471 & n13522 ;
  assign n16278 = n4466 & n12936 ;
  assign n16279 = n4468 & n13235 ;
  assign n16280 = n16278 | n16279 ;
  assign n16281 = n16277 | n16280 ;
  assign n16282 = n4475 & n13537 ;
  assign n16283 = n4475 & n13539 ;
  assign n16284 = ( ~n13248 & n16282 ) | ( ~n13248 & n16283 ) | ( n16282 & n16283 ) ;
  assign n16285 = n16281 | n16284 ;
  assign n16286 = n4475 | n16281 ;
  assign n16287 = ( n13530 & n16285 ) | ( n13530 & n16286 ) | ( n16285 & n16286 ) ;
  assign n16288 = x17 | n16287 ;
  assign n16289 = ~x17 & n16287 ;
  assign n16290 = ( ~n16287 & n16288 ) | ( ~n16287 & n16289 ) | ( n16288 & n16289 ) ;
  assign n16291 = n16276 & n16290 ;
  assign n16292 = n14976 & ~n14977 ;
  assign n16293 = n14812 & ~n14977 ;
  assign n16294 = n16292 | n16293 ;
  assign n16295 = n4471 & n13235 ;
  assign n16296 = n4466 & ~n12616 ;
  assign n16297 = n4468 & n12936 ;
  assign n16298 = n16296 | n16297 ;
  assign n16299 = n16295 | n16298 ;
  assign n16300 = n4475 | n16295 ;
  assign n16301 = n16298 | n16300 ;
  assign n16302 = ( n13561 & n16299 ) | ( n13561 & n16301 ) | ( n16299 & n16301 ) ;
  assign n16303 = x17 & n16301 ;
  assign n16304 = x17 & n16299 ;
  assign n16305 = ( n13561 & n16303 ) | ( n13561 & n16304 ) | ( n16303 & n16304 ) ;
  assign n16306 = x17 & ~n16304 ;
  assign n16307 = x17 & ~n16303 ;
  assign n16308 = ( ~n13561 & n16306 ) | ( ~n13561 & n16307 ) | ( n16306 & n16307 ) ;
  assign n16309 = ( n16302 & ~n16305 ) | ( n16302 & n16308 ) | ( ~n16305 & n16308 ) ;
  assign n16310 = n16294 & n16309 ;
  assign n16311 = n16294 & ~n16310 ;
  assign n16312 = ~n14832 & n14974 ;
  assign n16313 = n14832 & ~n14974 ;
  assign n16314 = n16312 | n16313 ;
  assign n16315 = n4471 & n12936 ;
  assign n16316 = n4466 & n12010 ;
  assign n16317 = n4468 & ~n12616 ;
  assign n16318 = n16316 | n16317 ;
  assign n16319 = n16315 | n16318 ;
  assign n16320 = n4475 | n16315 ;
  assign n16321 = n16318 | n16320 ;
  assign n16322 = ( ~n13591 & n16319 ) | ( ~n13591 & n16321 ) | ( n16319 & n16321 ) ;
  assign n16323 = ~x17 & n16321 ;
  assign n16324 = ~x17 & n16319 ;
  assign n16325 = ( ~n13591 & n16323 ) | ( ~n13591 & n16324 ) | ( n16323 & n16324 ) ;
  assign n16326 = x17 | n16324 ;
  assign n16327 = x17 | n16323 ;
  assign n16328 = ( ~n13591 & n16326 ) | ( ~n13591 & n16327 ) | ( n16326 & n16327 ) ;
  assign n16329 = ( ~n16322 & n16325 ) | ( ~n16322 & n16328 ) | ( n16325 & n16328 ) ;
  assign n16330 = n16314 & n16329 ;
  assign n16331 = n14970 & n14972 ;
  assign n16332 = n14970 | n14972 ;
  assign n16333 = ~n16331 & n16332 ;
  assign n16335 = n4466 & ~n11663 ;
  assign n16336 = n4468 & n12010 ;
  assign n16337 = n16335 | n16336 ;
  assign n16334 = n4471 & ~n12616 ;
  assign n16339 = n4475 | n16334 ;
  assign n16340 = n16337 | n16339 ;
  assign n16338 = n16334 | n16337 ;
  assign n16341 = n16338 & n16340 ;
  assign n16342 = ( ~n12626 & n16340 ) | ( ~n12626 & n16341 ) | ( n16340 & n16341 ) ;
  assign n16343 = ~x17 & n16341 ;
  assign n16344 = ~x17 & n16340 ;
  assign n16345 = ( ~n12626 & n16343 ) | ( ~n12626 & n16344 ) | ( n16343 & n16344 ) ;
  assign n16346 = x17 | n16343 ;
  assign n16347 = x17 | n16344 ;
  assign n16348 = ( ~n12626 & n16346 ) | ( ~n12626 & n16347 ) | ( n16346 & n16347 ) ;
  assign n16349 = ( ~n16342 & n16345 ) | ( ~n16342 & n16348 ) | ( n16345 & n16348 ) ;
  assign n16350 = n16333 & n16349 ;
  assign n16351 = n14871 | n14968 ;
  assign n16352 = ~n14969 & n16351 ;
  assign n16354 = n4466 & n11363 ;
  assign n16355 = n4468 & ~n11663 ;
  assign n16356 = n16354 | n16355 ;
  assign n16353 = n4471 & n12010 ;
  assign n16358 = n4475 | n16353 ;
  assign n16359 = n16356 | n16358 ;
  assign n16357 = n16353 | n16356 ;
  assign n16360 = n16357 & n16359 ;
  assign n16361 = ( ~n12028 & n16359 ) | ( ~n12028 & n16360 ) | ( n16359 & n16360 ) ;
  assign n16362 = n16359 | n16360 ;
  assign n16363 = ( n12017 & n16361 ) | ( n12017 & n16362 ) | ( n16361 & n16362 ) ;
  assign n16364 = ~x17 & n16363 ;
  assign n16365 = x17 | n16363 ;
  assign n16366 = ( ~n16363 & n16364 ) | ( ~n16363 & n16365 ) | ( n16364 & n16365 ) ;
  assign n16367 = n16352 & n16366 ;
  assign n16368 = n16352 & ~n16367 ;
  assign n16369 = ~n16352 & n16366 ;
  assign n16370 = n16368 | n16369 ;
  assign n16371 = n14895 | n14966 ;
  assign n16372 = ~n14967 & n16371 ;
  assign n16373 = n4466 & n10649 ;
  assign n16374 = n4468 & n11363 ;
  assign n16375 = n16373 | n16374 ;
  assign n16376 = n4471 & ~n11663 ;
  assign n16377 = n4475 | n16376 ;
  assign n16378 = n16375 | n16377 ;
  assign n16379 = n16375 | n16376 ;
  assign n16380 = n12048 & ~n16379 ;
  assign n16381 = ( n11672 & ~n16379 ) | ( n11672 & n16380 ) | ( ~n16379 & n16380 ) ;
  assign n16382 = n16378 & ~n16381 ;
  assign n16383 = ( n12040 & n16378 ) | ( n12040 & n16382 ) | ( n16378 & n16382 ) ;
  assign n16384 = x17 & n16383 ;
  assign n16385 = x17 & ~n16383 ;
  assign n16386 = ( n16383 & ~n16384 ) | ( n16383 & n16385 ) | ( ~n16384 & n16385 ) ;
  assign n16387 = n16372 & n16386 ;
  assign n16388 = n16372 & ~n16387 ;
  assign n16389 = ~n16372 & n16386 ;
  assign n16390 = n16388 | n16389 ;
  assign n16391 = n14962 & n14964 ;
  assign n16392 = n14962 | n14964 ;
  assign n16393 = ~n16391 & n16392 ;
  assign n16394 = n4471 & n11363 ;
  assign n16395 = n4466 & n10325 ;
  assign n16396 = n4468 & n10649 ;
  assign n16397 = n16395 | n16396 ;
  assign n16398 = n16394 | n16397 ;
  assign n16399 = n4475 | n16398 ;
  assign n16400 = ( n12059 & n16398 ) | ( n12059 & n16399 ) | ( n16398 & n16399 ) ;
  assign n16401 = x17 & n16399 ;
  assign n16402 = x17 & n16398 ;
  assign n16403 = ( n12059 & n16401 ) | ( n12059 & n16402 ) | ( n16401 & n16402 ) ;
  assign n16404 = x17 & ~n16401 ;
  assign n16405 = x17 & ~n16402 ;
  assign n16406 = ( ~n12059 & n16404 ) | ( ~n12059 & n16405 ) | ( n16404 & n16405 ) ;
  assign n16407 = ( n16400 & ~n16403 ) | ( n16400 & n16406 ) | ( ~n16403 & n16406 ) ;
  assign n16408 = n16393 & n16407 ;
  assign n16409 = n14949 & n14960 ;
  assign n16410 = n14949 & ~n16409 ;
  assign n16411 = n4471 & n10649 ;
  assign n16412 = n4466 & n10654 ;
  assign n16413 = n4468 & n10325 ;
  assign n16414 = n16412 | n16413 ;
  assign n16415 = n16411 | n16414 ;
  assign n16416 = n4475 | n16411 ;
  assign n16417 = n16414 | n16416 ;
  assign n16418 = ( n10702 & n16415 ) | ( n10702 & n16417 ) | ( n16415 & n16417 ) ;
  assign n16419 = n16415 | n16417 ;
  assign n16420 = ( n10695 & n16418 ) | ( n10695 & n16419 ) | ( n16418 & n16419 ) ;
  assign n16421 = x17 & n16420 ;
  assign n16422 = x17 & ~n16420 ;
  assign n16423 = ( n16420 & ~n16421 ) | ( n16420 & n16422 ) | ( ~n16421 & n16422 ) ;
  assign n16424 = ~n14949 & n14960 ;
  assign n16425 = n16423 & n16424 ;
  assign n16426 = ( n16410 & n16423 ) | ( n16410 & n16425 ) | ( n16423 & n16425 ) ;
  assign n16427 = n16423 | n16424 ;
  assign n16428 = n16410 | n16427 ;
  assign n16429 = ~n16426 & n16428 ;
  assign n16430 = n4471 & n10325 ;
  assign n16431 = n4466 & ~n10662 ;
  assign n16432 = n4468 & n10654 ;
  assign n16433 = n16431 | n16432 ;
  assign n16434 = n16430 | n16433 ;
  assign n16435 = n4475 | n16434 ;
  assign n16436 = ( ~n10957 & n16434 ) | ( ~n10957 & n16435 ) | ( n16434 & n16435 ) ;
  assign n16437 = n16434 | n16435 ;
  assign n16438 = ( n10949 & n16436 ) | ( n10949 & n16437 ) | ( n16436 & n16437 ) ;
  assign n16439 = ~x17 & n16438 ;
  assign n16440 = x17 & n16434 ;
  assign n16441 = x17 & n4475 ;
  assign n16442 = ( x17 & n16434 ) | ( x17 & n16441 ) | ( n16434 & n16441 ) ;
  assign n16443 = ( ~n10957 & n16440 ) | ( ~n10957 & n16442 ) | ( n16440 & n16442 ) ;
  assign n16444 = n16440 | n16442 ;
  assign n16445 = ( n10949 & n16443 ) | ( n10949 & n16444 ) | ( n16443 & n16444 ) ;
  assign n16446 = x17 & ~n16445 ;
  assign n16447 = n16439 | n16446 ;
  assign n16448 = n14928 & n14946 ;
  assign n16449 = n14928 | n14946 ;
  assign n16450 = ~n16448 & n16449 ;
  assign n16451 = n16447 & n16450 ;
  assign n16452 = n16447 | n16450 ;
  assign n16453 = ~n16451 & n16452 ;
  assign n16454 = n14921 | n14924 ;
  assign n16455 = ~n14924 & n14926 ;
  assign n16456 = ( n14922 & n16454 ) | ( n14922 & ~n16455 ) | ( n16454 & ~n16455 ) ;
  assign n16457 = ~n14928 & n16456 ;
  assign n16458 = n4471 & n10654 ;
  assign n16459 = n4466 & n10667 ;
  assign n16460 = n4468 & ~n10662 ;
  assign n16461 = n16459 | n16460 ;
  assign n16462 = n16458 | n16461 ;
  assign n16463 = n4475 | n16458 ;
  assign n16464 = n16461 | n16463 ;
  assign n16465 = ( n10978 & n16462 ) | ( n10978 & n16464 ) | ( n16462 & n16464 ) ;
  assign n16466 = x17 & n16464 ;
  assign n16467 = x17 & n16462 ;
  assign n16468 = ( n10978 & n16466 ) | ( n10978 & n16467 ) | ( n16466 & n16467 ) ;
  assign n16469 = x17 & ~n16467 ;
  assign n16470 = x17 & ~n16466 ;
  assign n16471 = ( ~n10978 & n16469 ) | ( ~n10978 & n16470 ) | ( n16469 & n16470 ) ;
  assign n16472 = ( n16465 & ~n16468 ) | ( n16465 & n16471 ) | ( ~n16468 & n16471 ) ;
  assign n16473 = n16457 & n16472 ;
  assign n16474 = n4475 & n10784 ;
  assign n16475 = n4468 & ~n10678 ;
  assign n16476 = n4471 & ~n10675 ;
  assign n16477 = n16475 | n16476 ;
  assign n16478 = x17 | n16477 ;
  assign n16479 = n16474 | n16478 ;
  assign n16480 = ~x17 & n16479 ;
  assign n16481 = x17 & ~n4461 ;
  assign n16482 = ( x17 & n10678 ) | ( x17 & n16481 ) | ( n10678 & n16481 ) ;
  assign n16483 = n16479 & n16482 ;
  assign n16484 = n16474 | n16477 ;
  assign n16485 = n16482 & ~n16484 ;
  assign n16486 = ( n16480 & n16483 ) | ( n16480 & n16485 ) | ( n16483 & n16485 ) ;
  assign n16487 = n4471 & n10667 ;
  assign n16488 = n4466 & ~n10678 ;
  assign n16489 = n4468 & ~n10675 ;
  assign n16490 = n16488 | n16489 ;
  assign n16491 = n16487 | n16490 ;
  assign n16492 = n10837 | n16491 ;
  assign n16493 = n4475 | n16487 ;
  assign n16494 = n16490 | n16493 ;
  assign n16495 = ~x17 & n16494 ;
  assign n16496 = n16492 & n16495 ;
  assign n16497 = x17 | n16496 ;
  assign n16498 = n3536 & ~n10678 ;
  assign n16499 = n16496 & n16498 ;
  assign n16500 = n16492 & n16494 ;
  assign n16501 = n16498 & ~n16500 ;
  assign n16502 = ( n16497 & n16499 ) | ( n16497 & n16501 ) | ( n16499 & n16501 ) ;
  assign n16503 = n16486 & n16502 ;
  assign n16504 = ( n16496 & n16497 ) | ( n16496 & ~n16500 ) | ( n16497 & ~n16500 ) ;
  assign n16505 = n16486 | n16498 ;
  assign n16506 = ( n16498 & n16504 ) | ( n16498 & n16505 ) | ( n16504 & n16505 ) ;
  assign n16507 = ~n16503 & n16506 ;
  assign n16508 = n4471 & ~n10662 ;
  assign n16509 = n4466 & ~n10675 ;
  assign n16510 = n4468 & n10667 ;
  assign n16511 = n16509 | n16510 ;
  assign n16512 = n16508 | n16511 ;
  assign n16513 = ( n4475 & n10850 ) | ( n4475 & n16512 ) | ( n10850 & n16512 ) ;
  assign n16514 = ( x17 & n4475 ) | ( x17 & ~n16512 ) | ( n4475 & ~n16512 ) ;
  assign n16515 = ( x17 & n10850 ) | ( x17 & n16514 ) | ( n10850 & n16514 ) ;
  assign n16516 = ~n16513 & n16515 ;
  assign n16517 = n16512 | n16515 ;
  assign n16518 = ( ~x17 & n16516 ) | ( ~x17 & n16517 ) | ( n16516 & n16517 ) ;
  assign n16519 = n16503 | n16518 ;
  assign n16520 = ( n16503 & n16507 ) | ( n16503 & n16519 ) | ( n16507 & n16519 ) ;
  assign n16521 = n16457 | n16472 ;
  assign n16522 = ~n16473 & n16521 ;
  assign n16523 = n16473 | n16522 ;
  assign n16524 = ( n16473 & n16520 ) | ( n16473 & n16523 ) | ( n16520 & n16523 ) ;
  assign n16525 = n16453 & n16524 ;
  assign n16526 = n16451 | n16525 ;
  assign n16527 = n16429 & n16526 ;
  assign n16528 = n16426 | n16527 ;
  assign n16529 = ~n16393 & n16407 ;
  assign n16530 = ( n16393 & ~n16408 ) | ( n16393 & n16529 ) | ( ~n16408 & n16529 ) ;
  assign n16531 = n16408 | n16530 ;
  assign n16532 = ( n16408 & n16528 ) | ( n16408 & n16531 ) | ( n16528 & n16531 ) ;
  assign n16533 = n16390 & n16532 ;
  assign n16534 = n16387 | n16533 ;
  assign n16535 = n16370 & n16534 ;
  assign n16536 = n16367 | n16535 ;
  assign n16537 = n16333 | n16349 ;
  assign n16538 = ~n16350 & n16537 ;
  assign n16539 = n16350 | n16538 ;
  assign n16540 = ( n16350 & n16536 ) | ( n16350 & n16539 ) | ( n16536 & n16539 ) ;
  assign n16541 = n16314 | n16329 ;
  assign n16542 = ~n16330 & n16541 ;
  assign n16543 = n16330 | n16542 ;
  assign n16544 = ( n16330 & n16540 ) | ( n16330 & n16543 ) | ( n16540 & n16543 ) ;
  assign n16545 = ~n16294 & n16309 ;
  assign n16546 = n16544 & n16545 ;
  assign n16547 = ( n16311 & n16544 ) | ( n16311 & n16546 ) | ( n16544 & n16546 ) ;
  assign n16548 = n16310 | n16547 ;
  assign n16549 = ~n16276 & n16290 ;
  assign n16550 = ( n16276 & ~n16291 ) | ( n16276 & n16549 ) | ( ~n16291 & n16549 ) ;
  assign n16551 = n16291 | n16550 ;
  assign n16552 = ( n16291 & n16548 ) | ( n16291 & n16551 ) | ( n16548 & n16551 ) ;
  assign n16553 = n16273 & n16552 ;
  assign n16554 = n16234 | n16250 ;
  assign n16555 = ~n16251 & n16554 ;
  assign n16556 = n16270 & n16555 ;
  assign n16557 = ( n16553 & n16555 ) | ( n16553 & n16556 ) | ( n16555 & n16556 ) ;
  assign n16558 = n16251 | n16557 ;
  assign n16559 = n16228 | n16558 ;
  assign n16560 = ( n16228 & ~n16232 ) | ( n16228 & n16559 ) | ( ~n16232 & n16559 ) ;
  assign n16561 = ~n16207 & n16560 ;
  assign n16562 = n16205 | n16561 ;
  assign n16563 = n16183 | n16562 ;
  assign n16564 = ( n16183 & n16186 ) | ( n16183 & n16563 ) | ( n16186 & n16563 ) ;
  assign n16565 = n16156 | n16564 ;
  assign n16566 = ( n16156 & ~n16159 ) | ( n16156 & n16565 ) | ( ~n16159 & n16565 ) ;
  assign n16567 = ~n16127 & n16566 ;
  assign n16568 = n16127 & ~n16566 ;
  assign n16569 = n16567 | n16568 ;
  assign n16570 = n3547 & ~n8982 ;
  assign n16571 = ( n3547 & n9051 ) | ( n3547 & n16570 ) | ( n9051 & n16570 ) ;
  assign n16572 = n3541 & n9022 ;
  assign n16573 = n16571 | n16572 ;
  assign n16574 = n3541 | n16571 ;
  assign n16575 = ( ~n9019 & n16573 ) | ( ~n9019 & n16574 ) | ( n16573 & n16574 ) ;
  assign n16576 = n3544 | n16575 ;
  assign n16577 = ( ~n8017 & n16575 ) | ( ~n8017 & n16576 ) | ( n16575 & n16576 ) ;
  assign n16578 = n3537 | n16577 ;
  assign n16579 = ( ~n10242 & n16577 ) | ( ~n10242 & n16578 ) | ( n16577 & n16578 ) ;
  assign n16580 = ~x20 & n16578 ;
  assign n16581 = ~x20 & n16577 ;
  assign n16582 = ( ~n10242 & n16580 ) | ( ~n10242 & n16581 ) | ( n16580 & n16581 ) ;
  assign n16583 = x20 | n16580 ;
  assign n16584 = x20 | n16581 ;
  assign n16585 = ( ~n10242 & n16583 ) | ( ~n10242 & n16584 ) | ( n16583 & n16584 ) ;
  assign n16586 = ( ~n16579 & n16582 ) | ( ~n16579 & n16585 ) | ( n16582 & n16585 ) ;
  assign n16587 = n16034 | n16053 ;
  assign n16588 = ( n16034 & ~n16036 ) | ( n16034 & n16587 ) | ( ~n16036 & n16587 ) ;
  assign n16589 = n16586 & n16588 ;
  assign n16590 = n16586 | n16588 ;
  assign n16591 = ~n16589 & n16590 ;
  assign n16592 = ( n4455 & n15952 ) | ( n4455 & n15954 ) | ( n15952 & n15954 ) ;
  assign n16593 = n9101 | n15048 ;
  assign n16594 = n555 | n606 ;
  assign n16595 = n16593 | n16594 ;
  assign n16596 = n6983 | n16595 ;
  assign n16597 = n6971 | n16596 ;
  assign n16598 = n1443 | n6807 ;
  assign n16599 = n1490 | n16598 ;
  assign n16600 = n16597 | n16599 ;
  assign n16601 = n728 | n1615 ;
  assign n16602 = n2040 | n16601 ;
  assign n16603 = n667 | n2696 ;
  assign n16604 = n296 | n16603 ;
  assign n16605 = n16602 | n16604 ;
  assign n16606 = n171 | n3389 ;
  assign n16607 = n16605 | n16606 ;
  assign n16608 = n16600 | n16607 ;
  assign n16609 = n183 | n343 ;
  assign n16610 = n3308 | n16609 ;
  assign n16611 = n280 | n16610 ;
  assign n16612 = n15931 | n16611 ;
  assign n16613 = n15927 & ~n16612 ;
  assign n16614 = ~n16608 & n16613 ;
  assign n16615 = n15931 & n16611 ;
  assign n16616 = ( ~n15927 & n16611 ) | ( ~n15927 & n16615 ) | ( n16611 & n16615 ) ;
  assign n16617 = ( ~n15932 & n16608 ) | ( ~n15932 & n16616 ) | ( n16608 & n16616 ) ;
  assign n16618 = n16614 | n16617 ;
  assign n16619 = x17 & ~n16617 ;
  assign n16620 = ( ~n16617 & n16618 ) | ( ~n16617 & n16619 ) | ( n16618 & n16619 ) ;
  assign n16621 = ~n16614 & n16620 ;
  assign n16622 = ~x17 & n16618 ;
  assign n16623 = n16621 | n16622 ;
  assign n16624 = n1065 & n5192 ;
  assign n16625 = ( n1065 & n5179 ) | ( n1065 & n16624 ) | ( n5179 & n16624 ) ;
  assign n16626 = n1060 & n4245 ;
  assign n16627 = ( n1060 & n4303 ) | ( n1060 & n16626 ) | ( n4303 & n16626 ) ;
  assign n16628 = n16625 | n16627 ;
  assign n16629 = n1057 & n5117 ;
  assign n16630 = ( n1057 & ~n5037 ) | ( n1057 & n16629 ) | ( ~n5037 & n16629 ) ;
  assign n16631 = n16628 | n16630 ;
  assign n16632 = n16623 & n16631 ;
  assign n16633 = n1062 | n16625 ;
  assign n16634 = n16627 | n16633 ;
  assign n16635 = n16630 | n16634 ;
  assign n16636 = n16623 & n16635 ;
  assign n16637 = ( ~n5270 & n16632 ) | ( ~n5270 & n16636 ) | ( n16632 & n16636 ) ;
  assign n16638 = n16623 | n16631 ;
  assign n16639 = n16623 | n16635 ;
  assign n16640 = ( ~n5270 & n16638 ) | ( ~n5270 & n16639 ) | ( n16638 & n16639 ) ;
  assign n16641 = ~n16637 & n16640 ;
  assign n16642 = n16592 & n16641 ;
  assign n16643 = n16592 | n16641 ;
  assign n16644 = ~n16642 & n16643 ;
  assign n16645 = n15958 | n15977 ;
  assign n16646 = ( n15958 & ~n15961 ) | ( n15958 & n16645 ) | ( ~n15961 & n16645 ) ;
  assign n16647 = n16644 & n16646 ;
  assign n16648 = n16644 | n16646 ;
  assign n16649 = ~n16647 & n16648 ;
  assign n16650 = n1826 & n5108 ;
  assign n16651 = n1823 & n5997 ;
  assign n16652 = ( n1823 & n5979 ) | ( n1823 & n16651 ) | ( n5979 & n16651 ) ;
  assign n16653 = n16650 | n16652 ;
  assign n16654 = n1829 & n5857 ;
  assign n16655 = ( n1829 & ~n5899 ) | ( n1829 & n16654 ) | ( ~n5899 & n16654 ) ;
  assign n16656 = n16653 | n16655 ;
  assign n16657 = n1821 | n16656 ;
  assign n16658 = ( ~n6151 & n16656 ) | ( ~n6151 & n16657 ) | ( n16656 & n16657 ) ;
  assign n16659 = ~x29 & n16657 ;
  assign n16660 = ~x29 & n16656 ;
  assign n16661 = ( ~n6151 & n16659 ) | ( ~n6151 & n16660 ) | ( n16659 & n16660 ) ;
  assign n16662 = x29 | n16659 ;
  assign n16663 = x29 | n16660 ;
  assign n16664 = ( ~n6151 & n16662 ) | ( ~n6151 & n16663 ) | ( n16662 & n16663 ) ;
  assign n16665 = ( ~n16658 & n16661 ) | ( ~n16658 & n16664 ) | ( n16661 & n16664 ) ;
  assign n16666 = n16649 & n16665 ;
  assign n16667 = n16649 & ~n16666 ;
  assign n16668 = n2312 & ~n6091 ;
  assign n16669 = n2308 & n7036 ;
  assign n16670 = ( n2308 & n7023 ) | ( n2308 & n16669 ) | ( n7023 & n16669 ) ;
  assign n16671 = n16668 | n16670 ;
  assign n16672 = n2315 & n6950 ;
  assign n16673 = n16671 | n16672 ;
  assign n16674 = n2306 | n16673 ;
  assign n16675 = n16673 & n16674 ;
  assign n16676 = ( ~n7107 & n16674 ) | ( ~n7107 & n16675 ) | ( n16674 & n16675 ) ;
  assign n16677 = ~x26 & n16675 ;
  assign n16678 = ~x26 & n16674 ;
  assign n16679 = ( ~n7107 & n16677 ) | ( ~n7107 & n16678 ) | ( n16677 & n16678 ) ;
  assign n16680 = x26 | n16677 ;
  assign n16681 = x26 | n16678 ;
  assign n16682 = ( ~n7107 & n16680 ) | ( ~n7107 & n16681 ) | ( n16680 & n16681 ) ;
  assign n16683 = ( ~n16676 & n16679 ) | ( ~n16676 & n16682 ) | ( n16679 & n16682 ) ;
  assign n16684 = n16665 & n16683 ;
  assign n16685 = ~n16649 & n16684 ;
  assign n16686 = ( n16667 & n16683 ) | ( n16667 & n16685 ) | ( n16683 & n16685 ) ;
  assign n16687 = n16665 | n16683 ;
  assign n16688 = ( ~n16649 & n16683 ) | ( ~n16649 & n16687 ) | ( n16683 & n16687 ) ;
  assign n16689 = n16667 | n16688 ;
  assign n16690 = ~n16686 & n16689 ;
  assign n16691 = n15984 | n16003 ;
  assign n16692 = ( n15984 & ~n15987 ) | ( n15984 & n16691 ) | ( ~n15987 & n16691 ) ;
  assign n16693 = n16690 & n16692 ;
  assign n16694 = n16690 | n16692 ;
  assign n16695 = ~n16693 & n16694 ;
  assign n16696 = n2925 & n6889 ;
  assign n16697 = ( n2925 & ~n6884 ) | ( n2925 & n16696 ) | ( ~n6884 & n16696 ) ;
  assign n16698 = n2928 & n7907 ;
  assign n16699 = ( n2928 & n7902 ) | ( n2928 & n16698 ) | ( n7902 & n16698 ) ;
  assign n16700 = n2932 & n8079 ;
  assign n16701 = ( n2932 & ~n8070 ) | ( n2932 & n16700 ) | ( ~n8070 & n16700 ) ;
  assign n16702 = n16699 | n16701 ;
  assign n16703 = n16697 | n16702 ;
  assign n16704 = n2936 | n16703 ;
  assign n16705 = ( ~n8156 & n16703 ) | ( ~n8156 & n16704 ) | ( n16703 & n16704 ) ;
  assign n16706 = ~x23 & n16704 ;
  assign n16707 = ~x23 & n16703 ;
  assign n16708 = ( ~n8156 & n16706 ) | ( ~n8156 & n16707 ) | ( n16706 & n16707 ) ;
  assign n16709 = x23 | n16706 ;
  assign n16710 = x23 | n16707 ;
  assign n16711 = ( ~n8156 & n16709 ) | ( ~n8156 & n16710 ) | ( n16709 & n16710 ) ;
  assign n16712 = ( ~n16705 & n16708 ) | ( ~n16705 & n16711 ) | ( n16708 & n16711 ) ;
  assign n16713 = n16695 & n16712 ;
  assign n16714 = n16695 & ~n16713 ;
  assign n16716 = n16009 | n16028 ;
  assign n16717 = ( n16009 & ~n16011 ) | ( n16009 & n16716 ) | ( ~n16011 & n16716 ) ;
  assign n16715 = ~n16695 & n16712 ;
  assign n16718 = n16715 & n16717 ;
  assign n16719 = ( n16714 & n16717 ) | ( n16714 & n16718 ) | ( n16717 & n16718 ) ;
  assign n16720 = n16715 | n16717 ;
  assign n16721 = n16714 | n16720 ;
  assign n16722 = ~n16719 & n16721 ;
  assign n16723 = n16591 & n16722 ;
  assign n16724 = n16591 | n16722 ;
  assign n16725 = ~n16723 & n16724 ;
  assign n16726 = ~n15906 & n16056 ;
  assign n16727 = ( n15906 & n15908 ) | ( n15906 & ~n16726 ) | ( n15908 & ~n16726 ) ;
  assign n16728 = n16725 & n16727 ;
  assign n16729 = n16725 | n16727 ;
  assign n16730 = ~n16728 & n16729 ;
  assign n16731 = n16062 & n16730 ;
  assign n16732 = n16728 | n16731 ;
  assign n16733 = n16728 | n16730 ;
  assign n16734 = ( n16065 & n16732 ) | ( n16065 & n16733 ) | ( n16732 & n16733 ) ;
  assign n16735 = n3544 & ~n8982 ;
  assign n16736 = ( n3544 & n9051 ) | ( n3544 & n16735 ) | ( n9051 & n16735 ) ;
  assign n16737 = n3537 | n16736 ;
  assign n16738 = n9442 & ~n16736 ;
  assign n16739 = n9074 & ~n16736 ;
  assign n16740 = ( ~n9440 & n16738 ) | ( ~n9440 & n16739 ) | ( n16738 & n16739 ) ;
  assign n16741 = n16737 & ~n16740 ;
  assign n16742 = n16736 & n16737 ;
  assign n16743 = ( ~n9442 & n16737 ) | ( ~n9442 & n16742 ) | ( n16737 & n16742 ) ;
  assign n16744 = ( ~n9072 & n16741 ) | ( ~n9072 & n16743 ) | ( n16741 & n16743 ) ;
  assign n16745 = ~x20 & n16741 ;
  assign n16746 = ~x20 & n16743 ;
  assign n16747 = ( ~n9072 & n16745 ) | ( ~n9072 & n16746 ) | ( n16745 & n16746 ) ;
  assign n16748 = x20 | n16745 ;
  assign n16749 = x20 | n16746 ;
  assign n16750 = ( ~n9072 & n16748 ) | ( ~n9072 & n16749 ) | ( n16748 & n16749 ) ;
  assign n16751 = ( ~n16744 & n16747 ) | ( ~n16744 & n16750 ) | ( n16747 & n16750 ) ;
  assign n16752 = n1065 & n5117 ;
  assign n16753 = ( n1065 & ~n5037 ) | ( n1065 & n16752 ) | ( ~n5037 & n16752 ) ;
  assign n16754 = n1057 & n5108 ;
  assign n16755 = n1060 & n5192 ;
  assign n16756 = ( n1060 & n5179 ) | ( n1060 & n16755 ) | ( n5179 & n16755 ) ;
  assign n16757 = n16754 | n16756 ;
  assign n16758 = n16753 | n16757 ;
  assign n16759 = n1062 | n16758 ;
  assign n16760 = ( ~n5220 & n16758 ) | ( ~n5220 & n16759 ) | ( n16758 & n16759 ) ;
  assign n16761 = n1384 | n3312 ;
  assign n16762 = n7948 | n16761 ;
  assign n16763 = n1447 | n5072 ;
  assign n16764 = n16762 | n16763 ;
  assign n16765 = n4357 | n16764 ;
  assign n16766 = n3370 | n16765 ;
  assign n16767 = n2129 | n16766 ;
  assign n16768 = n1125 | n2625 ;
  assign n16769 = n2248 | n14364 ;
  assign n16770 = n16768 | n16769 ;
  assign n16771 = n178 | n292 ;
  assign n16772 = n1165 | n16771 ;
  assign n16773 = n175 | n447 ;
  assign n16774 = n96 | n16773 ;
  assign n16775 = n16772 | n16774 ;
  assign n16776 = n1031 | n16775 ;
  assign n16777 = n16770 | n16776 ;
  assign n16778 = n1460 | n3431 ;
  assign n16779 = n914 | n16778 ;
  assign n16780 = n2117 | n16779 ;
  assign n16781 = n112 | n309 ;
  assign n16782 = n887 | n16781 ;
  assign n16783 = n16780 | n16782 ;
  assign n16784 = n16777 | n16783 ;
  assign n16785 = n16767 | n16784 ;
  assign n16786 = n967 | n980 ;
  assign n16787 = n153 | n806 ;
  assign n16788 = n16786 | n16787 ;
  assign n16789 = n369 | n510 ;
  assign n16790 = n206 | n16789 ;
  assign n16791 = n203 | n16790 ;
  assign n16792 = n16788 | n16791 ;
  assign n16793 = n126 | n16792 ;
  assign n16794 = n680 | n869 ;
  assign n16795 = n1663 | n16794 ;
  assign n16796 = n2683 | n16795 ;
  assign n16797 = n205 | n457 ;
  assign n16798 = n92 | n16797 ;
  assign n16799 = n5901 | n16798 ;
  assign n16800 = n13870 | n16799 ;
  assign n16801 = n16796 | n16800 ;
  assign n16802 = n456 | n594 ;
  assign n16803 = n5097 | n16802 ;
  assign n16804 = n355 | n616 ;
  assign n16805 = n1114 | n16804 ;
  assign n16806 = n16803 | n16805 ;
  assign n16807 = n517 | n16806 ;
  assign n16808 = n16801 | n16807 ;
  assign n16809 = n16793 | n16808 ;
  assign n16810 = n16785 | n16809 ;
  assign n16811 = n16620 | n16810 ;
  assign n16812 = n16620 & n16810 ;
  assign n16813 = n16811 & ~n16812 ;
  assign n16814 = n16758 & n16813 ;
  assign n16815 = n16759 & n16813 ;
  assign n16816 = ( ~n5220 & n16814 ) | ( ~n5220 & n16815 ) | ( n16814 & n16815 ) ;
  assign n16817 = n16813 & ~n16815 ;
  assign n16818 = n16813 & ~n16814 ;
  assign n16819 = ( n5220 & n16817 ) | ( n5220 & n16818 ) | ( n16817 & n16818 ) ;
  assign n16820 = ( n16760 & ~n16816 ) | ( n16760 & n16819 ) | ( ~n16816 & n16819 ) ;
  assign n16821 = n16592 | n16637 ;
  assign n16822 = ( n16637 & n16641 ) | ( n16637 & n16821 ) | ( n16641 & n16821 ) ;
  assign n16823 = n16820 & n16822 ;
  assign n16824 = n16820 | n16822 ;
  assign n16825 = ~n16823 & n16824 ;
  assign n16826 = n1823 & n5857 ;
  assign n16827 = ( n1823 & ~n5899 ) | ( n1823 & n16826 ) | ( ~n5899 & n16826 ) ;
  assign n16828 = n1829 & ~n6091 ;
  assign n16829 = n1826 & n5997 ;
  assign n16830 = ( n1826 & n5979 ) | ( n1826 & n16829 ) | ( n5979 & n16829 ) ;
  assign n16831 = n16828 | n16830 ;
  assign n16832 = n16827 | n16831 ;
  assign n16833 = n1821 | n16832 ;
  assign n16834 = n16832 & n16833 ;
  assign n16835 = ( n6108 & n16833 ) | ( n6108 & n16834 ) | ( n16833 & n16834 ) ;
  assign n16836 = x29 & n16834 ;
  assign n16837 = x29 & n16833 ;
  assign n16838 = ( n6108 & n16836 ) | ( n6108 & n16837 ) | ( n16836 & n16837 ) ;
  assign n16839 = x29 & ~n16836 ;
  assign n16840 = x29 & ~n16837 ;
  assign n16841 = ( ~n6108 & n16839 ) | ( ~n6108 & n16840 ) | ( n16839 & n16840 ) ;
  assign n16842 = ( n16835 & ~n16838 ) | ( n16835 & n16841 ) | ( ~n16838 & n16841 ) ;
  assign n16843 = n16825 & n16842 ;
  assign n16844 = n16825 | n16842 ;
  assign n16845 = ~n16843 & n16844 ;
  assign n16846 = n16647 | n16665 ;
  assign n16847 = ( n16647 & n16649 ) | ( n16647 & n16846 ) | ( n16649 & n16846 ) ;
  assign n16848 = n16845 & n16847 ;
  assign n16849 = n16845 | n16847 ;
  assign n16850 = ~n16848 & n16849 ;
  assign n16851 = n2308 & n6950 ;
  assign n16852 = n2312 & n7036 ;
  assign n16853 = ( n2312 & n7023 ) | ( n2312 & n16852 ) | ( n7023 & n16852 ) ;
  assign n16854 = n16851 | n16853 ;
  assign n16855 = n2315 & n6889 ;
  assign n16856 = ( n2315 & ~n6884 ) | ( n2315 & n16855 ) | ( ~n6884 & n16855 ) ;
  assign n16857 = n16854 | n16856 ;
  assign n16858 = n2306 | n16856 ;
  assign n16859 = n16854 | n16858 ;
  assign n16860 = ( ~n7061 & n16857 ) | ( ~n7061 & n16859 ) | ( n16857 & n16859 ) ;
  assign n16861 = ~x26 & n16859 ;
  assign n16862 = ~x26 & n16857 ;
  assign n16863 = ( ~n7061 & n16861 ) | ( ~n7061 & n16862 ) | ( n16861 & n16862 ) ;
  assign n16864 = x26 | n16862 ;
  assign n16865 = x26 | n16861 ;
  assign n16866 = ( ~n7061 & n16864 ) | ( ~n7061 & n16865 ) | ( n16864 & n16865 ) ;
  assign n16867 = ( ~n16860 & n16863 ) | ( ~n16860 & n16866 ) | ( n16863 & n16866 ) ;
  assign n16868 = n16850 & ~n16867 ;
  assign n16869 = n16850 | n16867 ;
  assign n16870 = ( ~n16850 & n16868 ) | ( ~n16850 & n16869 ) | ( n16868 & n16869 ) ;
  assign n16871 = n16686 | n16692 ;
  assign n16872 = ( n16686 & n16690 ) | ( n16686 & n16871 ) | ( n16690 & n16871 ) ;
  assign n16873 = n16870 & n16872 ;
  assign n16874 = n16870 | n16872 ;
  assign n16875 = ~n16873 & n16874 ;
  assign n16876 = n2925 & n7907 ;
  assign n16877 = ( n2925 & n7902 ) | ( n2925 & n16876 ) | ( n7902 & n16876 ) ;
  assign n16878 = n2928 & n8079 ;
  assign n16879 = ( n2928 & ~n8070 ) | ( n2928 & n16878 ) | ( ~n8070 & n16878 ) ;
  assign n16880 = n16877 | n16879 ;
  assign n16881 = n2932 & ~n8017 ;
  assign n16882 = n16880 | n16881 ;
  assign n16883 = n2936 | n16880 ;
  assign n16884 = n16881 | n16883 ;
  assign n16885 = ( n8104 & n16882 ) | ( n8104 & n16884 ) | ( n16882 & n16884 ) ;
  assign n16886 = x23 & n16884 ;
  assign n16887 = x23 & n16882 ;
  assign n16888 = ( n8104 & n16886 ) | ( n8104 & n16887 ) | ( n16886 & n16887 ) ;
  assign n16889 = x23 & ~n16887 ;
  assign n16890 = x23 & ~n16886 ;
  assign n16891 = ( ~n8104 & n16889 ) | ( ~n8104 & n16890 ) | ( n16889 & n16890 ) ;
  assign n16892 = ( n16885 & ~n16888 ) | ( n16885 & n16891 ) | ( ~n16888 & n16891 ) ;
  assign n16893 = n16873 | n16892 ;
  assign n16894 = ( n16873 & n16875 ) | ( n16873 & n16893 ) | ( n16875 & n16893 ) ;
  assign n16895 = n16751 & n16894 ;
  assign n16896 = n16751 | n16894 ;
  assign n16897 = ~n16895 & n16896 ;
  assign n16898 = n1060 & n5117 ;
  assign n16899 = ( n1060 & ~n5037 ) | ( n1060 & n16898 ) | ( ~n5037 & n16898 ) ;
  assign n16900 = n1065 & n5108 ;
  assign n16901 = n1057 & n5997 ;
  assign n16902 = ( n1057 & n5979 ) | ( n1057 & n16901 ) | ( n5979 & n16901 ) ;
  assign n16903 = n16900 | n16902 ;
  assign n16904 = n16899 | n16903 ;
  assign n16905 = n1062 | n16904 ;
  assign n16906 = ( n6181 & n16904 ) | ( n6181 & n16905 ) | ( n16904 & n16905 ) ;
  assign n16907 = n5931 | n5932 ;
  assign n16908 = n1281 | n4367 ;
  assign n16909 = n2145 & ~n16908 ;
  assign n16910 = ~n16907 & n16909 ;
  assign n16911 = n182 | n1247 ;
  assign n16912 = n16910 & ~n16911 ;
  assign n16913 = ~n12986 & n16912 ;
  assign n16914 = n6801 | n13003 ;
  assign n16915 = n6054 | n12962 ;
  assign n16916 = n16914 | n16915 ;
  assign n16917 = n53 | n503 ;
  assign n16918 = n834 | n16917 ;
  assign n16919 = n175 | n477 ;
  assign n16920 = n92 | n16919 ;
  assign n16921 = n16918 | n16920 ;
  assign n16922 = n310 | n349 ;
  assign n16923 = n16921 | n16922 ;
  assign n16924 = n281 | n318 ;
  assign n16925 = n3389 | n16924 ;
  assign n16926 = n372 | n2214 ;
  assign n16927 = n16925 | n16926 ;
  assign n16928 = n16923 | n16927 ;
  assign n16929 = n16916 | n16928 ;
  assign n16930 = n728 | n5860 ;
  assign n16931 = n205 | n451 ;
  assign n16932 = n450 | n16931 ;
  assign n16933 = n16930 | n16932 ;
  assign n16934 = n344 | n16933 ;
  assign n16935 = n487 | n676 ;
  assign n16936 = n16934 | n16935 ;
  assign n16937 = n16929 | n16936 ;
  assign n16938 = n16913 & ~n16937 ;
  assign n16939 = n783 | n11076 ;
  assign n16940 = n5183 | n16939 ;
  assign n16941 = n511 | n4249 ;
  assign n16942 = n189 | n16941 ;
  assign n16943 = n16940 | n16942 ;
  assign n16944 = n333 | n16943 ;
  assign n16945 = n16938 & ~n16944 ;
  assign n16946 = n16810 & n16945 ;
  assign n16947 = n16810 | n16945 ;
  assign n16948 = n1062 & n16947 ;
  assign n16949 = ( n16904 & n16947 ) | ( n16904 & n16948 ) | ( n16947 & n16948 ) ;
  assign n16950 = ~n16946 & n16949 ;
  assign n16951 = ~n16946 & n16947 ;
  assign n16952 = n16904 & n16951 ;
  assign n16953 = ( n6181 & n16950 ) | ( n6181 & n16952 ) | ( n16950 & n16952 ) ;
  assign n16954 = n16906 & ~n16953 ;
  assign n16955 = n16811 & ~n16815 ;
  assign n16956 = n16811 & ~n16814 ;
  assign n16957 = ( n5220 & n16955 ) | ( n5220 & n16956 ) | ( n16955 & n16956 ) ;
  assign n16958 = n16946 & n16947 ;
  assign n16959 = ( n16947 & ~n16949 ) | ( n16947 & n16958 ) | ( ~n16949 & n16958 ) ;
  assign n16960 = ~n16946 & n16959 ;
  assign n16961 = n16947 & ~n16952 ;
  assign n16962 = ~n16946 & n16961 ;
  assign n16963 = ( ~n6181 & n16960 ) | ( ~n6181 & n16962 ) | ( n16960 & n16962 ) ;
  assign n16964 = ~n16957 & n16963 ;
  assign n16965 = ( n16954 & ~n16957 ) | ( n16954 & n16964 ) | ( ~n16957 & n16964 ) ;
  assign n16966 = n16957 & ~n16963 ;
  assign n16967 = ~n16954 & n16966 ;
  assign n16968 = n16965 | n16967 ;
  assign n16969 = n16823 | n16842 ;
  assign n16970 = ( n16823 & n16825 ) | ( n16823 & n16969 ) | ( n16825 & n16969 ) ;
  assign n16971 = ~n16968 & n16970 ;
  assign n16972 = n16968 & ~n16970 ;
  assign n16973 = n16971 | n16972 ;
  assign n16974 = n1826 & n5857 ;
  assign n16975 = ( n1826 & ~n5899 ) | ( n1826 & n16974 ) | ( ~n5899 & n16974 ) ;
  assign n16976 = n1823 & ~n6091 ;
  assign n16977 = n1829 & n7036 ;
  assign n16978 = ( n1829 & n7023 ) | ( n1829 & n16977 ) | ( n7023 & n16977 ) ;
  assign n16979 = n16976 | n16978 ;
  assign n16980 = n16975 | n16979 ;
  assign n16981 = n1821 | n16980 ;
  assign n16982 = n16980 & n16981 ;
  assign n16983 = ( n7136 & n16981 ) | ( n7136 & n16982 ) | ( n16981 & n16982 ) ;
  assign n16984 = x29 & n16982 ;
  assign n16985 = x29 & n16981 ;
  assign n16986 = ( n7136 & n16984 ) | ( n7136 & n16985 ) | ( n16984 & n16985 ) ;
  assign n16987 = x29 & ~n16984 ;
  assign n16988 = x29 & ~n16985 ;
  assign n16989 = ( ~n7136 & n16987 ) | ( ~n7136 & n16988 ) | ( n16987 & n16988 ) ;
  assign n16990 = ( n16983 & ~n16986 ) | ( n16983 & n16989 ) | ( ~n16986 & n16989 ) ;
  assign n16991 = ~n16973 & n16990 ;
  assign n16992 = n16973 & ~n16990 ;
  assign n16993 = n16991 | n16992 ;
  assign n16994 = n2312 & n6950 ;
  assign n16995 = n2308 & n6889 ;
  assign n16996 = ( n2308 & ~n6884 ) | ( n2308 & n16995 ) | ( ~n6884 & n16995 ) ;
  assign n16997 = n16994 | n16996 ;
  assign n16998 = n2315 & n7907 ;
  assign n16999 = ( n2315 & n7902 ) | ( n2315 & n16998 ) | ( n7902 & n16998 ) ;
  assign n17000 = n16997 | n16999 ;
  assign n17001 = n2306 | n16999 ;
  assign n17002 = n16997 | n17001 ;
  assign n17003 = ( ~n8193 & n17000 ) | ( ~n8193 & n17002 ) | ( n17000 & n17002 ) ;
  assign n17004 = ~x26 & n17002 ;
  assign n17005 = ~x26 & n17000 ;
  assign n17006 = ( ~n8193 & n17004 ) | ( ~n8193 & n17005 ) | ( n17004 & n17005 ) ;
  assign n17007 = x26 | n17005 ;
  assign n17008 = x26 | n17004 ;
  assign n17009 = ( ~n8193 & n17007 ) | ( ~n8193 & n17008 ) | ( n17007 & n17008 ) ;
  assign n17010 = ( ~n17003 & n17006 ) | ( ~n17003 & n17009 ) | ( n17006 & n17009 ) ;
  assign n17011 = n16993 | n17010 ;
  assign n17012 = n16993 & ~n17010 ;
  assign n17013 = ( ~n16993 & n17011 ) | ( ~n16993 & n17012 ) | ( n17011 & n17012 ) ;
  assign n17014 = n16848 | n16867 ;
  assign n17015 = ( n16848 & n16850 ) | ( n16848 & n17014 ) | ( n16850 & n17014 ) ;
  assign n17016 = ~n17013 & n17015 ;
  assign n17017 = n17013 & ~n17015 ;
  assign n17018 = n17016 | n17017 ;
  assign n17019 = n2925 & n8079 ;
  assign n17020 = ( n2925 & ~n8070 ) | ( n2925 & n17019 ) | ( ~n8070 & n17019 ) ;
  assign n17021 = n2928 | n17020 ;
  assign n17022 = ( ~n8017 & n17020 ) | ( ~n8017 & n17021 ) | ( n17020 & n17021 ) ;
  assign n17023 = n2932 & n9022 ;
  assign n17024 = ( n2932 & ~n9019 ) | ( n2932 & n17023 ) | ( ~n9019 & n17023 ) ;
  assign n17025 = n17022 | n17024 ;
  assign n17026 = n2936 | n17024 ;
  assign n17027 = n17022 | n17026 ;
  assign n17028 = ( ~n9416 & n17025 ) | ( ~n9416 & n17027 ) | ( n17025 & n17027 ) ;
  assign n17029 = ~x23 & n17027 ;
  assign n17030 = ~x23 & n17025 ;
  assign n17031 = ( ~n9416 & n17029 ) | ( ~n9416 & n17030 ) | ( n17029 & n17030 ) ;
  assign n17032 = x23 | n17030 ;
  assign n17033 = x23 | n17029 ;
  assign n17034 = ( ~n9416 & n17032 ) | ( ~n9416 & n17033 ) | ( n17032 & n17033 ) ;
  assign n17035 = ( ~n17028 & n17031 ) | ( ~n17028 & n17034 ) | ( n17031 & n17034 ) ;
  assign n17036 = n17018 | n17035 ;
  assign n17037 = n17018 & ~n17035 ;
  assign n17038 = ( ~n17018 & n17036 ) | ( ~n17018 & n17037 ) | ( n17036 & n17037 ) ;
  assign n17039 = n16897 & ~n17038 ;
  assign n17040 = n16897 | n17038 ;
  assign n17041 = ( ~n16897 & n17039 ) | ( ~n16897 & n17040 ) | ( n17039 & n17040 ) ;
  assign n17042 = n16713 | n16719 ;
  assign n17043 = n16875 & ~n16892 ;
  assign n17044 = n16875 | n16892 ;
  assign n17045 = ( ~n16875 & n17043 ) | ( ~n16875 & n17044 ) | ( n17043 & n17044 ) ;
  assign n17046 = n17042 & n17045 ;
  assign n17047 = n17042 | n17045 ;
  assign n17048 = ~n17046 & n17047 ;
  assign n17049 = n3541 & ~n8982 ;
  assign n17050 = ( n3541 & n9051 ) | ( n3541 & n17049 ) | ( n9051 & n17049 ) ;
  assign n17051 = n3544 & ~n9022 ;
  assign n17052 = ( n3544 & n17050 ) | ( n3544 & ~n17051 ) | ( n17050 & ~n17051 ) ;
  assign n17053 = n3544 | n17050 ;
  assign n17054 = ( ~n9019 & n17052 ) | ( ~n9019 & n17053 ) | ( n17052 & n17053 ) ;
  assign n17055 = n3537 | n17054 ;
  assign n17056 = ( n9078 & n17054 ) | ( n9078 & n17055 ) | ( n17054 & n17055 ) ;
  assign n17057 = x20 & n17055 ;
  assign n17058 = x20 & n17054 ;
  assign n17059 = ( n9078 & n17057 ) | ( n9078 & n17058 ) | ( n17057 & n17058 ) ;
  assign n17060 = x20 & ~n17057 ;
  assign n17061 = x20 & ~n17058 ;
  assign n17062 = ( ~n9078 & n17060 ) | ( ~n9078 & n17061 ) | ( n17060 & n17061 ) ;
  assign n17063 = ( n17056 & ~n17059 ) | ( n17056 & n17062 ) | ( ~n17059 & n17062 ) ;
  assign n17064 = n17046 | n17063 ;
  assign n17065 = ( n17046 & n17048 ) | ( n17046 & n17064 ) | ( n17048 & n17064 ) ;
  assign n17066 = ~n17041 & n17065 ;
  assign n17067 = n17041 & ~n17065 ;
  assign n17068 = n17066 | n17067 ;
  assign n17069 = n17048 & ~n17063 ;
  assign n17070 = n17048 | n17063 ;
  assign n17071 = ( ~n17048 & n17069 ) | ( ~n17048 & n17070 ) | ( n17069 & n17070 ) ;
  assign n17072 = n16589 | n16722 ;
  assign n17073 = ( n16589 & n16591 ) | ( n16589 & n17072 ) | ( n16591 & n17072 ) ;
  assign n17074 = n17071 & n17073 ;
  assign n17075 = n17071 | n17073 ;
  assign n17076 = ~n17074 & n17075 ;
  assign n17077 = n17074 | n17076 ;
  assign n17078 = ~n17068 & n17077 ;
  assign n17079 = ~n17068 & n17074 ;
  assign n17080 = ( n16734 & n17078 ) | ( n16734 & n17079 ) | ( n17078 & n17079 ) ;
  assign n17081 = ( ~n16064 & n16730 ) | ( ~n16064 & n16731 ) | ( n16730 & n16731 ) ;
  assign n17082 = n16728 & n17076 ;
  assign n17083 = n17074 | n17082 ;
  assign n17084 = ~n17068 & n17083 ;
  assign n17085 = ( n17078 & n17081 ) | ( n17078 & n17084 ) | ( n17081 & n17084 ) ;
  assign n17086 = ( n15882 & n17080 ) | ( n15882 & n17085 ) | ( n17080 & n17085 ) ;
  assign n17087 = ( n16734 & n17074 ) | ( n16734 & n17077 ) | ( n17074 & n17077 ) ;
  assign n17088 = n17068 & ~n17087 ;
  assign n17089 = ( n17077 & n17081 ) | ( n17077 & n17083 ) | ( n17081 & n17083 ) ;
  assign n17090 = n17068 & ~n17089 ;
  assign n17091 = ( ~n15882 & n17088 ) | ( ~n15882 & n17090 ) | ( n17088 & n17090 ) ;
  assign n17092 = n17086 | n17091 ;
  assign n17093 = n16734 & n17076 ;
  assign n17094 = ( n17076 & n17081 ) | ( n17076 & n17082 ) | ( n17081 & n17082 ) ;
  assign n17095 = ( n15882 & n17093 ) | ( n15882 & n17094 ) | ( n17093 & n17094 ) ;
  assign n17096 = n16734 | n17076 ;
  assign n17097 = n16728 | n17081 ;
  assign n17098 = n17076 | n17097 ;
  assign n17099 = ( n15882 & n17096 ) | ( n15882 & n17098 ) | ( n17096 & n17098 ) ;
  assign n17100 = ~n17095 & n17099 ;
  assign n17101 = ~n17092 & n17100 ;
  assign n17102 = n17092 & ~n17100 ;
  assign n17103 = n17101 | n17102 ;
  assign n17104 = ( n16065 & n16730 ) | ( n16065 & n16731 ) | ( n16730 & n16731 ) ;
  assign n17105 = ( n15882 & n17081 ) | ( n15882 & n17104 ) | ( n17081 & n17104 ) ;
  assign n17106 = n16062 | n16065 ;
  assign n17107 = n16730 | n17106 ;
  assign n17108 = ~n16062 & n16064 ;
  assign n17109 = ~n16730 & n17108 ;
  assign n17110 = ( n15882 & n17107 ) | ( n15882 & ~n17109 ) | ( n17107 & ~n17109 ) ;
  assign n17111 = ~n17105 & n17110 ;
  assign n17112 = n17100 & n17111 ;
  assign n17113 = n17100 | n17111 ;
  assign n17114 = ~n17112 & n17113 ;
  assign n17115 = ~n16069 & n17111 ;
  assign n17116 = n17112 | n17115 ;
  assign n17117 = ( n17112 & n17114 ) | ( n17112 & n17116 ) | ( n17114 & n17116 ) ;
  assign n17118 = ~n17103 & n17117 ;
  assign n17119 = n17112 | n17114 ;
  assign n17120 = ~n17103 & n17119 ;
  assign n17121 = n16069 & ~n17111 ;
  assign n17122 = n16070 | n16098 ;
  assign n17123 = ~n16070 & n16072 ;
  assign n17124 = ( ~n16070 & n16094 ) | ( ~n16070 & n17123 ) | ( n16094 & n17123 ) ;
  assign n17125 = ~n17122 & n17124 ;
  assign n17126 = n17121 | n17125 ;
  assign n17127 = ( n15435 & n17122 ) | ( n15435 & ~n17124 ) | ( n17122 & ~n17124 ) ;
  assign n17128 = ~n17121 & n17127 ;
  assign n17129 = ( n15446 & ~n17126 ) | ( n15446 & n17128 ) | ( ~n17126 & n17128 ) ;
  assign n17130 = ( n17118 & n17120 ) | ( n17118 & n17129 ) | ( n17120 & n17129 ) ;
  assign n17131 = n17103 & ~n17117 ;
  assign n17132 = n17103 & ~n17119 ;
  assign n17133 = ( ~n17129 & n17131 ) | ( ~n17129 & n17132 ) | ( n17131 & n17132 ) ;
  assign n17134 = n17130 | n17133 ;
  assign n17136 = n5237 & n17111 ;
  assign n17137 = n5231 & n17100 ;
  assign n17138 = n17136 | n17137 ;
  assign n17135 = n5234 & ~n17092 ;
  assign n17140 = n5227 | n17135 ;
  assign n17141 = n17138 | n17140 ;
  assign n17139 = n17135 | n17138 ;
  assign n17142 = n17139 & n17141 ;
  assign n17143 = ( ~n17134 & n17141 ) | ( ~n17134 & n17142 ) | ( n17141 & n17142 ) ;
  assign n17144 = ~x14 & n17142 ;
  assign n17145 = ~x14 & n17141 ;
  assign n17146 = ( ~n17134 & n17144 ) | ( ~n17134 & n17145 ) | ( n17144 & n17145 ) ;
  assign n17147 = x14 | n17144 ;
  assign n17148 = x14 | n17145 ;
  assign n17149 = ( ~n17134 & n17147 ) | ( ~n17134 & n17148 ) | ( n17147 & n17148 ) ;
  assign n17150 = ( ~n17143 & n17146 ) | ( ~n17143 & n17149 ) | ( n17146 & n17149 ) ;
  assign n17151 = ~n16569 & n17150 ;
  assign n17152 = n16569 | n17151 ;
  assign n17153 = n16569 & n17150 ;
  assign n17154 = n17152 & ~n17153 ;
  assign n17155 = ~n16159 & n16564 ;
  assign n17156 = n16159 & ~n16564 ;
  assign n17157 = n17155 | n17156 ;
  assign n17158 = n17115 | n17129 ;
  assign n17159 = n17114 & n17115 ;
  assign n17160 = ( n17114 & n17129 ) | ( n17114 & n17159 ) | ( n17129 & n17159 ) ;
  assign n17161 = n17158 & ~n17160 ;
  assign n17162 = n5237 & ~n16069 ;
  assign n17163 = n5231 & n17111 ;
  assign n17164 = n17162 | n17163 ;
  assign n17165 = n5234 & n17100 ;
  assign n17166 = n5227 | n17165 ;
  assign n17167 = n17164 | n17166 ;
  assign n17168 = n17164 | n17165 ;
  assign n17169 = n17113 & ~n17117 ;
  assign n17170 = n17168 | n17169 ;
  assign n17171 = ( ~n17129 & n17168 ) | ( ~n17129 & n17170 ) | ( n17168 & n17170 ) ;
  assign n17172 = n17167 & n17171 ;
  assign n17173 = ( n17161 & n17167 ) | ( n17161 & n17172 ) | ( n17167 & n17172 ) ;
  assign n17174 = ~x14 & n17173 ;
  assign n17175 = x14 | n17173 ;
  assign n17176 = ( ~n17173 & n17174 ) | ( ~n17173 & n17175 ) | ( n17174 & n17175 ) ;
  assign n17177 = ~n17157 & n17176 ;
  assign n17178 = n17157 | n17177 ;
  assign n17179 = n17157 & n17176 ;
  assign n17180 = n17178 & ~n17179 ;
  assign n17181 = n16186 & n16562 ;
  assign n17182 = n16186 | n16562 ;
  assign n17183 = ~n17181 & n17182 ;
  assign n17184 = ~n17115 & n17129 ;
  assign n17185 = ( n15446 & ~n17125 ) | ( n15446 & n17127 ) | ( ~n17125 & n17127 ) ;
  assign n17186 = ~n17184 & n17185 ;
  assign n17187 = n5237 & n15886 ;
  assign n17188 = n5231 & ~n16069 ;
  assign n17189 = n17187 | n17188 ;
  assign n17190 = n5234 & n17111 ;
  assign n17191 = n5227 | n17190 ;
  assign n17192 = n17189 | n17191 ;
  assign n17193 = n17189 | n17190 ;
  assign n17194 = n17115 | n17121 ;
  assign n17195 = ~n17193 & n17194 ;
  assign n17196 = ( n17129 & ~n17193 ) | ( n17129 & n17195 ) | ( ~n17193 & n17195 ) ;
  assign n17197 = n17192 & ~n17196 ;
  assign n17198 = ( n17186 & n17192 ) | ( n17186 & n17197 ) | ( n17192 & n17197 ) ;
  assign n17199 = x14 & n17198 ;
  assign n17200 = x14 & ~n17198 ;
  assign n17201 = ( n17198 & ~n17199 ) | ( n17198 & n17200 ) | ( ~n17199 & n17200 ) ;
  assign n17202 = n17183 & n17201 ;
  assign n17203 = n17183 & ~n17202 ;
  assign n17204 = ~n17183 & n17201 ;
  assign n17205 = n17203 | n17204 ;
  assign n17206 = n16207 & ~n16560 ;
  assign n17207 = n16561 | n17206 ;
  assign n17208 = n5234 & ~n16069 ;
  assign n17209 = n5237 & ~n16085 ;
  assign n17210 = n5231 & n15886 ;
  assign n17211 = n17209 | n17210 ;
  assign n17212 = n17208 | n17211 ;
  assign n17213 = n5227 | n17212 ;
  assign n17214 = ( ~n16107 & n17212 ) | ( ~n16107 & n17213 ) | ( n17212 & n17213 ) ;
  assign n17215 = ~x14 & n17213 ;
  assign n17216 = ~x14 & n17212 ;
  assign n17217 = ( ~n16107 & n17215 ) | ( ~n16107 & n17216 ) | ( n17215 & n17216 ) ;
  assign n17218 = x14 | n17215 ;
  assign n17219 = x14 | n17216 ;
  assign n17220 = ( ~n16107 & n17218 ) | ( ~n16107 & n17219 ) | ( n17218 & n17219 ) ;
  assign n17221 = ( ~n17214 & n17217 ) | ( ~n17214 & n17220 ) | ( n17217 & n17220 ) ;
  assign n17222 = ~n17207 & n17221 ;
  assign n17223 = n17207 | n17222 ;
  assign n17224 = n17207 & n17221 ;
  assign n17225 = n17223 & ~n17224 ;
  assign n17226 = ~n16232 & n16558 ;
  assign n17227 = n16232 & ~n16558 ;
  assign n17228 = n17226 | n17227 ;
  assign n17230 = n5237 & n15434 ;
  assign n17231 = n5231 & ~n16085 ;
  assign n17232 = n17230 | n17231 ;
  assign n17229 = n5234 & n15886 ;
  assign n17234 = n5227 | n17229 ;
  assign n17235 = n17232 | n17234 ;
  assign n17233 = n17229 | n17232 ;
  assign n17236 = n17233 & n17235 ;
  assign n17237 = ( ~n16140 & n17235 ) | ( ~n16140 & n17236 ) | ( n17235 & n17236 ) ;
  assign n17238 = ~x14 & n17236 ;
  assign n17239 = ~x14 & n17235 ;
  assign n17240 = ( ~n16140 & n17238 ) | ( ~n16140 & n17239 ) | ( n17238 & n17239 ) ;
  assign n17241 = x14 | n17238 ;
  assign n17242 = x14 | n17239 ;
  assign n17243 = ( ~n16140 & n17241 ) | ( ~n16140 & n17242 ) | ( n17241 & n17242 ) ;
  assign n17244 = ( ~n17237 & n17240 ) | ( ~n17237 & n17243 ) | ( n17240 & n17243 ) ;
  assign n17245 = ~n17228 & n17244 ;
  assign n17246 = n17228 | n17245 ;
  assign n17247 = n17228 & n17244 ;
  assign n17248 = n17246 & ~n17247 ;
  assign n17249 = n16270 | n16555 ;
  assign n17250 = n16553 | n17249 ;
  assign n17251 = ~n16557 & n17250 ;
  assign n17252 = n5234 & ~n16085 ;
  assign n17253 = n5237 & n14591 ;
  assign n17254 = n5231 & n15434 ;
  assign n17255 = n17253 | n17254 ;
  assign n17256 = n17252 | n17255 ;
  assign n17257 = n5227 | n17252 ;
  assign n17258 = n17255 | n17257 ;
  assign n17259 = ( ~n16167 & n17256 ) | ( ~n16167 & n17258 ) | ( n17256 & n17258 ) ;
  assign n17260 = ~x14 & n17258 ;
  assign n17261 = ~x14 & n17256 ;
  assign n17262 = ( ~n16167 & n17260 ) | ( ~n16167 & n17261 ) | ( n17260 & n17261 ) ;
  assign n17263 = x14 | n17261 ;
  assign n17264 = x14 | n17260 ;
  assign n17265 = ( ~n16167 & n17263 ) | ( ~n16167 & n17264 ) | ( n17263 & n17264 ) ;
  assign n17266 = ( ~n17259 & n17262 ) | ( ~n17259 & n17265 ) | ( n17262 & n17265 ) ;
  assign n17267 = n17251 & n17266 ;
  assign n17268 = n16552 & ~n16553 ;
  assign n17269 = n16273 & ~n16553 ;
  assign n17270 = n17268 | n17269 ;
  assign n17271 = n5234 & n15434 ;
  assign n17272 = n5237 & n14329 ;
  assign n17273 = n5231 & n14591 ;
  assign n17274 = n17272 | n17273 ;
  assign n17275 = n17271 | n17274 ;
  assign n17276 = n5227 | n17271 ;
  assign n17277 = n17274 | n17276 ;
  assign n17278 = ( n15453 & n17275 ) | ( n15453 & n17277 ) | ( n17275 & n17277 ) ;
  assign n17279 = x14 & n17277 ;
  assign n17280 = x14 & n17275 ;
  assign n17281 = ( n15453 & n17279 ) | ( n15453 & n17280 ) | ( n17279 & n17280 ) ;
  assign n17282 = x14 & ~n17280 ;
  assign n17283 = x14 & ~n17279 ;
  assign n17284 = ( ~n15453 & n17282 ) | ( ~n15453 & n17283 ) | ( n17282 & n17283 ) ;
  assign n17285 = ( n17278 & ~n17281 ) | ( n17278 & n17284 ) | ( ~n17281 & n17284 ) ;
  assign n17286 = n17270 & n17285 ;
  assign n17287 = n17270 & ~n17286 ;
  assign n17288 = ~n17270 & n17285 ;
  assign n17289 = n17287 | n17288 ;
  assign n17290 = n16544 | n16545 ;
  assign n17291 = n16311 | n17290 ;
  assign n17292 = ~n16547 & n17291 ;
  assign n17294 = n5237 & n13522 ;
  assign n17295 = n5231 & n14607 ;
  assign n17296 = n17294 | n17295 ;
  assign n17293 = n5234 & n14329 ;
  assign n17298 = n5227 | n17293 ;
  assign n17299 = n17296 | n17298 ;
  assign n17297 = n17293 | n17296 ;
  assign n17300 = n17297 & n17299 ;
  assign n17301 = ( n14656 & n17299 ) | ( n14656 & n17300 ) | ( n17299 & n17300 ) ;
  assign n17302 = x14 & n17300 ;
  assign n17303 = x14 & n17299 ;
  assign n17304 = ( n14656 & n17302 ) | ( n14656 & n17303 ) | ( n17302 & n17303 ) ;
  assign n17305 = x14 & ~n17302 ;
  assign n17306 = x14 & ~n17303 ;
  assign n17307 = ( ~n14656 & n17305 ) | ( ~n14656 & n17306 ) | ( n17305 & n17306 ) ;
  assign n17308 = ( n17301 & ~n17304 ) | ( n17301 & n17307 ) | ( ~n17304 & n17307 ) ;
  assign n17309 = n17292 & n17308 ;
  assign n17310 = n16548 & n16550 ;
  assign n17311 = n16548 | n16550 ;
  assign n17312 = ~n17310 & n17311 ;
  assign n17314 = n5237 & n14607 ;
  assign n17315 = n5231 & n14329 ;
  assign n17316 = n17314 | n17315 ;
  assign n17313 = n5234 & n14591 ;
  assign n17318 = n5227 | n17313 ;
  assign n17319 = n17316 | n17318 ;
  assign n17317 = n17313 | n17316 ;
  assign n17320 = n17317 & n17319 ;
  assign n17321 = ( n14629 & n17319 ) | ( n14629 & n17320 ) | ( n17319 & n17320 ) ;
  assign n17322 = x14 & n17320 ;
  assign n17323 = x14 & n17319 ;
  assign n17324 = ( n14629 & n17322 ) | ( n14629 & n17323 ) | ( n17322 & n17323 ) ;
  assign n17325 = x14 & ~n17322 ;
  assign n17326 = x14 & ~n17323 ;
  assign n17327 = ( ~n14629 & n17325 ) | ( ~n14629 & n17326 ) | ( n17325 & n17326 ) ;
  assign n17328 = ( n17321 & ~n17324 ) | ( n17321 & n17327 ) | ( ~n17324 & n17327 ) ;
  assign n17329 = n17312 & n17328 ;
  assign n17330 = n17312 | n17328 ;
  assign n17331 = ~n17329 & n17330 ;
  assign n17332 = n17309 & n17331 ;
  assign n17333 = n17329 | n17331 ;
  assign n17334 = n16540 & n16542 ;
  assign n17335 = n16540 | n16542 ;
  assign n17336 = ~n17334 & n17335 ;
  assign n17337 = n5237 & n13235 ;
  assign n17338 = n5231 & n13522 ;
  assign n17339 = n17337 | n17338 ;
  assign n17340 = n5234 & n14607 ;
  assign n17341 = n5227 | n17340 ;
  assign n17342 = n17339 | n17341 ;
  assign n17343 = n17339 | n17340 ;
  assign n17344 = n14696 | n17343 ;
  assign n17345 = n14698 | n17343 ;
  assign n17346 = ( ~n13248 & n17344 ) | ( ~n13248 & n17345 ) | ( n17344 & n17345 ) ;
  assign n17347 = n17342 & n17346 ;
  assign n17348 = ( n14687 & n17342 ) | ( n14687 & n17347 ) | ( n17342 & n17347 ) ;
  assign n17349 = ~x14 & n17348 ;
  assign n17350 = x14 | n17348 ;
  assign n17351 = ( ~n17348 & n17349 ) | ( ~n17348 & n17350 ) | ( n17349 & n17350 ) ;
  assign n17352 = n17336 & n17351 ;
  assign n17353 = n17336 & ~n17352 ;
  assign n17354 = ~n17336 & n17351 ;
  assign n17355 = n17353 | n17354 ;
  assign n17356 = n16536 & n16538 ;
  assign n17357 = n16536 | n16538 ;
  assign n17358 = ~n17356 & n17357 ;
  assign n17359 = n5234 & n13522 ;
  assign n17360 = n5237 & n12936 ;
  assign n17361 = n5231 & n13235 ;
  assign n17362 = n17360 | n17361 ;
  assign n17363 = n17359 | n17362 ;
  assign n17364 = n5227 & n13537 ;
  assign n17365 = n5227 & n13539 ;
  assign n17366 = ( ~n13248 & n17364 ) | ( ~n13248 & n17365 ) | ( n17364 & n17365 ) ;
  assign n17367 = n17363 | n17366 ;
  assign n17368 = n5227 | n17363 ;
  assign n17369 = ( n13530 & n17367 ) | ( n13530 & n17368 ) | ( n17367 & n17368 ) ;
  assign n17370 = x14 | n17369 ;
  assign n17371 = ~x14 & n17369 ;
  assign n17372 = ( ~n17369 & n17370 ) | ( ~n17369 & n17371 ) | ( n17370 & n17371 ) ;
  assign n17373 = n17358 & n17372 ;
  assign n17374 = n16534 & ~n16535 ;
  assign n17375 = n16370 & ~n16535 ;
  assign n17376 = n17374 | n17375 ;
  assign n17377 = n5234 & n13235 ;
  assign n17378 = n5237 & ~n12616 ;
  assign n17379 = n5231 & n12936 ;
  assign n17380 = n17378 | n17379 ;
  assign n17381 = n17377 | n17380 ;
  assign n17382 = n5227 | n17377 ;
  assign n17383 = n17380 | n17382 ;
  assign n17384 = ( n13561 & n17381 ) | ( n13561 & n17383 ) | ( n17381 & n17383 ) ;
  assign n17385 = x14 & n17383 ;
  assign n17386 = x14 & n17381 ;
  assign n17387 = ( n13561 & n17385 ) | ( n13561 & n17386 ) | ( n17385 & n17386 ) ;
  assign n17388 = x14 & ~n17386 ;
  assign n17389 = x14 & ~n17385 ;
  assign n17390 = ( ~n13561 & n17388 ) | ( ~n13561 & n17389 ) | ( n17388 & n17389 ) ;
  assign n17391 = ( n17384 & ~n17387 ) | ( n17384 & n17390 ) | ( ~n17387 & n17390 ) ;
  assign n17392 = n17376 & n17391 ;
  assign n17393 = n17376 & ~n17392 ;
  assign n17394 = ~n16390 & n16532 ;
  assign n17395 = n16390 & ~n16532 ;
  assign n17396 = n17394 | n17395 ;
  assign n17397 = n5234 & n12936 ;
  assign n17398 = n5237 & n12010 ;
  assign n17399 = n5231 & ~n12616 ;
  assign n17400 = n17398 | n17399 ;
  assign n17401 = n17397 | n17400 ;
  assign n17402 = n5227 | n17397 ;
  assign n17403 = n17400 | n17402 ;
  assign n17404 = ( ~n13591 & n17401 ) | ( ~n13591 & n17403 ) | ( n17401 & n17403 ) ;
  assign n17405 = ~x14 & n17403 ;
  assign n17406 = ~x14 & n17401 ;
  assign n17407 = ( ~n13591 & n17405 ) | ( ~n13591 & n17406 ) | ( n17405 & n17406 ) ;
  assign n17408 = x14 | n17406 ;
  assign n17409 = x14 | n17405 ;
  assign n17410 = ( ~n13591 & n17408 ) | ( ~n13591 & n17409 ) | ( n17408 & n17409 ) ;
  assign n17411 = ( ~n17404 & n17407 ) | ( ~n17404 & n17410 ) | ( n17407 & n17410 ) ;
  assign n17412 = n17396 & n17411 ;
  assign n17413 = n16528 & n16530 ;
  assign n17414 = n16528 | n16530 ;
  assign n17415 = ~n17413 & n17414 ;
  assign n17417 = n5237 & ~n11663 ;
  assign n17418 = n5231 & n12010 ;
  assign n17419 = n17417 | n17418 ;
  assign n17416 = n5234 & ~n12616 ;
  assign n17421 = n5227 | n17416 ;
  assign n17422 = n17419 | n17421 ;
  assign n17420 = n17416 | n17419 ;
  assign n17423 = n17420 & n17422 ;
  assign n17424 = ( ~n12626 & n17422 ) | ( ~n12626 & n17423 ) | ( n17422 & n17423 ) ;
  assign n17425 = ~x14 & n17423 ;
  assign n17426 = ~x14 & n17422 ;
  assign n17427 = ( ~n12626 & n17425 ) | ( ~n12626 & n17426 ) | ( n17425 & n17426 ) ;
  assign n17428 = x14 | n17425 ;
  assign n17429 = x14 | n17426 ;
  assign n17430 = ( ~n12626 & n17428 ) | ( ~n12626 & n17429 ) | ( n17428 & n17429 ) ;
  assign n17431 = ( ~n17424 & n17427 ) | ( ~n17424 & n17430 ) | ( n17427 & n17430 ) ;
  assign n17432 = n17415 & n17431 ;
  assign n17433 = n16429 | n16526 ;
  assign n17434 = ~n16527 & n17433 ;
  assign n17436 = n5237 & n11363 ;
  assign n17437 = n5231 & ~n11663 ;
  assign n17438 = n17436 | n17437 ;
  assign n17435 = n5234 & n12010 ;
  assign n17440 = n5227 | n17435 ;
  assign n17441 = n17438 | n17440 ;
  assign n17439 = n17435 | n17438 ;
  assign n17442 = n17439 & n17441 ;
  assign n17443 = ( ~n12028 & n17441 ) | ( ~n12028 & n17442 ) | ( n17441 & n17442 ) ;
  assign n17444 = n17441 | n17442 ;
  assign n17445 = ( n12017 & n17443 ) | ( n12017 & n17444 ) | ( n17443 & n17444 ) ;
  assign n17446 = ~x14 & n17445 ;
  assign n17447 = x14 | n17445 ;
  assign n17448 = ( ~n17445 & n17446 ) | ( ~n17445 & n17447 ) | ( n17446 & n17447 ) ;
  assign n17449 = n17434 & n17448 ;
  assign n17450 = n17434 & ~n17449 ;
  assign n17451 = ~n17434 & n17448 ;
  assign n17452 = n17450 | n17451 ;
  assign n17453 = n16453 | n16524 ;
  assign n17454 = ~n16525 & n17453 ;
  assign n17455 = n5237 & n10649 ;
  assign n17456 = n5231 & n11363 ;
  assign n17457 = n17455 | n17456 ;
  assign n17458 = n5234 & ~n11663 ;
  assign n17459 = n5227 | n17458 ;
  assign n17460 = n17457 | n17459 ;
  assign n17461 = n17457 | n17458 ;
  assign n17462 = n12048 & ~n17461 ;
  assign n17463 = ( n11672 & ~n17461 ) | ( n11672 & n17462 ) | ( ~n17461 & n17462 ) ;
  assign n17464 = n17460 & ~n17463 ;
  assign n17465 = ( n12040 & n17460 ) | ( n12040 & n17464 ) | ( n17460 & n17464 ) ;
  assign n17466 = x14 & n17465 ;
  assign n17467 = x14 & ~n17465 ;
  assign n17468 = ( n17465 & ~n17466 ) | ( n17465 & n17467 ) | ( ~n17466 & n17467 ) ;
  assign n17469 = n17454 & n17468 ;
  assign n17470 = n17454 & ~n17469 ;
  assign n17471 = ~n17454 & n17468 ;
  assign n17472 = n17470 | n17471 ;
  assign n17473 = n16520 & n16522 ;
  assign n17474 = n16520 | n16522 ;
  assign n17475 = ~n17473 & n17474 ;
  assign n17476 = n5234 & n11363 ;
  assign n17477 = n5237 & n10325 ;
  assign n17478 = n5231 & n10649 ;
  assign n17479 = n17477 | n17478 ;
  assign n17480 = n17476 | n17479 ;
  assign n17481 = n5227 | n17480 ;
  assign n17482 = ( n12059 & n17480 ) | ( n12059 & n17481 ) | ( n17480 & n17481 ) ;
  assign n17483 = x14 & n17481 ;
  assign n17484 = x14 & n17480 ;
  assign n17485 = ( n12059 & n17483 ) | ( n12059 & n17484 ) | ( n17483 & n17484 ) ;
  assign n17486 = x14 & ~n17483 ;
  assign n17487 = x14 & ~n17484 ;
  assign n17488 = ( ~n12059 & n17486 ) | ( ~n12059 & n17487 ) | ( n17486 & n17487 ) ;
  assign n17489 = ( n17482 & ~n17485 ) | ( n17482 & n17488 ) | ( ~n17485 & n17488 ) ;
  assign n17490 = n17475 & n17489 ;
  assign n17491 = n16507 & n16518 ;
  assign n17492 = n16507 & ~n17491 ;
  assign n17493 = n5234 & n10649 ;
  assign n17494 = n5237 & n10654 ;
  assign n17495 = n5231 & n10325 ;
  assign n17496 = n17494 | n17495 ;
  assign n17497 = n17493 | n17496 ;
  assign n17498 = n5227 | n17493 ;
  assign n17499 = n17496 | n17498 ;
  assign n17500 = ( n10702 & n17497 ) | ( n10702 & n17499 ) | ( n17497 & n17499 ) ;
  assign n17501 = n17497 | n17499 ;
  assign n17502 = ( n10695 & n17500 ) | ( n10695 & n17501 ) | ( n17500 & n17501 ) ;
  assign n17503 = x14 & n17502 ;
  assign n17504 = x14 & ~n17502 ;
  assign n17505 = ( n17502 & ~n17503 ) | ( n17502 & n17504 ) | ( ~n17503 & n17504 ) ;
  assign n17506 = ~n16507 & n16518 ;
  assign n17507 = n17505 & n17506 ;
  assign n17508 = ( n17492 & n17505 ) | ( n17492 & n17507 ) | ( n17505 & n17507 ) ;
  assign n17509 = n17505 | n17506 ;
  assign n17510 = n17492 | n17509 ;
  assign n17511 = ~n17508 & n17510 ;
  assign n17512 = n5234 & n10325 ;
  assign n17513 = n5237 & ~n10662 ;
  assign n17514 = n5231 & n10654 ;
  assign n17515 = n17513 | n17514 ;
  assign n17516 = n17512 | n17515 ;
  assign n17517 = n5227 | n17516 ;
  assign n17518 = ( ~n10957 & n17516 ) | ( ~n10957 & n17517 ) | ( n17516 & n17517 ) ;
  assign n17519 = n17516 | n17517 ;
  assign n17520 = ( n10949 & n17518 ) | ( n10949 & n17519 ) | ( n17518 & n17519 ) ;
  assign n17521 = ~x14 & n17520 ;
  assign n17522 = x14 & n17516 ;
  assign n17523 = x14 & n5227 ;
  assign n17524 = ( x14 & n17516 ) | ( x14 & n17523 ) | ( n17516 & n17523 ) ;
  assign n17525 = ( ~n10957 & n17522 ) | ( ~n10957 & n17524 ) | ( n17522 & n17524 ) ;
  assign n17526 = n17522 | n17524 ;
  assign n17527 = ( n10949 & n17525 ) | ( n10949 & n17526 ) | ( n17525 & n17526 ) ;
  assign n17528 = x14 & ~n17527 ;
  assign n17529 = n17521 | n17528 ;
  assign n17530 = n16486 & n16504 ;
  assign n17531 = n16486 | n16504 ;
  assign n17532 = ~n17530 & n17531 ;
  assign n17533 = n17529 & n17532 ;
  assign n17534 = n17529 | n17532 ;
  assign n17535 = ~n17533 & n17534 ;
  assign n17536 = n16479 | n16482 ;
  assign n17537 = ~n16482 & n16484 ;
  assign n17538 = ( n16480 & n17536 ) | ( n16480 & ~n17537 ) | ( n17536 & ~n17537 ) ;
  assign n17539 = ~n16486 & n17538 ;
  assign n17540 = n5234 & n10654 ;
  assign n17541 = n5237 & n10667 ;
  assign n17542 = n5231 & ~n10662 ;
  assign n17543 = n17541 | n17542 ;
  assign n17544 = n17540 | n17543 ;
  assign n17545 = n5227 | n17540 ;
  assign n17546 = n17543 | n17545 ;
  assign n17547 = ( n10978 & n17544 ) | ( n10978 & n17546 ) | ( n17544 & n17546 ) ;
  assign n17548 = x14 & n17546 ;
  assign n17549 = x14 & n17544 ;
  assign n17550 = ( n10978 & n17548 ) | ( n10978 & n17549 ) | ( n17548 & n17549 ) ;
  assign n17551 = x14 & ~n17549 ;
  assign n17552 = x14 & ~n17548 ;
  assign n17553 = ( ~n10978 & n17551 ) | ( ~n10978 & n17552 ) | ( n17551 & n17552 ) ;
  assign n17554 = ( n17547 & ~n17550 ) | ( n17547 & n17553 ) | ( ~n17550 & n17553 ) ;
  assign n17555 = n17539 & n17554 ;
  assign n17556 = n5227 & n10784 ;
  assign n17557 = n5231 & ~n10678 ;
  assign n17558 = n5234 & ~n10675 ;
  assign n17559 = n17557 | n17558 ;
  assign n17560 = x14 | n17559 ;
  assign n17561 = n17556 | n17560 ;
  assign n17562 = ~x14 & n17561 ;
  assign n17563 = x14 & ~n5223 ;
  assign n17564 = ( x14 & n10678 ) | ( x14 & n17563 ) | ( n10678 & n17563 ) ;
  assign n17565 = n17561 & n17564 ;
  assign n17566 = n17556 | n17559 ;
  assign n17567 = n17564 & ~n17566 ;
  assign n17568 = ( n17562 & n17565 ) | ( n17562 & n17567 ) | ( n17565 & n17567 ) ;
  assign n17569 = n5234 & n10667 ;
  assign n17570 = n5237 & ~n10678 ;
  assign n17571 = n5231 & ~n10675 ;
  assign n17572 = n17570 | n17571 ;
  assign n17573 = n17569 | n17572 ;
  assign n17574 = n10837 | n17573 ;
  assign n17575 = n5227 | n17569 ;
  assign n17576 = n17572 | n17575 ;
  assign n17577 = ~x14 & n17576 ;
  assign n17578 = n17574 & n17577 ;
  assign n17579 = x14 | n17578 ;
  assign n17580 = n4461 & ~n10678 ;
  assign n17581 = n17578 & n17580 ;
  assign n17582 = n17574 & n17576 ;
  assign n17583 = n17580 & ~n17582 ;
  assign n17584 = ( n17579 & n17581 ) | ( n17579 & n17583 ) | ( n17581 & n17583 ) ;
  assign n17585 = n17568 & n17584 ;
  assign n17586 = ( n17578 & n17579 ) | ( n17578 & ~n17582 ) | ( n17579 & ~n17582 ) ;
  assign n17587 = n17568 | n17580 ;
  assign n17588 = ( n17580 & n17586 ) | ( n17580 & n17587 ) | ( n17586 & n17587 ) ;
  assign n17589 = ~n17585 & n17588 ;
  assign n17590 = n5234 & ~n10662 ;
  assign n17591 = n5237 & ~n10675 ;
  assign n17592 = n5231 & n10667 ;
  assign n17593 = n17591 | n17592 ;
  assign n17594 = n17590 | n17593 ;
  assign n17595 = ( n5227 & n10850 ) | ( n5227 & n17594 ) | ( n10850 & n17594 ) ;
  assign n17596 = ( x14 & n5227 ) | ( x14 & ~n17594 ) | ( n5227 & ~n17594 ) ;
  assign n17597 = ( x14 & n10850 ) | ( x14 & n17596 ) | ( n10850 & n17596 ) ;
  assign n17598 = ~n17595 & n17597 ;
  assign n17599 = n17594 | n17597 ;
  assign n17600 = ( ~x14 & n17598 ) | ( ~x14 & n17599 ) | ( n17598 & n17599 ) ;
  assign n17601 = n17585 | n17600 ;
  assign n17602 = ( n17585 & n17589 ) | ( n17585 & n17601 ) | ( n17589 & n17601 ) ;
  assign n17603 = n17539 | n17554 ;
  assign n17604 = ~n17555 & n17603 ;
  assign n17605 = n17555 | n17604 ;
  assign n17606 = ( n17555 & n17602 ) | ( n17555 & n17605 ) | ( n17602 & n17605 ) ;
  assign n17607 = n17535 & n17606 ;
  assign n17608 = n17533 | n17607 ;
  assign n17609 = n17511 & n17608 ;
  assign n17610 = n17508 | n17609 ;
  assign n17611 = ~n17475 & n17489 ;
  assign n17612 = ( n17475 & ~n17490 ) | ( n17475 & n17611 ) | ( ~n17490 & n17611 ) ;
  assign n17613 = n17490 | n17612 ;
  assign n17614 = ( n17490 & n17610 ) | ( n17490 & n17613 ) | ( n17610 & n17613 ) ;
  assign n17615 = n17472 & n17614 ;
  assign n17616 = n17469 | n17615 ;
  assign n17617 = n17452 & n17616 ;
  assign n17618 = n17449 | n17617 ;
  assign n17619 = n17415 | n17431 ;
  assign n17620 = ~n17432 & n17619 ;
  assign n17621 = n17432 | n17620 ;
  assign n17622 = ( n17432 & n17618 ) | ( n17432 & n17621 ) | ( n17618 & n17621 ) ;
  assign n17623 = n17396 | n17411 ;
  assign n17624 = ~n17412 & n17623 ;
  assign n17625 = n17412 | n17624 ;
  assign n17626 = ( n17412 & n17622 ) | ( n17412 & n17625 ) | ( n17622 & n17625 ) ;
  assign n17627 = ~n17376 & n17391 ;
  assign n17628 = n17626 & n17627 ;
  assign n17629 = ( n17393 & n17626 ) | ( n17393 & n17628 ) | ( n17626 & n17628 ) ;
  assign n17630 = n17392 | n17629 ;
  assign n17631 = ~n17358 & n17372 ;
  assign n17632 = ( n17358 & ~n17373 ) | ( n17358 & n17631 ) | ( ~n17373 & n17631 ) ;
  assign n17633 = n17373 | n17632 ;
  assign n17634 = ( n17373 & n17630 ) | ( n17373 & n17633 ) | ( n17630 & n17633 ) ;
  assign n17635 = n17355 & n17634 ;
  assign n17636 = n17352 | n17635 ;
  assign n17637 = n17292 & ~n17309 ;
  assign n17638 = ~n17292 & n17308 ;
  assign n17639 = n17637 | n17638 ;
  assign n17640 = n17636 & n17639 ;
  assign n17641 = n17329 | n17640 ;
  assign n17642 = ( n17332 & n17333 ) | ( n17332 & n17641 ) | ( n17333 & n17641 ) ;
  assign n17643 = n17286 | n17642 ;
  assign n17644 = ( n17286 & n17289 ) | ( n17286 & n17643 ) | ( n17289 & n17643 ) ;
  assign n17645 = ~n17251 & n17266 ;
  assign n17646 = ( n17251 & ~n17267 ) | ( n17251 & n17645 ) | ( ~n17267 & n17645 ) ;
  assign n17647 = n17267 | n17646 ;
  assign n17648 = ( n17267 & n17644 ) | ( n17267 & n17647 ) | ( n17644 & n17647 ) ;
  assign n17649 = n17245 | n17648 ;
  assign n17650 = ( n17245 & ~n17248 ) | ( n17245 & n17649 ) | ( ~n17248 & n17649 ) ;
  assign n17651 = ~n17225 & n17650 ;
  assign n17652 = n17222 | n17651 ;
  assign n17653 = n17202 | n17652 ;
  assign n17654 = ( n17202 & n17205 ) | ( n17202 & n17653 ) | ( n17205 & n17653 ) ;
  assign n17655 = n17177 | n17654 ;
  assign n17656 = ( n17177 & ~n17180 ) | ( n17177 & n17655 ) | ( ~n17180 & n17655 ) ;
  assign n17657 = ~n17154 & n17656 ;
  assign n17658 = n17151 | n17657 ;
  assign n17745 = ~n15088 & n15091 ;
  assign n17746 = ( n15088 & n15093 ) | ( n15088 & ~n17745 ) | ( n15093 & ~n17745 ) ;
  assign n17659 = n1057 & n10649 ;
  assign n17660 = n1065 & n10325 ;
  assign n17661 = n1060 & n10654 ;
  assign n17662 = n17660 | n17661 ;
  assign n17663 = n17659 | n17662 ;
  assign n17664 = n1062 | n17661 ;
  assign n17665 = n17660 | n17664 ;
  assign n17666 = n17659 | n17665 ;
  assign n17667 = ( n10702 & n17663 ) | ( n10702 & n17666 ) | ( n17663 & n17666 ) ;
  assign n17668 = n17663 | n17666 ;
  assign n17669 = ( n10695 & n17667 ) | ( n10695 & n17668 ) | ( n17667 & n17668 ) ;
  assign n17670 = n435 | n456 ;
  assign n17671 = n1615 | n17670 ;
  assign n17672 = n1692 | n17671 ;
  assign n17673 = n7917 | n10338 ;
  assign n17674 = n17672 | n17673 ;
  assign n17675 = n1418 | n17674 ;
  assign n17676 = n321 | n680 ;
  assign n17677 = n7931 | n17676 ;
  assign n17678 = n311 | n702 ;
  assign n17679 = n124 | n4249 ;
  assign n17680 = n17678 | n17679 ;
  assign n17681 = n527 | n887 ;
  assign n17682 = n17680 | n17681 ;
  assign n17683 = n17677 | n17682 ;
  assign n17684 = n17675 | n17683 ;
  assign n17685 = n443 | n17684 ;
  assign n17686 = n332 | n9120 ;
  assign n17687 = n1000 | n4182 ;
  assign n17688 = n179 | n295 ;
  assign n17689 = n465 | n568 ;
  assign n17690 = n17688 | n17689 ;
  assign n17691 = n17687 | n17690 ;
  assign n17692 = n17686 | n17691 ;
  assign n17693 = n390 | n437 ;
  assign n17694 = n12387 | n17693 ;
  assign n17695 = n207 | n449 ;
  assign n17696 = n17694 | n17695 ;
  assign n17697 = n779 | n857 ;
  assign n17698 = n839 | n17697 ;
  assign n17699 = n17696 | n17698 ;
  assign n17700 = n160 | n412 ;
  assign n17701 = n501 | n17700 ;
  assign n17702 = n17699 | n17701 ;
  assign n17703 = n17692 | n17702 ;
  assign n17704 = n235 | n7919 ;
  assign n17705 = n17703 | n17704 ;
  assign n17706 = n17685 | n17705 ;
  assign n17707 = n931 | n5123 ;
  assign n17708 = n190 | n720 ;
  assign n17709 = n223 | n17708 ;
  assign n17710 = n17707 | n17709 ;
  assign n17711 = n239 | n616 ;
  assign n17712 = n96 | n17711 ;
  assign n17713 = n3395 | n17712 ;
  assign n17714 = n5072 | n15243 ;
  assign n17715 = n17713 | n17714 ;
  assign n17716 = n17710 | n17715 ;
  assign n17717 = n330 | n387 ;
  assign n17718 = n3330 | n17717 ;
  assign n17719 = n269 | n644 ;
  assign n17720 = n155 | n17719 ;
  assign n17721 = n17718 | n17720 ;
  assign n17722 = n1176 | n17721 ;
  assign n17723 = n17716 | n17722 ;
  assign n17724 = n348 | n500 ;
  assign n17725 = n575 | n1380 ;
  assign n17726 = n282 | n17725 ;
  assign n17727 = n17724 | n17726 ;
  assign n17728 = n17723 | n17727 ;
  assign n17729 = n88 | n451 ;
  assign n17730 = n284 | n600 ;
  assign n17731 = n17729 | n17730 ;
  assign n17732 = n675 | n895 ;
  assign n17733 = n17731 | n17732 ;
  assign n17734 = n17728 | n17733 ;
  assign n17735 = n17706 | n17734 ;
  assign n17736 = n17659 & n17735 ;
  assign n17737 = ( n17665 & n17735 ) | ( n17665 & n17736 ) | ( n17735 & n17736 ) ;
  assign n17738 = ( n17662 & n17735 ) | ( n17662 & n17736 ) | ( n17735 & n17736 ) ;
  assign n17739 = ( n10702 & n17737 ) | ( n10702 & n17738 ) | ( n17737 & n17738 ) ;
  assign n17740 = n17737 | n17738 ;
  assign n17741 = ( n10695 & n17739 ) | ( n10695 & n17740 ) | ( n17739 & n17740 ) ;
  assign n17742 = n17669 & ~n17741 ;
  assign n17743 = ~n17669 & n17735 ;
  assign n17744 = n17742 | n17743 ;
  assign n17747 = n17744 & n17746 ;
  assign n17748 = n17746 & ~n17747 ;
  assign n17750 = n1826 & n11363 ;
  assign n17751 = n1823 & ~n11663 ;
  assign n17752 = n17750 | n17751 ;
  assign n17749 = n1829 & n12010 ;
  assign n17754 = n1821 | n17749 ;
  assign n17755 = n17752 | n17754 ;
  assign n17753 = n17749 | n17752 ;
  assign n17756 = n17753 & n17755 ;
  assign n17757 = ( ~n12028 & n17755 ) | ( ~n12028 & n17756 ) | ( n17755 & n17756 ) ;
  assign n17758 = n17755 | n17756 ;
  assign n17759 = ( n12017 & n17757 ) | ( n12017 & n17758 ) | ( n17757 & n17758 ) ;
  assign n17760 = ~x29 & n17759 ;
  assign n17761 = x29 | n17759 ;
  assign n17762 = ( ~n17759 & n17760 ) | ( ~n17759 & n17761 ) | ( n17760 & n17761 ) ;
  assign n17763 = n17744 & ~n17746 ;
  assign n17764 = n17762 & n17763 ;
  assign n17765 = ( n17748 & n17762 ) | ( n17748 & n17764 ) | ( n17762 & n17764 ) ;
  assign n17766 = n17762 | n17763 ;
  assign n17767 = n17748 | n17766 ;
  assign n17768 = ~n17765 & n17767 ;
  assign n17769 = n15097 & n17768 ;
  assign n17770 = ( n15103 & n17768 ) | ( n15103 & n17769 ) | ( n17768 & n17769 ) ;
  assign n17771 = n15097 | n17768 ;
  assign n17772 = n15103 | n17771 ;
  assign n17773 = ~n17770 & n17772 ;
  assign n17775 = n2312 & ~n12616 ;
  assign n17776 = n2308 & n12936 ;
  assign n17777 = n17775 | n17776 ;
  assign n17774 = n2315 & n13235 ;
  assign n17779 = n2306 | n17774 ;
  assign n17780 = n17777 | n17779 ;
  assign n17778 = n17774 | n17777 ;
  assign n17781 = n17778 & n17780 ;
  assign n17782 = ( n13561 & n17780 ) | ( n13561 & n17781 ) | ( n17780 & n17781 ) ;
  assign n17783 = x26 & n17781 ;
  assign n17784 = x26 & n17780 ;
  assign n17785 = ( n13561 & n17783 ) | ( n13561 & n17784 ) | ( n17783 & n17784 ) ;
  assign n17786 = x26 & ~n17783 ;
  assign n17787 = x26 & ~n17784 ;
  assign n17788 = ( ~n13561 & n17786 ) | ( ~n13561 & n17787 ) | ( n17786 & n17787 ) ;
  assign n17789 = ( n17782 & ~n17785 ) | ( n17782 & n17788 ) | ( ~n17785 & n17788 ) ;
  assign n17790 = n17773 & n17789 ;
  assign n17791 = n17773 & ~n17790 ;
  assign n17792 = ~n17773 & n17789 ;
  assign n17793 = n17791 | n17792 ;
  assign n17794 = ~n15121 & n15124 ;
  assign n17795 = ( n15121 & n15126 ) | ( n15121 & ~n17794 ) | ( n15126 & ~n17794 ) ;
  assign n17796 = n17793 & ~n17795 ;
  assign n17797 = ~n17793 & n17795 ;
  assign n17798 = n17796 | n17797 ;
  assign n17799 = n2932 & n14329 ;
  assign n17800 = n2925 & n13522 ;
  assign n17801 = n2928 & n14607 ;
  assign n17802 = n17800 | n17801 ;
  assign n17803 = n17799 | n17802 ;
  assign n17804 = n2936 | n17799 ;
  assign n17805 = n17802 | n17804 ;
  assign n17806 = ( n14656 & n17803 ) | ( n14656 & n17805 ) | ( n17803 & n17805 ) ;
  assign n17807 = x23 & n17805 ;
  assign n17808 = x23 & n17803 ;
  assign n17809 = ( n14656 & n17807 ) | ( n14656 & n17808 ) | ( n17807 & n17808 ) ;
  assign n17810 = x23 & ~n17808 ;
  assign n17811 = x23 & ~n17807 ;
  assign n17812 = ( ~n14656 & n17810 ) | ( ~n14656 & n17811 ) | ( n17810 & n17811 ) ;
  assign n17813 = ( n17806 & ~n17809 ) | ( n17806 & n17812 ) | ( ~n17809 & n17812 ) ;
  assign n17814 = n17798 & n17813 ;
  assign n17815 = n17798 | n17813 ;
  assign n17816 = ~n17814 & n17815 ;
  assign n17817 = ~n15144 & n15146 ;
  assign n17818 = ( n15144 & n15148 ) | ( n15144 & ~n17817 ) | ( n15148 & ~n17817 ) ;
  assign n17819 = n17816 & n17818 ;
  assign n17820 = n17816 | n17818 ;
  assign n17821 = ~n17819 & n17820 ;
  assign n17823 = n3544 & n14591 ;
  assign n17824 = n3541 & n15434 ;
  assign n17825 = n17823 | n17824 ;
  assign n17822 = n3547 & ~n16085 ;
  assign n17827 = n3537 | n17822 ;
  assign n17828 = n17825 | n17827 ;
  assign n17826 = n17822 | n17825 ;
  assign n17829 = n17826 & n17828 ;
  assign n17830 = ( ~n16167 & n17828 ) | ( ~n16167 & n17829 ) | ( n17828 & n17829 ) ;
  assign n17831 = ~x20 & n17829 ;
  assign n17832 = ~x20 & n17828 ;
  assign n17833 = ( ~n16167 & n17831 ) | ( ~n16167 & n17832 ) | ( n17831 & n17832 ) ;
  assign n17834 = x20 | n17831 ;
  assign n17835 = x20 | n17832 ;
  assign n17836 = ( ~n16167 & n17834 ) | ( ~n16167 & n17835 ) | ( n17834 & n17835 ) ;
  assign n17837 = ( ~n17830 & n17833 ) | ( ~n17830 & n17836 ) | ( n17833 & n17836 ) ;
  assign n17838 = n17821 & n17837 ;
  assign n17839 = n17821 & ~n17838 ;
  assign n17840 = ~n17821 & n17837 ;
  assign n17841 = n17839 | n17840 ;
  assign n17842 = ~n15470 & n15473 ;
  assign n17843 = ( n14999 & n15470 ) | ( n14999 & ~n17842 ) | ( n15470 & ~n17842 ) ;
  assign n17844 = n17841 & ~n17843 ;
  assign n17845 = ~n17841 & n17843 ;
  assign n17846 = n17844 | n17845 ;
  assign n17847 = n4471 & n17111 ;
  assign n17848 = n4466 & n15886 ;
  assign n17849 = n4468 & ~n16069 ;
  assign n17850 = n17848 | n17849 ;
  assign n17851 = n17847 | n17850 ;
  assign n17852 = n4475 & ~n17194 ;
  assign n17853 = ~n17129 & n17852 ;
  assign n17854 = n17851 | n17853 ;
  assign n17855 = n4475 | n17851 ;
  assign n17856 = ( n17186 & n17854 ) | ( n17186 & n17855 ) | ( n17854 & n17855 ) ;
  assign n17857 = x17 | n17856 ;
  assign n17858 = ~x17 & n17856 ;
  assign n17859 = ( ~n17856 & n17857 ) | ( ~n17856 & n17858 ) | ( n17857 & n17858 ) ;
  assign n17860 = n17846 & n17859 ;
  assign n17861 = n17846 | n17859 ;
  assign n17862 = ~n17860 & n17861 ;
  assign n17863 = n16123 & n17862 ;
  assign n17864 = ( n16567 & n17862 ) | ( n16567 & n17863 ) | ( n17862 & n17863 ) ;
  assign n17865 = n16123 | n17862 ;
  assign n17866 = n16567 | n17865 ;
  assign n17867 = ~n17864 & n17866 ;
  assign n17868 = n2932 & ~n8982 ;
  assign n17869 = ( n2932 & n9051 ) | ( n2932 & n17868 ) | ( n9051 & n17868 ) ;
  assign n17870 = n2928 & n9022 ;
  assign n17871 = n17869 | n17870 ;
  assign n17872 = n2928 | n17869 ;
  assign n17873 = ( ~n9019 & n17871 ) | ( ~n9019 & n17872 ) | ( n17871 & n17872 ) ;
  assign n17874 = n2925 | n17873 ;
  assign n17875 = ( ~n8017 & n17873 ) | ( ~n8017 & n17874 ) | ( n17873 & n17874 ) ;
  assign n17876 = n2936 | n17875 ;
  assign n17877 = ( ~n10242 & n17875 ) | ( ~n10242 & n17876 ) | ( n17875 & n17876 ) ;
  assign n17878 = ~x23 & n17876 ;
  assign n17879 = ~x23 & n17875 ;
  assign n17880 = ( ~n10242 & n17878 ) | ( ~n10242 & n17879 ) | ( n17878 & n17879 ) ;
  assign n17881 = x23 | n17878 ;
  assign n17882 = x23 | n17879 ;
  assign n17883 = ( ~n10242 & n17881 ) | ( ~n10242 & n17882 ) | ( n17881 & n17882 ) ;
  assign n17884 = ( ~n17877 & n17880 ) | ( ~n17877 & n17883 ) | ( n17880 & n17883 ) ;
  assign n17885 = n17016 | n17035 ;
  assign n17886 = ( n17016 & ~n17018 ) | ( n17016 & n17885 ) | ( ~n17018 & n17885 ) ;
  assign n17887 = n17884 & n17886 ;
  assign n17888 = n17884 | n17886 ;
  assign n17889 = ~n17887 & n17888 ;
  assign n17890 = n1739 | n6985 ;
  assign n17891 = n6835 | n17890 ;
  assign n17892 = n114 | n317 ;
  assign n17893 = n8983 | n17892 ;
  assign n17894 = n209 | n13343 ;
  assign n17895 = n17893 | n17894 ;
  assign n17896 = n64 | n666 ;
  assign n17897 = n133 | n269 ;
  assign n17898 = n17896 | n17897 ;
  assign n17899 = n155 | n349 ;
  assign n17900 = n104 | n676 ;
  assign n17901 = n17899 | n17900 ;
  assign n17902 = n17898 | n17901 ;
  assign n17903 = n17895 | n17902 ;
  assign n17904 = ( ~n497 & n17891 ) | ( ~n497 & n17903 ) | ( n17891 & n17903 ) ;
  assign n17905 = n17891 & n17903 ;
  assign n17906 = ( ~n10875 & n17904 ) | ( ~n10875 & n17905 ) | ( n17904 & n17905 ) ;
  assign n17907 = n10876 | n17906 ;
  assign n17908 = n314 | n888 ;
  assign n17909 = n10887 | n17908 ;
  assign n17910 = n278 | n616 ;
  assign n17911 = n212 | n273 ;
  assign n17912 = n17910 | n17911 ;
  assign n17913 = n229 | n17912 ;
  assign n17914 = n17909 | n17913 ;
  assign n17915 = n554 | n17694 ;
  assign n17916 = n697 | n7027 ;
  assign n17917 = n12274 | n17916 ;
  assign n17918 = n17915 | n17917 ;
  assign n17919 = n382 | n661 ;
  assign n17920 = n1349 | n1355 ;
  assign n17921 = n17919 | n17920 ;
  assign n17922 = n17918 | n17921 ;
  assign n17923 = n748 | n783 ;
  assign n17924 = n17710 | n17923 ;
  assign n17925 = n289 | n318 ;
  assign n17926 = n153 | n17925 ;
  assign n17927 = n341 | n477 ;
  assign n17928 = n17926 | n17927 ;
  assign n17929 = n17924 | n17928 ;
  assign n17930 = n17922 | n17929 ;
  assign n17931 = n17914 | n17930 ;
  assign n17932 = n259 | n2050 ;
  assign n17933 = n178 | n2192 ;
  assign n17934 = n17932 | n17933 ;
  assign n17935 = n333 | n443 ;
  assign n17936 = n500 | n17935 ;
  assign n17937 = n17934 | n17936 ;
  assign n17938 = n17931 | n17937 ;
  assign n17939 = n17907 | n17938 ;
  assign n17940 = ( ~x20 & n16810 ) | ( ~x20 & n17939 ) | ( n16810 & n17939 ) ;
  assign n17941 = n16810 | n17939 ;
  assign n17942 = ~n17940 & n17941 ;
  assign n17943 = n16810 & n17939 ;
  assign n17944 = n17941 & ~n17943 ;
  assign n17945 = x20 | n17944 ;
  assign n17946 = ~n17942 & n17945 ;
  assign n17947 = n16959 | n17946 ;
  assign n17948 = n16961 | n17946 ;
  assign n17949 = ( ~n6181 & n17947 ) | ( ~n6181 & n17948 ) | ( n17947 & n17948 ) ;
  assign n17950 = n16959 & n17946 ;
  assign n17951 = n16961 & n17946 ;
  assign n17952 = ( ~n6181 & n17950 ) | ( ~n6181 & n17951 ) | ( n17950 & n17951 ) ;
  assign n17953 = n17949 & ~n17952 ;
  assign n17954 = n1060 & n5108 ;
  assign n17955 = n1065 & n5997 ;
  assign n17956 = ( n1065 & n5979 ) | ( n1065 & n17955 ) | ( n5979 & n17955 ) ;
  assign n17957 = n17954 | n17956 ;
  assign n17958 = n1057 & n5857 ;
  assign n17959 = ( n1057 & ~n5899 ) | ( n1057 & n17958 ) | ( ~n5899 & n17958 ) ;
  assign n17960 = n17957 | n17959 ;
  assign n17961 = n1062 | n17960 ;
  assign n17962 = ( ~n6151 & n17960 ) | ( ~n6151 & n17961 ) | ( n17960 & n17961 ) ;
  assign n17963 = ~n17953 & n17962 ;
  assign n17964 = n17953 & ~n17962 ;
  assign n17965 = n17963 | n17964 ;
  assign n17966 = n1826 & ~n6091 ;
  assign n17967 = n1823 & n7036 ;
  assign n17968 = ( n1823 & n7023 ) | ( n1823 & n17967 ) | ( n7023 & n17967 ) ;
  assign n17969 = n17966 | n17968 ;
  assign n17970 = n1829 & n6950 ;
  assign n17971 = n17969 | n17970 ;
  assign n17972 = n1821 | n17971 ;
  assign n17973 = ( ~n7107 & n17971 ) | ( ~n7107 & n17972 ) | ( n17971 & n17972 ) ;
  assign n17974 = ~x29 & n17972 ;
  assign n17975 = ~x29 & n17971 ;
  assign n17976 = ( ~n7107 & n17974 ) | ( ~n7107 & n17975 ) | ( n17974 & n17975 ) ;
  assign n17977 = x29 | n17974 ;
  assign n17978 = x29 | n17975 ;
  assign n17979 = ( ~n7107 & n17977 ) | ( ~n7107 & n17978 ) | ( n17977 & n17978 ) ;
  assign n17980 = ( ~n17973 & n17976 ) | ( ~n17973 & n17979 ) | ( n17976 & n17979 ) ;
  assign n17981 = n17965 & n17980 ;
  assign n17982 = n17965 | n17980 ;
  assign n17983 = ~n17981 & n17982 ;
  assign n17984 = ~n16965 & n16968 ;
  assign n17985 = ( n16965 & n16970 ) | ( n16965 & ~n17984 ) | ( n16970 & ~n17984 ) ;
  assign n17986 = n17983 & n17985 ;
  assign n17987 = n17983 | n17985 ;
  assign n17988 = ~n17986 & n17987 ;
  assign n17989 = n2312 & n6889 ;
  assign n17990 = ( n2312 & ~n6884 ) | ( n2312 & n17989 ) | ( ~n6884 & n17989 ) ;
  assign n17991 = n2308 & n7907 ;
  assign n17992 = ( n2308 & n7902 ) | ( n2308 & n17991 ) | ( n7902 & n17991 ) ;
  assign n17993 = n2315 & n8079 ;
  assign n17994 = ( n2315 & ~n8070 ) | ( n2315 & n17993 ) | ( ~n8070 & n17993 ) ;
  assign n17995 = n17992 | n17994 ;
  assign n17996 = n17990 | n17995 ;
  assign n17997 = n2306 | n17996 ;
  assign n17998 = n17996 & n17997 ;
  assign n17999 = ( ~n8156 & n17997 ) | ( ~n8156 & n17998 ) | ( n17997 & n17998 ) ;
  assign n18000 = ~x26 & n17998 ;
  assign n18001 = ~x26 & n17997 ;
  assign n18002 = ( ~n8156 & n18000 ) | ( ~n8156 & n18001 ) | ( n18000 & n18001 ) ;
  assign n18003 = x26 | n18000 ;
  assign n18004 = x26 | n18001 ;
  assign n18005 = ( ~n8156 & n18003 ) | ( ~n8156 & n18004 ) | ( n18003 & n18004 ) ;
  assign n18006 = ( ~n17999 & n18002 ) | ( ~n17999 & n18005 ) | ( n18002 & n18005 ) ;
  assign n18007 = n17988 & n18006 ;
  assign n18008 = n17988 & ~n18007 ;
  assign n18009 = ~n17988 & n18006 ;
  assign n18010 = n18008 | n18009 ;
  assign n18011 = n16991 | n17010 ;
  assign n18012 = ( n16991 & ~n16993 ) | ( n16991 & n18011 ) | ( ~n16993 & n18011 ) ;
  assign n18013 = n18010 & n18012 ;
  assign n18014 = n18010 | n18012 ;
  assign n18015 = ~n18013 & n18014 ;
  assign n18016 = n17889 & ~n18015 ;
  assign n18017 = n17889 | n18015 ;
  assign n18018 = ( ~n17889 & n18016 ) | ( ~n17889 & n18017 ) | ( n18016 & n18017 ) ;
  assign n18019 = ~n16895 & n17038 ;
  assign n18020 = ( n16895 & n16897 ) | ( n16895 & ~n18019 ) | ( n16897 & ~n18019 ) ;
  assign n18021 = n18018 & n18020 ;
  assign n18022 = n18018 | n18020 ;
  assign n18023 = ~n18021 & n18022 ;
  assign n18024 = n17066 | n17078 ;
  assign n18025 = n17066 | n17084 ;
  assign n18026 = ( n17081 & n18024 ) | ( n17081 & n18025 ) | ( n18024 & n18025 ) ;
  assign n18027 = n18023 & n18026 ;
  assign n18028 = n18023 & n18024 ;
  assign n18029 = n17066 | n17079 ;
  assign n18030 = n18023 & n18029 ;
  assign n18031 = ( n16734 & n18028 ) | ( n16734 & n18030 ) | ( n18028 & n18030 ) ;
  assign n18032 = ( n15882 & n18027 ) | ( n15882 & n18031 ) | ( n18027 & n18031 ) ;
  assign n18033 = ( n16734 & n18024 ) | ( n16734 & n18029 ) | ( n18024 & n18029 ) ;
  assign n18034 = n18023 | n18033 ;
  assign n18035 = n18023 | n18026 ;
  assign n18036 = ( n15882 & n18034 ) | ( n15882 & n18035 ) | ( n18034 & n18035 ) ;
  assign n18037 = ~n18032 & n18036 ;
  assign n18038 = ~n17092 & n18037 ;
  assign n18039 = n17092 & ~n18037 ;
  assign n18040 = n18038 | n18039 ;
  assign n18041 = ~n17101 & n17103 ;
  assign n18042 = ( n17101 & n17117 ) | ( n17101 & ~n18041 ) | ( n17117 & ~n18041 ) ;
  assign n18043 = ~n18040 & n18042 ;
  assign n18044 = ( n17101 & n17119 ) | ( n17101 & ~n18041 ) | ( n17119 & ~n18041 ) ;
  assign n18045 = ~n18040 & n18044 ;
  assign n18046 = ( n17129 & n18043 ) | ( n17129 & n18045 ) | ( n18043 & n18045 ) ;
  assign n18047 = n18040 & ~n18044 ;
  assign n18048 = n18040 & ~n18042 ;
  assign n18049 = ( ~n17129 & n18047 ) | ( ~n17129 & n18048 ) | ( n18047 & n18048 ) ;
  assign n18050 = n18046 | n18049 ;
  assign n18052 = n5237 & n17100 ;
  assign n18053 = n5231 & ~n17092 ;
  assign n18054 = n18052 | n18053 ;
  assign n18051 = n5234 & n18037 ;
  assign n18056 = n5227 | n18051 ;
  assign n18057 = n18054 | n18056 ;
  assign n18055 = n18051 | n18054 ;
  assign n18058 = n18055 & n18057 ;
  assign n18059 = ( ~n18050 & n18057 ) | ( ~n18050 & n18058 ) | ( n18057 & n18058 ) ;
  assign n18060 = ~x14 & n18058 ;
  assign n18061 = ~x14 & n18057 ;
  assign n18062 = ( ~n18050 & n18060 ) | ( ~n18050 & n18061 ) | ( n18060 & n18061 ) ;
  assign n18063 = x14 | n18060 ;
  assign n18064 = x14 | n18061 ;
  assign n18065 = ( ~n18050 & n18063 ) | ( ~n18050 & n18064 ) | ( n18063 & n18064 ) ;
  assign n18066 = ( ~n18059 & n18062 ) | ( ~n18059 & n18065 ) | ( n18062 & n18065 ) ;
  assign n18067 = n17867 & n18066 ;
  assign n18068 = n17867 & ~n18067 ;
  assign n18069 = ~n17867 & n18066 ;
  assign n18070 = n18068 | n18069 ;
  assign n18071 = n17658 & n18070 ;
  assign n18072 = n17658 & ~n18071 ;
  assign n18073 = ~n17658 & n18070 ;
  assign n18074 = n18072 | n18073 ;
  assign n18075 = n18021 | n18028 ;
  assign n18076 = n18021 | n18030 ;
  assign n18077 = ( n16734 & n18075 ) | ( n16734 & n18076 ) | ( n18075 & n18076 ) ;
  assign n18078 = n17981 | n17986 ;
  assign n18079 = n1065 & n5857 ;
  assign n18080 = ( n1065 & ~n5899 ) | ( n1065 & n18079 ) | ( ~n5899 & n18079 ) ;
  assign n18081 = n1057 & ~n6091 ;
  assign n18082 = n1060 & n5997 ;
  assign n18083 = ( n1060 & n5979 ) | ( n1060 & n18082 ) | ( n5979 & n18082 ) ;
  assign n18084 = n18081 | n18083 ;
  assign n18085 = n18080 | n18084 ;
  assign n18086 = n1062 | n18085 ;
  assign n18087 = ( n6108 & n18085 ) | ( n6108 & n18086 ) | ( n18085 & n18086 ) ;
  assign n18088 = n661 | n13866 ;
  assign n18089 = n624 | n18088 ;
  assign n18090 = ~n1336 & n5878 ;
  assign n18091 = ~n5909 & n18090 ;
  assign n18092 = ~n18089 & n18091 ;
  assign n18093 = ~n995 & n18092 ;
  assign n18094 = ~n5150 & n18093 ;
  assign n18095 = ~n617 & n18094 ;
  assign n18096 = ~n1782 & n18095 ;
  assign n18097 = n94 | n820 ;
  assign n18098 = n5052 | n18097 ;
  assign n18099 = n142 | n18098 ;
  assign n18100 = n178 | n841 ;
  assign n18101 = n309 | n18100 ;
  assign n18102 = n477 | n676 ;
  assign n18103 = n4016 | n18102 ;
  assign n18104 = n18101 | n18103 ;
  assign n18105 = n7880 | n8052 ;
  assign n18106 = n1460 | n18105 ;
  assign n18107 = n18104 | n18106 ;
  assign n18108 = n4197 | n18107 ;
  assign n18109 = n901 | n991 ;
  assign n18110 = n993 | n18109 ;
  assign n18111 = n254 | n513 ;
  assign n18112 = n214 | n444 ;
  assign n18113 = n139 | n555 ;
  assign n18114 = n18112 | n18113 ;
  assign n18115 = n18111 | n18114 ;
  assign n18116 = n18110 | n18115 ;
  assign n18117 = n1030 | n1303 ;
  assign n18118 = n574 | n648 ;
  assign n18119 = n344 | n18118 ;
  assign n18120 = n18117 | n18119 ;
  assign n18121 = n18116 | n18120 ;
  assign n18122 = n18108 | n18121 ;
  assign n18123 = n237 | n667 ;
  assign n18124 = n281 | n18123 ;
  assign n18125 = n92 | n938 ;
  assign n18126 = n16797 | n18125 ;
  assign n18127 = n18124 | n18126 ;
  assign n18128 = n198 | n250 ;
  assign n18129 = n18127 | n18128 ;
  assign n18130 = n783 | n18129 ;
  assign n18131 = n18122 | n18130 ;
  assign n18132 = n18099 | n18131 ;
  assign n18133 = n18096 & ~n18132 ;
  assign n18134 = n17940 | n18133 ;
  assign n18135 = n17940 & n18133 ;
  assign n18136 = n18134 & ~n18135 ;
  assign n18137 = n18086 & n18136 ;
  assign n18138 = n18085 & n18136 ;
  assign n18139 = ( n6108 & n18137 ) | ( n6108 & n18138 ) | ( n18137 & n18138 ) ;
  assign n18140 = n18136 & ~n18138 ;
  assign n18141 = n18136 & ~n18137 ;
  assign n18142 = ( ~n6108 & n18140 ) | ( ~n6108 & n18141 ) | ( n18140 & n18141 ) ;
  assign n18143 = ( n18087 & ~n18139 ) | ( n18087 & n18142 ) | ( ~n18139 & n18142 ) ;
  assign n18144 = n17949 & ~n17962 ;
  assign n18145 = ( n17949 & ~n17953 ) | ( n17949 & n18144 ) | ( ~n17953 & n18144 ) ;
  assign n18146 = n18143 & ~n18145 ;
  assign n18147 = ~n18143 & n18145 ;
  assign n18148 = n18146 | n18147 ;
  assign n18149 = n1823 & n6950 ;
  assign n18150 = n1826 & n7036 ;
  assign n18151 = ( n1826 & n7023 ) | ( n1826 & n18150 ) | ( n7023 & n18150 ) ;
  assign n18152 = n18149 | n18151 ;
  assign n18153 = n1829 & n6889 ;
  assign n18154 = ( n1829 & ~n6884 ) | ( n1829 & n18153 ) | ( ~n6884 & n18153 ) ;
  assign n18156 = n1821 | n18154 ;
  assign n18157 = n18152 | n18156 ;
  assign n18155 = n18152 | n18154 ;
  assign n18158 = n18155 & n18157 ;
  assign n18159 = ( ~n7061 & n18157 ) | ( ~n7061 & n18158 ) | ( n18157 & n18158 ) ;
  assign n18160 = ~x29 & n18158 ;
  assign n18161 = ~x29 & n18157 ;
  assign n18162 = ( ~n7061 & n18160 ) | ( ~n7061 & n18161 ) | ( n18160 & n18161 ) ;
  assign n18163 = x29 | n18160 ;
  assign n18164 = x29 | n18161 ;
  assign n18165 = ( ~n7061 & n18163 ) | ( ~n7061 & n18164 ) | ( n18163 & n18164 ) ;
  assign n18166 = ( ~n18159 & n18162 ) | ( ~n18159 & n18165 ) | ( n18162 & n18165 ) ;
  assign n18167 = ~n18148 & n18166 ;
  assign n18168 = n18148 & ~n18166 ;
  assign n18169 = n18167 | n18168 ;
  assign n18170 = n18078 & ~n18169 ;
  assign n18171 = n18078 & ~n18170 ;
  assign n18172 = n2925 & ~n8982 ;
  assign n18173 = ( n2925 & n9051 ) | ( n2925 & n18172 ) | ( n9051 & n18172 ) ;
  assign n18174 = n2936 | n18173 ;
  assign n18175 = n9442 & ~n18173 ;
  assign n18176 = n9074 & ~n18173 ;
  assign n18177 = ( ~n9440 & n18175 ) | ( ~n9440 & n18176 ) | ( n18175 & n18176 ) ;
  assign n18178 = n18174 & ~n18177 ;
  assign n18179 = n18173 & n18174 ;
  assign n18180 = ( ~n9442 & n18174 ) | ( ~n9442 & n18179 ) | ( n18174 & n18179 ) ;
  assign n18181 = ( ~n9072 & n18178 ) | ( ~n9072 & n18180 ) | ( n18178 & n18180 ) ;
  assign n18182 = ~x23 & n18178 ;
  assign n18183 = ~x23 & n18180 ;
  assign n18184 = ( ~n9072 & n18182 ) | ( ~n9072 & n18183 ) | ( n18182 & n18183 ) ;
  assign n18185 = x23 | n18182 ;
  assign n18186 = x23 | n18183 ;
  assign n18187 = ( ~n9072 & n18185 ) | ( ~n9072 & n18186 ) | ( n18185 & n18186 ) ;
  assign n18188 = ( ~n18181 & n18184 ) | ( ~n18181 & n18187 ) | ( n18184 & n18187 ) ;
  assign n18189 = n2312 & n7907 ;
  assign n18190 = ( n2312 & n7902 ) | ( n2312 & n18189 ) | ( n7902 & n18189 ) ;
  assign n18191 = n2308 & n8079 ;
  assign n18192 = ( n2308 & ~n8070 ) | ( n2308 & n18191 ) | ( ~n8070 & n18191 ) ;
  assign n18193 = n18190 | n18192 ;
  assign n18194 = n2315 & ~n8017 ;
  assign n18195 = n18193 | n18194 ;
  assign n18196 = n2306 | n18193 ;
  assign n18197 = n18194 | n18196 ;
  assign n18198 = ( n8104 & n18195 ) | ( n8104 & n18197 ) | ( n18195 & n18197 ) ;
  assign n18199 = x26 & n18197 ;
  assign n18200 = x26 & n18195 ;
  assign n18201 = ( n8104 & n18199 ) | ( n8104 & n18200 ) | ( n18199 & n18200 ) ;
  assign n18202 = x26 & ~n18200 ;
  assign n18203 = x26 & ~n18199 ;
  assign n18204 = ( ~n8104 & n18202 ) | ( ~n8104 & n18203 ) | ( n18202 & n18203 ) ;
  assign n18205 = ( n18198 & ~n18201 ) | ( n18198 & n18204 ) | ( ~n18201 & n18204 ) ;
  assign n18206 = ~n18169 & n18205 ;
  assign n18207 = ~n18078 & n18206 ;
  assign n18208 = ~n18169 & n18188 ;
  assign n18209 = n18078 & n18208 ;
  assign n18210 = ( n18188 & n18207 ) | ( n18188 & n18209 ) | ( n18207 & n18209 ) ;
  assign n18211 = ( n18188 & n18205 ) | ( n18188 & n18209 ) | ( n18205 & n18209 ) ;
  assign n18212 = ( n18171 & n18210 ) | ( n18171 & n18211 ) | ( n18210 & n18211 ) ;
  assign n18213 = n18169 & ~n18188 ;
  assign n18214 = ( n18078 & n18188 ) | ( n18078 & ~n18213 ) | ( n18188 & ~n18213 ) ;
  assign n18215 = n18207 | n18214 ;
  assign n18216 = n18205 | n18214 ;
  assign n18217 = ( n18171 & n18215 ) | ( n18171 & n18216 ) | ( n18215 & n18216 ) ;
  assign n18218 = ~n18212 & n18217 ;
  assign n18302 = n18146 | n18166 ;
  assign n18303 = ( n18146 & ~n18148 ) | ( n18146 & n18302 ) | ( ~n18148 & n18302 ) ;
  assign n18219 = n18135 | n18137 ;
  assign n18220 = n18085 | n18135 ;
  assign n18221 = ( n18135 & n18136 ) | ( n18135 & n18220 ) | ( n18136 & n18220 ) ;
  assign n18222 = ( n6108 & n18219 ) | ( n6108 & n18221 ) | ( n18219 & n18221 ) ;
  assign n18223 = n13857 | n13917 ;
  assign n18224 = n13916 | n18223 ;
  assign n18225 = n13853 | n18224 ;
  assign n18226 = n461 | n574 ;
  assign n18227 = n6985 | n18226 ;
  assign n18228 = n67 | n477 ;
  assign n18229 = n388 | n18228 ;
  assign n18230 = n18227 | n18229 ;
  assign n18231 = n291 | n555 ;
  assign n18232 = n568 | n18231 ;
  assign n18233 = n18230 | n18232 ;
  assign n18234 = n599 | n18233 ;
  assign n18235 = n1725 | n18234 ;
  assign n18236 = n18225 | n18235 ;
  assign n18237 = n257 | n289 ;
  assign n18238 = n1301 | n18237 ;
  assign n18239 = n139 | n255 ;
  assign n18240 = n278 | n18239 ;
  assign n18241 = n18238 | n18240 ;
  assign n18242 = n395 | n18241 ;
  assign n18243 = n18236 | n18242 ;
  assign n18244 = n155 | n332 ;
  assign n18245 = n205 | n208 ;
  assign n18246 = n468 | n801 ;
  assign n18247 = n18245 | n18246 ;
  assign n18248 = n390 | n18247 ;
  assign n18249 = n55 | n12690 ;
  assign n18250 = n3313 | n18249 ;
  assign n18251 = n18248 | n18250 ;
  assign n18252 = n261 | n602 ;
  assign n18253 = n510 | n901 ;
  assign n18254 = n18252 | n18253 ;
  assign n18255 = n96 | n725 ;
  assign n18256 = n283 | n18255 ;
  assign n18257 = n18254 | n18256 ;
  assign n18258 = n2638 | n18257 ;
  assign n18259 = n18251 | n18258 ;
  assign n18260 = n18244 | n18259 ;
  assign n18261 = n235 | n4246 ;
  assign n18262 = n399 | n3431 ;
  assign n18263 = n18261 | n18262 ;
  assign n18264 = n88 | n412 ;
  assign n18265 = n456 | n18264 ;
  assign n18266 = n193 | n18265 ;
  assign n18267 = n18263 | n18266 ;
  assign n18268 = n434 | n18267 ;
  assign n18269 = n18260 | n18268 ;
  assign n18270 = n18243 | n18269 ;
  assign n18271 = n18133 & n18270 ;
  assign n18272 = n18133 | n18270 ;
  assign n18273 = n18135 & n18272 ;
  assign n18274 = ~n18271 & n18273 ;
  assign n18275 = ~n18271 & n18272 ;
  assign n18276 = ( n18137 & n18274 ) | ( n18137 & n18275 ) | ( n18274 & n18275 ) ;
  assign n18277 = n18221 & n18275 ;
  assign n18278 = ( n6108 & n18276 ) | ( n6108 & n18277 ) | ( n18276 & n18277 ) ;
  assign n18279 = n18222 & ~n18278 ;
  assign n18280 = n1057 & n7036 ;
  assign n18281 = ( n1057 & n7023 ) | ( n1057 & n18280 ) | ( n7023 & n18280 ) ;
  assign n18282 = n1060 & n5857 ;
  assign n18283 = ( n1060 & ~n5899 ) | ( n1060 & n18282 ) | ( ~n5899 & n18282 ) ;
  assign n18284 = n1065 & ~n6091 ;
  assign n18285 = n1062 | n18284 ;
  assign n18286 = n18283 | n18285 ;
  assign n18287 = n18281 | n18286 ;
  assign n18288 = n18283 | n18284 ;
  assign n18289 = n18281 | n18288 ;
  assign n18290 = ( n7136 & n18287 ) | ( n7136 & n18289 ) | ( n18287 & n18289 ) ;
  assign n18291 = n18272 & ~n18276 ;
  assign n18292 = ~n18271 & n18291 ;
  assign n18293 = n18272 & ~n18275 ;
  assign n18294 = ( ~n18221 & n18272 ) | ( ~n18221 & n18293 ) | ( n18272 & n18293 ) ;
  assign n18295 = ~n18271 & n18294 ;
  assign n18296 = ( ~n6108 & n18292 ) | ( ~n6108 & n18295 ) | ( n18292 & n18295 ) ;
  assign n18297 = n18290 & n18296 ;
  assign n18298 = ( n18279 & n18290 ) | ( n18279 & n18297 ) | ( n18290 & n18297 ) ;
  assign n18299 = n18290 | n18296 ;
  assign n18300 = n18279 | n18299 ;
  assign n18301 = ~n18298 & n18300 ;
  assign n18304 = n18301 & n18303 ;
  assign n18305 = n18303 & ~n18304 ;
  assign n18306 = n1826 & n6950 ;
  assign n18307 = n1823 & n6889 ;
  assign n18308 = ( n1823 & ~n6884 ) | ( n1823 & n18307 ) | ( ~n6884 & n18307 ) ;
  assign n18309 = n18306 | n18308 ;
  assign n18310 = n1829 & n7907 ;
  assign n18311 = ( n1829 & n7902 ) | ( n1829 & n18310 ) | ( n7902 & n18310 ) ;
  assign n18313 = n1821 | n18311 ;
  assign n18314 = n18309 | n18313 ;
  assign n18312 = n18309 | n18311 ;
  assign n18315 = n18312 & n18314 ;
  assign n18316 = ( ~n8193 & n18314 ) | ( ~n8193 & n18315 ) | ( n18314 & n18315 ) ;
  assign n18317 = ~x29 & n18315 ;
  assign n18318 = ~x29 & n18314 ;
  assign n18319 = ( ~n8193 & n18317 ) | ( ~n8193 & n18318 ) | ( n18317 & n18318 ) ;
  assign n18320 = x29 | n18317 ;
  assign n18321 = x29 | n18318 ;
  assign n18322 = ( ~n8193 & n18320 ) | ( ~n8193 & n18321 ) | ( n18320 & n18321 ) ;
  assign n18323 = ( ~n18316 & n18319 ) | ( ~n18316 & n18322 ) | ( n18319 & n18322 ) ;
  assign n18324 = n18301 & n18323 ;
  assign n18325 = ~n18303 & n18324 ;
  assign n18326 = ( n18305 & n18323 ) | ( n18305 & n18325 ) | ( n18323 & n18325 ) ;
  assign n18327 = n18301 | n18323 ;
  assign n18328 = ( ~n18303 & n18323 ) | ( ~n18303 & n18327 ) | ( n18323 & n18327 ) ;
  assign n18329 = n18305 | n18328 ;
  assign n18330 = ~n18326 & n18329 ;
  assign n18331 = n2312 & n8079 ;
  assign n18332 = ( n2312 & ~n8070 ) | ( n2312 & n18331 ) | ( ~n8070 & n18331 ) ;
  assign n18333 = n2308 | n18332 ;
  assign n18334 = ( ~n8017 & n18332 ) | ( ~n8017 & n18333 ) | ( n18332 & n18333 ) ;
  assign n18335 = n2315 & n9022 ;
  assign n18336 = ( n2315 & ~n9019 ) | ( n2315 & n18335 ) | ( ~n9019 & n18335 ) ;
  assign n18337 = n18334 | n18336 ;
  assign n18338 = n2306 | n18336 ;
  assign n18339 = n18334 | n18338 ;
  assign n18340 = ( ~n9416 & n18337 ) | ( ~n9416 & n18339 ) | ( n18337 & n18339 ) ;
  assign n18341 = ~x26 & n18339 ;
  assign n18342 = ~x26 & n18337 ;
  assign n18343 = ( ~n9416 & n18341 ) | ( ~n9416 & n18342 ) | ( n18341 & n18342 ) ;
  assign n18344 = x26 | n18342 ;
  assign n18345 = x26 | n18341 ;
  assign n18346 = ( ~n9416 & n18344 ) | ( ~n9416 & n18345 ) | ( n18344 & n18345 ) ;
  assign n18347 = ( ~n18340 & n18343 ) | ( ~n18340 & n18346 ) | ( n18343 & n18346 ) ;
  assign n18348 = n18330 & ~n18347 ;
  assign n18349 = n18330 | n18347 ;
  assign n18350 = ( ~n18330 & n18348 ) | ( ~n18330 & n18349 ) | ( n18348 & n18349 ) ;
  assign n18351 = n18218 & n18350 ;
  assign n18352 = n18350 & ~n18351 ;
  assign n18353 = ( n18218 & ~n18351 ) | ( n18218 & n18352 ) | ( ~n18351 & n18352 ) ;
  assign n18354 = ( n18171 & n18205 ) | ( n18171 & n18207 ) | ( n18205 & n18207 ) ;
  assign n18355 = n18169 & ~n18205 ;
  assign n18356 = ( n18078 & ~n18205 ) | ( n18078 & n18355 ) | ( ~n18205 & n18355 ) ;
  assign n18357 = ~n18171 & n18356 ;
  assign n18358 = n18354 | n18357 ;
  assign n18359 = n18007 | n18012 ;
  assign n18360 = ( n18007 & n18010 ) | ( n18007 & n18359 ) | ( n18010 & n18359 ) ;
  assign n18361 = ~n18358 & n18360 ;
  assign n18362 = n18358 & ~n18360 ;
  assign n18363 = n18361 | n18362 ;
  assign n18364 = n2928 & ~n8982 ;
  assign n18365 = ( n2928 & n9051 ) | ( n2928 & n18364 ) | ( n9051 & n18364 ) ;
  assign n18366 = n2925 & ~n9022 ;
  assign n18367 = ( n2925 & n18365 ) | ( n2925 & ~n18366 ) | ( n18365 & ~n18366 ) ;
  assign n18368 = n2925 | n18365 ;
  assign n18369 = ( ~n9019 & n18367 ) | ( ~n9019 & n18368 ) | ( n18367 & n18368 ) ;
  assign n18370 = n2936 | n18369 ;
  assign n18371 = ( n9078 & n18369 ) | ( n9078 & n18370 ) | ( n18369 & n18370 ) ;
  assign n18372 = x23 & n18370 ;
  assign n18373 = x23 & n18369 ;
  assign n18374 = ( n9078 & n18372 ) | ( n9078 & n18373 ) | ( n18372 & n18373 ) ;
  assign n18375 = x23 & ~n18372 ;
  assign n18376 = x23 & ~n18373 ;
  assign n18377 = ( ~n9078 & n18375 ) | ( ~n9078 & n18376 ) | ( n18375 & n18376 ) ;
  assign n18378 = ( n18371 & ~n18374 ) | ( n18371 & n18377 ) | ( ~n18374 & n18377 ) ;
  assign n18379 = n18361 | n18378 ;
  assign n18380 = ( n18361 & ~n18363 ) | ( n18361 & n18379 ) | ( ~n18363 & n18379 ) ;
  assign n18381 = n18353 & n18380 ;
  assign n18382 = n18353 | n18380 ;
  assign n18383 = ~n18381 & n18382 ;
  assign n18384 = ~n18363 & n18378 ;
  assign n18385 = n18363 & ~n18378 ;
  assign n18386 = n18384 | n18385 ;
  assign n18387 = n17887 | n18015 ;
  assign n18388 = ( n17887 & n17889 ) | ( n17887 & n18387 ) | ( n17889 & n18387 ) ;
  assign n18389 = ~n18386 & n18388 ;
  assign n18390 = n18386 & ~n18388 ;
  assign n18391 = n18389 | n18390 ;
  assign n18392 = ~n18389 & n18391 ;
  assign n18393 = n18383 & ~n18392 ;
  assign n18394 = n18383 & n18389 ;
  assign n18395 = ( n18077 & n18393 ) | ( n18077 & n18394 ) | ( n18393 & n18394 ) ;
  assign n18396 = n18021 | n18023 ;
  assign n18397 = ~n18391 & n18396 ;
  assign n18398 = n18389 | n18397 ;
  assign n18399 = n18383 & n18398 ;
  assign n18400 = n18021 & ~n18391 ;
  assign n18401 = n18389 | n18400 ;
  assign n18402 = n18383 & n18401 ;
  assign n18403 = ( n18026 & n18399 ) | ( n18026 & n18402 ) | ( n18399 & n18402 ) ;
  assign n18404 = ( n15882 & n18395 ) | ( n15882 & n18403 ) | ( n18395 & n18403 ) ;
  assign n18405 = ( n18077 & n18389 ) | ( n18077 & ~n18392 ) | ( n18389 & ~n18392 ) ;
  assign n18406 = n18383 | n18405 ;
  assign n18407 = ( n18026 & n18398 ) | ( n18026 & n18401 ) | ( n18398 & n18401 ) ;
  assign n18408 = n18383 | n18407 ;
  assign n18409 = ( n15882 & n18406 ) | ( n15882 & n18408 ) | ( n18406 & n18408 ) ;
  assign n18410 = ~n18404 & n18409 ;
  assign n18411 = n18212 | n18351 ;
  assign n18429 = n18326 | n18347 ;
  assign n18430 = ( n18326 & n18330 ) | ( n18326 & n18429 ) | ( n18330 & n18429 ) ;
  assign n18412 = n2315 & ~n8982 ;
  assign n18413 = ( n2315 & n9051 ) | ( n2315 & n18412 ) | ( n9051 & n18412 ) ;
  assign n18414 = n2308 & n9022 ;
  assign n18415 = n18413 | n18414 ;
  assign n18416 = n2308 | n18413 ;
  assign n18417 = ( ~n9019 & n18415 ) | ( ~n9019 & n18416 ) | ( n18415 & n18416 ) ;
  assign n18418 = n2312 | n18417 ;
  assign n18419 = ( ~n8017 & n18417 ) | ( ~n8017 & n18418 ) | ( n18417 & n18418 ) ;
  assign n18420 = n2306 | n18419 ;
  assign n18421 = ( ~n10242 & n18419 ) | ( ~n10242 & n18420 ) | ( n18419 & n18420 ) ;
  assign n18422 = ~x26 & n18420 ;
  assign n18423 = ~x26 & n18419 ;
  assign n18424 = ( ~n10242 & n18422 ) | ( ~n10242 & n18423 ) | ( n18422 & n18423 ) ;
  assign n18425 = x26 | n18422 ;
  assign n18426 = x26 | n18423 ;
  assign n18427 = ( ~n10242 & n18425 ) | ( ~n10242 & n18426 ) | ( n18425 & n18426 ) ;
  assign n18428 = ( ~n18421 & n18424 ) | ( ~n18421 & n18427 ) | ( n18424 & n18427 ) ;
  assign n18431 = n18428 & n18430 ;
  assign n18432 = n18430 & ~n18431 ;
  assign n18433 = ( ~n6108 & n18291 ) | ( ~n6108 & n18294 ) | ( n18291 & n18294 ) ;
  assign n18434 = n96 | n841 ;
  assign n18435 = n1678 | n18434 ;
  assign n18436 = n246 | n1172 ;
  assign n18437 = n959 | n18436 ;
  assign n18438 = n18435 | n18437 ;
  assign n18439 = n103 | n126 ;
  assign n18440 = n39 | n18439 ;
  assign n18441 = n18438 | n18440 ;
  assign n18442 = n4333 | n4334 ;
  assign n18443 = n3362 | n5011 ;
  assign n18444 = n18442 | n18443 ;
  assign n18445 = n71 | n364 ;
  assign n18446 = n448 | n487 ;
  assign n18447 = n18445 | n18446 ;
  assign n18448 = n412 | n441 ;
  assign n18449 = n416 | n432 ;
  assign n18450 = n18448 | n18449 ;
  assign n18451 = n312 | n568 ;
  assign n18452 = n18450 | n18451 ;
  assign n18453 = n18447 | n18452 ;
  assign n18454 = n18444 | n18453 ;
  assign n18455 = n18441 | n18454 ;
  assign n18456 = n3356 | n11101 ;
  assign n18457 = n320 | n434 ;
  assign n18458 = n1723 | n18457 ;
  assign n18459 = n801 | n3444 ;
  assign n18460 = n18458 | n18459 ;
  assign n18461 = n1030 | n4367 ;
  assign n18462 = n483 | n820 ;
  assign n18463 = n7928 | n18462 ;
  assign n18464 = n18461 | n18463 ;
  assign n18465 = n18460 | n18464 ;
  assign n18466 = n660 | n721 ;
  assign n18467 = n980 | n1013 ;
  assign n18468 = n18466 | n18467 ;
  assign n18469 = n264 | n938 ;
  assign n18470 = n18468 | n18469 ;
  assign n18471 = n18465 | n18470 ;
  assign n18472 = n18456 | n18471 ;
  assign n18473 = n18455 | n18472 ;
  assign n18474 = n357 | n1034 ;
  assign n18475 = n7834 | n18474 ;
  assign n18476 = n284 | n291 ;
  assign n18477 = n1631 | n18476 ;
  assign n18478 = n99 | n540 ;
  assign n18479 = n18477 | n18478 ;
  assign n18480 = n18475 | n18479 ;
  assign n18481 = n249 | n458 ;
  assign n18482 = n578 | n18481 ;
  assign n18483 = n203 | n18482 ;
  assign n18484 = n18480 | n18483 ;
  assign n18485 = n1505 | n1518 ;
  assign n18486 = n18484 | n18485 ;
  assign n18487 = n18473 | n18486 ;
  assign n18488 = n179 | n806 ;
  assign n18489 = n12387 | n18488 ;
  assign n18490 = n477 | n775 ;
  assign n18491 = n444 | n18490 ;
  assign n18492 = n18489 | n18491 ;
  assign n18493 = n75 | n2736 ;
  assign n18494 = n18492 | n18493 ;
  assign n18495 = n354 | n18494 ;
  assign n18496 = n18487 | n18495 ;
  assign n18497 = n18270 | n18496 ;
  assign n18498 = ( ~x23 & n18270 ) | ( ~x23 & n18496 ) | ( n18270 & n18496 ) ;
  assign n18499 = n18497 & ~n18498 ;
  assign n18500 = n18270 & n18496 ;
  assign n18501 = n18497 & ~n18500 ;
  assign n18502 = x23 | n18501 ;
  assign n18503 = ~n18499 & n18502 ;
  assign n18504 = n1057 & n6950 ;
  assign n18505 = n1060 & ~n6091 ;
  assign n18506 = n1065 & n7036 ;
  assign n18507 = ( n1065 & n7023 ) | ( n1065 & n18506 ) | ( n7023 & n18506 ) ;
  assign n18508 = n18505 | n18507 ;
  assign n18509 = n1062 | n18508 ;
  assign n18510 = n18504 | n18509 ;
  assign n18511 = ~n18503 & n18510 ;
  assign n18512 = n18504 | n18508 ;
  assign n18513 = ~n18503 & n18512 ;
  assign n18514 = ( ~n7107 & n18511 ) | ( ~n7107 & n18513 ) | ( n18511 & n18513 ) ;
  assign n18515 = n18503 & ~n18510 ;
  assign n18516 = n18503 & ~n18512 ;
  assign n18517 = ( n7107 & n18515 ) | ( n7107 & n18516 ) | ( n18515 & n18516 ) ;
  assign n18518 = n18514 | n18517 ;
  assign n18519 = n18433 | n18518 ;
  assign n18520 = n18433 & n18518 ;
  assign n18521 = n18519 & ~n18520 ;
  assign n18522 = n18298 | n18301 ;
  assign n18523 = n18521 & n18522 ;
  assign n18524 = n18298 & n18521 ;
  assign n18525 = ( n18303 & n18523 ) | ( n18303 & n18524 ) | ( n18523 & n18524 ) ;
  assign n18526 = n18521 | n18522 ;
  assign n18527 = n18298 | n18521 ;
  assign n18528 = ( n18303 & n18526 ) | ( n18303 & n18527 ) | ( n18526 & n18527 ) ;
  assign n18529 = ~n18525 & n18528 ;
  assign n18530 = n1826 & n6889 ;
  assign n18531 = ( n1826 & ~n6884 ) | ( n1826 & n18530 ) | ( ~n6884 & n18530 ) ;
  assign n18532 = n1823 & n7907 ;
  assign n18533 = ( n1823 & n7902 ) | ( n1823 & n18532 ) | ( n7902 & n18532 ) ;
  assign n18534 = n1829 & n8079 ;
  assign n18535 = ( n1829 & ~n8070 ) | ( n1829 & n18534 ) | ( ~n8070 & n18534 ) ;
  assign n18536 = n18533 | n18535 ;
  assign n18537 = n18531 | n18536 ;
  assign n18538 = n1821 | n18537 ;
  assign n18539 = ( ~n8156 & n18537 ) | ( ~n8156 & n18538 ) | ( n18537 & n18538 ) ;
  assign n18540 = ~x29 & n18538 ;
  assign n18541 = ~x29 & n18537 ;
  assign n18542 = ( ~n8156 & n18540 ) | ( ~n8156 & n18541 ) | ( n18540 & n18541 ) ;
  assign n18543 = x29 | n18540 ;
  assign n18544 = x29 | n18541 ;
  assign n18545 = ( ~n8156 & n18543 ) | ( ~n8156 & n18544 ) | ( n18543 & n18544 ) ;
  assign n18546 = ( ~n18539 & n18542 ) | ( ~n18539 & n18545 ) | ( n18542 & n18545 ) ;
  assign n18547 = n18529 & ~n18546 ;
  assign n18548 = n18529 | n18546 ;
  assign n18549 = ( ~n18529 & n18547 ) | ( ~n18529 & n18548 ) | ( n18547 & n18548 ) ;
  assign n18550 = n18428 & n18549 ;
  assign n18551 = ~n18430 & n18550 ;
  assign n18552 = ( n18432 & n18549 ) | ( n18432 & n18551 ) | ( n18549 & n18551 ) ;
  assign n18553 = n18428 | n18549 ;
  assign n18554 = ( ~n18430 & n18549 ) | ( ~n18430 & n18553 ) | ( n18549 & n18553 ) ;
  assign n18555 = n18432 | n18554 ;
  assign n18556 = ~n18552 & n18555 ;
  assign n18557 = n18411 & n18556 ;
  assign n18558 = n18411 | n18556 ;
  assign n18559 = ~n18557 & n18558 ;
  assign n18560 = n18381 | n18393 ;
  assign n18561 = n18559 & n18560 ;
  assign n18562 = n18381 | n18394 ;
  assign n18563 = n18559 & n18562 ;
  assign n18564 = ( n18077 & n18561 ) | ( n18077 & n18563 ) | ( n18561 & n18563 ) ;
  assign n18565 = n18381 | n18399 ;
  assign n18566 = n18559 & n18565 ;
  assign n18567 = n18381 | n18402 ;
  assign n18568 = n18559 & n18567 ;
  assign n18569 = ( n18026 & n18566 ) | ( n18026 & n18568 ) | ( n18566 & n18568 ) ;
  assign n18570 = ( n15882 & n18564 ) | ( n15882 & n18569 ) | ( n18564 & n18569 ) ;
  assign n18571 = ( n18077 & n18560 ) | ( n18077 & n18562 ) | ( n18560 & n18562 ) ;
  assign n18572 = n18559 | n18571 ;
  assign n18573 = ( n18026 & n18565 ) | ( n18026 & n18567 ) | ( n18565 & n18567 ) ;
  assign n18574 = n18559 | n18573 ;
  assign n18575 = ( n15882 & n18572 ) | ( n15882 & n18574 ) | ( n18572 & n18574 ) ;
  assign n18576 = ~n18570 & n18575 ;
  assign n18577 = n18410 & n18576 ;
  assign n18578 = n18077 & ~n18391 ;
  assign n18579 = ( n18026 & n18397 ) | ( n18026 & n18400 ) | ( n18397 & n18400 ) ;
  assign n18580 = ( n15882 & n18578 ) | ( n15882 & n18579 ) | ( n18578 & n18579 ) ;
  assign n18581 = ( n18021 & n18026 ) | ( n18021 & n18396 ) | ( n18026 & n18396 ) ;
  assign n18582 = n18391 & ~n18581 ;
  assign n18583 = ~n18077 & n18391 ;
  assign n18584 = ( ~n15882 & n18582 ) | ( ~n15882 & n18583 ) | ( n18582 & n18583 ) ;
  assign n18585 = n18580 | n18584 ;
  assign n18586 = ~n18410 & n18585 ;
  assign n18587 = n18037 & ~n18585 ;
  assign n18588 = ~n18586 & n18587 ;
  assign n18589 = n18410 | n18576 ;
  assign n18590 = n18410 & ~n18585 ;
  assign n18591 = n18589 & n18590 ;
  assign n18592 = ( n18588 & n18589 ) | ( n18588 & n18591 ) | ( n18589 & n18591 ) ;
  assign n18593 = ~n18577 & n18592 ;
  assign n18594 = n18038 | n18043 ;
  assign n18595 = ~n18037 & n18585 ;
  assign n18596 = n18587 | n18595 ;
  assign n18597 = ( n18586 & ~n18588 ) | ( n18586 & n18596 ) | ( ~n18588 & n18596 ) ;
  assign n18598 = ~n18577 & n18591 ;
  assign n18599 = ~n18577 & n18589 ;
  assign n18600 = ( ~n18597 & n18598 ) | ( ~n18597 & n18599 ) | ( n18598 & n18599 ) ;
  assign n18601 = ( n18593 & n18594 ) | ( n18593 & n18600 ) | ( n18594 & n18600 ) ;
  assign n18602 = n18038 | n18045 ;
  assign n18603 = ( n18593 & n18600 ) | ( n18593 & n18602 ) | ( n18600 & n18602 ) ;
  assign n18604 = ( n17129 & n18601 ) | ( n17129 & n18603 ) | ( n18601 & n18603 ) ;
  assign n18605 = ~n18590 & n18597 ;
  assign n18606 = n18588 | n18590 ;
  assign n18607 = ( n18594 & ~n18605 ) | ( n18594 & n18606 ) | ( ~n18605 & n18606 ) ;
  assign n18608 = ( n18602 & ~n18605 ) | ( n18602 & n18606 ) | ( ~n18605 & n18606 ) ;
  assign n18609 = ( n17129 & n18607 ) | ( n17129 & n18608 ) | ( n18607 & n18608 ) ;
  assign n18610 = ~n18604 & n18609 ;
  assign n18611 = n18599 & ~n18604 ;
  assign n18612 = n18610 | n18611 ;
  assign n18613 = n6122 & n18576 ;
  assign n18614 = n6125 & ~n18585 ;
  assign n18615 = n6119 & n18410 ;
  assign n18616 = n18614 | n18615 ;
  assign n18617 = n18613 | n18616 ;
  assign n18618 = n6115 | n18613 ;
  assign n18619 = n18616 | n18618 ;
  assign n18620 = ( n18612 & n18617 ) | ( n18612 & n18619 ) | ( n18617 & n18619 ) ;
  assign n18621 = x11 & n18619 ;
  assign n18622 = x11 & n18617 ;
  assign n18623 = ( n18612 & n18621 ) | ( n18612 & n18622 ) | ( n18621 & n18622 ) ;
  assign n18624 = x11 & ~n18622 ;
  assign n18625 = x11 & ~n18621 ;
  assign n18626 = ( ~n18612 & n18624 ) | ( ~n18612 & n18625 ) | ( n18624 & n18625 ) ;
  assign n18627 = ( n18620 & ~n18623 ) | ( n18620 & n18626 ) | ( ~n18623 & n18626 ) ;
  assign n18628 = n18073 & n18627 ;
  assign n18629 = ( n18072 & n18627 ) | ( n18072 & n18628 ) | ( n18627 & n18628 ) ;
  assign n18630 = n18074 & ~n18629 ;
  assign n18631 = ~n18073 & n18627 ;
  assign n18632 = ~n18072 & n18631 ;
  assign n18633 = n18630 | n18632 ;
  assign n18634 = n17154 & n17656 ;
  assign n18635 = n17154 | n17656 ;
  assign n18636 = ~n18634 & n18635 ;
  assign n18637 = n6122 & n18410 ;
  assign n18638 = n6125 & n18037 ;
  assign n18639 = n6119 & ~n18585 ;
  assign n18640 = n18638 | n18639 ;
  assign n18641 = n18637 | n18640 ;
  assign n18642 = n18594 & ~n18596 ;
  assign n18643 = ~n18596 & n18602 ;
  assign n18644 = ( n17129 & n18642 ) | ( n17129 & n18643 ) | ( n18642 & n18643 ) ;
  assign n18645 = n18590 | n18597 ;
  assign n18646 = n18588 & ~n18590 ;
  assign n18647 = ( n18594 & ~n18645 ) | ( n18594 & n18646 ) | ( ~n18645 & n18646 ) ;
  assign n18648 = ( n18602 & ~n18645 ) | ( n18602 & n18646 ) | ( ~n18645 & n18646 ) ;
  assign n18649 = ( n17129 & n18647 ) | ( n17129 & n18648 ) | ( n18647 & n18648 ) ;
  assign n18650 = ( n18587 & n18644 ) | ( n18587 & ~n18649 ) | ( n18644 & ~n18649 ) ;
  assign n18651 = n6115 & ~n18586 ;
  assign n18652 = ~n18609 & n18651 ;
  assign n18653 = ( n6115 & n18650 ) | ( n6115 & n18652 ) | ( n18650 & n18652 ) ;
  assign n18654 = n18641 | n18653 ;
  assign n18655 = x11 | n18641 ;
  assign n18656 = n18653 | n18655 ;
  assign n18657 = ~x11 & n18655 ;
  assign n18658 = ( ~x11 & n18653 ) | ( ~x11 & n18657 ) | ( n18653 & n18657 ) ;
  assign n18659 = ( ~n18654 & n18656 ) | ( ~n18654 & n18658 ) | ( n18656 & n18658 ) ;
  assign n18660 = ~n18636 & n18659 ;
  assign n18661 = n18636 & ~n18659 ;
  assign n18662 = n18660 | n18661 ;
  assign n18663 = n17180 & n17654 ;
  assign n18664 = n17180 | n17654 ;
  assign n18665 = ~n18663 & n18664 ;
  assign n18666 = n6122 & ~n18585 ;
  assign n18667 = n6125 & ~n17092 ;
  assign n18668 = n6119 & n18037 ;
  assign n18669 = n18667 | n18668 ;
  assign n18670 = n18666 | n18669 ;
  assign n18671 = ( n17129 & n18594 ) | ( n17129 & n18602 ) | ( n18594 & n18602 ) ;
  assign n18672 = ~n18644 & n18671 ;
  assign n18673 = n18594 | n18596 ;
  assign n18674 = n18596 | n18602 ;
  assign n18675 = ( n17129 & n18673 ) | ( n17129 & n18674 ) | ( n18673 & n18674 ) ;
  assign n18676 = n6115 & ~n18675 ;
  assign n18677 = ( n6115 & n18672 ) | ( n6115 & n18676 ) | ( n18672 & n18676 ) ;
  assign n18678 = n18670 | n18677 ;
  assign n18679 = x11 | n18670 ;
  assign n18680 = n18677 | n18679 ;
  assign n18681 = ~x11 & n18679 ;
  assign n18682 = ( ~x11 & n18677 ) | ( ~x11 & n18681 ) | ( n18677 & n18681 ) ;
  assign n18683 = ( ~n18678 & n18680 ) | ( ~n18678 & n18682 ) | ( n18680 & n18682 ) ;
  assign n18684 = ~n18665 & n18683 ;
  assign n18685 = n18665 & ~n18683 ;
  assign n18686 = n18684 | n18685 ;
  assign n18687 = ~n17205 & n17652 ;
  assign n18688 = n17205 & ~n17652 ;
  assign n18689 = n18687 | n18688 ;
  assign n18690 = n6122 & n18037 ;
  assign n18691 = n6125 & n17100 ;
  assign n18692 = n6119 & ~n17092 ;
  assign n18693 = n18691 | n18692 ;
  assign n18694 = n18690 | n18693 ;
  assign n18695 = n6115 | n18690 ;
  assign n18696 = n18693 | n18695 ;
  assign n18697 = ( ~n18050 & n18694 ) | ( ~n18050 & n18696 ) | ( n18694 & n18696 ) ;
  assign n18698 = ~x11 & n18696 ;
  assign n18699 = ~x11 & n18694 ;
  assign n18700 = ( ~n18050 & n18698 ) | ( ~n18050 & n18699 ) | ( n18698 & n18699 ) ;
  assign n18701 = x11 | n18699 ;
  assign n18702 = x11 | n18698 ;
  assign n18703 = ( ~n18050 & n18701 ) | ( ~n18050 & n18702 ) | ( n18701 & n18702 ) ;
  assign n18704 = ( ~n18697 & n18700 ) | ( ~n18697 & n18703 ) | ( n18700 & n18703 ) ;
  assign n18705 = n18689 & n18704 ;
  assign n18706 = n18689 | n18704 ;
  assign n18707 = ~n18705 & n18706 ;
  assign n18708 = n17225 & n17650 ;
  assign n18709 = n17225 | n17650 ;
  assign n18710 = ~n18708 & n18709 ;
  assign n18711 = n6122 & ~n17092 ;
  assign n18712 = n6125 & n17111 ;
  assign n18713 = n6119 & n17100 ;
  assign n18714 = n18712 | n18713 ;
  assign n18715 = n18711 | n18714 ;
  assign n18716 = n6115 | n18711 ;
  assign n18717 = n18714 | n18716 ;
  assign n18718 = ( ~n17134 & n18715 ) | ( ~n17134 & n18717 ) | ( n18715 & n18717 ) ;
  assign n18719 = ~x11 & n18717 ;
  assign n18720 = ~x11 & n18715 ;
  assign n18721 = ( ~n17134 & n18719 ) | ( ~n17134 & n18720 ) | ( n18719 & n18720 ) ;
  assign n18722 = x11 | n18720 ;
  assign n18723 = x11 | n18719 ;
  assign n18724 = ( ~n17134 & n18722 ) | ( ~n17134 & n18723 ) | ( n18722 & n18723 ) ;
  assign n18725 = ( ~n18718 & n18721 ) | ( ~n18718 & n18724 ) | ( n18721 & n18724 ) ;
  assign n18726 = ~n18710 & n18725 ;
  assign n18727 = n17248 & n17648 ;
  assign n18728 = n17248 | n17648 ;
  assign n18729 = ~n18727 & n18728 ;
  assign n18730 = n6122 & n17100 ;
  assign n18731 = n6125 & ~n16069 ;
  assign n18732 = n6119 & n17111 ;
  assign n18733 = n18731 | n18732 ;
  assign n18734 = n18730 | n18733 ;
  assign n18735 = n6115 & n17169 ;
  assign n18736 = ~n17129 & n18735 ;
  assign n18737 = n18734 | n18736 ;
  assign n18738 = n6115 | n18734 ;
  assign n18739 = ( n17161 & n18737 ) | ( n17161 & n18738 ) | ( n18737 & n18738 ) ;
  assign n18740 = x11 | n18739 ;
  assign n18741 = ~x11 & n18739 ;
  assign n18742 = ( ~n18739 & n18740 ) | ( ~n18739 & n18741 ) | ( n18740 & n18741 ) ;
  assign n18743 = ~n18729 & n18742 ;
  assign n18744 = n18729 & ~n18742 ;
  assign n18745 = n18743 | n18744 ;
  assign n18746 = n17644 & n17646 ;
  assign n18747 = n17644 | n17646 ;
  assign n18748 = ~n18746 & n18747 ;
  assign n18749 = n6125 & n15886 ;
  assign n18750 = n6119 & ~n16069 ;
  assign n18751 = n18749 | n18750 ;
  assign n18752 = n6122 & n17111 ;
  assign n18753 = n6115 | n18752 ;
  assign n18754 = n18751 | n18753 ;
  assign n18755 = n18751 | n18752 ;
  assign n18756 = n17194 & ~n18755 ;
  assign n18757 = ( n17129 & ~n18755 ) | ( n17129 & n18756 ) | ( ~n18755 & n18756 ) ;
  assign n18758 = n18754 & ~n18757 ;
  assign n18759 = ( n17186 & n18754 ) | ( n17186 & n18758 ) | ( n18754 & n18758 ) ;
  assign n18760 = x11 & n18759 ;
  assign n18761 = x11 & ~n18759 ;
  assign n18762 = ( n18759 & ~n18760 ) | ( n18759 & n18761 ) | ( ~n18760 & n18761 ) ;
  assign n18763 = n18748 & n18762 ;
  assign n18764 = n17289 & n17642 ;
  assign n18765 = n17289 | n17642 ;
  assign n18766 = ~n18764 & n18765 ;
  assign n18767 = n6122 & ~n16069 ;
  assign n18768 = n6125 & ~n16085 ;
  assign n18769 = n6119 & n15886 ;
  assign n18770 = n18768 | n18769 ;
  assign n18771 = n18767 | n18770 ;
  assign n18772 = n6115 | n18771 ;
  assign n18773 = ( ~n16107 & n18771 ) | ( ~n16107 & n18772 ) | ( n18771 & n18772 ) ;
  assign n18774 = ~x11 & n18772 ;
  assign n18775 = ~x11 & n18771 ;
  assign n18776 = ( ~n16107 & n18774 ) | ( ~n16107 & n18775 ) | ( n18774 & n18775 ) ;
  assign n18777 = x11 | n18774 ;
  assign n18778 = x11 | n18775 ;
  assign n18779 = ( ~n16107 & n18777 ) | ( ~n16107 & n18778 ) | ( n18777 & n18778 ) ;
  assign n18780 = ( ~n18773 & n18776 ) | ( ~n18773 & n18779 ) | ( n18776 & n18779 ) ;
  assign n18781 = n18766 & n18780 ;
  assign n18782 = n18766 & ~n18781 ;
  assign n18783 = ~n18766 & n18780 ;
  assign n18784 = n18782 | n18783 ;
  assign n18785 = ( n17331 & n17332 ) | ( n17331 & n17640 ) | ( n17332 & n17640 ) ;
  assign n18786 = n17309 | n17331 ;
  assign n18787 = n17640 | n18786 ;
  assign n18788 = ~n18785 & n18787 ;
  assign n18789 = n6122 & n15886 ;
  assign n18790 = n6125 & n15434 ;
  assign n18791 = n6119 & ~n16085 ;
  assign n18792 = n18790 | n18791 ;
  assign n18793 = n18789 | n18792 ;
  assign n18794 = n6115 | n18789 ;
  assign n18795 = n18792 | n18794 ;
  assign n18796 = ( ~n16140 & n18793 ) | ( ~n16140 & n18795 ) | ( n18793 & n18795 ) ;
  assign n18797 = ~x11 & n18795 ;
  assign n18798 = ~x11 & n18793 ;
  assign n18799 = ( ~n16140 & n18797 ) | ( ~n16140 & n18798 ) | ( n18797 & n18798 ) ;
  assign n18800 = x11 | n18798 ;
  assign n18801 = x11 | n18797 ;
  assign n18802 = ( ~n16140 & n18800 ) | ( ~n16140 & n18801 ) | ( n18800 & n18801 ) ;
  assign n18803 = ( ~n18796 & n18799 ) | ( ~n18796 & n18802 ) | ( n18799 & n18802 ) ;
  assign n18804 = n18788 & n18803 ;
  assign n18805 = n17636 & ~n17640 ;
  assign n18806 = n17639 & ~n17640 ;
  assign n18807 = n18805 | n18806 ;
  assign n18808 = n6122 & ~n16085 ;
  assign n18809 = n6125 & n14591 ;
  assign n18810 = n6119 & n15434 ;
  assign n18811 = n18809 | n18810 ;
  assign n18812 = n18808 | n18811 ;
  assign n18813 = n6115 | n18808 ;
  assign n18814 = n18811 | n18813 ;
  assign n18815 = ( ~n16167 & n18812 ) | ( ~n16167 & n18814 ) | ( n18812 & n18814 ) ;
  assign n18816 = ~x11 & n18814 ;
  assign n18817 = ~x11 & n18812 ;
  assign n18818 = ( ~n16167 & n18816 ) | ( ~n16167 & n18817 ) | ( n18816 & n18817 ) ;
  assign n18819 = x11 | n18817 ;
  assign n18820 = x11 | n18816 ;
  assign n18821 = ( ~n16167 & n18819 ) | ( ~n16167 & n18820 ) | ( n18819 & n18820 ) ;
  assign n18822 = ( ~n18815 & n18818 ) | ( ~n18815 & n18821 ) | ( n18818 & n18821 ) ;
  assign n18823 = n18807 & n18822 ;
  assign n18824 = n18807 & ~n18823 ;
  assign n18825 = ~n18807 & n18822 ;
  assign n18826 = n18824 | n18825 ;
  assign n18827 = n17634 & ~n17635 ;
  assign n18828 = n17355 & ~n17635 ;
  assign n18829 = n18827 | n18828 ;
  assign n18830 = n6122 & n15434 ;
  assign n18831 = n6125 & n14329 ;
  assign n18832 = n6119 & n14591 ;
  assign n18833 = n18831 | n18832 ;
  assign n18834 = n18830 | n18833 ;
  assign n18835 = n6115 | n18830 ;
  assign n18836 = n18833 | n18835 ;
  assign n18837 = ( n15453 & n18834 ) | ( n15453 & n18836 ) | ( n18834 & n18836 ) ;
  assign n18838 = x11 & n18836 ;
  assign n18839 = x11 & n18834 ;
  assign n18840 = ( n15453 & n18838 ) | ( n15453 & n18839 ) | ( n18838 & n18839 ) ;
  assign n18841 = x11 & ~n18839 ;
  assign n18842 = x11 & ~n18838 ;
  assign n18843 = ( ~n15453 & n18841 ) | ( ~n15453 & n18842 ) | ( n18841 & n18842 ) ;
  assign n18844 = ( n18837 & ~n18840 ) | ( n18837 & n18843 ) | ( ~n18840 & n18843 ) ;
  assign n18845 = n18829 & n18844 ;
  assign n18846 = n18829 & ~n18845 ;
  assign n18847 = ~n18829 & n18844 ;
  assign n18848 = n18846 | n18847 ;
  assign n18849 = n17626 | n17627 ;
  assign n18850 = n17393 | n18849 ;
  assign n18851 = ~n17629 & n18850 ;
  assign n18853 = n6125 & n13522 ;
  assign n18854 = n6119 & n14607 ;
  assign n18855 = n18853 | n18854 ;
  assign n18852 = n6122 & n14329 ;
  assign n18857 = n6115 | n18852 ;
  assign n18858 = n18855 | n18857 ;
  assign n18856 = n18852 | n18855 ;
  assign n18859 = n18856 & n18858 ;
  assign n18860 = ( n14656 & n18858 ) | ( n14656 & n18859 ) | ( n18858 & n18859 ) ;
  assign n18861 = x11 & n18859 ;
  assign n18862 = x11 & n18858 ;
  assign n18863 = ( n14656 & n18861 ) | ( n14656 & n18862 ) | ( n18861 & n18862 ) ;
  assign n18864 = x11 & ~n18861 ;
  assign n18865 = x11 & ~n18862 ;
  assign n18866 = ( ~n14656 & n18864 ) | ( ~n14656 & n18865 ) | ( n18864 & n18865 ) ;
  assign n18867 = ( n18860 & ~n18863 ) | ( n18860 & n18866 ) | ( ~n18863 & n18866 ) ;
  assign n18868 = n18851 & n18867 ;
  assign n18869 = n17630 & n17632 ;
  assign n18870 = n17630 | n17632 ;
  assign n18871 = ~n18869 & n18870 ;
  assign n18873 = n6125 & n14607 ;
  assign n18874 = n6119 & n14329 ;
  assign n18875 = n18873 | n18874 ;
  assign n18872 = n6122 & n14591 ;
  assign n18877 = n6115 | n18872 ;
  assign n18878 = n18875 | n18877 ;
  assign n18876 = n18872 | n18875 ;
  assign n18879 = n18876 & n18878 ;
  assign n18880 = ( n14629 & n18878 ) | ( n14629 & n18879 ) | ( n18878 & n18879 ) ;
  assign n18881 = x11 & n18879 ;
  assign n18882 = x11 & n18878 ;
  assign n18883 = ( n14629 & n18881 ) | ( n14629 & n18882 ) | ( n18881 & n18882 ) ;
  assign n18884 = x11 & ~n18881 ;
  assign n18885 = x11 & ~n18882 ;
  assign n18886 = ( ~n14629 & n18884 ) | ( ~n14629 & n18885 ) | ( n18884 & n18885 ) ;
  assign n18887 = ( n18880 & ~n18883 ) | ( n18880 & n18886 ) | ( ~n18883 & n18886 ) ;
  assign n18888 = n18871 & n18887 ;
  assign n18889 = n18871 | n18887 ;
  assign n18890 = ~n18888 & n18889 ;
  assign n18891 = n18868 & n18890 ;
  assign n18892 = n18888 | n18890 ;
  assign n18893 = n17622 & n17624 ;
  assign n18894 = n17622 | n17624 ;
  assign n18895 = ~n18893 & n18894 ;
  assign n18896 = n6125 & n13235 ;
  assign n18897 = n6119 & n13522 ;
  assign n18898 = n18896 | n18897 ;
  assign n18899 = n6122 & n14607 ;
  assign n18900 = n6115 | n18899 ;
  assign n18901 = n18898 | n18900 ;
  assign n18902 = n18898 | n18899 ;
  assign n18903 = n14696 | n18902 ;
  assign n18904 = n14698 | n18902 ;
  assign n18905 = ( ~n13248 & n18903 ) | ( ~n13248 & n18904 ) | ( n18903 & n18904 ) ;
  assign n18906 = n18901 & n18905 ;
  assign n18907 = ( n14687 & n18901 ) | ( n14687 & n18906 ) | ( n18901 & n18906 ) ;
  assign n18908 = ~x11 & n18907 ;
  assign n18909 = x11 | n18907 ;
  assign n18910 = ( ~n18907 & n18908 ) | ( ~n18907 & n18909 ) | ( n18908 & n18909 ) ;
  assign n18911 = n18895 & n18910 ;
  assign n18912 = n18895 & ~n18911 ;
  assign n18913 = ~n18895 & n18910 ;
  assign n18914 = n18912 | n18913 ;
  assign n18915 = n17618 & n17620 ;
  assign n18916 = n17618 | n17620 ;
  assign n18917 = ~n18915 & n18916 ;
  assign n18918 = n6122 & n13522 ;
  assign n18919 = n6125 & n12936 ;
  assign n18920 = n6119 & n13235 ;
  assign n18921 = n18919 | n18920 ;
  assign n18922 = n18918 | n18921 ;
  assign n18923 = n6115 & n13537 ;
  assign n18924 = n6115 & n13539 ;
  assign n18925 = ( ~n13248 & n18923 ) | ( ~n13248 & n18924 ) | ( n18923 & n18924 ) ;
  assign n18926 = n18922 | n18925 ;
  assign n18927 = n6115 | n18922 ;
  assign n18928 = ( n13530 & n18926 ) | ( n13530 & n18927 ) | ( n18926 & n18927 ) ;
  assign n18929 = x11 | n18928 ;
  assign n18930 = ~x11 & n18928 ;
  assign n18931 = ( ~n18928 & n18929 ) | ( ~n18928 & n18930 ) | ( n18929 & n18930 ) ;
  assign n18932 = n18917 & n18931 ;
  assign n18933 = n17616 & ~n17617 ;
  assign n18934 = n17452 & ~n17617 ;
  assign n18935 = n18933 | n18934 ;
  assign n18936 = n6122 & n13235 ;
  assign n18937 = n6125 & ~n12616 ;
  assign n18938 = n6119 & n12936 ;
  assign n18939 = n18937 | n18938 ;
  assign n18940 = n18936 | n18939 ;
  assign n18941 = n6115 | n18936 ;
  assign n18942 = n18939 | n18941 ;
  assign n18943 = ( n13561 & n18940 ) | ( n13561 & n18942 ) | ( n18940 & n18942 ) ;
  assign n18944 = x11 & n18942 ;
  assign n18945 = x11 & n18940 ;
  assign n18946 = ( n13561 & n18944 ) | ( n13561 & n18945 ) | ( n18944 & n18945 ) ;
  assign n18947 = x11 & ~n18945 ;
  assign n18948 = x11 & ~n18944 ;
  assign n18949 = ( ~n13561 & n18947 ) | ( ~n13561 & n18948 ) | ( n18947 & n18948 ) ;
  assign n18950 = ( n18943 & ~n18946 ) | ( n18943 & n18949 ) | ( ~n18946 & n18949 ) ;
  assign n18951 = n18935 & n18950 ;
  assign n18952 = n18935 & ~n18951 ;
  assign n18953 = ~n17472 & n17614 ;
  assign n18954 = n17472 & ~n17614 ;
  assign n18955 = n18953 | n18954 ;
  assign n18956 = n6122 & n12936 ;
  assign n18957 = n6125 & n12010 ;
  assign n18958 = n6119 & ~n12616 ;
  assign n18959 = n18957 | n18958 ;
  assign n18960 = n18956 | n18959 ;
  assign n18961 = n6115 | n18956 ;
  assign n18962 = n18959 | n18961 ;
  assign n18963 = ( ~n13591 & n18960 ) | ( ~n13591 & n18962 ) | ( n18960 & n18962 ) ;
  assign n18964 = ~x11 & n18962 ;
  assign n18965 = ~x11 & n18960 ;
  assign n18966 = ( ~n13591 & n18964 ) | ( ~n13591 & n18965 ) | ( n18964 & n18965 ) ;
  assign n18967 = x11 | n18965 ;
  assign n18968 = x11 | n18964 ;
  assign n18969 = ( ~n13591 & n18967 ) | ( ~n13591 & n18968 ) | ( n18967 & n18968 ) ;
  assign n18970 = ( ~n18963 & n18966 ) | ( ~n18963 & n18969 ) | ( n18966 & n18969 ) ;
  assign n18971 = n18955 & n18970 ;
  assign n18972 = n17610 & n17612 ;
  assign n18973 = n17610 | n17612 ;
  assign n18974 = ~n18972 & n18973 ;
  assign n18976 = n6125 & ~n11663 ;
  assign n18977 = n6119 & n12010 ;
  assign n18978 = n18976 | n18977 ;
  assign n18975 = n6122 & ~n12616 ;
  assign n18980 = n6115 | n18975 ;
  assign n18981 = n18978 | n18980 ;
  assign n18979 = n18975 | n18978 ;
  assign n18982 = n18979 & n18981 ;
  assign n18983 = ( ~n12626 & n18981 ) | ( ~n12626 & n18982 ) | ( n18981 & n18982 ) ;
  assign n18984 = ~x11 & n18982 ;
  assign n18985 = ~x11 & n18981 ;
  assign n18986 = ( ~n12626 & n18984 ) | ( ~n12626 & n18985 ) | ( n18984 & n18985 ) ;
  assign n18987 = x11 | n18984 ;
  assign n18988 = x11 | n18985 ;
  assign n18989 = ( ~n12626 & n18987 ) | ( ~n12626 & n18988 ) | ( n18987 & n18988 ) ;
  assign n18990 = ( ~n18983 & n18986 ) | ( ~n18983 & n18989 ) | ( n18986 & n18989 ) ;
  assign n18991 = n18974 & n18990 ;
  assign n18992 = n17511 | n17608 ;
  assign n18993 = ~n17609 & n18992 ;
  assign n18995 = n6125 & n11363 ;
  assign n18996 = n6119 & ~n11663 ;
  assign n18997 = n18995 | n18996 ;
  assign n18994 = n6122 & n12010 ;
  assign n18999 = n6115 | n18994 ;
  assign n19000 = n18997 | n18999 ;
  assign n18998 = n18994 | n18997 ;
  assign n19001 = n18998 & n19000 ;
  assign n19002 = ( ~n12028 & n19000 ) | ( ~n12028 & n19001 ) | ( n19000 & n19001 ) ;
  assign n19003 = n19000 | n19001 ;
  assign n19004 = ( n12017 & n19002 ) | ( n12017 & n19003 ) | ( n19002 & n19003 ) ;
  assign n19005 = ~x11 & n19004 ;
  assign n19006 = x11 | n19004 ;
  assign n19007 = ( ~n19004 & n19005 ) | ( ~n19004 & n19006 ) | ( n19005 & n19006 ) ;
  assign n19008 = n18993 & n19007 ;
  assign n19009 = n18993 & ~n19008 ;
  assign n19010 = ~n18993 & n19007 ;
  assign n19011 = n19009 | n19010 ;
  assign n19012 = n17535 | n17606 ;
  assign n19013 = ~n17607 & n19012 ;
  assign n19014 = n6125 & n10649 ;
  assign n19015 = n6119 & n11363 ;
  assign n19016 = n19014 | n19015 ;
  assign n19017 = n6122 & ~n11663 ;
  assign n19018 = n6115 | n19017 ;
  assign n19019 = n19016 | n19018 ;
  assign n19020 = n19016 | n19017 ;
  assign n19021 = n12048 & ~n19020 ;
  assign n19022 = ( n11672 & ~n19020 ) | ( n11672 & n19021 ) | ( ~n19020 & n19021 ) ;
  assign n19023 = n19019 & ~n19022 ;
  assign n19024 = ( n12040 & n19019 ) | ( n12040 & n19023 ) | ( n19019 & n19023 ) ;
  assign n19025 = x11 & n19024 ;
  assign n19026 = x11 & ~n19024 ;
  assign n19027 = ( n19024 & ~n19025 ) | ( n19024 & n19026 ) | ( ~n19025 & n19026 ) ;
  assign n19028 = n19013 & n19027 ;
  assign n19029 = n19013 & ~n19028 ;
  assign n19030 = ~n19013 & n19027 ;
  assign n19031 = n19029 | n19030 ;
  assign n19032 = n17602 & n17604 ;
  assign n19033 = n17602 | n17604 ;
  assign n19034 = ~n19032 & n19033 ;
  assign n19035 = n6122 & n11363 ;
  assign n19036 = n6125 & n10325 ;
  assign n19037 = n6119 & n10649 ;
  assign n19038 = n19036 | n19037 ;
  assign n19039 = n19035 | n19038 ;
  assign n19040 = n6115 | n19039 ;
  assign n19041 = ( n12059 & n19039 ) | ( n12059 & n19040 ) | ( n19039 & n19040 ) ;
  assign n19042 = x11 & n19040 ;
  assign n19043 = x11 & n19039 ;
  assign n19044 = ( n12059 & n19042 ) | ( n12059 & n19043 ) | ( n19042 & n19043 ) ;
  assign n19045 = x11 & ~n19042 ;
  assign n19046 = x11 & ~n19043 ;
  assign n19047 = ( ~n12059 & n19045 ) | ( ~n12059 & n19046 ) | ( n19045 & n19046 ) ;
  assign n19048 = ( n19041 & ~n19044 ) | ( n19041 & n19047 ) | ( ~n19044 & n19047 ) ;
  assign n19049 = n19034 & n19048 ;
  assign n19050 = n17589 & n17600 ;
  assign n19051 = n17589 & ~n19050 ;
  assign n19052 = n6122 & n10649 ;
  assign n19053 = n6125 & n10654 ;
  assign n19054 = n6119 & n10325 ;
  assign n19055 = n19053 | n19054 ;
  assign n19056 = n19052 | n19055 ;
  assign n19057 = n6115 | n19052 ;
  assign n19058 = n19055 | n19057 ;
  assign n19059 = ( n10702 & n19056 ) | ( n10702 & n19058 ) | ( n19056 & n19058 ) ;
  assign n19060 = n19056 | n19058 ;
  assign n19061 = ( n10695 & n19059 ) | ( n10695 & n19060 ) | ( n19059 & n19060 ) ;
  assign n19062 = x11 & n19061 ;
  assign n19063 = x11 & ~n19061 ;
  assign n19064 = ( n19061 & ~n19062 ) | ( n19061 & n19063 ) | ( ~n19062 & n19063 ) ;
  assign n19065 = ~n17589 & n17600 ;
  assign n19066 = n19064 & n19065 ;
  assign n19067 = ( n19051 & n19064 ) | ( n19051 & n19066 ) | ( n19064 & n19066 ) ;
  assign n19068 = n19064 | n19065 ;
  assign n19069 = n19051 | n19068 ;
  assign n19070 = ~n19067 & n19069 ;
  assign n19071 = n6122 & n10325 ;
  assign n19072 = n6125 & ~n10662 ;
  assign n19073 = n6119 & n10654 ;
  assign n19074 = n19072 | n19073 ;
  assign n19075 = n19071 | n19074 ;
  assign n19076 = n6115 | n19075 ;
  assign n19077 = ( ~n10957 & n19075 ) | ( ~n10957 & n19076 ) | ( n19075 & n19076 ) ;
  assign n19078 = n19075 | n19076 ;
  assign n19079 = ( n10949 & n19077 ) | ( n10949 & n19078 ) | ( n19077 & n19078 ) ;
  assign n19080 = ~x11 & n19079 ;
  assign n19081 = x11 & n19075 ;
  assign n19082 = x11 & n6115 ;
  assign n19083 = ( x11 & n19075 ) | ( x11 & n19082 ) | ( n19075 & n19082 ) ;
  assign n19084 = ( ~n10957 & n19081 ) | ( ~n10957 & n19083 ) | ( n19081 & n19083 ) ;
  assign n19085 = n19081 | n19083 ;
  assign n19086 = ( n10949 & n19084 ) | ( n10949 & n19085 ) | ( n19084 & n19085 ) ;
  assign n19087 = x11 & ~n19086 ;
  assign n19088 = n19080 | n19087 ;
  assign n19089 = n17568 & n17586 ;
  assign n19090 = n17568 | n17586 ;
  assign n19091 = ~n19089 & n19090 ;
  assign n19092 = n19088 & n19091 ;
  assign n19093 = n19088 | n19091 ;
  assign n19094 = ~n19092 & n19093 ;
  assign n19095 = n17561 | n17564 ;
  assign n19096 = ~n17564 & n17566 ;
  assign n19097 = ( n17562 & n19095 ) | ( n17562 & ~n19096 ) | ( n19095 & ~n19096 ) ;
  assign n19098 = ~n17568 & n19097 ;
  assign n19099 = n6122 & n10654 ;
  assign n19100 = n6125 & n10667 ;
  assign n19101 = n6119 & ~n10662 ;
  assign n19102 = n19100 | n19101 ;
  assign n19103 = n19099 | n19102 ;
  assign n19104 = n6115 | n19099 ;
  assign n19105 = n19102 | n19104 ;
  assign n19106 = ( n10978 & n19103 ) | ( n10978 & n19105 ) | ( n19103 & n19105 ) ;
  assign n19107 = x11 & n19105 ;
  assign n19108 = x11 & n19103 ;
  assign n19109 = ( n10978 & n19107 ) | ( n10978 & n19108 ) | ( n19107 & n19108 ) ;
  assign n19110 = x11 & ~n19108 ;
  assign n19111 = x11 & ~n19107 ;
  assign n19112 = ( ~n10978 & n19110 ) | ( ~n10978 & n19111 ) | ( n19110 & n19111 ) ;
  assign n19113 = ( n19106 & ~n19109 ) | ( n19106 & n19112 ) | ( ~n19109 & n19112 ) ;
  assign n19114 = n19098 & n19113 ;
  assign n19115 = n6115 & n10784 ;
  assign n19116 = n6119 & ~n10678 ;
  assign n19117 = n6122 & ~n10675 ;
  assign n19118 = n19116 | n19117 ;
  assign n19119 = x11 | n19118 ;
  assign n19120 = n19115 | n19119 ;
  assign n19121 = ~x11 & n19120 ;
  assign n19122 = x11 & ~n6114 ;
  assign n19123 = ( x11 & n10678 ) | ( x11 & n19122 ) | ( n10678 & n19122 ) ;
  assign n19124 = n19120 & n19123 ;
  assign n19125 = n19115 | n19118 ;
  assign n19126 = n19123 & ~n19125 ;
  assign n19127 = ( n19121 & n19124 ) | ( n19121 & n19126 ) | ( n19124 & n19126 ) ;
  assign n19128 = n6122 & n10667 ;
  assign n19129 = n6125 & ~n10678 ;
  assign n19130 = n6119 & ~n10675 ;
  assign n19131 = n19129 | n19130 ;
  assign n19132 = n19128 | n19131 ;
  assign n19133 = n10837 | n19132 ;
  assign n19134 = n6115 | n19128 ;
  assign n19135 = n19131 | n19134 ;
  assign n19136 = ~x11 & n19135 ;
  assign n19137 = n19133 & n19136 ;
  assign n19138 = x11 | n19137 ;
  assign n19139 = n5223 & ~n10678 ;
  assign n19140 = n19137 & n19139 ;
  assign n19141 = n19133 & n19135 ;
  assign n19142 = n19139 & ~n19141 ;
  assign n19143 = ( n19138 & n19140 ) | ( n19138 & n19142 ) | ( n19140 & n19142 ) ;
  assign n19144 = n19127 & n19143 ;
  assign n19145 = ( n19137 & n19138 ) | ( n19137 & ~n19141 ) | ( n19138 & ~n19141 ) ;
  assign n19146 = n19127 | n19139 ;
  assign n19147 = ( n19139 & n19145 ) | ( n19139 & n19146 ) | ( n19145 & n19146 ) ;
  assign n19148 = ~n19144 & n19147 ;
  assign n19149 = n6122 & ~n10662 ;
  assign n19150 = n6125 & ~n10675 ;
  assign n19151 = n6119 & n10667 ;
  assign n19152 = n19150 | n19151 ;
  assign n19153 = n19149 | n19152 ;
  assign n19154 = ( n6115 & n10850 ) | ( n6115 & n19153 ) | ( n10850 & n19153 ) ;
  assign n19155 = ( x11 & n6115 ) | ( x11 & ~n19153 ) | ( n6115 & ~n19153 ) ;
  assign n19156 = ( x11 & n10850 ) | ( x11 & n19155 ) | ( n10850 & n19155 ) ;
  assign n19157 = ~n19154 & n19156 ;
  assign n19158 = n19153 | n19156 ;
  assign n19159 = ( ~x11 & n19157 ) | ( ~x11 & n19158 ) | ( n19157 & n19158 ) ;
  assign n19160 = n19144 | n19159 ;
  assign n19161 = ( n19144 & n19148 ) | ( n19144 & n19160 ) | ( n19148 & n19160 ) ;
  assign n19162 = n19098 | n19113 ;
  assign n19163 = ~n19114 & n19162 ;
  assign n19164 = n19114 | n19163 ;
  assign n19165 = ( n19114 & n19161 ) | ( n19114 & n19164 ) | ( n19161 & n19164 ) ;
  assign n19166 = n19094 & n19165 ;
  assign n19167 = n19092 | n19166 ;
  assign n19168 = n19070 & n19167 ;
  assign n19169 = n19067 | n19168 ;
  assign n19170 = ~n19034 & n19048 ;
  assign n19171 = ( n19034 & ~n19049 ) | ( n19034 & n19170 ) | ( ~n19049 & n19170 ) ;
  assign n19172 = n19049 | n19171 ;
  assign n19173 = ( n19049 & n19169 ) | ( n19049 & n19172 ) | ( n19169 & n19172 ) ;
  assign n19174 = n19031 & n19173 ;
  assign n19175 = n19028 | n19174 ;
  assign n19176 = n19011 & n19175 ;
  assign n19177 = n19008 | n19176 ;
  assign n19178 = n18974 | n18990 ;
  assign n19179 = ~n18991 & n19178 ;
  assign n19180 = n18991 | n19179 ;
  assign n19181 = ( n18991 & n19177 ) | ( n18991 & n19180 ) | ( n19177 & n19180 ) ;
  assign n19182 = n18955 | n18970 ;
  assign n19183 = ~n18971 & n19182 ;
  assign n19184 = n18971 | n19183 ;
  assign n19185 = ( n18971 & n19181 ) | ( n18971 & n19184 ) | ( n19181 & n19184 ) ;
  assign n19186 = ~n18935 & n18950 ;
  assign n19187 = n19185 & n19186 ;
  assign n19188 = ( n18952 & n19185 ) | ( n18952 & n19187 ) | ( n19185 & n19187 ) ;
  assign n19189 = n18951 | n19188 ;
  assign n19190 = ~n18917 & n18931 ;
  assign n19191 = ( n18917 & ~n18932 ) | ( n18917 & n19190 ) | ( ~n18932 & n19190 ) ;
  assign n19192 = n18932 | n19191 ;
  assign n19193 = ( n18932 & n19189 ) | ( n18932 & n19192 ) | ( n19189 & n19192 ) ;
  assign n19194 = n18914 & n19193 ;
  assign n19195 = n18911 | n19194 ;
  assign n19196 = n18851 & ~n18868 ;
  assign n19197 = ~n18851 & n18867 ;
  assign n19198 = n19196 | n19197 ;
  assign n19199 = n19195 & n19198 ;
  assign n19200 = n18888 | n19199 ;
  assign n19201 = ( n18891 & n18892 ) | ( n18891 & n19200 ) | ( n18892 & n19200 ) ;
  assign n19202 = n18845 | n19201 ;
  assign n19203 = ( n18845 & n18848 ) | ( n18845 & n19202 ) | ( n18848 & n19202 ) ;
  assign n19204 = n18823 | n19203 ;
  assign n19205 = ( n18823 & n18826 ) | ( n18823 & n19204 ) | ( n18826 & n19204 ) ;
  assign n19206 = ~n18788 & n18803 ;
  assign n19207 = ( n18788 & ~n18804 ) | ( n18788 & n19206 ) | ( ~n18804 & n19206 ) ;
  assign n19208 = n18804 | n19207 ;
  assign n19209 = ( n18804 & n19205 ) | ( n18804 & n19208 ) | ( n19205 & n19208 ) ;
  assign n19210 = n18781 | n19209 ;
  assign n19211 = ( n18781 & n18784 ) | ( n18781 & n19210 ) | ( n18784 & n19210 ) ;
  assign n19212 = n18748 | n18762 ;
  assign n19213 = ~n18763 & n19212 ;
  assign n19214 = n18763 | n19213 ;
  assign n19215 = ( n18763 & n19211 ) | ( n18763 & n19214 ) | ( n19211 & n19214 ) ;
  assign n19216 = ~n18745 & n19215 ;
  assign n19217 = n18743 | n19216 ;
  assign n19218 = n18710 & ~n18725 ;
  assign n19219 = n18726 | n19218 ;
  assign n19220 = ~n18726 & n19219 ;
  assign n19221 = ( n18726 & n19217 ) | ( n18726 & ~n19220 ) | ( n19217 & ~n19220 ) ;
  assign n19222 = n18705 | n19221 ;
  assign n19223 = ( n18705 & n18707 ) | ( n18705 & n19222 ) | ( n18707 & n19222 ) ;
  assign n19224 = n18684 | n19223 ;
  assign n19225 = ( n18684 & ~n18686 ) | ( n18684 & n19224 ) | ( ~n18686 & n19224 ) ;
  assign n19226 = ~n18662 & n19225 ;
  assign n19227 = n18660 | n19226 ;
  assign n19228 = n18633 & n19227 ;
  assign n19229 = n18633 | n19227 ;
  assign n19230 = ~n19228 & n19229 ;
  assign n19304 = n18525 | n18546 ;
  assign n19305 = ( n18525 & n18529 ) | ( n18525 & n19304 ) | ( n18529 & n19304 ) ;
  assign n19231 = n1065 & n6950 ;
  assign n19232 = n1060 & n7036 ;
  assign n19233 = ( n1060 & n7023 ) | ( n1060 & n19232 ) | ( n7023 & n19232 ) ;
  assign n19234 = n19231 | n19233 ;
  assign n19235 = n1057 & n6889 ;
  assign n19236 = ( n1057 & ~n6884 ) | ( n1057 & n19235 ) | ( ~n6884 & n19235 ) ;
  assign n19237 = n19234 | n19236 ;
  assign n19238 = n1062 | n19236 ;
  assign n19239 = n19234 | n19238 ;
  assign n19240 = ( ~n7061 & n19237 ) | ( ~n7061 & n19239 ) | ( n19237 & n19239 ) ;
  assign n19241 = n324 | n3337 ;
  assign n19242 = n11753 | n11758 ;
  assign n19243 = n280 | n17688 ;
  assign n19244 = n436 | n1136 ;
  assign n19245 = ( ~n11091 & n19243 ) | ( ~n11091 & n19244 ) | ( n19243 & n19244 ) ;
  assign n19246 = n11091 | n11763 ;
  assign n19247 = n19245 | n19246 ;
  assign n19248 = n19242 | n19247 ;
  assign n19249 = n204 | n19248 ;
  assign n19250 = n19241 | n19249 ;
  assign n19251 = n399 | n483 ;
  assign n19252 = n590 | n638 ;
  assign n19253 = n19251 | n19252 ;
  assign n19254 = n79 | n560 ;
  assign n19255 = n199 | n19254 ;
  assign n19256 = n19253 | n19255 ;
  assign n19257 = n680 | n1028 ;
  assign n19258 = n2050 | n19257 ;
  assign n19259 = n19256 | n19258 ;
  assign n19260 = n442 | n10379 ;
  assign n19261 = n1251 | n19260 ;
  assign n19262 = n53 | n19261 ;
  assign n19263 = n19259 | n19262 ;
  assign n19264 = n689 | n758 ;
  assign n19265 = n8001 | n19264 ;
  assign n19266 = n19263 | n19265 ;
  assign n19267 = n19250 | n19266 ;
  assign n19268 = n18498 & ~n19267 ;
  assign n19269 = ~n18498 & n19267 ;
  assign n19270 = n19268 | n19269 ;
  assign n19271 = n19239 & n19270 ;
  assign n19272 = n19237 & n19270 ;
  assign n19273 = ( ~n7061 & n19271 ) | ( ~n7061 & n19272 ) | ( n19271 & n19272 ) ;
  assign n19274 = n19270 & ~n19272 ;
  assign n19275 = n19270 & ~n19271 ;
  assign n19276 = ( n7061 & n19274 ) | ( n7061 & n19275 ) | ( n19274 & n19275 ) ;
  assign n19277 = ( n19240 & ~n19273 ) | ( n19240 & n19276 ) | ( ~n19273 & n19276 ) ;
  assign n19278 = n18433 & ~n18514 ;
  assign n19279 = ( ~n18514 & n18518 ) | ( ~n18514 & n19278 ) | ( n18518 & n19278 ) ;
  assign n19280 = n19277 | n19279 ;
  assign n19281 = n19277 & n19279 ;
  assign n19282 = n19280 & ~n19281 ;
  assign n19288 = n1829 & ~n8017 ;
  assign n19283 = n1826 & n7907 ;
  assign n19284 = ( n1826 & n7902 ) | ( n1826 & n19283 ) | ( n7902 & n19283 ) ;
  assign n19285 = n1823 & n8079 ;
  assign n19286 = ( n1823 & ~n8070 ) | ( n1823 & n19285 ) | ( ~n8070 & n19285 ) ;
  assign n19287 = n19284 | n19286 ;
  assign n19290 = n1821 | n19287 ;
  assign n19291 = n19288 | n19290 ;
  assign n19289 = n19287 | n19288 ;
  assign n19292 = n19289 & n19291 ;
  assign n19293 = ( n8104 & n19291 ) | ( n8104 & n19292 ) | ( n19291 & n19292 ) ;
  assign n19294 = x29 & n19292 ;
  assign n19295 = x29 & n19291 ;
  assign n19296 = ( n8104 & n19294 ) | ( n8104 & n19295 ) | ( n19294 & n19295 ) ;
  assign n19297 = x29 & ~n19294 ;
  assign n19298 = x29 & ~n19295 ;
  assign n19299 = ( ~n8104 & n19297 ) | ( ~n8104 & n19298 ) | ( n19297 & n19298 ) ;
  assign n19300 = ( n19293 & ~n19296 ) | ( n19293 & n19299 ) | ( ~n19296 & n19299 ) ;
  assign n19301 = n19282 & n19300 ;
  assign n19302 = n19282 | n19300 ;
  assign n19303 = ~n19301 & n19302 ;
  assign n19306 = n19303 & n19305 ;
  assign n19307 = n19305 & ~n19306 ;
  assign n19308 = n2308 & ~n8982 ;
  assign n19309 = ( n2308 & n9051 ) | ( n2308 & n19308 ) | ( n9051 & n19308 ) ;
  assign n19310 = n2312 & ~n9022 ;
  assign n19311 = ( n2312 & n19309 ) | ( n2312 & ~n19310 ) | ( n19309 & ~n19310 ) ;
  assign n19312 = n2312 | n19309 ;
  assign n19313 = ( ~n9019 & n19311 ) | ( ~n9019 & n19312 ) | ( n19311 & n19312 ) ;
  assign n19314 = n2306 | n19313 ;
  assign n19315 = ( n9078 & n19313 ) | ( n9078 & n19314 ) | ( n19313 & n19314 ) ;
  assign n19316 = x26 & n19314 ;
  assign n19317 = x26 & n19313 ;
  assign n19318 = ( n9078 & n19316 ) | ( n9078 & n19317 ) | ( n19316 & n19317 ) ;
  assign n19319 = x26 & ~n19316 ;
  assign n19320 = x26 & ~n19317 ;
  assign n19321 = ( ~n9078 & n19319 ) | ( ~n9078 & n19320 ) | ( n19319 & n19320 ) ;
  assign n19322 = ( n19315 & ~n19318 ) | ( n19315 & n19321 ) | ( ~n19318 & n19321 ) ;
  assign n19323 = n19303 & n19322 ;
  assign n19324 = ~n19305 & n19323 ;
  assign n19325 = ( n19307 & n19322 ) | ( n19307 & n19324 ) | ( n19322 & n19324 ) ;
  assign n19326 = n19303 | n19322 ;
  assign n19327 = ( ~n19305 & n19322 ) | ( ~n19305 & n19326 ) | ( n19322 & n19326 ) ;
  assign n19328 = n19307 | n19327 ;
  assign n19329 = ~n19325 & n19328 ;
  assign n19330 = n18431 | n18551 ;
  assign n19331 = n18431 | n18549 ;
  assign n19332 = ( n18432 & n19330 ) | ( n18432 & n19331 ) | ( n19330 & n19331 ) ;
  assign n19333 = n19329 & n19332 ;
  assign n19334 = n19329 | n19332 ;
  assign n19335 = ~n19333 & n19334 ;
  assign n19336 = n18557 | n18561 ;
  assign n19337 = n19335 & n19336 ;
  assign n19338 = n18557 | n18563 ;
  assign n19339 = n19335 & n19338 ;
  assign n19340 = ( n18077 & n19337 ) | ( n18077 & n19339 ) | ( n19337 & n19339 ) ;
  assign n19341 = n18557 | n18566 ;
  assign n19342 = n19335 & n19341 ;
  assign n19343 = n18557 | n18568 ;
  assign n19344 = n19335 & n19343 ;
  assign n19345 = ( n18026 & n19342 ) | ( n18026 & n19344 ) | ( n19342 & n19344 ) ;
  assign n19346 = ( n15882 & n19340 ) | ( n15882 & n19345 ) | ( n19340 & n19345 ) ;
  assign n19347 = ( n18077 & n19336 ) | ( n18077 & n19338 ) | ( n19336 & n19338 ) ;
  assign n19348 = n19335 | n19347 ;
  assign n19349 = ( n18026 & n19341 ) | ( n18026 & n19343 ) | ( n19341 & n19343 ) ;
  assign n19350 = n19335 | n19349 ;
  assign n19351 = ( n15882 & n19348 ) | ( n15882 & n19350 ) | ( n19348 & n19350 ) ;
  assign n19352 = ~n19346 & n19351 ;
  assign n19353 = n1060 & n6950 ;
  assign n19354 = n1065 & n6889 ;
  assign n19355 = ( n1065 & ~n6884 ) | ( n1065 & n19354 ) | ( ~n6884 & n19354 ) ;
  assign n19356 = n19353 | n19355 ;
  assign n19357 = n1057 & n7907 ;
  assign n19358 = ( n1057 & n7902 ) | ( n1057 & n19357 ) | ( n7902 & n19357 ) ;
  assign n19359 = n19356 | n19358 ;
  assign n19360 = n1062 | n19358 ;
  assign n19361 = n19356 | n19360 ;
  assign n19362 = ( ~n8193 & n19359 ) | ( ~n8193 & n19361 ) | ( n19359 & n19361 ) ;
  assign n19363 = n126 | n212 ;
  assign n19364 = n5982 | n19363 ;
  assign n19365 = n354 | n19364 ;
  assign n19366 = n163 | n213 ;
  assign n19367 = n283 | n19366 ;
  assign n19368 = n8971 | n10344 ;
  assign n19369 = n19367 | n19368 ;
  assign n19370 = n19365 | n19369 ;
  assign n19371 = n15198 | n15201 ;
  assign n19372 = n3311 | n15030 ;
  assign n19373 = n292 | n648 ;
  assign n19374 = n67 | n88 ;
  assign n19375 = n19373 | n19374 ;
  assign n19376 = n312 | n886 ;
  assign n19377 = n19375 | n19376 ;
  assign n19378 = n19372 | n19377 ;
  assign n19379 = n19371 | n19378 ;
  assign n19380 = ( n282 & n318 ) | ( n282 & ~n10369 ) | ( n318 & ~n10369 ) ;
  assign n19381 = n249 | n10369 ;
  assign n19382 = n19380 | n19381 ;
  assign n19383 = n355 | n720 ;
  assign n19384 = n19382 | n19383 ;
  assign n19385 = n15070 | n19384 ;
  assign n19386 = n19379 | n19385 ;
  assign n19387 = n19370 | n19386 ;
  assign n19388 = n77 | n607 ;
  assign n19389 = n10732 | n19388 ;
  assign n19390 = n578 | n680 ;
  assign n19391 = n19389 | n19390 ;
  assign n19392 = n938 | n19391 ;
  assign n19393 = n5049 | n19392 ;
  assign n19394 = n5045 | n19393 ;
  assign n19395 = n39 | n190 ;
  assign n19396 = ( n566 & ~n2220 ) | ( n566 & n19395 ) | ( ~n2220 & n19395 ) ;
  assign n19397 = n182 | n2220 ;
  assign n19398 = n19396 | n19397 ;
  assign n19399 = n3376 | n19398 ;
  assign n19400 = n19394 | n19399 ;
  assign n19401 = n502 | n679 ;
  assign n19402 = n117 | n4249 ;
  assign n19403 = n19401 | n19402 ;
  assign n19404 = n309 | n434 ;
  assign n19405 = n437 | n19404 ;
  assign n19406 = n19403 | n19405 ;
  assign n19407 = n19400 | n19406 ;
  assign n19408 = n19387 | n19407 ;
  assign n19409 = n19267 & ~n19408 ;
  assign n19410 = ~n19267 & n19408 ;
  assign n19411 = n19409 | n19410 ;
  assign n19412 = n19361 & ~n19411 ;
  assign n19413 = n19359 & ~n19411 ;
  assign n19414 = ( ~n8193 & n19412 ) | ( ~n8193 & n19413 ) | ( n19412 & n19413 ) ;
  assign n19415 = n19362 & ~n19414 ;
  assign n19416 = n19239 & ~n19270 ;
  assign n19417 = n19268 | n19416 ;
  assign n19418 = n19237 & ~n19270 ;
  assign n19419 = n19268 | n19418 ;
  assign n19420 = ( ~n7061 & n19417 ) | ( ~n7061 & n19419 ) | ( n19417 & n19419 ) ;
  assign n19421 = n19410 | n19413 ;
  assign n19422 = n19409 | n19421 ;
  assign n19423 = n19410 | n19412 ;
  assign n19424 = n19409 | n19423 ;
  assign n19425 = ( ~n8193 & n19422 ) | ( ~n8193 & n19424 ) | ( n19422 & n19424 ) ;
  assign n19426 = n19420 & ~n19425 ;
  assign n19427 = ( n19415 & n19420 ) | ( n19415 & n19426 ) | ( n19420 & n19426 ) ;
  assign n19428 = ~n19420 & n19425 ;
  assign n19429 = ~n19415 & n19428 ;
  assign n19430 = n19427 | n19429 ;
  assign n19431 = n19280 & ~n19300 ;
  assign n19432 = ( n19280 & ~n19282 ) | ( n19280 & n19431 ) | ( ~n19282 & n19431 ) ;
  assign n19433 = n19430 | n19432 ;
  assign n19434 = n19430 & n19432 ;
  assign n19435 = n19433 & ~n19434 ;
  assign n19436 = n1826 & n8079 ;
  assign n19437 = ( n1826 & ~n8070 ) | ( n1826 & n19436 ) | ( ~n8070 & n19436 ) ;
  assign n19438 = n1823 | n19437 ;
  assign n19439 = ( ~n8017 & n19437 ) | ( ~n8017 & n19438 ) | ( n19437 & n19438 ) ;
  assign n19440 = n1829 & n9022 ;
  assign n19441 = ( n1829 & ~n9019 ) | ( n1829 & n19440 ) | ( ~n9019 & n19440 ) ;
  assign n19442 = n19439 | n19441 ;
  assign n19443 = n1821 | n19441 ;
  assign n19444 = n19439 | n19443 ;
  assign n19445 = ( ~n9416 & n19442 ) | ( ~n9416 & n19444 ) | ( n19442 & n19444 ) ;
  assign n19446 = ~x29 & n19444 ;
  assign n19447 = ~x29 & n19442 ;
  assign n19448 = ( ~n9416 & n19446 ) | ( ~n9416 & n19447 ) | ( n19446 & n19447 ) ;
  assign n19449 = x29 | n19447 ;
  assign n19450 = x29 | n19446 ;
  assign n19451 = ( ~n9416 & n19449 ) | ( ~n9416 & n19450 ) | ( n19449 & n19450 ) ;
  assign n19452 = ( ~n19445 & n19448 ) | ( ~n19445 & n19451 ) | ( n19448 & n19451 ) ;
  assign n19453 = n2306 & ~n9442 ;
  assign n19454 = n2306 & ~n9074 ;
  assign n19455 = ( n9440 & n19453 ) | ( n9440 & n19454 ) | ( n19453 & n19454 ) ;
  assign n19456 = n2312 & ~n8982 ;
  assign n19457 = ( n2312 & n9051 ) | ( n2312 & n19456 ) | ( n9051 & n19456 ) ;
  assign n19458 = n19455 | n19457 ;
  assign n19459 = n2306 | n19457 ;
  assign n19460 = ( ~n9442 & n19457 ) | ( ~n9442 & n19459 ) | ( n19457 & n19459 ) ;
  assign n19461 = ( ~n9072 & n19458 ) | ( ~n9072 & n19460 ) | ( n19458 & n19460 ) ;
  assign n19462 = ~x26 & n19458 ;
  assign n19463 = ~x26 & n19460 ;
  assign n19464 = ( ~n9072 & n19462 ) | ( ~n9072 & n19463 ) | ( n19462 & n19463 ) ;
  assign n19465 = x26 | n19462 ;
  assign n19466 = x26 | n19463 ;
  assign n19467 = ( ~n9072 & n19465 ) | ( ~n9072 & n19466 ) | ( n19465 & n19466 ) ;
  assign n19468 = ( ~n19461 & n19464 ) | ( ~n19461 & n19467 ) | ( n19464 & n19467 ) ;
  assign n19469 = n19452 & n19468 ;
  assign n19470 = n19452 & ~n19469 ;
  assign n19471 = ~n19452 & n19468 ;
  assign n19472 = n19470 | n19471 ;
  assign n19473 = n19435 & n19472 ;
  assign n19474 = n19435 | n19472 ;
  assign n19475 = ~n19473 & n19474 ;
  assign n19476 = n19306 & n19475 ;
  assign n19477 = ( n19325 & n19475 ) | ( n19325 & n19476 ) | ( n19475 & n19476 ) ;
  assign n19478 = n19306 | n19475 ;
  assign n19479 = n19325 | n19478 ;
  assign n19480 = ~n19477 & n19479 ;
  assign n19481 = n19333 | n19337 ;
  assign n19482 = n19480 & n19481 ;
  assign n19483 = n19333 | n19339 ;
  assign n19484 = n19480 & n19483 ;
  assign n19485 = ( n18077 & n19482 ) | ( n18077 & n19484 ) | ( n19482 & n19484 ) ;
  assign n19486 = n19333 & n19480 ;
  assign n19487 = ( n19345 & n19480 ) | ( n19345 & n19486 ) | ( n19480 & n19486 ) ;
  assign n19488 = ( n15882 & n19485 ) | ( n15882 & n19487 ) | ( n19485 & n19487 ) ;
  assign n19489 = ( n18077 & n19481 ) | ( n18077 & n19483 ) | ( n19481 & n19483 ) ;
  assign n19490 = n19480 | n19489 ;
  assign n19491 = n19333 | n19345 ;
  assign n19492 = n19480 | n19491 ;
  assign n19493 = ( n15882 & n19490 ) | ( n15882 & n19492 ) | ( n19490 & n19492 ) ;
  assign n19494 = ~n19488 & n19493 ;
  assign n19495 = n19352 & n19494 ;
  assign n19496 = n18576 & n19352 ;
  assign n19497 = n18576 | n19352 ;
  assign n19498 = ~n19496 & n19497 ;
  assign n19499 = n19496 | n19498 ;
  assign n19500 = n19352 | n19494 ;
  assign n19501 = ~n19495 & n19500 ;
  assign n19502 = n19495 | n19501 ;
  assign n19503 = ( n19495 & n19499 ) | ( n19495 & n19502 ) | ( n19499 & n19502 ) ;
  assign n19504 = n19495 | n19496 ;
  assign n19505 = ( n19495 & n19501 ) | ( n19495 & n19504 ) | ( n19501 & n19504 ) ;
  assign n19506 = ( n18577 & n19503 ) | ( n18577 & n19505 ) | ( n19503 & n19505 ) ;
  assign n19507 = n19503 | n19505 ;
  assign n19508 = ( n18604 & n19506 ) | ( n18604 & n19507 ) | ( n19506 & n19507 ) ;
  assign n19509 = ~n19427 & n19430 ;
  assign n19510 = n19250 | n19263 ;
  assign n19511 = n2146 | n13912 ;
  assign n19512 = n10358 | n19511 ;
  assign n19513 = ( ~n1025 & n10793 ) | ( ~n1025 & n19512 ) | ( n10793 & n19512 ) ;
  assign n19514 = n10793 & n19512 ;
  assign n19515 = ( ~n1022 & n19513 ) | ( ~n1022 & n19514 ) | ( n19513 & n19514 ) ;
  assign n19516 = n1026 | n19515 ;
  assign n19517 = n801 | n18458 ;
  assign n19518 = n2748 | n15191 ;
  assign n19519 = n19517 | n19518 ;
  assign n19520 = n450 | n491 ;
  assign n19521 = n952 | n19520 ;
  assign n19522 = n184 | n19521 ;
  assign n19523 = n110 | n19522 ;
  assign n19524 = n19519 | n19523 ;
  assign n19525 = n5069 | n10344 ;
  assign n19526 = n15032 | n19525 ;
  assign n19527 = n4142 | n19526 ;
  assign n19528 = n10374 | n19527 ;
  assign n19529 = n4197 | n6932 ;
  assign n19530 = n1675 | n3431 ;
  assign n19531 = n19529 | n19530 ;
  assign n19532 = n114 | n19531 ;
  assign n19533 = n94 | n806 ;
  assign n19534 = n237 | n355 ;
  assign n19535 = n19533 | n19534 ;
  assign n19536 = n310 | n762 ;
  assign n19537 = n517 | n19536 ;
  assign n19538 = n19535 | n19537 ;
  assign n19539 = n19532 | n19538 ;
  assign n19540 = n19528 | n19539 ;
  assign n19541 = n19524 | n19540 ;
  assign n19542 = n414 | n539 ;
  assign n19543 = n54 | n498 ;
  assign n19544 = n19542 | n19543 ;
  assign n19545 = n179 | n1166 ;
  assign n19546 = n171 | n19545 ;
  assign n19547 = n19544 | n19546 ;
  assign n19548 = n131 | n435 ;
  assign n19549 = n19547 | n19548 ;
  assign n19550 = n19541 | n19549 ;
  assign n19551 = n19516 | n19550 ;
  assign n19552 = n19265 | n19551 ;
  assign n19553 = n19510 | n19552 ;
  assign n19554 = n19267 & n19551 ;
  assign n19555 = n19553 & ~n19554 ;
  assign n19556 = x26 | n19555 ;
  assign n19557 = x26 & ~n19551 ;
  assign n19558 = ( x26 & ~n19267 ) | ( x26 & n19557 ) | ( ~n19267 & n19557 ) ;
  assign n19559 = n19553 & n19558 ;
  assign n19560 = n19556 & ~n19559 ;
  assign n19561 = n19421 & ~n19560 ;
  assign n19562 = n19423 & ~n19560 ;
  assign n19563 = ( ~n8193 & n19561 ) | ( ~n8193 & n19562 ) | ( n19561 & n19562 ) ;
  assign n19564 = ~n19421 & n19560 ;
  assign n19565 = ~n19423 & n19560 ;
  assign n19566 = ( n8193 & n19564 ) | ( n8193 & n19565 ) | ( n19564 & n19565 ) ;
  assign n19567 = n19563 | n19566 ;
  assign n19568 = n1060 & n6889 ;
  assign n19569 = ( n1060 & ~n6884 ) | ( n1060 & n19568 ) | ( ~n6884 & n19568 ) ;
  assign n19570 = n1065 & n7907 ;
  assign n19571 = ( n1065 & n7902 ) | ( n1065 & n19570 ) | ( n7902 & n19570 ) ;
  assign n19572 = n1057 & n8079 ;
  assign n19573 = ( n1057 & ~n8070 ) | ( n1057 & n19572 ) | ( ~n8070 & n19572 ) ;
  assign n19574 = n19571 | n19573 ;
  assign n19575 = n19569 | n19574 ;
  assign n19576 = n1062 | n19575 ;
  assign n19577 = ( ~n8156 & n19575 ) | ( ~n8156 & n19576 ) | ( n19575 & n19576 ) ;
  assign n19578 = n19567 & n19577 ;
  assign n19579 = n19567 | n19577 ;
  assign n19580 = ~n19578 & n19579 ;
  assign n19581 = n19509 | n19580 ;
  assign n19582 = n19427 & ~n19580 ;
  assign n19583 = ( n19432 & n19581 ) | ( n19432 & ~n19582 ) | ( n19581 & ~n19582 ) ;
  assign n19584 = n19509 & n19580 ;
  assign n19585 = ~n19427 & n19580 ;
  assign n19586 = ( n19432 & n19584 ) | ( n19432 & n19585 ) | ( n19584 & n19585 ) ;
  assign n19587 = n19583 & ~n19586 ;
  assign n19588 = n1829 & ~n8982 ;
  assign n19589 = ( n1829 & n9051 ) | ( n1829 & n19588 ) | ( n9051 & n19588 ) ;
  assign n19590 = n1823 & n9022 ;
  assign n19591 = n19589 | n19590 ;
  assign n19592 = n1823 | n19589 ;
  assign n19593 = ( ~n9019 & n19591 ) | ( ~n9019 & n19592 ) | ( n19591 & n19592 ) ;
  assign n19594 = n1826 | n19593 ;
  assign n19595 = ( ~n8017 & n19593 ) | ( ~n8017 & n19594 ) | ( n19593 & n19594 ) ;
  assign n19596 = n1821 | n19595 ;
  assign n19597 = ( ~n10242 & n19595 ) | ( ~n10242 & n19596 ) | ( n19595 & n19596 ) ;
  assign n19598 = ~x29 & n19596 ;
  assign n19599 = ~x29 & n19595 ;
  assign n19600 = ( ~n10242 & n19598 ) | ( ~n10242 & n19599 ) | ( n19598 & n19599 ) ;
  assign n19601 = x29 | n19598 ;
  assign n19602 = x29 | n19599 ;
  assign n19603 = ( ~n10242 & n19601 ) | ( ~n10242 & n19602 ) | ( n19601 & n19602 ) ;
  assign n19604 = ( ~n19597 & n19600 ) | ( ~n19597 & n19603 ) | ( n19600 & n19603 ) ;
  assign n19605 = n19587 & n19604 ;
  assign n19606 = n19587 & ~n19605 ;
  assign n19607 = n19469 | n19472 ;
  assign n19608 = ( n19435 & n19469 ) | ( n19435 & n19607 ) | ( n19469 & n19607 ) ;
  assign n19609 = ~n19587 & n19604 ;
  assign n19610 = n19608 & n19609 ;
  assign n19611 = ( n19606 & n19608 ) | ( n19606 & n19610 ) | ( n19608 & n19610 ) ;
  assign n19612 = n19608 | n19609 ;
  assign n19613 = n19606 | n19612 ;
  assign n19614 = ~n19611 & n19613 ;
  assign n19615 = n19477 | n19482 ;
  assign n19616 = n19614 & n19615 ;
  assign n19617 = n19477 | n19484 ;
  assign n19618 = n19614 & n19617 ;
  assign n19619 = ( n18077 & n19616 ) | ( n18077 & n19618 ) | ( n19616 & n19618 ) ;
  assign n19620 = n19477 | n19486 ;
  assign n19621 = n19614 & n19620 ;
  assign n19622 = n19477 | n19480 ;
  assign n19623 = n19614 & n19622 ;
  assign n19624 = ( n19345 & n19621 ) | ( n19345 & n19623 ) | ( n19621 & n19623 ) ;
  assign n19625 = ( n15882 & n19619 ) | ( n15882 & n19624 ) | ( n19619 & n19624 ) ;
  assign n19626 = ( n19345 & n19620 ) | ( n19345 & n19622 ) | ( n19620 & n19622 ) ;
  assign n19627 = n19614 | n19626 ;
  assign n19628 = ( n18077 & n19615 ) | ( n18077 & n19617 ) | ( n19615 & n19617 ) ;
  assign n19629 = n19614 | n19628 ;
  assign n19630 = ( n15882 & n19627 ) | ( n15882 & n19629 ) | ( n19627 & n19629 ) ;
  assign n19631 = ~n19625 & n19630 ;
  assign n19632 = n19494 & n19631 ;
  assign n19633 = n19494 | n19631 ;
  assign n19634 = ~n19632 & n19633 ;
  assign n19635 = n19503 & n19634 ;
  assign n19636 = n19505 & n19634 ;
  assign n19637 = ( n18577 & n19635 ) | ( n18577 & n19636 ) | ( n19635 & n19636 ) ;
  assign n19638 = n19635 | n19636 ;
  assign n19639 = ( n18604 & n19637 ) | ( n18604 & n19638 ) | ( n19637 & n19638 ) ;
  assign n19640 = n19508 & ~n19639 ;
  assign n19641 = n7074 & n19352 ;
  assign n19642 = n7068 & n19494 ;
  assign n19643 = n19641 | n19642 ;
  assign n19644 = n7079 & n19631 ;
  assign n19645 = n7078 | n19644 ;
  assign n19646 = n19643 | n19645 ;
  assign n19647 = n19643 | n19644 ;
  assign n19648 = n19632 | n19634 ;
  assign n19649 = ( n19503 & n19632 ) | ( n19503 & n19648 ) | ( n19632 & n19648 ) ;
  assign n19650 = ( n19505 & n19632 ) | ( n19505 & n19648 ) | ( n19632 & n19648 ) ;
  assign n19651 = ( n18577 & n19649 ) | ( n18577 & n19650 ) | ( n19649 & n19650 ) ;
  assign n19652 = n19633 & ~n19651 ;
  assign n19653 = n19647 | n19652 ;
  assign n19654 = n19649 | n19650 ;
  assign n19655 = n19633 & ~n19654 ;
  assign n19656 = n19647 | n19655 ;
  assign n19657 = ( ~n18604 & n19653 ) | ( ~n18604 & n19656 ) | ( n19653 & n19656 ) ;
  assign n19658 = n19646 & n19657 ;
  assign n19659 = ( n19640 & n19646 ) | ( n19640 & n19658 ) | ( n19646 & n19658 ) ;
  assign n19660 = ~x8 & n19659 ;
  assign n19661 = x8 | n19659 ;
  assign n19662 = ( ~n19659 & n19660 ) | ( ~n19659 & n19661 ) | ( n19660 & n19661 ) ;
  assign n19663 = n19230 & n19662 ;
  assign n19664 = n19230 & ~n19663 ;
  assign n19665 = ~n19230 & n19662 ;
  assign n19666 = n19664 | n19665 ;
  assign n19667 = ~n18686 & n19223 ;
  assign n19668 = n18686 & ~n19223 ;
  assign n19669 = n19667 | n19668 ;
  assign n19670 = n18577 & n19498 ;
  assign n19671 = ( n18604 & n19498 ) | ( n18604 & n19670 ) | ( n19498 & n19670 ) ;
  assign n19672 = n18577 | n19498 ;
  assign n19673 = n18604 | n19672 ;
  assign n19674 = ~n19671 & n19673 ;
  assign n19676 = n7074 & n18410 ;
  assign n19677 = n7068 & n18576 ;
  assign n19678 = n19676 | n19677 ;
  assign n19675 = n7079 & n19352 ;
  assign n19680 = n7078 | n19675 ;
  assign n19681 = n19678 | n19680 ;
  assign n19679 = n19675 | n19678 ;
  assign n19682 = n19679 & n19681 ;
  assign n19683 = ( n19674 & n19681 ) | ( n19674 & n19682 ) | ( n19681 & n19682 ) ;
  assign n19684 = x8 & n19682 ;
  assign n19685 = x8 & n19681 ;
  assign n19686 = ( n19674 & n19684 ) | ( n19674 & n19685 ) | ( n19684 & n19685 ) ;
  assign n19687 = x8 & ~n19684 ;
  assign n19688 = x8 & ~n19685 ;
  assign n19689 = ( ~n19674 & n19687 ) | ( ~n19674 & n19688 ) | ( n19687 & n19688 ) ;
  assign n19690 = ( n19683 & ~n19686 ) | ( n19683 & n19689 ) | ( ~n19686 & n19689 ) ;
  assign n19691 = ~n19669 & n19690 ;
  assign n19692 = n18707 & n19221 ;
  assign n19693 = n18707 | n19221 ;
  assign n19694 = ~n19692 & n19693 ;
  assign n19696 = n7074 & ~n18585 ;
  assign n19697 = n7068 & n18410 ;
  assign n19698 = n19696 | n19697 ;
  assign n19695 = n7079 & n18576 ;
  assign n19700 = n7078 | n19695 ;
  assign n19701 = n19698 | n19700 ;
  assign n19699 = n19695 | n19698 ;
  assign n19702 = n19699 & n19701 ;
  assign n19703 = ( n18612 & n19701 ) | ( n18612 & n19702 ) | ( n19701 & n19702 ) ;
  assign n19704 = x8 & n19702 ;
  assign n19705 = x8 & n19701 ;
  assign n19706 = ( n18612 & n19704 ) | ( n18612 & n19705 ) | ( n19704 & n19705 ) ;
  assign n19707 = x8 & ~n19704 ;
  assign n19708 = x8 & ~n19705 ;
  assign n19709 = ( ~n18612 & n19707 ) | ( ~n18612 & n19708 ) | ( n19707 & n19708 ) ;
  assign n19710 = ( n19703 & ~n19706 ) | ( n19703 & n19709 ) | ( ~n19706 & n19709 ) ;
  assign n19711 = n19694 & n19710 ;
  assign n19712 = n19217 & ~n19219 ;
  assign n19713 = ~n19217 & n19219 ;
  assign n19714 = n19712 | n19713 ;
  assign n19715 = n7079 & n18410 ;
  assign n19716 = n7074 & n18037 ;
  assign n19717 = n7068 & ~n18585 ;
  assign n19718 = n19716 | n19717 ;
  assign n19719 = n19715 | n19718 ;
  assign n19720 = n18586 & ~n19719 ;
  assign n19721 = ( n18609 & ~n19719 ) | ( n18609 & n19720 ) | ( ~n19719 & n19720 ) ;
  assign n19722 = ~n18650 & n19721 ;
  assign n19723 = n7078 | n19715 ;
  assign n19724 = n19718 | n19723 ;
  assign n19725 = ~n19722 & n19724 ;
  assign n19726 = x8 & n19724 ;
  assign n19727 = ~n19722 & n19726 ;
  assign n19728 = x8 & ~n19726 ;
  assign n19729 = ( x8 & n19722 ) | ( x8 & n19728 ) | ( n19722 & n19728 ) ;
  assign n19730 = ( n19725 & ~n19727 ) | ( n19725 & n19729 ) | ( ~n19727 & n19729 ) ;
  assign n19731 = ~n19714 & n19730 ;
  assign n19732 = n18745 & ~n19215 ;
  assign n19733 = n19216 | n19732 ;
  assign n19734 = n7079 & ~n18585 ;
  assign n19735 = n7074 & ~n17092 ;
  assign n19736 = n7068 & n18037 ;
  assign n19737 = n19735 | n19736 ;
  assign n19738 = n19734 | n19737 ;
  assign n19739 = n18675 & ~n19738 ;
  assign n19740 = ~n18672 & n19739 ;
  assign n19741 = n7078 | n19734 ;
  assign n19742 = n19737 | n19741 ;
  assign n19743 = ~n19740 & n19742 ;
  assign n19744 = x8 & n19742 ;
  assign n19745 = ~n19740 & n19744 ;
  assign n19746 = x8 & ~n19744 ;
  assign n19747 = ( x8 & n19740 ) | ( x8 & n19746 ) | ( n19740 & n19746 ) ;
  assign n19748 = ( n19743 & ~n19745 ) | ( n19743 & n19747 ) | ( ~n19745 & n19747 ) ;
  assign n19749 = ~n19733 & n19748 ;
  assign n19750 = n19733 | n19749 ;
  assign n19751 = n19733 & n19748 ;
  assign n19752 = n19750 & ~n19751 ;
  assign n19753 = n19211 & n19213 ;
  assign n19754 = n19211 | n19213 ;
  assign n19755 = ~n19753 & n19754 ;
  assign n19756 = n7079 & n18037 ;
  assign n19757 = n7074 & n17100 ;
  assign n19758 = n7068 & ~n17092 ;
  assign n19759 = n19757 | n19758 ;
  assign n19760 = n19756 | n19759 ;
  assign n19761 = n7078 | n19756 ;
  assign n19762 = n19759 | n19761 ;
  assign n19763 = ( ~n18050 & n19760 ) | ( ~n18050 & n19762 ) | ( n19760 & n19762 ) ;
  assign n19764 = ~x8 & n19762 ;
  assign n19765 = ~x8 & n19760 ;
  assign n19766 = ( ~n18050 & n19764 ) | ( ~n18050 & n19765 ) | ( n19764 & n19765 ) ;
  assign n19767 = x8 | n19765 ;
  assign n19768 = x8 | n19764 ;
  assign n19769 = ( ~n18050 & n19767 ) | ( ~n18050 & n19768 ) | ( n19767 & n19768 ) ;
  assign n19770 = ( ~n19763 & n19766 ) | ( ~n19763 & n19769 ) | ( n19766 & n19769 ) ;
  assign n19771 = n19755 & n19770 ;
  assign n19772 = ~n18784 & n19209 ;
  assign n19773 = n18784 & ~n19209 ;
  assign n19774 = n19772 | n19773 ;
  assign n19775 = n7079 & ~n17092 ;
  assign n19776 = n7074 & n17111 ;
  assign n19777 = n7068 & n17100 ;
  assign n19778 = n19776 | n19777 ;
  assign n19779 = n19775 | n19778 ;
  assign n19780 = n7078 | n19775 ;
  assign n19781 = n19778 | n19780 ;
  assign n19782 = ( ~n17134 & n19779 ) | ( ~n17134 & n19781 ) | ( n19779 & n19781 ) ;
  assign n19783 = ~x8 & n19781 ;
  assign n19784 = ~x8 & n19779 ;
  assign n19785 = ( ~n17134 & n19783 ) | ( ~n17134 & n19784 ) | ( n19783 & n19784 ) ;
  assign n19786 = x8 | n19784 ;
  assign n19787 = x8 | n19783 ;
  assign n19788 = ( ~n17134 & n19786 ) | ( ~n17134 & n19787 ) | ( n19786 & n19787 ) ;
  assign n19789 = ( ~n19782 & n19785 ) | ( ~n19782 & n19788 ) | ( n19785 & n19788 ) ;
  assign n19790 = n19774 & n19789 ;
  assign n19791 = n19774 | n19789 ;
  assign n19792 = ~n19790 & n19791 ;
  assign n19793 = n19205 & n19207 ;
  assign n19794 = n19205 | n19207 ;
  assign n19795 = ~n19793 & n19794 ;
  assign n19796 = n7074 & ~n16069 ;
  assign n19797 = n7068 & n17111 ;
  assign n19798 = n19796 | n19797 ;
  assign n19799 = n7079 & n17100 ;
  assign n19800 = n7078 | n19799 ;
  assign n19801 = n19798 | n19800 ;
  assign n19802 = n19798 | n19799 ;
  assign n19803 = n17169 | n19802 ;
  assign n19804 = ( ~n17129 & n19802 ) | ( ~n17129 & n19803 ) | ( n19802 & n19803 ) ;
  assign n19805 = n19801 & n19804 ;
  assign n19806 = ( n17161 & n19801 ) | ( n17161 & n19805 ) | ( n19801 & n19805 ) ;
  assign n19807 = ~x8 & n19806 ;
  assign n19808 = x8 | n19806 ;
  assign n19809 = ( ~n19806 & n19807 ) | ( ~n19806 & n19808 ) | ( n19807 & n19808 ) ;
  assign n19810 = n19795 & n19809 ;
  assign n19811 = n18826 & n19203 ;
  assign n19812 = n18826 | n19203 ;
  assign n19813 = ~n19811 & n19812 ;
  assign n19814 = n7074 & n15886 ;
  assign n19815 = n7068 & ~n16069 ;
  assign n19816 = n19814 | n19815 ;
  assign n19817 = n7079 & n17111 ;
  assign n19818 = n7078 | n19817 ;
  assign n19819 = n19816 | n19818 ;
  assign n19820 = n19816 | n19817 ;
  assign n19821 = n17194 & ~n19820 ;
  assign n19822 = ( n17129 & ~n19820 ) | ( n17129 & n19821 ) | ( ~n19820 & n19821 ) ;
  assign n19823 = n19819 & ~n19822 ;
  assign n19824 = ( n17186 & n19819 ) | ( n17186 & n19823 ) | ( n19819 & n19823 ) ;
  assign n19825 = x8 & n19824 ;
  assign n19826 = x8 & ~n19824 ;
  assign n19827 = ( n19824 & ~n19825 ) | ( n19824 & n19826 ) | ( ~n19825 & n19826 ) ;
  assign n19828 = n19813 & n19827 ;
  assign n19829 = n19813 & ~n19828 ;
  assign n19830 = ~n19813 & n19827 ;
  assign n19831 = n19829 | n19830 ;
  assign n19832 = n18848 & n19201 ;
  assign n19833 = n18848 | n19201 ;
  assign n19834 = ~n19832 & n19833 ;
  assign n19835 = n7079 & ~n16069 ;
  assign n19836 = n7074 & ~n16085 ;
  assign n19837 = n7068 & n15886 ;
  assign n19838 = n19836 | n19837 ;
  assign n19839 = n19835 | n19838 ;
  assign n19840 = n7078 | n19839 ;
  assign n19841 = ( ~n16107 & n19839 ) | ( ~n16107 & n19840 ) | ( n19839 & n19840 ) ;
  assign n19842 = ~x8 & n19840 ;
  assign n19843 = ~x8 & n19839 ;
  assign n19844 = ( ~n16107 & n19842 ) | ( ~n16107 & n19843 ) | ( n19842 & n19843 ) ;
  assign n19845 = x8 | n19842 ;
  assign n19846 = x8 | n19843 ;
  assign n19847 = ( ~n16107 & n19845 ) | ( ~n16107 & n19846 ) | ( n19845 & n19846 ) ;
  assign n19848 = ( ~n19841 & n19844 ) | ( ~n19841 & n19847 ) | ( n19844 & n19847 ) ;
  assign n19849 = n19834 & n19848 ;
  assign n19850 = n19834 & ~n19849 ;
  assign n19851 = ~n19834 & n19848 ;
  assign n19852 = n19850 | n19851 ;
  assign n19853 = ( n18890 & n18891 ) | ( n18890 & n19199 ) | ( n18891 & n19199 ) ;
  assign n19854 = n18868 | n18890 ;
  assign n19855 = n19199 | n19854 ;
  assign n19856 = ~n19853 & n19855 ;
  assign n19857 = n7079 & n15886 ;
  assign n19858 = n7074 & n15434 ;
  assign n19859 = n7068 & ~n16085 ;
  assign n19860 = n19858 | n19859 ;
  assign n19861 = n19857 | n19860 ;
  assign n19862 = n7078 | n19857 ;
  assign n19863 = n19860 | n19862 ;
  assign n19864 = ( ~n16140 & n19861 ) | ( ~n16140 & n19863 ) | ( n19861 & n19863 ) ;
  assign n19865 = ~x8 & n19863 ;
  assign n19866 = ~x8 & n19861 ;
  assign n19867 = ( ~n16140 & n19865 ) | ( ~n16140 & n19866 ) | ( n19865 & n19866 ) ;
  assign n19868 = x8 | n19866 ;
  assign n19869 = x8 | n19865 ;
  assign n19870 = ( ~n16140 & n19868 ) | ( ~n16140 & n19869 ) | ( n19868 & n19869 ) ;
  assign n19871 = ( ~n19864 & n19867 ) | ( ~n19864 & n19870 ) | ( n19867 & n19870 ) ;
  assign n19872 = n19856 & n19871 ;
  assign n19873 = n19195 & ~n19199 ;
  assign n19874 = n19198 & ~n19199 ;
  assign n19875 = n19873 | n19874 ;
  assign n19876 = n7079 & ~n16085 ;
  assign n19877 = n7074 & n14591 ;
  assign n19878 = n7068 & n15434 ;
  assign n19879 = n19877 | n19878 ;
  assign n19880 = n19876 | n19879 ;
  assign n19881 = n7078 | n19876 ;
  assign n19882 = n19879 | n19881 ;
  assign n19883 = ( ~n16167 & n19880 ) | ( ~n16167 & n19882 ) | ( n19880 & n19882 ) ;
  assign n19884 = ~x8 & n19882 ;
  assign n19885 = ~x8 & n19880 ;
  assign n19886 = ( ~n16167 & n19884 ) | ( ~n16167 & n19885 ) | ( n19884 & n19885 ) ;
  assign n19887 = x8 | n19885 ;
  assign n19888 = x8 | n19884 ;
  assign n19889 = ( ~n16167 & n19887 ) | ( ~n16167 & n19888 ) | ( n19887 & n19888 ) ;
  assign n19890 = ( ~n19883 & n19886 ) | ( ~n19883 & n19889 ) | ( n19886 & n19889 ) ;
  assign n19891 = n19875 & n19890 ;
  assign n19892 = n19875 & ~n19891 ;
  assign n19893 = ~n19875 & n19890 ;
  assign n19894 = n19892 | n19893 ;
  assign n19895 = n19193 & ~n19194 ;
  assign n19896 = n18914 & ~n19194 ;
  assign n19897 = n19895 | n19896 ;
  assign n19898 = n7079 & n15434 ;
  assign n19899 = n7074 & n14329 ;
  assign n19900 = n7068 & n14591 ;
  assign n19901 = n19899 | n19900 ;
  assign n19902 = n19898 | n19901 ;
  assign n19903 = n7078 | n19898 ;
  assign n19904 = n19901 | n19903 ;
  assign n19905 = ( n15453 & n19902 ) | ( n15453 & n19904 ) | ( n19902 & n19904 ) ;
  assign n19906 = x8 & n19904 ;
  assign n19907 = x8 & n19902 ;
  assign n19908 = ( n15453 & n19906 ) | ( n15453 & n19907 ) | ( n19906 & n19907 ) ;
  assign n19909 = x8 & ~n19907 ;
  assign n19910 = x8 & ~n19906 ;
  assign n19911 = ( ~n15453 & n19909 ) | ( ~n15453 & n19910 ) | ( n19909 & n19910 ) ;
  assign n19912 = ( n19905 & ~n19908 ) | ( n19905 & n19911 ) | ( ~n19908 & n19911 ) ;
  assign n19913 = n19897 & n19912 ;
  assign n19914 = n19897 & ~n19913 ;
  assign n19915 = ~n19897 & n19912 ;
  assign n19916 = n19914 | n19915 ;
  assign n19917 = n19185 | n19186 ;
  assign n19918 = n18952 | n19917 ;
  assign n19919 = ~n19188 & n19918 ;
  assign n19921 = n7074 & n13522 ;
  assign n19922 = n7068 & n14607 ;
  assign n19923 = n19921 | n19922 ;
  assign n19920 = n7079 & n14329 ;
  assign n19925 = n7078 | n19920 ;
  assign n19926 = n19923 | n19925 ;
  assign n19924 = n19920 | n19923 ;
  assign n19927 = n19924 & n19926 ;
  assign n19928 = ( n14656 & n19926 ) | ( n14656 & n19927 ) | ( n19926 & n19927 ) ;
  assign n19929 = x8 & n19927 ;
  assign n19930 = x8 & n19926 ;
  assign n19931 = ( n14656 & n19929 ) | ( n14656 & n19930 ) | ( n19929 & n19930 ) ;
  assign n19932 = x8 & ~n19929 ;
  assign n19933 = x8 & ~n19930 ;
  assign n19934 = ( ~n14656 & n19932 ) | ( ~n14656 & n19933 ) | ( n19932 & n19933 ) ;
  assign n19935 = ( n19928 & ~n19931 ) | ( n19928 & n19934 ) | ( ~n19931 & n19934 ) ;
  assign n19936 = n19919 & n19935 ;
  assign n19937 = n19189 & n19191 ;
  assign n19938 = n19189 | n19191 ;
  assign n19939 = ~n19937 & n19938 ;
  assign n19941 = n7074 & n14607 ;
  assign n19942 = n7068 & n14329 ;
  assign n19943 = n19941 | n19942 ;
  assign n19940 = n7079 & n14591 ;
  assign n19945 = n7078 | n19940 ;
  assign n19946 = n19943 | n19945 ;
  assign n19944 = n19940 | n19943 ;
  assign n19947 = n19944 & n19946 ;
  assign n19948 = ( n14629 & n19946 ) | ( n14629 & n19947 ) | ( n19946 & n19947 ) ;
  assign n19949 = x8 & n19947 ;
  assign n19950 = x8 & n19946 ;
  assign n19951 = ( n14629 & n19949 ) | ( n14629 & n19950 ) | ( n19949 & n19950 ) ;
  assign n19952 = x8 & ~n19949 ;
  assign n19953 = x8 & ~n19950 ;
  assign n19954 = ( ~n14629 & n19952 ) | ( ~n14629 & n19953 ) | ( n19952 & n19953 ) ;
  assign n19955 = ( n19948 & ~n19951 ) | ( n19948 & n19954 ) | ( ~n19951 & n19954 ) ;
  assign n19956 = n19939 & n19955 ;
  assign n19957 = n19939 | n19955 ;
  assign n19958 = ~n19956 & n19957 ;
  assign n19959 = n19936 & n19958 ;
  assign n19960 = n19956 | n19958 ;
  assign n19961 = n19181 & n19183 ;
  assign n19962 = n19181 | n19183 ;
  assign n19963 = ~n19961 & n19962 ;
  assign n19964 = n7074 & n13235 ;
  assign n19965 = n7068 & n13522 ;
  assign n19966 = n19964 | n19965 ;
  assign n19967 = n7079 & n14607 ;
  assign n19968 = n7078 | n19967 ;
  assign n19969 = n19966 | n19968 ;
  assign n19970 = n19966 | n19967 ;
  assign n19971 = n14696 | n19970 ;
  assign n19972 = n14698 | n19970 ;
  assign n19973 = ( ~n13248 & n19971 ) | ( ~n13248 & n19972 ) | ( n19971 & n19972 ) ;
  assign n19974 = n19969 & n19973 ;
  assign n19975 = ( n14687 & n19969 ) | ( n14687 & n19974 ) | ( n19969 & n19974 ) ;
  assign n19976 = ~x8 & n19975 ;
  assign n19977 = x8 | n19975 ;
  assign n19978 = ( ~n19975 & n19976 ) | ( ~n19975 & n19977 ) | ( n19976 & n19977 ) ;
  assign n19979 = n19963 & n19978 ;
  assign n19980 = n19963 & ~n19979 ;
  assign n19981 = ~n19963 & n19978 ;
  assign n19982 = n19980 | n19981 ;
  assign n19983 = n19177 & n19179 ;
  assign n19984 = n19177 | n19179 ;
  assign n19985 = ~n19983 & n19984 ;
  assign n19986 = n7079 & n13522 ;
  assign n19987 = n7074 & n12936 ;
  assign n19988 = n7068 & n13235 ;
  assign n19989 = n19987 | n19988 ;
  assign n19990 = n19986 | n19989 ;
  assign n19991 = n7078 & n13537 ;
  assign n19992 = n7078 & n13539 ;
  assign n19993 = ( ~n13248 & n19991 ) | ( ~n13248 & n19992 ) | ( n19991 & n19992 ) ;
  assign n19994 = n19990 | n19993 ;
  assign n19995 = n7078 | n19990 ;
  assign n19996 = ( n13530 & n19994 ) | ( n13530 & n19995 ) | ( n19994 & n19995 ) ;
  assign n19997 = x8 | n19996 ;
  assign n19998 = ~x8 & n19996 ;
  assign n19999 = ( ~n19996 & n19997 ) | ( ~n19996 & n19998 ) | ( n19997 & n19998 ) ;
  assign n20000 = n19985 & n19999 ;
  assign n20001 = n19175 & ~n19176 ;
  assign n20002 = n19011 & ~n19176 ;
  assign n20003 = n20001 | n20002 ;
  assign n20004 = n7079 & n13235 ;
  assign n20005 = n7074 & ~n12616 ;
  assign n20006 = n7068 & n12936 ;
  assign n20007 = n20005 | n20006 ;
  assign n20008 = n20004 | n20007 ;
  assign n20009 = n7078 | n20004 ;
  assign n20010 = n20007 | n20009 ;
  assign n20011 = ( n13561 & n20008 ) | ( n13561 & n20010 ) | ( n20008 & n20010 ) ;
  assign n20012 = x8 & n20010 ;
  assign n20013 = x8 & n20008 ;
  assign n20014 = ( n13561 & n20012 ) | ( n13561 & n20013 ) | ( n20012 & n20013 ) ;
  assign n20015 = x8 & ~n20013 ;
  assign n20016 = x8 & ~n20012 ;
  assign n20017 = ( ~n13561 & n20015 ) | ( ~n13561 & n20016 ) | ( n20015 & n20016 ) ;
  assign n20018 = ( n20011 & ~n20014 ) | ( n20011 & n20017 ) | ( ~n20014 & n20017 ) ;
  assign n20019 = n20003 & n20018 ;
  assign n20020 = n20003 & ~n20019 ;
  assign n20021 = ~n19031 & n19173 ;
  assign n20022 = n19031 & ~n19173 ;
  assign n20023 = n20021 | n20022 ;
  assign n20024 = n7079 & n12936 ;
  assign n20025 = n7074 & n12010 ;
  assign n20026 = n7068 & ~n12616 ;
  assign n20027 = n20025 | n20026 ;
  assign n20028 = n20024 | n20027 ;
  assign n20029 = n7078 | n20024 ;
  assign n20030 = n20027 | n20029 ;
  assign n20031 = ( ~n13591 & n20028 ) | ( ~n13591 & n20030 ) | ( n20028 & n20030 ) ;
  assign n20032 = ~x8 & n20030 ;
  assign n20033 = ~x8 & n20028 ;
  assign n20034 = ( ~n13591 & n20032 ) | ( ~n13591 & n20033 ) | ( n20032 & n20033 ) ;
  assign n20035 = x8 | n20033 ;
  assign n20036 = x8 | n20032 ;
  assign n20037 = ( ~n13591 & n20035 ) | ( ~n13591 & n20036 ) | ( n20035 & n20036 ) ;
  assign n20038 = ( ~n20031 & n20034 ) | ( ~n20031 & n20037 ) | ( n20034 & n20037 ) ;
  assign n20039 = n20023 & n20038 ;
  assign n20040 = n19169 & n19171 ;
  assign n20041 = n19169 | n19171 ;
  assign n20042 = ~n20040 & n20041 ;
  assign n20044 = n7074 & ~n11663 ;
  assign n20045 = n7068 & n12010 ;
  assign n20046 = n20044 | n20045 ;
  assign n20043 = n7079 & ~n12616 ;
  assign n20048 = n7078 | n20043 ;
  assign n20049 = n20046 | n20048 ;
  assign n20047 = n20043 | n20046 ;
  assign n20050 = n20047 & n20049 ;
  assign n20051 = ( ~n12626 & n20049 ) | ( ~n12626 & n20050 ) | ( n20049 & n20050 ) ;
  assign n20052 = ~x8 & n20050 ;
  assign n20053 = ~x8 & n20049 ;
  assign n20054 = ( ~n12626 & n20052 ) | ( ~n12626 & n20053 ) | ( n20052 & n20053 ) ;
  assign n20055 = x8 | n20052 ;
  assign n20056 = x8 | n20053 ;
  assign n20057 = ( ~n12626 & n20055 ) | ( ~n12626 & n20056 ) | ( n20055 & n20056 ) ;
  assign n20058 = ( ~n20051 & n20054 ) | ( ~n20051 & n20057 ) | ( n20054 & n20057 ) ;
  assign n20059 = n20042 & n20058 ;
  assign n20060 = n19070 | n19167 ;
  assign n20061 = ~n19168 & n20060 ;
  assign n20063 = n7074 & n11363 ;
  assign n20064 = n7068 & ~n11663 ;
  assign n20065 = n20063 | n20064 ;
  assign n20062 = n7079 & n12010 ;
  assign n20067 = n7078 | n20062 ;
  assign n20068 = n20065 | n20067 ;
  assign n20066 = n20062 | n20065 ;
  assign n20069 = n20066 & n20068 ;
  assign n20070 = ( ~n12028 & n20068 ) | ( ~n12028 & n20069 ) | ( n20068 & n20069 ) ;
  assign n20071 = n20068 | n20069 ;
  assign n20072 = ( n12017 & n20070 ) | ( n12017 & n20071 ) | ( n20070 & n20071 ) ;
  assign n20073 = ~x8 & n20072 ;
  assign n20074 = x8 | n20072 ;
  assign n20075 = ( ~n20072 & n20073 ) | ( ~n20072 & n20074 ) | ( n20073 & n20074 ) ;
  assign n20076 = n20061 & n20075 ;
  assign n20077 = n20061 & ~n20076 ;
  assign n20078 = ~n20061 & n20075 ;
  assign n20079 = n20077 | n20078 ;
  assign n20080 = n19094 | n19165 ;
  assign n20081 = ~n19166 & n20080 ;
  assign n20082 = n7074 & n10649 ;
  assign n20083 = n7068 & n11363 ;
  assign n20084 = n20082 | n20083 ;
  assign n20085 = n7079 & ~n11663 ;
  assign n20086 = n7078 | n20085 ;
  assign n20087 = n20084 | n20086 ;
  assign n20088 = n20084 | n20085 ;
  assign n20089 = n12048 & ~n20088 ;
  assign n20090 = ( n11672 & ~n20088 ) | ( n11672 & n20089 ) | ( ~n20088 & n20089 ) ;
  assign n20091 = n20087 & ~n20090 ;
  assign n20092 = ( n12040 & n20087 ) | ( n12040 & n20091 ) | ( n20087 & n20091 ) ;
  assign n20093 = x8 & n20092 ;
  assign n20094 = x8 & ~n20092 ;
  assign n20095 = ( n20092 & ~n20093 ) | ( n20092 & n20094 ) | ( ~n20093 & n20094 ) ;
  assign n20096 = n20081 & n20095 ;
  assign n20097 = n20081 & ~n20096 ;
  assign n20098 = ~n20081 & n20095 ;
  assign n20099 = n20097 | n20098 ;
  assign n20100 = n19161 & n19163 ;
  assign n20101 = n19161 | n19163 ;
  assign n20102 = ~n20100 & n20101 ;
  assign n20103 = n7079 & n11363 ;
  assign n20104 = n7074 & n10325 ;
  assign n20105 = n7068 & n10649 ;
  assign n20106 = n20104 | n20105 ;
  assign n20107 = n20103 | n20106 ;
  assign n20108 = n7078 | n20107 ;
  assign n20109 = ( n12059 & n20107 ) | ( n12059 & n20108 ) | ( n20107 & n20108 ) ;
  assign n20110 = x8 & n20108 ;
  assign n20111 = x8 & n20107 ;
  assign n20112 = ( n12059 & n20110 ) | ( n12059 & n20111 ) | ( n20110 & n20111 ) ;
  assign n20113 = x8 & ~n20110 ;
  assign n20114 = x8 & ~n20111 ;
  assign n20115 = ( ~n12059 & n20113 ) | ( ~n12059 & n20114 ) | ( n20113 & n20114 ) ;
  assign n20116 = ( n20109 & ~n20112 ) | ( n20109 & n20115 ) | ( ~n20112 & n20115 ) ;
  assign n20117 = n20102 & n20116 ;
  assign n20118 = n19148 & n19159 ;
  assign n20119 = n19148 & ~n20118 ;
  assign n20120 = n7079 & n10649 ;
  assign n20121 = n7074 & n10654 ;
  assign n20122 = n7068 & n10325 ;
  assign n20123 = n20121 | n20122 ;
  assign n20124 = n20120 | n20123 ;
  assign n20125 = n7078 | n20120 ;
  assign n20126 = n20123 | n20125 ;
  assign n20127 = ( n10702 & n20124 ) | ( n10702 & n20126 ) | ( n20124 & n20126 ) ;
  assign n20128 = n20124 | n20126 ;
  assign n20129 = ( n10695 & n20127 ) | ( n10695 & n20128 ) | ( n20127 & n20128 ) ;
  assign n20130 = x8 & n20129 ;
  assign n20131 = x8 & ~n20129 ;
  assign n20132 = ( n20129 & ~n20130 ) | ( n20129 & n20131 ) | ( ~n20130 & n20131 ) ;
  assign n20133 = ~n19148 & n19159 ;
  assign n20134 = n20132 & n20133 ;
  assign n20135 = ( n20119 & n20132 ) | ( n20119 & n20134 ) | ( n20132 & n20134 ) ;
  assign n20136 = n20132 | n20133 ;
  assign n20137 = n20119 | n20136 ;
  assign n20138 = ~n20135 & n20137 ;
  assign n20139 = n7079 & n10325 ;
  assign n20140 = n7074 & ~n10662 ;
  assign n20141 = n7068 & n10654 ;
  assign n20142 = n20140 | n20141 ;
  assign n20143 = n20139 | n20142 ;
  assign n20144 = n7078 | n20143 ;
  assign n20145 = ( ~n10957 & n20143 ) | ( ~n10957 & n20144 ) | ( n20143 & n20144 ) ;
  assign n20146 = n20143 | n20144 ;
  assign n20147 = ( n10949 & n20145 ) | ( n10949 & n20146 ) | ( n20145 & n20146 ) ;
  assign n20148 = ~x8 & n20147 ;
  assign n20149 = x8 & n20143 ;
  assign n20150 = x8 & n7078 ;
  assign n20151 = ( x8 & n20143 ) | ( x8 & n20150 ) | ( n20143 & n20150 ) ;
  assign n20152 = ( ~n10957 & n20149 ) | ( ~n10957 & n20151 ) | ( n20149 & n20151 ) ;
  assign n20153 = n20149 | n20151 ;
  assign n20154 = ( n10949 & n20152 ) | ( n10949 & n20153 ) | ( n20152 & n20153 ) ;
  assign n20155 = x8 & ~n20154 ;
  assign n20156 = n20148 | n20155 ;
  assign n20157 = n19127 & n19145 ;
  assign n20158 = n19127 | n19145 ;
  assign n20159 = ~n20157 & n20158 ;
  assign n20160 = n20156 & n20159 ;
  assign n20161 = n20156 | n20159 ;
  assign n20162 = ~n20160 & n20161 ;
  assign n20163 = n19120 | n19123 ;
  assign n20164 = ~n19123 & n19125 ;
  assign n20165 = ( n19121 & n20163 ) | ( n19121 & ~n20164 ) | ( n20163 & ~n20164 ) ;
  assign n20166 = ~n19127 & n20165 ;
  assign n20167 = n7079 & n10654 ;
  assign n20168 = n7074 & n10667 ;
  assign n20169 = n7068 & ~n10662 ;
  assign n20170 = n20168 | n20169 ;
  assign n20171 = n20167 | n20170 ;
  assign n20172 = n7078 | n20167 ;
  assign n20173 = n20170 | n20172 ;
  assign n20174 = ( n10978 & n20171 ) | ( n10978 & n20173 ) | ( n20171 & n20173 ) ;
  assign n20175 = x8 & n20173 ;
  assign n20176 = x8 & n20171 ;
  assign n20177 = ( n10978 & n20175 ) | ( n10978 & n20176 ) | ( n20175 & n20176 ) ;
  assign n20178 = x8 & ~n20176 ;
  assign n20179 = x8 & ~n20175 ;
  assign n20180 = ( ~n10978 & n20178 ) | ( ~n10978 & n20179 ) | ( n20178 & n20179 ) ;
  assign n20181 = ( n20174 & ~n20177 ) | ( n20174 & n20180 ) | ( ~n20177 & n20180 ) ;
  assign n20182 = n20166 & n20181 ;
  assign n20183 = n7078 & n10784 ;
  assign n20184 = n7068 & ~n10678 ;
  assign n20185 = n7079 & ~n10675 ;
  assign n20186 = n20184 | n20185 ;
  assign n20187 = x8 | n20186 ;
  assign n20188 = n20183 | n20187 ;
  assign n20189 = ~x8 & n20188 ;
  assign n20190 = x8 & ~n7067 ;
  assign n20191 = ( x8 & n10678 ) | ( x8 & n20190 ) | ( n10678 & n20190 ) ;
  assign n20192 = n20188 & n20191 ;
  assign n20193 = n20183 | n20186 ;
  assign n20194 = n20191 & ~n20193 ;
  assign n20195 = ( n20189 & n20192 ) | ( n20189 & n20194 ) | ( n20192 & n20194 ) ;
  assign n20196 = n7079 & n10667 ;
  assign n20197 = n7074 & ~n10678 ;
  assign n20198 = n7068 & ~n10675 ;
  assign n20199 = n20197 | n20198 ;
  assign n20200 = n20196 | n20199 ;
  assign n20201 = n10837 | n20200 ;
  assign n20202 = n7078 | n20196 ;
  assign n20203 = n20199 | n20202 ;
  assign n20204 = ~x8 & n20203 ;
  assign n20205 = n20201 & n20204 ;
  assign n20206 = x8 | n20205 ;
  assign n20207 = n6114 & ~n10678 ;
  assign n20208 = n20205 & n20207 ;
  assign n20209 = n20201 & n20203 ;
  assign n20210 = n20207 & ~n20209 ;
  assign n20211 = ( n20206 & n20208 ) | ( n20206 & n20210 ) | ( n20208 & n20210 ) ;
  assign n20212 = n20195 & n20211 ;
  assign n20213 = ( n20205 & n20206 ) | ( n20205 & ~n20209 ) | ( n20206 & ~n20209 ) ;
  assign n20214 = n20195 | n20207 ;
  assign n20215 = ( n20207 & n20213 ) | ( n20207 & n20214 ) | ( n20213 & n20214 ) ;
  assign n20216 = ~n20212 & n20215 ;
  assign n20217 = n7079 & ~n10662 ;
  assign n20218 = n7074 & ~n10675 ;
  assign n20219 = n7068 & n10667 ;
  assign n20220 = n20218 | n20219 ;
  assign n20221 = n20217 | n20220 ;
  assign n20222 = ( n7078 & n10850 ) | ( n7078 & n20221 ) | ( n10850 & n20221 ) ;
  assign n20223 = ( x8 & n7078 ) | ( x8 & ~n20221 ) | ( n7078 & ~n20221 ) ;
  assign n20224 = ( x8 & n10850 ) | ( x8 & n20223 ) | ( n10850 & n20223 ) ;
  assign n20225 = ~n20222 & n20224 ;
  assign n20226 = n20221 | n20224 ;
  assign n20227 = ( ~x8 & n20225 ) | ( ~x8 & n20226 ) | ( n20225 & n20226 ) ;
  assign n20228 = n20212 | n20227 ;
  assign n20229 = ( n20212 & n20216 ) | ( n20212 & n20228 ) | ( n20216 & n20228 ) ;
  assign n20230 = n20166 | n20181 ;
  assign n20231 = ~n20182 & n20230 ;
  assign n20232 = n20182 | n20231 ;
  assign n20233 = ( n20182 & n20229 ) | ( n20182 & n20232 ) | ( n20229 & n20232 ) ;
  assign n20234 = n20162 & n20233 ;
  assign n20235 = n20160 | n20234 ;
  assign n20236 = n20138 & n20235 ;
  assign n20237 = n20135 | n20236 ;
  assign n20238 = ~n20102 & n20116 ;
  assign n20239 = ( n20102 & ~n20117 ) | ( n20102 & n20238 ) | ( ~n20117 & n20238 ) ;
  assign n20240 = n20117 | n20239 ;
  assign n20241 = ( n20117 & n20237 ) | ( n20117 & n20240 ) | ( n20237 & n20240 ) ;
  assign n20242 = n20099 & n20241 ;
  assign n20243 = n20096 | n20242 ;
  assign n20244 = n20079 & n20243 ;
  assign n20245 = n20076 | n20244 ;
  assign n20246 = n20042 | n20058 ;
  assign n20247 = ~n20059 & n20246 ;
  assign n20248 = n20059 | n20247 ;
  assign n20249 = ( n20059 & n20245 ) | ( n20059 & n20248 ) | ( n20245 & n20248 ) ;
  assign n20250 = n20023 | n20038 ;
  assign n20251 = ~n20039 & n20250 ;
  assign n20252 = n20039 | n20251 ;
  assign n20253 = ( n20039 & n20249 ) | ( n20039 & n20252 ) | ( n20249 & n20252 ) ;
  assign n20254 = ~n20003 & n20018 ;
  assign n20255 = n20253 & n20254 ;
  assign n20256 = ( n20020 & n20253 ) | ( n20020 & n20255 ) | ( n20253 & n20255 ) ;
  assign n20257 = n20019 | n20256 ;
  assign n20258 = ~n19985 & n19999 ;
  assign n20259 = ( n19985 & ~n20000 ) | ( n19985 & n20258 ) | ( ~n20000 & n20258 ) ;
  assign n20260 = n20000 | n20259 ;
  assign n20261 = ( n20000 & n20257 ) | ( n20000 & n20260 ) | ( n20257 & n20260 ) ;
  assign n20262 = n19982 & n20261 ;
  assign n20263 = n19979 | n20262 ;
  assign n20264 = n19919 & ~n19936 ;
  assign n20265 = ~n19919 & n19935 ;
  assign n20266 = n20264 | n20265 ;
  assign n20267 = n20263 & n20266 ;
  assign n20268 = n19956 | n20267 ;
  assign n20269 = ( n19959 & n19960 ) | ( n19959 & n20268 ) | ( n19960 & n20268 ) ;
  assign n20270 = n19913 | n20269 ;
  assign n20271 = ( n19913 & n19916 ) | ( n19913 & n20270 ) | ( n19916 & n20270 ) ;
  assign n20272 = n19891 | n20271 ;
  assign n20273 = ( n19891 & n19894 ) | ( n19891 & n20272 ) | ( n19894 & n20272 ) ;
  assign n20274 = ~n19856 & n19871 ;
  assign n20275 = ( n19856 & ~n19872 ) | ( n19856 & n20274 ) | ( ~n19872 & n20274 ) ;
  assign n20276 = n19872 | n20275 ;
  assign n20277 = ( n19872 & n20273 ) | ( n19872 & n20276 ) | ( n20273 & n20276 ) ;
  assign n20278 = n19849 | n20277 ;
  assign n20279 = ( n19849 & n19852 ) | ( n19849 & n20278 ) | ( n19852 & n20278 ) ;
  assign n20280 = n19828 | n20279 ;
  assign n20281 = ( n19828 & n19831 ) | ( n19828 & n20280 ) | ( n19831 & n20280 ) ;
  assign n20282 = n19795 | n19809 ;
  assign n20283 = ~n19810 & n20282 ;
  assign n20284 = n19810 | n20283 ;
  assign n20285 = ( n19810 & n20281 ) | ( n19810 & n20284 ) | ( n20281 & n20284 ) ;
  assign n20286 = n19792 & n20285 ;
  assign n20287 = n19790 | n20286 ;
  assign n20288 = ~n19755 & n19770 ;
  assign n20289 = ( n19755 & ~n19771 ) | ( n19755 & n20288 ) | ( ~n19771 & n20288 ) ;
  assign n20290 = n19771 | n20289 ;
  assign n20291 = ( n19771 & n20287 ) | ( n19771 & n20290 ) | ( n20287 & n20290 ) ;
  assign n20292 = ~n19752 & n20291 ;
  assign n20293 = n19749 | n20292 ;
  assign n20294 = n19714 | n19731 ;
  assign n20295 = n19714 & n19730 ;
  assign n20296 = n20294 & ~n20295 ;
  assign n20297 = n20293 & ~n20296 ;
  assign n20298 = n19731 | n20297 ;
  assign n20299 = n19694 & ~n19711 ;
  assign n20300 = ~n19694 & n19710 ;
  assign n20301 = n20299 | n20300 ;
  assign n20302 = n20298 & n20301 ;
  assign n20303 = n19711 | n20302 ;
  assign n20304 = n19669 | n19691 ;
  assign n20305 = n19669 & n19690 ;
  assign n20306 = n20304 & ~n20305 ;
  assign n20307 = n20303 & ~n20306 ;
  assign n20308 = n19691 | n20307 ;
  assign n20309 = n18662 & ~n19225 ;
  assign n20310 = n19226 | n20309 ;
  assign n20311 = n19499 & n19501 ;
  assign n20312 = n19496 & n19501 ;
  assign n20313 = ( n18577 & n20311 ) | ( n18577 & n20312 ) | ( n20311 & n20312 ) ;
  assign n20314 = n20311 | n20312 ;
  assign n20315 = ( n18604 & n20313 ) | ( n18604 & n20314 ) | ( n20313 & n20314 ) ;
  assign n20316 = ( n18576 & n18577 ) | ( n18576 & n19352 ) | ( n18577 & n19352 ) ;
  assign n20317 = n19501 | n20316 ;
  assign n20318 = n19497 | n19501 ;
  assign n20319 = ( n18604 & n20317 ) | ( n18604 & n20318 ) | ( n20317 & n20318 ) ;
  assign n20320 = ~n20315 & n20319 ;
  assign n20322 = n7074 & n18576 ;
  assign n20323 = n7068 & n19352 ;
  assign n20324 = n20322 | n20323 ;
  assign n20321 = n7079 & n19494 ;
  assign n20326 = n7078 | n20321 ;
  assign n20327 = n20324 | n20326 ;
  assign n20325 = n20321 | n20324 ;
  assign n20328 = n20325 & n20327 ;
  assign n20329 = ( n20320 & n20327 ) | ( n20320 & n20328 ) | ( n20327 & n20328 ) ;
  assign n20330 = x8 & n20328 ;
  assign n20331 = x8 & n20327 ;
  assign n20332 = ( n20320 & n20330 ) | ( n20320 & n20331 ) | ( n20330 & n20331 ) ;
  assign n20333 = x8 & ~n20330 ;
  assign n20334 = x8 & ~n20331 ;
  assign n20335 = ( ~n20320 & n20333 ) | ( ~n20320 & n20334 ) | ( n20333 & n20334 ) ;
  assign n20336 = ( n20329 & ~n20332 ) | ( n20329 & n20335 ) | ( ~n20332 & n20335 ) ;
  assign n20337 = ~n20310 & n20336 ;
  assign n20338 = n20310 | n20337 ;
  assign n20339 = n20310 & n20336 ;
  assign n20340 = n20338 & ~n20339 ;
  assign n20341 = ~n20337 & n20340 ;
  assign n20342 = ( n20308 & n20337 ) | ( n20308 & ~n20341 ) | ( n20337 & ~n20341 ) ;
  assign n20343 = n19666 & n20342 ;
  assign n20344 = n19666 & ~n20343 ;
  assign n20345 = ~n19666 & n20342 ;
  assign n20346 = n20344 | n20345 ;
  assign n20347 = n6891 | n7982 ;
  assign n20348 = n1124 | n5154 ;
  assign n20349 = n20347 | n20348 ;
  assign n20350 = n858 | n20349 ;
  assign n20351 = n1340 | n2835 ;
  assign n20352 = n1483 | n20351 ;
  assign n20353 = n225 | n13826 ;
  assign n20354 = n264 | n491 ;
  assign n20355 = n20353 | n20354 ;
  assign n20356 = n20352 | n20355 ;
  assign n20357 = n20350 | n20356 ;
  assign n20358 = n1460 | n4170 ;
  assign n20359 = n110 | n141 ;
  assign n20360 = n20358 | n20359 ;
  assign n20361 = n8004 | n20360 ;
  assign n20362 = n7969 | n20361 ;
  assign n20363 = n20357 | n20362 ;
  assign n20364 = n8069 | n20363 ;
  assign n20365 = n381 | n4246 ;
  assign n20366 = n324 | n20365 ;
  assign n20367 = n347 | n20366 ;
  assign n20368 = n7925 | n20367 ;
  assign n20369 = n20364 | n20368 ;
  assign n20370 = n10913 | n10916 ;
  assign n20371 = n795 | n4330 ;
  assign n20372 = n245 | n269 ;
  assign n20373 = n333 | n435 ;
  assign n20374 = n20372 | n20373 ;
  assign n20375 = n20371 | n20374 ;
  assign n20376 = n2849 | n20375 ;
  assign n20377 = ( ~n741 & n20370 ) | ( ~n741 & n20376 ) | ( n20370 & n20376 ) ;
  assign n20378 = n20370 & n20376 ;
  assign n20379 = ( n734 & n20377 ) | ( n734 & n20378 ) | ( n20377 & n20378 ) ;
  assign n20380 = n742 & ~n20379 ;
  assign n20381 = n325 | n806 ;
  assign n20382 = n500 | n20381 ;
  assign n20383 = n13288 | n18434 ;
  assign n20384 = n20382 | n20383 ;
  assign n20385 = n313 | n369 ;
  assign n20386 = n2188 | n20385 ;
  assign n20387 = n212 | n762 ;
  assign n20388 = n347 | n886 ;
  assign n20389 = n20387 | n20388 ;
  assign n20390 = n20386 | n20389 ;
  assign n20391 = n20384 | n20390 ;
  assign n20392 = n10772 | n15602 ;
  assign n20393 = n3431 | n20392 ;
  assign n20394 = n20391 | n20393 ;
  assign n20395 = n319 | n1785 ;
  assign n20396 = n1304 | n20395 ;
  assign n20397 = n460 | n20396 ;
  assign n20398 = n5017 | n20397 ;
  assign n20399 = n20394 | n20398 ;
  assign n20400 = n117 | n412 ;
  assign n20401 = n214 | n291 ;
  assign n20402 = n20400 | n20401 ;
  assign n20403 = n139 | n324 ;
  assign n20404 = n196 | n20403 ;
  assign n20405 = n20402 | n20404 ;
  assign n20406 = n20399 | n20405 ;
  assign n20407 = n20380 & ~n20406 ;
  assign n20408 = ~n20369 & n20407 ;
  assign n20409 = ( x29 & ~n20369 ) | ( x29 & n20407 ) | ( ~n20369 & n20407 ) ;
  assign n20410 = ~n20408 & n20409 ;
  assign n20411 = n20369 & ~n20407 ;
  assign n20412 = n20408 | n20411 ;
  assign n20413 = ~x29 & n20412 ;
  assign n20414 = n20410 | n20413 ;
  assign n20415 = n229 | n11747 ;
  assign n20416 = n1125 | n20415 ;
  assign n20417 = n811 | n995 ;
  assign n20418 = n20416 | n20417 ;
  assign n20419 = n6048 & ~n20418 ;
  assign n20420 = n259 | n7024 ;
  assign n20421 = n178 | n763 ;
  assign n20422 = n20420 | n20421 ;
  assign n20423 = n88 | n170 ;
  assign n20424 = n291 | n341 ;
  assign n20425 = n20423 | n20424 ;
  assign n20426 = n20422 | n20425 ;
  assign n20427 = ( n281 & n416 ) | ( n281 & ~n4334 ) | ( n416 & ~n4334 ) ;
  assign n20428 = n4334 | n20427 ;
  assign n20429 = n20426 | n20428 ;
  assign n20430 = n20419 & ~n20429 ;
  assign n20431 = n1418 | n10907 ;
  assign n20432 = n20430 & ~n20431 ;
  assign n20433 = ~n15600 & n20432 ;
  assign n20434 = n1301 | n3445 ;
  assign n20435 = n233 | n644 ;
  assign n20436 = n123 | n20435 ;
  assign n20437 = n20434 | n20436 ;
  assign n20438 = n206 | n208 ;
  assign n20439 = n858 | n20438 ;
  assign n20440 = n1114 | n20439 ;
  assign n20441 = n20437 | n20440 ;
  assign n20442 = n20433 & ~n20441 ;
  assign n20443 = n20407 & ~n20442 ;
  assign n20444 = ~n19558 & n20442 ;
  assign n20445 = n19554 & n20442 ;
  assign n20446 = ( n19555 & n20444 ) | ( n19555 & n20445 ) | ( n20444 & n20445 ) ;
  assign n20447 = n19558 & ~n20442 ;
  assign n20448 = n19554 | n20442 ;
  assign n20449 = ( n19555 & ~n20447 ) | ( n19555 & n20448 ) | ( ~n20447 & n20448 ) ;
  assign n20450 = ~n20446 & n20449 ;
  assign n20451 = n1057 & ~n8017 ;
  assign n20452 = n1060 & n7907 ;
  assign n20453 = ( n1060 & n7902 ) | ( n1060 & n20452 ) | ( n7902 & n20452 ) ;
  assign n20454 = n1065 & n8079 ;
  assign n20455 = ( n1065 & ~n8070 ) | ( n1065 & n20454 ) | ( ~n8070 & n20454 ) ;
  assign n20456 = n20453 | n20455 ;
  assign n20457 = n1062 | n20456 ;
  assign n20458 = n20451 | n20457 ;
  assign n20459 = n20446 | n20458 ;
  assign n20460 = ( n20446 & n20450 ) | ( n20446 & n20459 ) | ( n20450 & n20459 ) ;
  assign n20461 = ~n20407 & n20442 ;
  assign n20462 = n20443 | n20461 ;
  assign n20463 = ~n20443 & n20462 ;
  assign n20464 = ( n20443 & n20460 ) | ( n20443 & ~n20463 ) | ( n20460 & ~n20463 ) ;
  assign n20465 = n20414 & n20464 ;
  assign n20466 = n20451 | n20456 ;
  assign n20467 = n20446 | n20466 ;
  assign n20468 = ( n20446 & n20450 ) | ( n20446 & n20467 ) | ( n20450 & n20467 ) ;
  assign n20469 = ( n20443 & ~n20463 ) | ( n20443 & n20468 ) | ( ~n20463 & n20468 ) ;
  assign n20470 = n20414 & n20469 ;
  assign n20471 = ( n8104 & n20465 ) | ( n8104 & n20470 ) | ( n20465 & n20470 ) ;
  assign n20472 = n20414 | n20464 ;
  assign n20473 = n20414 | n20469 ;
  assign n20474 = ( n8104 & n20472 ) | ( n8104 & n20473 ) | ( n20472 & n20473 ) ;
  assign n20475 = ~n20471 & n20474 ;
  assign n20476 = n1057 & ~n8982 ;
  assign n20477 = ( n1057 & n9051 ) | ( n1057 & n20476 ) | ( n9051 & n20476 ) ;
  assign n20478 = n1065 & n9022 ;
  assign n20479 = n20477 | n20478 ;
  assign n20480 = n1065 | n20477 ;
  assign n20481 = ( ~n9019 & n20479 ) | ( ~n9019 & n20480 ) | ( n20479 & n20480 ) ;
  assign n20482 = n1060 | n20481 ;
  assign n20483 = ( ~n8017 & n20481 ) | ( ~n8017 & n20482 ) | ( n20481 & n20482 ) ;
  assign n20484 = n1062 | n20483 ;
  assign n20485 = ( ~n10242 & n20483 ) | ( ~n10242 & n20484 ) | ( n20483 & n20484 ) ;
  assign n20486 = n20475 & n20485 ;
  assign n20487 = n20475 | n20485 ;
  assign n20488 = ~n20486 & n20487 ;
  assign n20489 = n1821 & ~n9442 ;
  assign n20490 = n1821 & ~n9074 ;
  assign n20491 = ( n9440 & n20489 ) | ( n9440 & n20490 ) | ( n20489 & n20490 ) ;
  assign n20492 = n1826 & ~n8982 ;
  assign n20493 = ( n1826 & n9051 ) | ( n1826 & n20492 ) | ( n9051 & n20492 ) ;
  assign n20494 = n20491 | n20493 ;
  assign n20495 = n1821 | n20493 ;
  assign n20496 = ( ~n9442 & n20493 ) | ( ~n9442 & n20495 ) | ( n20493 & n20495 ) ;
  assign n20497 = ( ~n9072 & n20494 ) | ( ~n9072 & n20496 ) | ( n20494 & n20496 ) ;
  assign n20498 = ~x29 & n20494 ;
  assign n20499 = ~x29 & n20496 ;
  assign n20500 = ( ~n9072 & n20498 ) | ( ~n9072 & n20499 ) | ( n20498 & n20499 ) ;
  assign n20501 = x29 | n20498 ;
  assign n20502 = x29 | n20499 ;
  assign n20503 = ( ~n9072 & n20501 ) | ( ~n9072 & n20502 ) | ( n20501 & n20502 ) ;
  assign n20504 = ( ~n20497 & n20500 ) | ( ~n20497 & n20503 ) | ( n20500 & n20503 ) ;
  assign n20505 = n1060 & n8079 ;
  assign n20506 = ( n1060 & ~n8070 ) | ( n1060 & n20505 ) | ( ~n8070 & n20505 ) ;
  assign n20507 = n1065 | n20506 ;
  assign n20508 = ( ~n8017 & n20506 ) | ( ~n8017 & n20507 ) | ( n20506 & n20507 ) ;
  assign n20509 = n1057 & n9022 ;
  assign n20510 = ( n1057 & ~n9019 ) | ( n1057 & n20509 ) | ( ~n9019 & n20509 ) ;
  assign n20511 = n20508 | n20510 ;
  assign n20512 = n1062 | n20510 ;
  assign n20513 = n20508 | n20512 ;
  assign n20514 = ( ~n9416 & n20511 ) | ( ~n9416 & n20513 ) | ( n20511 & n20513 ) ;
  assign n20515 = n20504 & n20514 ;
  assign n20516 = n20504 & ~n20515 ;
  assign n20517 = ( n8104 & n20460 ) | ( n8104 & n20468 ) | ( n20460 & n20468 ) ;
  assign n20518 = ~n20462 & n20468 ;
  assign n20519 = n20460 & ~n20462 ;
  assign n20520 = ( n8104 & n20518 ) | ( n8104 & n20519 ) | ( n20518 & n20519 ) ;
  assign n20521 = n20517 & ~n20520 ;
  assign n20522 = n20461 | n20464 ;
  assign n20523 = n20461 | n20469 ;
  assign n20524 = ( n8104 & n20522 ) | ( n8104 & n20523 ) | ( n20522 & n20523 ) ;
  assign n20525 = ~n20521 & n20524 ;
  assign n20526 = ~n20504 & n20514 ;
  assign n20527 = ~n20525 & n20526 ;
  assign n20528 = ( n20516 & ~n20525 ) | ( n20516 & n20527 ) | ( ~n20525 & n20527 ) ;
  assign n20529 = n20488 & n20515 ;
  assign n20530 = ( n20488 & n20528 ) | ( n20488 & n20529 ) | ( n20528 & n20529 ) ;
  assign n20531 = n20488 | n20515 ;
  assign n20532 = n20528 | n20531 ;
  assign n20533 = ~n20530 & n20532 ;
  assign n20534 = ( n20504 & ~n20514 ) | ( n20504 & n20524 ) | ( ~n20514 & n20524 ) ;
  assign n20535 = n20504 & ~n20514 ;
  assign n20536 = ( ~n20521 & n20534 ) | ( ~n20521 & n20535 ) | ( n20534 & n20535 ) ;
  assign n20537 = ( ~n20504 & n20514 ) | ( ~n20504 & n20536 ) | ( n20514 & n20536 ) ;
  assign n20538 = ( ~n20525 & n20536 ) | ( ~n20525 & n20537 ) | ( n20536 & n20537 ) ;
  assign n20539 = ( n8104 & n20458 ) | ( n8104 & n20466 ) | ( n20458 & n20466 ) ;
  assign n20540 = n20450 & n20458 ;
  assign n20541 = n20450 & n20466 ;
  assign n20542 = ( n8104 & n20540 ) | ( n8104 & n20541 ) | ( n20540 & n20541 ) ;
  assign n20543 = n20450 & ~n20541 ;
  assign n20544 = n20450 & ~n20540 ;
  assign n20545 = ( ~n8104 & n20543 ) | ( ~n8104 & n20544 ) | ( n20543 & n20544 ) ;
  assign n20546 = ( n20539 & ~n20542 ) | ( n20539 & n20545 ) | ( ~n20542 & n20545 ) ;
  assign n20547 = n19563 | n19577 ;
  assign n20548 = ( n19563 & ~n19567 ) | ( n19563 & n20547 ) | ( ~n19567 & n20547 ) ;
  assign n20549 = n20546 & n20548 ;
  assign n20550 = n20546 | n20548 ;
  assign n20551 = ~n20549 & n20550 ;
  assign n20552 = n1823 & ~n8982 ;
  assign n20553 = ( n1823 & n9051 ) | ( n1823 & n20552 ) | ( n9051 & n20552 ) ;
  assign n20554 = n1826 & ~n9022 ;
  assign n20555 = ( n1826 & n20553 ) | ( n1826 & ~n20554 ) | ( n20553 & ~n20554 ) ;
  assign n20556 = n1826 | n20553 ;
  assign n20557 = ( ~n9019 & n20555 ) | ( ~n9019 & n20556 ) | ( n20555 & n20556 ) ;
  assign n20558 = n1821 | n20557 ;
  assign n20559 = ( n9078 & n20557 ) | ( n9078 & n20558 ) | ( n20557 & n20558 ) ;
  assign n20560 = x29 & n20558 ;
  assign n20561 = x29 & n20557 ;
  assign n20562 = ( n9078 & n20560 ) | ( n9078 & n20561 ) | ( n20560 & n20561 ) ;
  assign n20563 = x29 & ~n20560 ;
  assign n20564 = x29 & ~n20561 ;
  assign n20565 = ( ~n9078 & n20563 ) | ( ~n9078 & n20564 ) | ( n20563 & n20564 ) ;
  assign n20566 = ( n20559 & ~n20562 ) | ( n20559 & n20565 ) | ( ~n20562 & n20565 ) ;
  assign n20567 = n20549 | n20566 ;
  assign n20568 = ( n20549 & n20551 ) | ( n20549 & n20567 ) | ( n20551 & n20567 ) ;
  assign n20569 = ~n20538 & n20568 ;
  assign n20570 = n20538 & ~n20568 ;
  assign n20571 = n20569 | n20570 ;
  assign n20572 = n20551 & ~n20566 ;
  assign n20573 = n20551 | n20566 ;
  assign n20574 = ( ~n20551 & n20572 ) | ( ~n20551 & n20573 ) | ( n20572 & n20573 ) ;
  assign n20575 = n19583 & ~n19604 ;
  assign n20576 = ( n19583 & ~n19587 ) | ( n19583 & n20575 ) | ( ~n19587 & n20575 ) ;
  assign n20577 = n20574 & ~n20576 ;
  assign n20578 = ~n20574 & n20576 ;
  assign n20579 = n20577 | n20578 ;
  assign n20580 = n19611 & ~n20579 ;
  assign n20581 = n20577 | n20580 ;
  assign n20582 = ~n20571 & n20581 ;
  assign n20583 = n20569 | n20582 ;
  assign n20584 = n20533 & n20583 ;
  assign n20585 = ~n20577 & n20579 ;
  assign n20586 = n20571 | n20585 ;
  assign n20587 = ~n20569 & n20586 ;
  assign n20588 = n20533 & ~n20587 ;
  assign n20589 = ( n19619 & n20584 ) | ( n19619 & n20588 ) | ( n20584 & n20588 ) ;
  assign n20590 = n19611 | n19621 ;
  assign n20591 = ~n20579 & n20590 ;
  assign n20592 = n20577 | n20591 ;
  assign n20593 = ~n20571 & n20592 ;
  assign n20594 = n20569 | n20593 ;
  assign n20595 = n20533 & n20594 ;
  assign n20596 = n19611 | n19623 ;
  assign n20597 = ~n20579 & n20596 ;
  assign n20598 = n20577 | n20597 ;
  assign n20599 = ~n20571 & n20598 ;
  assign n20600 = n20569 | n20599 ;
  assign n20601 = n20533 & n20600 ;
  assign n20602 = ( n19345 & n20595 ) | ( n19345 & n20601 ) | ( n20595 & n20601 ) ;
  assign n20603 = ( n15882 & n20589 ) | ( n15882 & n20602 ) | ( n20589 & n20602 ) ;
  assign n20604 = ( n19619 & n20583 ) | ( n19619 & ~n20587 ) | ( n20583 & ~n20587 ) ;
  assign n20605 = n20533 | n20604 ;
  assign n20606 = ( n19345 & n20594 ) | ( n19345 & n20600 ) | ( n20594 & n20600 ) ;
  assign n20607 = n20533 | n20606 ;
  assign n20608 = ( n15882 & n20605 ) | ( n15882 & n20607 ) | ( n20605 & n20607 ) ;
  assign n20609 = ~n20603 & n20608 ;
  assign n20610 = ( n19619 & n20582 ) | ( n19619 & ~n20586 ) | ( n20582 & ~n20586 ) ;
  assign n20611 = ( n19345 & n20593 ) | ( n19345 & n20599 ) | ( n20593 & n20599 ) ;
  assign n20612 = ( n15882 & n20610 ) | ( n15882 & n20611 ) | ( n20610 & n20611 ) ;
  assign n20613 = ( n19619 & n20581 ) | ( n19619 & ~n20585 ) | ( n20581 & ~n20585 ) ;
  assign n20614 = n20571 & ~n20613 ;
  assign n20615 = ( n19345 & n20592 ) | ( n19345 & n20598 ) | ( n20592 & n20598 ) ;
  assign n20616 = n20571 & ~n20615 ;
  assign n20617 = ( ~n15882 & n20614 ) | ( ~n15882 & n20616 ) | ( n20614 & n20616 ) ;
  assign n20618 = n20612 | n20617 ;
  assign n20619 = ~n20609 & n20618 ;
  assign n20620 = n20609 & ~n20618 ;
  assign n20621 = n20619 | n20620 ;
  assign n20622 = ( n19619 & ~n20579 ) | ( n19619 & n20580 ) | ( ~n20579 & n20580 ) ;
  assign n20623 = ( n19345 & n20591 ) | ( n19345 & n20597 ) | ( n20591 & n20597 ) ;
  assign n20624 = ( n15882 & n20622 ) | ( n15882 & n20623 ) | ( n20622 & n20623 ) ;
  assign n20625 = n19611 | n19619 ;
  assign n20626 = n20579 & ~n20625 ;
  assign n20627 = ( n19345 & n20590 ) | ( n19345 & n20596 ) | ( n20590 & n20596 ) ;
  assign n20628 = n20579 & ~n20627 ;
  assign n20629 = ( ~n15882 & n20626 ) | ( ~n15882 & n20628 ) | ( n20626 & n20628 ) ;
  assign n20630 = n20624 | n20629 ;
  assign n20631 = n20618 | n20630 ;
  assign n20632 = n20618 & n20630 ;
  assign n20633 = n20631 & ~n20632 ;
  assign n20634 = n20631 & ~n20633 ;
  assign n20635 = n19631 & ~n20630 ;
  assign n20636 = ~n19631 & n20630 ;
  assign n20637 = n20635 | n20636 ;
  assign n20638 = n19650 & ~n20637 ;
  assign n20639 = n19648 & ~n20637 ;
  assign n20640 = n19632 & ~n20637 ;
  assign n20641 = ( n19503 & n20639 ) | ( n19503 & n20640 ) | ( n20639 & n20640 ) ;
  assign n20642 = ( n18577 & n20638 ) | ( n18577 & n20641 ) | ( n20638 & n20641 ) ;
  assign n20643 = n20635 | n20642 ;
  assign n20644 = ( n20631 & n20634 ) | ( n20631 & ~n20643 ) | ( n20634 & ~n20643 ) ;
  assign n20645 = n20638 | n20641 ;
  assign n20646 = n20635 | n20645 ;
  assign n20647 = ( n20631 & n20634 ) | ( n20631 & ~n20646 ) | ( n20634 & ~n20646 ) ;
  assign n20648 = ( ~n18604 & n20644 ) | ( ~n18604 & n20647 ) | ( n20644 & n20647 ) ;
  assign n20649 = n20621 & n20648 ;
  assign n20650 = n8122 & n20609 ;
  assign n20651 = n8115 & ~n20630 ;
  assign n20652 = n8118 & ~n20618 ;
  assign n20653 = n20651 | n20652 ;
  assign n20654 = n20650 | n20653 ;
  assign n20655 = n20621 | n20634 ;
  assign n20656 = n20621 | n20631 ;
  assign n20657 = ( ~n20643 & n20655 ) | ( ~n20643 & n20656 ) | ( n20655 & n20656 ) ;
  assign n20658 = ( ~n20646 & n20655 ) | ( ~n20646 & n20656 ) | ( n20655 & n20656 ) ;
  assign n20659 = ( ~n18604 & n20657 ) | ( ~n18604 & n20658 ) | ( n20657 & n20658 ) ;
  assign n20660 = n8125 | n20650 ;
  assign n20661 = n20653 | n20660 ;
  assign n20662 = ( n20654 & n20659 ) | ( n20654 & n20661 ) | ( n20659 & n20661 ) ;
  assign n20663 = n20654 & n20661 ;
  assign n20664 = ( ~n20649 & n20662 ) | ( ~n20649 & n20663 ) | ( n20662 & n20663 ) ;
  assign n20665 = x5 & n20664 ;
  assign n20666 = x5 & ~n20664 ;
  assign n20667 = ( n20664 & ~n20665 ) | ( n20664 & n20666 ) | ( ~n20665 & n20666 ) ;
  assign n20668 = n20345 & n20667 ;
  assign n20669 = ( n20344 & n20667 ) | ( n20344 & n20668 ) | ( n20667 & n20668 ) ;
  assign n20670 = n20346 & ~n20669 ;
  assign n20671 = ~n20345 & n20667 ;
  assign n20672 = ~n20344 & n20671 ;
  assign n20673 = n20670 | n20672 ;
  assign n20674 = n20308 & ~n20340 ;
  assign n20675 = n20308 & ~n20674 ;
  assign n20678 = n20633 & ~n20643 ;
  assign n20679 = n20633 & ~n20646 ;
  assign n20680 = ( ~n18604 & n20678 ) | ( ~n18604 & n20679 ) | ( n20678 & n20679 ) ;
  assign n20681 = n8125 & n20680 ;
  assign n20682 = n8122 & ~n20618 ;
  assign n20683 = n8115 & n19631 ;
  assign n20684 = n8118 & ~n20630 ;
  assign n20685 = n20683 | n20684 ;
  assign n20686 = n20682 | n20685 ;
  assign n20687 = ~n20633 & n20643 ;
  assign n20688 = ~n20633 & n20646 ;
  assign n20689 = ( n18604 & n20687 ) | ( n18604 & n20688 ) | ( n20687 & n20688 ) ;
  assign n20690 = n20686 | n20689 ;
  assign n20691 = n8125 | n20686 ;
  assign n20692 = ( n20681 & n20690 ) | ( n20681 & n20691 ) | ( n20690 & n20691 ) ;
  assign n20693 = x5 | n20692 ;
  assign n20694 = ~x5 & n20692 ;
  assign n20695 = ( ~n20692 & n20693 ) | ( ~n20692 & n20694 ) | ( n20693 & n20694 ) ;
  assign n20676 = n20308 | n20340 ;
  assign n20696 = ~n20676 & n20695 ;
  assign n20697 = ( n20675 & n20695 ) | ( n20675 & n20696 ) | ( n20695 & n20696 ) ;
  assign n20677 = ~n20675 & n20676 ;
  assign n20698 = n20677 | n20697 ;
  assign n20699 = n20676 & n20695 ;
  assign n20700 = ~n20675 & n20699 ;
  assign n20701 = n20698 & ~n20700 ;
  assign n20702 = n20303 & ~n20307 ;
  assign n20703 = n20306 | n20307 ;
  assign n20704 = ~n20702 & n20703 ;
  assign n20705 = ( n18604 & n20642 ) | ( n18604 & n20645 ) | ( n20642 & n20645 ) ;
  assign n20706 = ~n19654 & n20637 ;
  assign n20707 = ~n19651 & n20637 ;
  assign n20708 = ( ~n18604 & n20706 ) | ( ~n18604 & n20707 ) | ( n20706 & n20707 ) ;
  assign n20709 = n20705 | n20708 ;
  assign n20710 = n8122 & ~n20630 ;
  assign n20711 = n8115 & n19494 ;
  assign n20712 = n8118 & n19631 ;
  assign n20713 = n20711 | n20712 ;
  assign n20714 = n20710 | n20713 ;
  assign n20715 = n8125 | n20710 ;
  assign n20716 = n20713 | n20715 ;
  assign n20717 = ( ~n20709 & n20714 ) | ( ~n20709 & n20716 ) | ( n20714 & n20716 ) ;
  assign n20718 = ~x5 & n20716 ;
  assign n20719 = ~x5 & n20714 ;
  assign n20720 = ( ~n20709 & n20718 ) | ( ~n20709 & n20719 ) | ( n20718 & n20719 ) ;
  assign n20721 = x5 | n20719 ;
  assign n20722 = x5 | n20718 ;
  assign n20723 = ( ~n20709 & n20721 ) | ( ~n20709 & n20722 ) | ( n20721 & n20722 ) ;
  assign n20724 = ( ~n20717 & n20720 ) | ( ~n20717 & n20723 ) | ( n20720 & n20723 ) ;
  assign n20725 = ~n20704 & n20724 ;
  assign n20726 = n20704 | n20725 ;
  assign n20727 = n20704 & n20724 ;
  assign n20728 = n20726 & ~n20727 ;
  assign n20729 = n20298 & ~n20302 ;
  assign n20730 = n20301 & ~n20302 ;
  assign n20731 = n20729 | n20730 ;
  assign n20732 = n8122 & n19631 ;
  assign n20733 = n8115 & n19352 ;
  assign n20734 = n8118 & n19494 ;
  assign n20735 = n20733 | n20734 ;
  assign n20736 = n20732 | n20735 ;
  assign n20737 = n8125 & n19652 ;
  assign n20738 = n8125 & n19655 ;
  assign n20739 = ( ~n18604 & n20737 ) | ( ~n18604 & n20738 ) | ( n20737 & n20738 ) ;
  assign n20740 = n20736 | n20739 ;
  assign n20741 = n8125 | n20736 ;
  assign n20742 = ( n19640 & n20740 ) | ( n19640 & n20741 ) | ( n20740 & n20741 ) ;
  assign n20743 = x5 | n20742 ;
  assign n20744 = ~x5 & n20742 ;
  assign n20745 = ( ~n20742 & n20743 ) | ( ~n20742 & n20744 ) | ( n20743 & n20744 ) ;
  assign n20746 = n20731 & n20745 ;
  assign n20747 = n20731 & ~n20746 ;
  assign n20748 = ~n20731 & n20745 ;
  assign n20749 = n20747 | n20748 ;
  assign n20750 = n20293 & ~n20297 ;
  assign n20751 = n20296 | n20297 ;
  assign n20752 = ~n20750 & n20751 ;
  assign n20753 = n8122 & n19494 ;
  assign n20754 = n8115 & n18576 ;
  assign n20755 = n8118 & n19352 ;
  assign n20756 = n20754 | n20755 ;
  assign n20757 = n20753 | n20756 ;
  assign n20758 = n8125 | n20753 ;
  assign n20759 = n20756 | n20758 ;
  assign n20760 = ( n20320 & n20757 ) | ( n20320 & n20759 ) | ( n20757 & n20759 ) ;
  assign n20761 = x5 & n20759 ;
  assign n20762 = x5 & n20757 ;
  assign n20763 = ( n20320 & n20761 ) | ( n20320 & n20762 ) | ( n20761 & n20762 ) ;
  assign n20764 = x5 & ~n20762 ;
  assign n20765 = x5 & ~n20761 ;
  assign n20766 = ( ~n20320 & n20764 ) | ( ~n20320 & n20765 ) | ( n20764 & n20765 ) ;
  assign n20767 = ( n20760 & ~n20763 ) | ( n20760 & n20766 ) | ( ~n20763 & n20766 ) ;
  assign n20768 = ~n20752 & n20767 ;
  assign n20769 = n20752 | n20768 ;
  assign n20770 = n20752 & n20767 ;
  assign n20771 = n20769 & ~n20770 ;
  assign n20772 = n20291 & ~n20292 ;
  assign n20773 = n19752 | n20292 ;
  assign n20774 = ~n20772 & n20773 ;
  assign n20775 = n8122 & n19352 ;
  assign n20776 = n8115 & n18410 ;
  assign n20777 = n8118 & n18576 ;
  assign n20778 = n20776 | n20777 ;
  assign n20779 = n20775 | n20778 ;
  assign n20780 = n8125 | n20775 ;
  assign n20781 = n20778 | n20780 ;
  assign n20782 = ( n19674 & n20779 ) | ( n19674 & n20781 ) | ( n20779 & n20781 ) ;
  assign n20783 = x5 & n20781 ;
  assign n20784 = x5 & n20779 ;
  assign n20785 = ( n19674 & n20783 ) | ( n19674 & n20784 ) | ( n20783 & n20784 ) ;
  assign n20786 = x5 & ~n20784 ;
  assign n20787 = x5 & ~n20783 ;
  assign n20788 = ( ~n19674 & n20786 ) | ( ~n19674 & n20787 ) | ( n20786 & n20787 ) ;
  assign n20789 = ( n20782 & ~n20785 ) | ( n20782 & n20788 ) | ( ~n20785 & n20788 ) ;
  assign n20790 = ~n20774 & n20789 ;
  assign n20791 = n20774 | n20790 ;
  assign n20792 = n20774 & n20789 ;
  assign n20793 = n20791 & ~n20792 ;
  assign n20794 = n19792 | n20285 ;
  assign n20795 = ~n20286 & n20794 ;
  assign n20796 = n8122 & n18410 ;
  assign n20797 = n8115 & n18037 ;
  assign n20798 = n8118 & ~n18585 ;
  assign n20799 = n20797 | n20798 ;
  assign n20800 = n20796 | n20799 ;
  assign n20801 = n18586 & ~n20800 ;
  assign n20802 = ( n18609 & ~n20800 ) | ( n18609 & n20801 ) | ( ~n20800 & n20801 ) ;
  assign n20803 = ~n18650 & n20802 ;
  assign n20804 = n8125 | n20796 ;
  assign n20805 = n20799 | n20804 ;
  assign n20806 = ~n20803 & n20805 ;
  assign n20807 = x5 & n20805 ;
  assign n20808 = ~n20803 & n20807 ;
  assign n20809 = x5 & ~n20807 ;
  assign n20810 = ( x5 & n20803 ) | ( x5 & n20809 ) | ( n20803 & n20809 ) ;
  assign n20811 = ( n20806 & ~n20808 ) | ( n20806 & n20810 ) | ( ~n20808 & n20810 ) ;
  assign n20812 = n20795 & n20811 ;
  assign n20813 = n20287 & n20289 ;
  assign n20814 = n20287 | n20289 ;
  assign n20815 = ~n20813 & n20814 ;
  assign n20817 = n8115 & ~n18585 ;
  assign n20818 = n8118 & n18410 ;
  assign n20819 = n20817 | n20818 ;
  assign n20816 = n8122 & n18576 ;
  assign n20821 = n8125 | n20816 ;
  assign n20822 = n20819 | n20821 ;
  assign n20820 = n20816 | n20819 ;
  assign n20823 = n20820 & n20822 ;
  assign n20824 = ( n18612 & n20822 ) | ( n18612 & n20823 ) | ( n20822 & n20823 ) ;
  assign n20825 = x5 & n20823 ;
  assign n20826 = x5 & n20822 ;
  assign n20827 = ( n18612 & n20825 ) | ( n18612 & n20826 ) | ( n20825 & n20826 ) ;
  assign n20828 = x5 & ~n20825 ;
  assign n20829 = x5 & ~n20826 ;
  assign n20830 = ( ~n18612 & n20828 ) | ( ~n18612 & n20829 ) | ( n20828 & n20829 ) ;
  assign n20831 = ( n20824 & ~n20827 ) | ( n20824 & n20830 ) | ( ~n20827 & n20830 ) ;
  assign n20832 = n20815 & n20831 ;
  assign n20833 = n20815 | n20831 ;
  assign n20834 = ~n20832 & n20833 ;
  assign n20835 = n20812 & n20834 ;
  assign n20836 = n20832 | n20834 ;
  assign n20837 = n20795 & ~n20812 ;
  assign n20838 = ~n20795 & n20811 ;
  assign n20839 = n20837 | n20838 ;
  assign n20840 = n20281 & n20283 ;
  assign n20841 = n20281 | n20283 ;
  assign n20842 = ~n20840 & n20841 ;
  assign n20843 = n8122 & ~n18585 ;
  assign n20844 = n8115 & ~n17092 ;
  assign n20845 = n8118 & n18037 ;
  assign n20846 = n20844 | n20845 ;
  assign n20847 = n20843 | n20846 ;
  assign n20848 = n8125 & ~n18675 ;
  assign n20849 = ( n8125 & n18672 ) | ( n8125 & n20848 ) | ( n18672 & n20848 ) ;
  assign n20850 = n20847 | n20849 ;
  assign n20851 = x5 | n20847 ;
  assign n20852 = n20849 | n20851 ;
  assign n20853 = ~x5 & n20851 ;
  assign n20854 = ( ~x5 & n20849 ) | ( ~x5 & n20853 ) | ( n20849 & n20853 ) ;
  assign n20855 = ( ~n20850 & n20852 ) | ( ~n20850 & n20854 ) | ( n20852 & n20854 ) ;
  assign n20856 = n20842 & n20855 ;
  assign n20857 = ~n19831 & n20279 ;
  assign n20858 = n19831 & ~n20279 ;
  assign n20859 = n20857 | n20858 ;
  assign n20860 = n8122 & n18037 ;
  assign n20861 = n8115 & n17100 ;
  assign n20862 = n8118 & ~n17092 ;
  assign n20863 = n20861 | n20862 ;
  assign n20864 = n20860 | n20863 ;
  assign n20865 = n8125 | n20860 ;
  assign n20866 = n20863 | n20865 ;
  assign n20867 = ( ~n18050 & n20864 ) | ( ~n18050 & n20866 ) | ( n20864 & n20866 ) ;
  assign n20868 = ~x5 & n20866 ;
  assign n20869 = ~x5 & n20864 ;
  assign n20870 = ( ~n18050 & n20868 ) | ( ~n18050 & n20869 ) | ( n20868 & n20869 ) ;
  assign n20871 = x5 | n20869 ;
  assign n20872 = x5 | n20868 ;
  assign n20873 = ( ~n18050 & n20871 ) | ( ~n18050 & n20872 ) | ( n20871 & n20872 ) ;
  assign n20874 = ( ~n20867 & n20870 ) | ( ~n20867 & n20873 ) | ( n20870 & n20873 ) ;
  assign n20875 = n20859 & n20874 ;
  assign n20876 = n20859 | n20874 ;
  assign n20877 = ~n20875 & n20876 ;
  assign n20878 = ~n19852 & n20277 ;
  assign n20879 = n19852 & ~n20277 ;
  assign n20880 = n20878 | n20879 ;
  assign n20881 = n8122 & ~n17092 ;
  assign n20882 = n8115 & n17111 ;
  assign n20883 = n8118 & n17100 ;
  assign n20884 = n20882 | n20883 ;
  assign n20885 = n20881 | n20884 ;
  assign n20886 = n8125 | n20881 ;
  assign n20887 = n20884 | n20886 ;
  assign n20888 = ( ~n17134 & n20885 ) | ( ~n17134 & n20887 ) | ( n20885 & n20887 ) ;
  assign n20889 = ~x5 & n20887 ;
  assign n20890 = ~x5 & n20885 ;
  assign n20891 = ( ~n17134 & n20889 ) | ( ~n17134 & n20890 ) | ( n20889 & n20890 ) ;
  assign n20892 = x5 | n20890 ;
  assign n20893 = x5 | n20889 ;
  assign n20894 = ( ~n17134 & n20892 ) | ( ~n17134 & n20893 ) | ( n20892 & n20893 ) ;
  assign n20895 = ( ~n20888 & n20891 ) | ( ~n20888 & n20894 ) | ( n20891 & n20894 ) ;
  assign n20896 = n20880 & n20895 ;
  assign n20897 = n20880 | n20895 ;
  assign n20898 = ~n20896 & n20897 ;
  assign n20899 = n20273 & n20275 ;
  assign n20900 = n20273 | n20275 ;
  assign n20901 = ~n20899 & n20900 ;
  assign n20902 = n8115 & ~n16069 ;
  assign n20903 = n8118 & n17111 ;
  assign n20904 = n20902 | n20903 ;
  assign n20905 = n8122 & n17100 ;
  assign n20906 = n8125 | n20905 ;
  assign n20907 = n20904 | n20906 ;
  assign n20908 = n20904 | n20905 ;
  assign n20909 = n17169 | n20908 ;
  assign n20910 = ( ~n17129 & n20908 ) | ( ~n17129 & n20909 ) | ( n20908 & n20909 ) ;
  assign n20911 = n20907 & n20910 ;
  assign n20912 = ( n17161 & n20907 ) | ( n17161 & n20911 ) | ( n20907 & n20911 ) ;
  assign n20913 = ~x5 & n20912 ;
  assign n20914 = x5 | n20912 ;
  assign n20915 = ( ~n20912 & n20913 ) | ( ~n20912 & n20914 ) | ( n20913 & n20914 ) ;
  assign n20916 = n20901 & n20915 ;
  assign n20917 = n19894 & n20271 ;
  assign n20918 = n19894 | n20271 ;
  assign n20919 = ~n20917 & n20918 ;
  assign n20920 = n8115 & n15886 ;
  assign n20921 = n8118 & ~n16069 ;
  assign n20922 = n20920 | n20921 ;
  assign n20923 = n8122 & n17111 ;
  assign n20924 = n8125 | n20923 ;
  assign n20925 = n20922 | n20924 ;
  assign n20926 = n20922 | n20923 ;
  assign n20927 = n17194 & ~n20926 ;
  assign n20928 = ( n17129 & ~n20926 ) | ( n17129 & n20927 ) | ( ~n20926 & n20927 ) ;
  assign n20929 = n20925 & ~n20928 ;
  assign n20930 = ( n17186 & n20925 ) | ( n17186 & n20929 ) | ( n20925 & n20929 ) ;
  assign n20931 = x5 & n20930 ;
  assign n20932 = x5 & ~n20930 ;
  assign n20933 = ( n20930 & ~n20931 ) | ( n20930 & n20932 ) | ( ~n20931 & n20932 ) ;
  assign n20934 = n20919 & n20933 ;
  assign n20935 = n20919 & ~n20934 ;
  assign n20936 = ~n20919 & n20933 ;
  assign n20937 = n20935 | n20936 ;
  assign n20938 = n19916 & n20269 ;
  assign n20939 = n19916 | n20269 ;
  assign n20940 = ~n20938 & n20939 ;
  assign n20941 = n8122 & ~n16069 ;
  assign n20942 = n8115 & ~n16085 ;
  assign n20943 = n8118 & n15886 ;
  assign n20944 = n20942 | n20943 ;
  assign n20945 = n20941 | n20944 ;
  assign n20946 = n8125 | n20945 ;
  assign n20947 = ( ~n16107 & n20945 ) | ( ~n16107 & n20946 ) | ( n20945 & n20946 ) ;
  assign n20948 = ~x5 & n20946 ;
  assign n20949 = ~x5 & n20945 ;
  assign n20950 = ( ~n16107 & n20948 ) | ( ~n16107 & n20949 ) | ( n20948 & n20949 ) ;
  assign n20951 = x5 | n20948 ;
  assign n20952 = x5 | n20949 ;
  assign n20953 = ( ~n16107 & n20951 ) | ( ~n16107 & n20952 ) | ( n20951 & n20952 ) ;
  assign n20954 = ( ~n20947 & n20950 ) | ( ~n20947 & n20953 ) | ( n20950 & n20953 ) ;
  assign n20955 = n20940 & n20954 ;
  assign n20956 = n20940 & ~n20955 ;
  assign n20957 = ~n20940 & n20954 ;
  assign n20958 = n20956 | n20957 ;
  assign n20959 = ( n19958 & n19959 ) | ( n19958 & n20267 ) | ( n19959 & n20267 ) ;
  assign n20960 = n19936 | n19958 ;
  assign n20961 = n20267 | n20960 ;
  assign n20962 = ~n20959 & n20961 ;
  assign n20963 = n8122 & n15886 ;
  assign n20964 = n8115 & n15434 ;
  assign n20965 = n8118 & ~n16085 ;
  assign n20966 = n20964 | n20965 ;
  assign n20967 = n20963 | n20966 ;
  assign n20968 = n8125 | n20963 ;
  assign n20969 = n20966 | n20968 ;
  assign n20970 = ( ~n16140 & n20967 ) | ( ~n16140 & n20969 ) | ( n20967 & n20969 ) ;
  assign n20971 = ~x5 & n20969 ;
  assign n20972 = ~x5 & n20967 ;
  assign n20973 = ( ~n16140 & n20971 ) | ( ~n16140 & n20972 ) | ( n20971 & n20972 ) ;
  assign n20974 = x5 | n20972 ;
  assign n20975 = x5 | n20971 ;
  assign n20976 = ( ~n16140 & n20974 ) | ( ~n16140 & n20975 ) | ( n20974 & n20975 ) ;
  assign n20977 = ( ~n20970 & n20973 ) | ( ~n20970 & n20976 ) | ( n20973 & n20976 ) ;
  assign n20978 = n20962 & n20977 ;
  assign n20979 = n20263 & ~n20267 ;
  assign n20980 = n20266 & ~n20267 ;
  assign n20981 = n20979 | n20980 ;
  assign n20982 = n8122 & ~n16085 ;
  assign n20983 = n8115 & n14591 ;
  assign n20984 = n8118 & n15434 ;
  assign n20985 = n20983 | n20984 ;
  assign n20986 = n20982 | n20985 ;
  assign n20987 = n8125 | n20982 ;
  assign n20988 = n20985 | n20987 ;
  assign n20989 = ( ~n16167 & n20986 ) | ( ~n16167 & n20988 ) | ( n20986 & n20988 ) ;
  assign n20990 = ~x5 & n20988 ;
  assign n20991 = ~x5 & n20986 ;
  assign n20992 = ( ~n16167 & n20990 ) | ( ~n16167 & n20991 ) | ( n20990 & n20991 ) ;
  assign n20993 = x5 | n20991 ;
  assign n20994 = x5 | n20990 ;
  assign n20995 = ( ~n16167 & n20993 ) | ( ~n16167 & n20994 ) | ( n20993 & n20994 ) ;
  assign n20996 = ( ~n20989 & n20992 ) | ( ~n20989 & n20995 ) | ( n20992 & n20995 ) ;
  assign n20997 = n20981 & n20996 ;
  assign n20998 = n20981 & ~n20997 ;
  assign n20999 = ~n20981 & n20996 ;
  assign n21000 = n20998 | n20999 ;
  assign n21001 = n20261 & ~n20262 ;
  assign n21002 = n19982 & ~n20262 ;
  assign n21003 = n21001 | n21002 ;
  assign n21004 = n8122 & n15434 ;
  assign n21005 = n8115 & n14329 ;
  assign n21006 = n8118 & n14591 ;
  assign n21007 = n21005 | n21006 ;
  assign n21008 = n21004 | n21007 ;
  assign n21009 = n8125 | n21004 ;
  assign n21010 = n21007 | n21009 ;
  assign n21011 = ( n15453 & n21008 ) | ( n15453 & n21010 ) | ( n21008 & n21010 ) ;
  assign n21012 = x5 & n21010 ;
  assign n21013 = x5 & n21008 ;
  assign n21014 = ( n15453 & n21012 ) | ( n15453 & n21013 ) | ( n21012 & n21013 ) ;
  assign n21015 = x5 & ~n21013 ;
  assign n21016 = x5 & ~n21012 ;
  assign n21017 = ( ~n15453 & n21015 ) | ( ~n15453 & n21016 ) | ( n21015 & n21016 ) ;
  assign n21018 = ( n21011 & ~n21014 ) | ( n21011 & n21017 ) | ( ~n21014 & n21017 ) ;
  assign n21019 = n21003 & n21018 ;
  assign n21020 = n21003 & ~n21019 ;
  assign n21021 = ~n21003 & n21018 ;
  assign n21022 = n21020 | n21021 ;
  assign n21023 = n20253 | n20254 ;
  assign n21024 = n20020 | n21023 ;
  assign n21025 = ~n20256 & n21024 ;
  assign n21027 = n8115 & n13522 ;
  assign n21028 = n8118 & n14607 ;
  assign n21029 = n21027 | n21028 ;
  assign n21026 = n8122 & n14329 ;
  assign n21031 = n8125 | n21026 ;
  assign n21032 = n21029 | n21031 ;
  assign n21030 = n21026 | n21029 ;
  assign n21033 = n21030 & n21032 ;
  assign n21034 = ( n14656 & n21032 ) | ( n14656 & n21033 ) | ( n21032 & n21033 ) ;
  assign n21035 = x5 & n21033 ;
  assign n21036 = x5 & n21032 ;
  assign n21037 = ( n14656 & n21035 ) | ( n14656 & n21036 ) | ( n21035 & n21036 ) ;
  assign n21038 = x5 & ~n21035 ;
  assign n21039 = x5 & ~n21036 ;
  assign n21040 = ( ~n14656 & n21038 ) | ( ~n14656 & n21039 ) | ( n21038 & n21039 ) ;
  assign n21041 = ( n21034 & ~n21037 ) | ( n21034 & n21040 ) | ( ~n21037 & n21040 ) ;
  assign n21042 = n21025 & n21041 ;
  assign n21043 = n20257 & n20259 ;
  assign n21044 = n20257 | n20259 ;
  assign n21045 = ~n21043 & n21044 ;
  assign n21047 = n8115 & n14607 ;
  assign n21048 = n8118 & n14329 ;
  assign n21049 = n21047 | n21048 ;
  assign n21046 = n8122 & n14591 ;
  assign n21051 = n8125 | n21046 ;
  assign n21052 = n21049 | n21051 ;
  assign n21050 = n21046 | n21049 ;
  assign n21053 = n21050 & n21052 ;
  assign n21054 = ( n14629 & n21052 ) | ( n14629 & n21053 ) | ( n21052 & n21053 ) ;
  assign n21055 = x5 & n21053 ;
  assign n21056 = x5 & n21052 ;
  assign n21057 = ( n14629 & n21055 ) | ( n14629 & n21056 ) | ( n21055 & n21056 ) ;
  assign n21058 = x5 & ~n21055 ;
  assign n21059 = x5 & ~n21056 ;
  assign n21060 = ( ~n14629 & n21058 ) | ( ~n14629 & n21059 ) | ( n21058 & n21059 ) ;
  assign n21061 = ( n21054 & ~n21057 ) | ( n21054 & n21060 ) | ( ~n21057 & n21060 ) ;
  assign n21062 = n21045 & n21061 ;
  assign n21063 = n21045 | n21061 ;
  assign n21064 = ~n21062 & n21063 ;
  assign n21065 = n21042 & n21064 ;
  assign n21066 = n21062 | n21064 ;
  assign n21067 = n20249 & n20251 ;
  assign n21068 = n20249 | n20251 ;
  assign n21069 = ~n21067 & n21068 ;
  assign n21070 = n8115 & n13235 ;
  assign n21071 = n8118 & n13522 ;
  assign n21072 = n21070 | n21071 ;
  assign n21073 = n8122 & n14607 ;
  assign n21074 = n8125 | n21073 ;
  assign n21075 = n21072 | n21074 ;
  assign n21076 = n21072 | n21073 ;
  assign n21077 = n14696 | n21076 ;
  assign n21078 = n14698 | n21076 ;
  assign n21079 = ( ~n13248 & n21077 ) | ( ~n13248 & n21078 ) | ( n21077 & n21078 ) ;
  assign n21080 = n21075 & n21079 ;
  assign n21081 = ( n14687 & n21075 ) | ( n14687 & n21080 ) | ( n21075 & n21080 ) ;
  assign n21082 = ~x5 & n21081 ;
  assign n21083 = x5 | n21081 ;
  assign n21084 = ( ~n21081 & n21082 ) | ( ~n21081 & n21083 ) | ( n21082 & n21083 ) ;
  assign n21085 = n21069 & n21084 ;
  assign n21086 = n21069 & ~n21085 ;
  assign n21087 = ~n21069 & n21084 ;
  assign n21088 = n21086 | n21087 ;
  assign n21089 = n20245 & n20247 ;
  assign n21090 = n20245 | n20247 ;
  assign n21091 = ~n21089 & n21090 ;
  assign n21092 = n8122 & n13522 ;
  assign n21093 = n8115 & n12936 ;
  assign n21094 = n8118 & n13235 ;
  assign n21095 = n21093 | n21094 ;
  assign n21096 = n21092 | n21095 ;
  assign n21097 = n8125 & n13537 ;
  assign n21098 = n8125 & n13539 ;
  assign n21099 = ( ~n13248 & n21097 ) | ( ~n13248 & n21098 ) | ( n21097 & n21098 ) ;
  assign n21100 = n21096 | n21099 ;
  assign n21101 = n8125 | n21096 ;
  assign n21102 = ( n13530 & n21100 ) | ( n13530 & n21101 ) | ( n21100 & n21101 ) ;
  assign n21103 = x5 | n21102 ;
  assign n21104 = ~x5 & n21102 ;
  assign n21105 = ( ~n21102 & n21103 ) | ( ~n21102 & n21104 ) | ( n21103 & n21104 ) ;
  assign n21106 = n21091 & n21105 ;
  assign n21107 = n20243 & ~n20244 ;
  assign n21108 = n20079 & ~n20244 ;
  assign n21109 = n21107 | n21108 ;
  assign n21110 = n8122 & n13235 ;
  assign n21111 = n8115 & ~n12616 ;
  assign n21112 = n8118 & n12936 ;
  assign n21113 = n21111 | n21112 ;
  assign n21114 = n21110 | n21113 ;
  assign n21115 = n8125 | n21110 ;
  assign n21116 = n21113 | n21115 ;
  assign n21117 = ( n13561 & n21114 ) | ( n13561 & n21116 ) | ( n21114 & n21116 ) ;
  assign n21118 = x5 & n21116 ;
  assign n21119 = x5 & n21114 ;
  assign n21120 = ( n13561 & n21118 ) | ( n13561 & n21119 ) | ( n21118 & n21119 ) ;
  assign n21121 = x5 & ~n21119 ;
  assign n21122 = x5 & ~n21118 ;
  assign n21123 = ( ~n13561 & n21121 ) | ( ~n13561 & n21122 ) | ( n21121 & n21122 ) ;
  assign n21124 = ( n21117 & ~n21120 ) | ( n21117 & n21123 ) | ( ~n21120 & n21123 ) ;
  assign n21125 = n21109 & n21124 ;
  assign n21126 = n21109 & ~n21125 ;
  assign n21127 = ~n20099 & n20241 ;
  assign n21128 = n20099 & ~n20241 ;
  assign n21129 = n21127 | n21128 ;
  assign n21130 = n8122 & n12936 ;
  assign n21131 = n8115 & n12010 ;
  assign n21132 = n8118 & ~n12616 ;
  assign n21133 = n21131 | n21132 ;
  assign n21134 = n21130 | n21133 ;
  assign n21135 = n8125 | n21130 ;
  assign n21136 = n21133 | n21135 ;
  assign n21137 = ( ~n13591 & n21134 ) | ( ~n13591 & n21136 ) | ( n21134 & n21136 ) ;
  assign n21138 = ~x5 & n21136 ;
  assign n21139 = ~x5 & n21134 ;
  assign n21140 = ( ~n13591 & n21138 ) | ( ~n13591 & n21139 ) | ( n21138 & n21139 ) ;
  assign n21141 = x5 | n21139 ;
  assign n21142 = x5 | n21138 ;
  assign n21143 = ( ~n13591 & n21141 ) | ( ~n13591 & n21142 ) | ( n21141 & n21142 ) ;
  assign n21144 = ( ~n21137 & n21140 ) | ( ~n21137 & n21143 ) | ( n21140 & n21143 ) ;
  assign n21145 = n21129 & n21144 ;
  assign n21146 = n20237 & n20239 ;
  assign n21147 = n20237 | n20239 ;
  assign n21148 = ~n21146 & n21147 ;
  assign n21150 = n8115 & ~n11663 ;
  assign n21151 = n8118 & n12010 ;
  assign n21152 = n21150 | n21151 ;
  assign n21149 = n8122 & ~n12616 ;
  assign n21154 = n8125 | n21149 ;
  assign n21155 = n21152 | n21154 ;
  assign n21153 = n21149 | n21152 ;
  assign n21156 = n21153 & n21155 ;
  assign n21157 = ( ~n12626 & n21155 ) | ( ~n12626 & n21156 ) | ( n21155 & n21156 ) ;
  assign n21158 = ~x5 & n21156 ;
  assign n21159 = ~x5 & n21155 ;
  assign n21160 = ( ~n12626 & n21158 ) | ( ~n12626 & n21159 ) | ( n21158 & n21159 ) ;
  assign n21161 = x5 | n21158 ;
  assign n21162 = x5 | n21159 ;
  assign n21163 = ( ~n12626 & n21161 ) | ( ~n12626 & n21162 ) | ( n21161 & n21162 ) ;
  assign n21164 = ( ~n21157 & n21160 ) | ( ~n21157 & n21163 ) | ( n21160 & n21163 ) ;
  assign n21165 = n21148 & n21164 ;
  assign n21166 = n20138 | n20235 ;
  assign n21167 = ~n20236 & n21166 ;
  assign n21169 = n8115 & n11363 ;
  assign n21170 = n8118 & ~n11663 ;
  assign n21171 = n21169 | n21170 ;
  assign n21168 = n8122 & n12010 ;
  assign n21173 = n8125 | n21168 ;
  assign n21174 = n21171 | n21173 ;
  assign n21172 = n21168 | n21171 ;
  assign n21175 = n21172 & n21174 ;
  assign n21176 = ( ~n12028 & n21174 ) | ( ~n12028 & n21175 ) | ( n21174 & n21175 ) ;
  assign n21177 = n21174 | n21175 ;
  assign n21178 = ( n12017 & n21176 ) | ( n12017 & n21177 ) | ( n21176 & n21177 ) ;
  assign n21179 = ~x5 & n21178 ;
  assign n21180 = x5 | n21178 ;
  assign n21181 = ( ~n21178 & n21179 ) | ( ~n21178 & n21180 ) | ( n21179 & n21180 ) ;
  assign n21182 = n21167 & n21181 ;
  assign n21183 = n21167 & ~n21182 ;
  assign n21184 = ~n21167 & n21181 ;
  assign n21185 = n21183 | n21184 ;
  assign n21186 = n20162 | n20233 ;
  assign n21187 = ~n20234 & n21186 ;
  assign n21188 = n8115 & n10649 ;
  assign n21189 = n8118 & n11363 ;
  assign n21190 = n21188 | n21189 ;
  assign n21191 = n8122 & ~n11663 ;
  assign n21192 = n8125 | n21191 ;
  assign n21193 = n21190 | n21192 ;
  assign n21194 = n21190 | n21191 ;
  assign n21195 = n12048 & ~n21194 ;
  assign n21196 = ( n11672 & ~n21194 ) | ( n11672 & n21195 ) | ( ~n21194 & n21195 ) ;
  assign n21197 = n21193 & ~n21196 ;
  assign n21198 = ( n12040 & n21193 ) | ( n12040 & n21197 ) | ( n21193 & n21197 ) ;
  assign n21199 = x5 & n21198 ;
  assign n21200 = x5 & ~n21198 ;
  assign n21201 = ( n21198 & ~n21199 ) | ( n21198 & n21200 ) | ( ~n21199 & n21200 ) ;
  assign n21202 = n21187 & n21201 ;
  assign n21203 = n21187 & ~n21202 ;
  assign n21204 = ~n21187 & n21201 ;
  assign n21205 = n21203 | n21204 ;
  assign n21206 = n20229 & n20231 ;
  assign n21207 = n20229 | n20231 ;
  assign n21208 = ~n21206 & n21207 ;
  assign n21209 = n8122 & n11363 ;
  assign n21210 = n8115 & n10325 ;
  assign n21211 = n8118 & n10649 ;
  assign n21212 = n21210 | n21211 ;
  assign n21213 = n21209 | n21212 ;
  assign n21214 = n8125 | n21213 ;
  assign n21215 = ( n12059 & n21213 ) | ( n12059 & n21214 ) | ( n21213 & n21214 ) ;
  assign n21216 = x5 & n21214 ;
  assign n21217 = x5 & n21213 ;
  assign n21218 = ( n12059 & n21216 ) | ( n12059 & n21217 ) | ( n21216 & n21217 ) ;
  assign n21219 = x5 & ~n21216 ;
  assign n21220 = x5 & ~n21217 ;
  assign n21221 = ( ~n12059 & n21219 ) | ( ~n12059 & n21220 ) | ( n21219 & n21220 ) ;
  assign n21222 = ( n21215 & ~n21218 ) | ( n21215 & n21221 ) | ( ~n21218 & n21221 ) ;
  assign n21223 = n21208 & n21222 ;
  assign n21224 = n20216 & n20227 ;
  assign n21225 = n20216 & ~n21224 ;
  assign n21226 = n8122 & n10649 ;
  assign n21227 = n8115 & n10654 ;
  assign n21228 = n8118 & n10325 ;
  assign n21229 = n21227 | n21228 ;
  assign n21230 = n21226 | n21229 ;
  assign n21231 = n8125 | n21226 ;
  assign n21232 = n21229 | n21231 ;
  assign n21233 = ( n10702 & n21230 ) | ( n10702 & n21232 ) | ( n21230 & n21232 ) ;
  assign n21234 = n21230 | n21232 ;
  assign n21235 = ( n10695 & n21233 ) | ( n10695 & n21234 ) | ( n21233 & n21234 ) ;
  assign n21236 = x5 & n21235 ;
  assign n21237 = x5 & ~n21235 ;
  assign n21238 = ( n21235 & ~n21236 ) | ( n21235 & n21237 ) | ( ~n21236 & n21237 ) ;
  assign n21239 = ~n20216 & n20227 ;
  assign n21240 = n21238 & n21239 ;
  assign n21241 = ( n21225 & n21238 ) | ( n21225 & n21240 ) | ( n21238 & n21240 ) ;
  assign n21242 = n21238 | n21239 ;
  assign n21243 = n21225 | n21242 ;
  assign n21244 = ~n21241 & n21243 ;
  assign n21245 = n8122 & n10325 ;
  assign n21246 = n8115 & ~n10662 ;
  assign n21247 = n8118 & n10654 ;
  assign n21248 = n21246 | n21247 ;
  assign n21249 = n21245 | n21248 ;
  assign n21250 = n8125 | n21249 ;
  assign n21251 = ( ~n10957 & n21249 ) | ( ~n10957 & n21250 ) | ( n21249 & n21250 ) ;
  assign n21252 = n21249 | n21250 ;
  assign n21253 = ( n10949 & n21251 ) | ( n10949 & n21252 ) | ( n21251 & n21252 ) ;
  assign n21254 = ~x5 & n21253 ;
  assign n21255 = x5 & n21249 ;
  assign n21256 = x5 & n8125 ;
  assign n21257 = ( x5 & n21249 ) | ( x5 & n21256 ) | ( n21249 & n21256 ) ;
  assign n21258 = ( ~n10957 & n21255 ) | ( ~n10957 & n21257 ) | ( n21255 & n21257 ) ;
  assign n21259 = n21255 | n21257 ;
  assign n21260 = ( n10949 & n21258 ) | ( n10949 & n21259 ) | ( n21258 & n21259 ) ;
  assign n21261 = x5 & ~n21260 ;
  assign n21262 = n21254 | n21261 ;
  assign n21263 = n20195 & n20213 ;
  assign n21264 = n20195 | n20213 ;
  assign n21265 = ~n21263 & n21264 ;
  assign n21266 = n21262 & n21265 ;
  assign n21267 = n21262 | n21265 ;
  assign n21268 = ~n21266 & n21267 ;
  assign n21269 = n20188 | n20191 ;
  assign n21270 = ~n20191 & n20193 ;
  assign n21271 = ( n20189 & n21269 ) | ( n20189 & ~n21270 ) | ( n21269 & ~n21270 ) ;
  assign n21272 = ~n20195 & n21271 ;
  assign n21273 = n8122 & n10654 ;
  assign n21274 = n8115 & n10667 ;
  assign n21275 = n8118 & ~n10662 ;
  assign n21276 = n21274 | n21275 ;
  assign n21277 = n21273 | n21276 ;
  assign n21278 = n8125 | n21273 ;
  assign n21279 = n21276 | n21278 ;
  assign n21280 = ( n10978 & n21277 ) | ( n10978 & n21279 ) | ( n21277 & n21279 ) ;
  assign n21281 = x5 & n21279 ;
  assign n21282 = x5 & n21277 ;
  assign n21283 = ( n10978 & n21281 ) | ( n10978 & n21282 ) | ( n21281 & n21282 ) ;
  assign n21284 = x5 & ~n21282 ;
  assign n21285 = x5 & ~n21281 ;
  assign n21286 = ( ~n10978 & n21284 ) | ( ~n10978 & n21285 ) | ( n21284 & n21285 ) ;
  assign n21287 = ( n21280 & ~n21283 ) | ( n21280 & n21286 ) | ( ~n21283 & n21286 ) ;
  assign n21288 = n21272 & n21287 ;
  assign n21289 = n8125 & n10784 ;
  assign n21290 = n8118 & ~n10678 ;
  assign n21291 = n8122 & ~n10675 ;
  assign n21292 = n21290 | n21291 ;
  assign n21293 = x5 | n21292 ;
  assign n21294 = n21289 | n21293 ;
  assign n21295 = ~x5 & n21294 ;
  assign n21296 = x5 & ~n8113 ;
  assign n21297 = ( x5 & n10678 ) | ( x5 & n21296 ) | ( n10678 & n21296 ) ;
  assign n21298 = n21294 & n21297 ;
  assign n21299 = n21289 | n21292 ;
  assign n21300 = n21297 & ~n21299 ;
  assign n21301 = ( n21295 & n21298 ) | ( n21295 & n21300 ) | ( n21298 & n21300 ) ;
  assign n21302 = n8122 & n10667 ;
  assign n21303 = n8115 & ~n10678 ;
  assign n21304 = n8118 & ~n10675 ;
  assign n21305 = n21303 | n21304 ;
  assign n21306 = n21302 | n21305 ;
  assign n21307 = n10837 | n21306 ;
  assign n21308 = n8125 | n21302 ;
  assign n21309 = n21305 | n21308 ;
  assign n21310 = ~x5 & n21309 ;
  assign n21311 = n21307 & n21310 ;
  assign n21312 = x5 | n21311 ;
  assign n21313 = n7067 & ~n10678 ;
  assign n21314 = n21311 & n21313 ;
  assign n21315 = n21307 & n21309 ;
  assign n21316 = n21313 & ~n21315 ;
  assign n21317 = ( n21312 & n21314 ) | ( n21312 & n21316 ) | ( n21314 & n21316 ) ;
  assign n21318 = n21301 & n21317 ;
  assign n21319 = ( n21311 & n21312 ) | ( n21311 & ~n21315 ) | ( n21312 & ~n21315 ) ;
  assign n21320 = n21301 | n21313 ;
  assign n21321 = ( n21313 & n21319 ) | ( n21313 & n21320 ) | ( n21319 & n21320 ) ;
  assign n21322 = ~n21318 & n21321 ;
  assign n21323 = n8122 & ~n10662 ;
  assign n21324 = n8115 & ~n10675 ;
  assign n21325 = n8118 & n10667 ;
  assign n21326 = n21324 | n21325 ;
  assign n21327 = n21323 | n21326 ;
  assign n21328 = ( n8125 & n10850 ) | ( n8125 & n21327 ) | ( n10850 & n21327 ) ;
  assign n21329 = ( x5 & n8125 ) | ( x5 & ~n21327 ) | ( n8125 & ~n21327 ) ;
  assign n21330 = ( x5 & n10850 ) | ( x5 & n21329 ) | ( n10850 & n21329 ) ;
  assign n21331 = ~n21328 & n21330 ;
  assign n21332 = n21327 | n21330 ;
  assign n21333 = ( ~x5 & n21331 ) | ( ~x5 & n21332 ) | ( n21331 & n21332 ) ;
  assign n21334 = n21318 | n21333 ;
  assign n21335 = ( n21318 & n21322 ) | ( n21318 & n21334 ) | ( n21322 & n21334 ) ;
  assign n21336 = n21272 | n21287 ;
  assign n21337 = ~n21288 & n21336 ;
  assign n21338 = n21288 | n21337 ;
  assign n21339 = ( n21288 & n21335 ) | ( n21288 & n21338 ) | ( n21335 & n21338 ) ;
  assign n21340 = n21268 & n21339 ;
  assign n21341 = n21266 | n21340 ;
  assign n21342 = n21244 & n21341 ;
  assign n21343 = n21241 | n21342 ;
  assign n21344 = ~n21208 & n21222 ;
  assign n21345 = ( n21208 & ~n21223 ) | ( n21208 & n21344 ) | ( ~n21223 & n21344 ) ;
  assign n21346 = n21223 | n21345 ;
  assign n21347 = ( n21223 & n21343 ) | ( n21223 & n21346 ) | ( n21343 & n21346 ) ;
  assign n21348 = n21205 & n21347 ;
  assign n21349 = n21202 | n21348 ;
  assign n21350 = n21185 & n21349 ;
  assign n21351 = n21182 | n21350 ;
  assign n21352 = n21148 | n21164 ;
  assign n21353 = ~n21165 & n21352 ;
  assign n21354 = n21165 | n21353 ;
  assign n21355 = ( n21165 & n21351 ) | ( n21165 & n21354 ) | ( n21351 & n21354 ) ;
  assign n21356 = n21129 | n21144 ;
  assign n21357 = ~n21145 & n21356 ;
  assign n21358 = n21145 | n21357 ;
  assign n21359 = ( n21145 & n21355 ) | ( n21145 & n21358 ) | ( n21355 & n21358 ) ;
  assign n21360 = ~n21109 & n21124 ;
  assign n21361 = n21359 & n21360 ;
  assign n21362 = ( n21126 & n21359 ) | ( n21126 & n21361 ) | ( n21359 & n21361 ) ;
  assign n21363 = n21125 | n21362 ;
  assign n21364 = ~n21091 & n21105 ;
  assign n21365 = ( n21091 & ~n21106 ) | ( n21091 & n21364 ) | ( ~n21106 & n21364 ) ;
  assign n21366 = n21106 | n21365 ;
  assign n21367 = ( n21106 & n21363 ) | ( n21106 & n21366 ) | ( n21363 & n21366 ) ;
  assign n21368 = n21088 & n21367 ;
  assign n21369 = n21085 | n21368 ;
  assign n21370 = n21025 & ~n21042 ;
  assign n21371 = ~n21025 & n21041 ;
  assign n21372 = n21370 | n21371 ;
  assign n21373 = n21369 & n21372 ;
  assign n21374 = n21062 | n21373 ;
  assign n21375 = ( n21065 & n21066 ) | ( n21065 & n21374 ) | ( n21066 & n21374 ) ;
  assign n21376 = n21019 | n21375 ;
  assign n21377 = ( n21019 & n21022 ) | ( n21019 & n21376 ) | ( n21022 & n21376 ) ;
  assign n21378 = n20997 | n21377 ;
  assign n21379 = ( n20997 & n21000 ) | ( n20997 & n21378 ) | ( n21000 & n21378 ) ;
  assign n21380 = ~n20962 & n20977 ;
  assign n21381 = ( n20962 & ~n20978 ) | ( n20962 & n21380 ) | ( ~n20978 & n21380 ) ;
  assign n21382 = n20978 | n21381 ;
  assign n21383 = ( n20978 & n21379 ) | ( n20978 & n21382 ) | ( n21379 & n21382 ) ;
  assign n21384 = n20955 | n21383 ;
  assign n21385 = ( n20955 & n20958 ) | ( n20955 & n21384 ) | ( n20958 & n21384 ) ;
  assign n21386 = n20934 | n21385 ;
  assign n21387 = ( n20934 & n20937 ) | ( n20934 & n21386 ) | ( n20937 & n21386 ) ;
  assign n21388 = n20901 | n20915 ;
  assign n21389 = ~n20916 & n21388 ;
  assign n21390 = n20916 | n21389 ;
  assign n21391 = ( n20916 & n21387 ) | ( n20916 & n21390 ) | ( n21387 & n21390 ) ;
  assign n21392 = n20898 & n21391 ;
  assign n21393 = n20896 | n21392 ;
  assign n21394 = n20877 & n21393 ;
  assign n21395 = n20875 | n21394 ;
  assign n21396 = ~n20842 & n20855 ;
  assign n21397 = ( n20842 & ~n20856 ) | ( n20842 & n21396 ) | ( ~n20856 & n21396 ) ;
  assign n21398 = n20856 | n21397 ;
  assign n21399 = ( n20856 & n21395 ) | ( n20856 & n21398 ) | ( n21395 & n21398 ) ;
  assign n21400 = n20839 & n21399 ;
  assign n21401 = n20832 | n21400 ;
  assign n21402 = ( n20835 & n20836 ) | ( n20835 & n21401 ) | ( n20836 & n21401 ) ;
  assign n21403 = n20790 | n21402 ;
  assign n21404 = ( n20790 & ~n20793 ) | ( n20790 & n21403 ) | ( ~n20793 & n21403 ) ;
  assign n21405 = n20768 | n21404 ;
  assign n21406 = ( n20768 & ~n20771 ) | ( n20768 & n21405 ) | ( ~n20771 & n21405 ) ;
  assign n21407 = n20746 | n21406 ;
  assign n21408 = ( n20746 & n20749 ) | ( n20746 & n21407 ) | ( n20749 & n21407 ) ;
  assign n21409 = n20725 | n21408 ;
  assign n21410 = ( n20725 & ~n20728 ) | ( n20725 & n21409 ) | ( ~n20728 & n21409 ) ;
  assign n21411 = ~n20701 & n21410 ;
  assign n21412 = n20697 | n21411 ;
  assign n21413 = n20673 & n21412 ;
  assign n21414 = n20673 | n21412 ;
  assign n21415 = ~n21413 & n21414 ;
  assign n21416 = n1062 & ~n9442 ;
  assign n21417 = n1062 & ~n9074 ;
  assign n21418 = ( n9440 & n21416 ) | ( n9440 & n21417 ) | ( n21416 & n21417 ) ;
  assign n21419 = n1060 & ~n8982 ;
  assign n21420 = ( n1060 & n9051 ) | ( n1060 & n21419 ) | ( n9051 & n21419 ) ;
  assign n21421 = n21418 | n21420 ;
  assign n21422 = n1062 | n21420 ;
  assign n21423 = ( ~n9442 & n21420 ) | ( ~n9442 & n21422 ) | ( n21420 & n21422 ) ;
  assign n21424 = ( ~n9072 & n21421 ) | ( ~n9072 & n21423 ) | ( n21421 & n21423 ) ;
  assign n21425 = n1641 | n8040 ;
  assign n21426 = n12372 | n21425 ;
  assign n21427 = n20361 | n21426 ;
  assign n21428 = n6905 | n21427 ;
  assign n21429 = n9030 | n9037 ;
  assign n21430 = n9027 | n21429 ;
  assign n21431 = n9012 | n21430 ;
  assign n21432 = n575 | n1014 ;
  assign n21433 = n112 | n21432 ;
  assign n21434 = n21431 | n21433 ;
  assign n21435 = n21428 | n21434 ;
  assign n21436 = n7947 & ~n21435 ;
  assign n21437 = ~n124 & n21436 ;
  assign n21438 = ~n858 & n8019 ;
  assign n21439 = ~n20349 & n21438 ;
  assign n21440 = ( n9018 & ~n9036 ) | ( n9018 & n21439 ) | ( ~n9036 & n21439 ) ;
  assign n21441 = n382 | n433 ;
  assign n21442 = n401 | n527 ;
  assign n21443 = n497 | n21442 ;
  assign n21444 = n21441 | n21443 ;
  assign n21445 = n9018 | n21444 ;
  assign n21446 = n21440 & ~n21445 ;
  assign n21447 = ~n21437 & n21446 ;
  assign n21448 = n124 | n21446 ;
  assign n21449 = n21436 & ~n21448 ;
  assign n21450 = n21423 & ~n21449 ;
  assign n21451 = ~n21447 & n21450 ;
  assign n21452 = n21447 | n21449 ;
  assign n21453 = n21421 & ~n21452 ;
  assign n21454 = ( ~n9072 & n21451 ) | ( ~n9072 & n21453 ) | ( n21451 & n21453 ) ;
  assign n21455 = n21424 & ~n21454 ;
  assign n21456 = n21449 | n21453 ;
  assign n21457 = n21447 | n21456 ;
  assign n21458 = n21447 & ~n21449 ;
  assign n21459 = ( n21449 & n21450 ) | ( n21449 & ~n21458 ) | ( n21450 & ~n21458 ) ;
  assign n21460 = n21447 | n21459 ;
  assign n21461 = ( ~n9072 & n21457 ) | ( ~n9072 & n21460 ) | ( n21457 & n21460 ) ;
  assign n21462 = ~n21455 & n21461 ;
  assign n21463 = ~n20409 & n21437 ;
  assign n21464 = n20409 & ~n21437 ;
  assign n21465 = n21463 | n21464 ;
  assign n21466 = n1065 & ~n8982 ;
  assign n21467 = ( n1065 & n9051 ) | ( n1065 & n21466 ) | ( n9051 & n21466 ) ;
  assign n21468 = n1060 & ~n9022 ;
  assign n21469 = ( n1060 & n21467 ) | ( n1060 & ~n21468 ) | ( n21467 & ~n21468 ) ;
  assign n21470 = n1060 | n21467 ;
  assign n21471 = ( ~n9019 & n21469 ) | ( ~n9019 & n21470 ) | ( n21469 & n21470 ) ;
  assign n21472 = n1062 | n21471 ;
  assign n21473 = ~n21465 & n21472 ;
  assign n21474 = n21463 | n21473 ;
  assign n21475 = ~n21465 & n21471 ;
  assign n21476 = n21463 | n21475 ;
  assign n21477 = ( n9078 & n21474 ) | ( n9078 & n21476 ) | ( n21474 & n21476 ) ;
  assign n21478 = ~n21462 & n21477 ;
  assign n21479 = n21462 & ~n21477 ;
  assign n21480 = n21478 | n21479 ;
  assign n21481 = n20471 | n20486 ;
  assign n21482 = ( n9078 & n21471 ) | ( n9078 & n21472 ) | ( n21471 & n21472 ) ;
  assign n21483 = n21465 & n21472 ;
  assign n21484 = n21465 & n21471 ;
  assign n21485 = ( n9078 & n21483 ) | ( n9078 & n21484 ) | ( n21483 & n21484 ) ;
  assign n21486 = n21465 & ~n21484 ;
  assign n21487 = n21465 & ~n21483 ;
  assign n21488 = ( ~n9078 & n21486 ) | ( ~n9078 & n21487 ) | ( n21486 & n21487 ) ;
  assign n21489 = ( n21482 & ~n21485 ) | ( n21482 & n21488 ) | ( ~n21485 & n21488 ) ;
  assign n21490 = n21481 & ~n21489 ;
  assign n21491 = ~n21481 & n21489 ;
  assign n21492 = n21490 | n21491 ;
  assign n21493 = n20530 | n20584 ;
  assign n21494 = ~n21492 & n21493 ;
  assign n21495 = n21490 | n21494 ;
  assign n21496 = ~n21480 & n21495 ;
  assign n21497 = n20530 | n20588 ;
  assign n21498 = ~n21492 & n21497 ;
  assign n21499 = n21490 | n21498 ;
  assign n21500 = ~n21480 & n21499 ;
  assign n21501 = ( n19619 & n21496 ) | ( n19619 & n21500 ) | ( n21496 & n21500 ) ;
  assign n21502 = n20530 | n20595 ;
  assign n21503 = ~n21492 & n21502 ;
  assign n21504 = n21490 | n21503 ;
  assign n21505 = ~n21480 & n21504 ;
  assign n21506 = n20530 | n20601 ;
  assign n21507 = ~n21492 & n21506 ;
  assign n21508 = n21490 | n21507 ;
  assign n21509 = ~n21480 & n21508 ;
  assign n21510 = ( n19345 & n21505 ) | ( n19345 & n21509 ) | ( n21505 & n21509 ) ;
  assign n21511 = ( n15882 & n21501 ) | ( n15882 & n21510 ) | ( n21501 & n21510 ) ;
  assign n21512 = ( n19619 & n21495 ) | ( n19619 & n21499 ) | ( n21495 & n21499 ) ;
  assign n21513 = n21480 & ~n21512 ;
  assign n21514 = ( n19345 & n21504 ) | ( n19345 & n21508 ) | ( n21504 & n21508 ) ;
  assign n21515 = n21480 & ~n21514 ;
  assign n21516 = ( ~n15882 & n21513 ) | ( ~n15882 & n21515 ) | ( n21513 & n21515 ) ;
  assign n21517 = n21511 | n21516 ;
  assign n21518 = ( ~n9072 & n21456 ) | ( ~n9072 & n21459 ) | ( n21456 & n21459 ) ;
  assign n21519 = n170 | n476 ;
  assign n21520 = n381 | n21519 ;
  assign n21521 = n758 | n8995 ;
  assign n21522 = n237 | n6896 ;
  assign n21523 = n8040 | n21522 ;
  assign n21524 = n7982 | n8005 ;
  assign n21525 = n8004 | n21524 ;
  assign n21526 = n21523 | n21525 ;
  assign n21527 = n21521 | n21526 ;
  assign n21528 = n7980 | n21527 ;
  assign n21529 = n7947 & ~n21528 ;
  assign n21530 = ~n21520 & n21529 ;
  assign n21531 = n21437 & n21530 ;
  assign n21532 = n21437 | n21530 ;
  assign n21533 = ~n21531 & n21532 ;
  assign n21534 = n21459 & ~n21533 ;
  assign n21535 = n21449 & ~n21533 ;
  assign n21536 = ( n21453 & ~n21533 ) | ( n21453 & n21535 ) | ( ~n21533 & n21535 ) ;
  assign n21537 = ( ~n9072 & n21534 ) | ( ~n9072 & n21536 ) | ( n21534 & n21536 ) ;
  assign n21538 = n21518 & ~n21537 ;
  assign n21539 = n21456 | n21533 ;
  assign n21540 = n21459 | n21533 ;
  assign n21541 = ( ~n9072 & n21539 ) | ( ~n9072 & n21540 ) | ( n21539 & n21540 ) ;
  assign n21542 = ~n21538 & n21541 ;
  assign n21543 = n21478 | n21501 ;
  assign n21544 = ~n21542 & n21543 ;
  assign n21545 = n21478 | n21510 ;
  assign n21546 = ~n21542 & n21545 ;
  assign n21547 = ( n15882 & n21544 ) | ( n15882 & n21546 ) | ( n21544 & n21546 ) ;
  assign n21548 = n21542 & ~n21543 ;
  assign n21549 = n21542 & ~n21545 ;
  assign n21550 = ( ~n15882 & n21548 ) | ( ~n15882 & n21549 ) | ( n21548 & n21549 ) ;
  assign n21551 = n21547 | n21550 ;
  assign n21552 = n21517 | n21551 ;
  assign n21553 = n21517 & n21551 ;
  assign n21554 = n21552 & ~n21553 ;
  assign n21555 = ( n19619 & n21494 ) | ( n19619 & n21498 ) | ( n21494 & n21498 ) ;
  assign n21556 = ( n19345 & n21503 ) | ( n19345 & n21507 ) | ( n21503 & n21507 ) ;
  assign n21557 = ( n15882 & n21555 ) | ( n15882 & n21556 ) | ( n21555 & n21556 ) ;
  assign n21558 = ( n19619 & n21493 ) | ( n19619 & n21497 ) | ( n21493 & n21497 ) ;
  assign n21559 = n21492 & ~n21558 ;
  assign n21560 = ( n19345 & n21502 ) | ( n19345 & n21506 ) | ( n21502 & n21506 ) ;
  assign n21561 = n21492 & ~n21560 ;
  assign n21562 = ( ~n15882 & n21559 ) | ( ~n15882 & n21561 ) | ( n21559 & n21561 ) ;
  assign n21563 = n21557 | n21562 ;
  assign n21564 = n21517 | n21563 ;
  assign n21565 = ~n20620 & n20621 ;
  assign n21566 = ( ~n20620 & n20634 ) | ( ~n20620 & n21565 ) | ( n20634 & n21565 ) ;
  assign n21567 = n21517 & n21563 ;
  assign n21568 = n21564 & ~n21567 ;
  assign n21569 = n20609 & ~n21563 ;
  assign n21570 = ~n20609 & n21563 ;
  assign n21571 = n21569 | n21570 ;
  assign n21572 = ~n21569 & n21571 ;
  assign n21573 = n21568 & ~n21572 ;
  assign n21574 = n21568 & n21569 ;
  assign n21575 = ( ~n21566 & n21573 ) | ( ~n21566 & n21574 ) | ( n21573 & n21574 ) ;
  assign n21576 = n21564 & ~n21575 ;
  assign n21577 = ~n20620 & n20631 ;
  assign n21578 = ( ~n20620 & n20621 ) | ( ~n20620 & n21577 ) | ( n20621 & n21577 ) ;
  assign n21579 = ( ~n21569 & n21572 ) | ( ~n21569 & n21578 ) | ( n21572 & n21578 ) ;
  assign n21580 = n21564 & ~n21568 ;
  assign n21581 = ( n21564 & n21579 ) | ( n21564 & n21580 ) | ( n21579 & n21580 ) ;
  assign n21582 = ( ~n20643 & n21576 ) | ( ~n20643 & n21581 ) | ( n21576 & n21581 ) ;
  assign n21583 = ( ~n20646 & n21576 ) | ( ~n20646 & n21581 ) | ( n21576 & n21581 ) ;
  assign n21584 = ( ~n18604 & n21582 ) | ( ~n18604 & n21583 ) | ( n21582 & n21583 ) ;
  assign n21585 = n21554 & ~n21584 ;
  assign n21586 = ~n21554 & n21584 ;
  assign n21587 = n21585 | n21586 ;
  assign n21588 = n9475 & ~n21551 ;
  assign n21589 = n9021 & ~n21563 ;
  assign n21590 = n9024 & ~n21517 ;
  assign n21591 = n21589 | n21590 ;
  assign n21592 = n21588 | n21591 ;
  assign n21593 = n8970 | n21588 ;
  assign n21594 = n21591 | n21593 ;
  assign n21595 = ( ~n21587 & n21592 ) | ( ~n21587 & n21594 ) | ( n21592 & n21594 ) ;
  assign n21596 = ~x2 & n21594 ;
  assign n21597 = ~x2 & n21592 ;
  assign n21598 = ( ~n21587 & n21596 ) | ( ~n21587 & n21597 ) | ( n21596 & n21597 ) ;
  assign n21599 = x2 | n21597 ;
  assign n21600 = x2 | n21596 ;
  assign n21601 = ( ~n21587 & n21599 ) | ( ~n21587 & n21600 ) | ( n21599 & n21600 ) ;
  assign n21602 = ( ~n21595 & n21598 ) | ( ~n21595 & n21601 ) | ( n21598 & n21601 ) ;
  assign n21603 = n21415 & n21602 ;
  assign n21604 = n21415 | n21602 ;
  assign n21605 = ~n21603 & n21604 ;
  assign n21606 = ~n20793 & n21402 ;
  assign n21607 = n20793 & ~n21402 ;
  assign n21608 = n21606 | n21607 ;
  assign n21610 = n9021 & n19494 ;
  assign n21611 = n9024 & n19631 ;
  assign n21612 = n21610 | n21611 ;
  assign n21609 = n9475 & ~n20630 ;
  assign n21614 = n8970 | n21609 ;
  assign n21615 = n21612 | n21614 ;
  assign n21613 = n21609 | n21612 ;
  assign n21616 = n21613 & n21615 ;
  assign n21617 = ( ~n20709 & n21615 ) | ( ~n20709 & n21616 ) | ( n21615 & n21616 ) ;
  assign n21618 = ~x2 & n21616 ;
  assign n21619 = ~x2 & n21615 ;
  assign n21620 = ( ~n20709 & n21618 ) | ( ~n20709 & n21619 ) | ( n21618 & n21619 ) ;
  assign n21621 = x2 | n21618 ;
  assign n21622 = x2 | n21619 ;
  assign n21623 = ( ~n20709 & n21621 ) | ( ~n20709 & n21622 ) | ( n21621 & n21622 ) ;
  assign n21624 = ( ~n21617 & n21620 ) | ( ~n21617 & n21623 ) | ( n21620 & n21623 ) ;
  assign n21625 = ~n21608 & n21624 ;
  assign n21626 = n21608 | n21625 ;
  assign n21627 = n21608 & n21624 ;
  assign n21628 = n21626 & ~n21627 ;
  assign n21629 = n21395 & n21397 ;
  assign n21630 = n21395 | n21397 ;
  assign n21631 = ~n21629 & n21630 ;
  assign n21633 = n9021 & ~n18585 ;
  assign n21634 = n9024 & n18410 ;
  assign n21635 = n21633 | n21634 ;
  assign n21632 = n9475 & n18576 ;
  assign n21637 = n8970 | n21632 ;
  assign n21638 = n21635 | n21637 ;
  assign n21636 = n21632 | n21635 ;
  assign n21639 = n21636 & n21638 ;
  assign n21640 = ( n18612 & n21638 ) | ( n18612 & n21639 ) | ( n21638 & n21639 ) ;
  assign n21641 = x2 & n21639 ;
  assign n21642 = x2 & n21638 ;
  assign n21643 = ( n18612 & n21641 ) | ( n18612 & n21642 ) | ( n21641 & n21642 ) ;
  assign n21644 = x2 & ~n21641 ;
  assign n21645 = x2 & ~n21642 ;
  assign n21646 = ( ~n18612 & n21644 ) | ( ~n18612 & n21645 ) | ( n21644 & n21645 ) ;
  assign n21647 = ( n21640 & ~n21643 ) | ( n21640 & n21646 ) | ( ~n21643 & n21646 ) ;
  assign n21648 = n9475 & n18410 ;
  assign n21649 = n9021 & n18037 ;
  assign n21650 = n9024 & ~n18585 ;
  assign n21651 = n21649 | n21650 ;
  assign n21652 = n21648 | n21651 ;
  assign n21653 = n18586 & ~n21652 ;
  assign n21654 = ( n18609 & ~n21652 ) | ( n18609 & n21653 ) | ( ~n21652 & n21653 ) ;
  assign n21655 = ~n18650 & n21654 ;
  assign n21656 = n8970 | n21648 ;
  assign n21657 = n21651 | n21656 ;
  assign n21658 = ~n21655 & n21657 ;
  assign n21659 = x2 & n21657 ;
  assign n21660 = ~n21655 & n21659 ;
  assign n21661 = x2 & ~n21659 ;
  assign n21662 = ( x2 & n21655 ) | ( x2 & n21661 ) | ( n21655 & n21661 ) ;
  assign n21663 = ( n21658 & ~n21660 ) | ( n21658 & n21662 ) | ( ~n21660 & n21662 ) ;
  assign n21664 = n9021 & ~n16069 ;
  assign n21665 = n9024 & n17111 ;
  assign n21666 = n21664 | n21665 ;
  assign n21667 = n9475 & n17100 ;
  assign n21668 = n8970 | n21667 ;
  assign n21669 = n21666 | n21668 ;
  assign n21670 = n21666 | n21667 ;
  assign n21671 = n17169 | n21670 ;
  assign n21672 = ( ~n17129 & n21670 ) | ( ~n17129 & n21671 ) | ( n21670 & n21671 ) ;
  assign n21673 = n21669 & n21672 ;
  assign n21674 = ( n17161 & n21669 ) | ( n17161 & n21673 ) | ( n21669 & n21673 ) ;
  assign n21675 = ~x2 & n21674 ;
  assign n21676 = x2 | n21674 ;
  assign n21677 = ( ~n21674 & n21675 ) | ( ~n21674 & n21676 ) | ( n21675 & n21676 ) ;
  assign n21678 = n9021 & n15886 ;
  assign n21679 = n9024 & ~n16069 ;
  assign n21680 = n21678 | n21679 ;
  assign n21681 = n9475 & n17111 ;
  assign n21682 = n8970 | n21681 ;
  assign n21683 = n21680 | n21682 ;
  assign n21684 = n21680 | n21681 ;
  assign n21685 = n17194 & ~n21684 ;
  assign n21686 = ( n17129 & ~n21684 ) | ( n17129 & n21685 ) | ( ~n21684 & n21685 ) ;
  assign n21687 = n21683 & ~n21686 ;
  assign n21688 = ( n17186 & n21683 ) | ( n17186 & n21687 ) | ( n21683 & n21687 ) ;
  assign n21689 = x2 & n21688 ;
  assign n21690 = x2 & ~n21688 ;
  assign n21691 = ( n21688 & ~n21689 ) | ( n21688 & n21690 ) | ( ~n21689 & n21690 ) ;
  assign n21692 = n21363 & n21365 ;
  assign n21693 = n21363 | n21365 ;
  assign n21694 = ~n21692 & n21693 ;
  assign n21696 = n9021 & n13522 ;
  assign n21697 = n9024 & n14607 ;
  assign n21698 = n21696 | n21697 ;
  assign n21695 = n9475 & n14329 ;
  assign n21700 = n8970 | n21695 ;
  assign n21701 = n21698 | n21700 ;
  assign n21699 = n21695 | n21698 ;
  assign n21702 = n21699 & n21701 ;
  assign n21703 = ( n14656 & n21701 ) | ( n14656 & n21702 ) | ( n21701 & n21702 ) ;
  assign n21704 = x2 & n21702 ;
  assign n21705 = x2 & n21701 ;
  assign n21706 = ( n14656 & n21704 ) | ( n14656 & n21705 ) | ( n21704 & n21705 ) ;
  assign n21707 = x2 & ~n21704 ;
  assign n21708 = x2 & ~n21705 ;
  assign n21709 = ( ~n14656 & n21707 ) | ( ~n14656 & n21708 ) | ( n21707 & n21708 ) ;
  assign n21710 = ( n21703 & ~n21706 ) | ( n21703 & n21709 ) | ( ~n21706 & n21709 ) ;
  assign n21711 = n9021 & n13235 ;
  assign n21712 = n9024 & n13522 ;
  assign n21713 = n21711 | n21712 ;
  assign n21714 = n9475 & n14607 ;
  assign n21715 = n8970 | n21714 ;
  assign n21716 = n21713 | n21715 ;
  assign n21717 = n21713 | n21714 ;
  assign n21718 = n14696 | n21717 ;
  assign n21719 = n14698 | n21717 ;
  assign n21720 = ( ~n13248 & n21718 ) | ( ~n13248 & n21719 ) | ( n21718 & n21719 ) ;
  assign n21721 = n21716 & n21720 ;
  assign n21722 = ( n14687 & n21716 ) | ( n14687 & n21721 ) | ( n21716 & n21721 ) ;
  assign n21723 = ~x2 & n21722 ;
  assign n21724 = x2 | n21722 ;
  assign n21725 = ( ~n21722 & n21723 ) | ( ~n21722 & n21724 ) | ( n21723 & n21724 ) ;
  assign n21726 = n21244 | n21341 ;
  assign n21727 = ~n21342 & n21726 ;
  assign n21728 = n21335 & n21337 ;
  assign n21729 = n21335 | n21337 ;
  assign n21730 = ~n21728 & n21729 ;
  assign n21731 = n9475 & n10649 ;
  assign n21732 = n9021 & n10654 ;
  assign n21733 = n9024 & n10325 ;
  assign n21734 = n21732 | n21733 ;
  assign n21735 = n21731 | n21734 ;
  assign n21736 = n8970 | n21731 ;
  assign n21737 = n21734 | n21736 ;
  assign n21738 = ( n10702 & n21735 ) | ( n10702 & n21737 ) | ( n21735 & n21737 ) ;
  assign n21739 = n21735 | n21737 ;
  assign n21740 = ( n10695 & n21738 ) | ( n10695 & n21739 ) | ( n21738 & n21739 ) ;
  assign n21741 = x2 & n21740 ;
  assign n21742 = x2 & ~n21740 ;
  assign n21743 = ( n21740 & ~n21741 ) | ( n21740 & n21742 ) | ( ~n21741 & n21742 ) ;
  assign n21744 = n21301 & n21319 ;
  assign n21745 = n21301 | n21319 ;
  assign n21746 = ~n21744 & n21745 ;
  assign n21747 = n8113 & ~n10678 ;
  assign n21748 = n9633 & n10784 ;
  assign n21749 = n9644 & ~n10678 ;
  assign n21750 = ( x2 & n9640 ) | ( x2 & n10675 ) | ( n9640 & n10675 ) ;
  assign n21751 = ~n21749 & n21750 ;
  assign n21752 = ~n21748 & n21751 ;
  assign n21753 = n9021 & ~n10678 ;
  assign n21754 = n9024 & ~n10675 ;
  assign n21755 = n21753 | n21754 ;
  assign n21756 = x2 & n9475 ;
  assign n21757 = n10667 & n21756 ;
  assign n21758 = ( x2 & n21755 ) | ( x2 & n21757 ) | ( n21755 & n21757 ) ;
  assign n21759 = n21752 & ~n21758 ;
  assign n21760 = n9660 & ~n10678 ;
  assign n21761 = n9633 | n21760 ;
  assign n21762 = ( n10837 & n21760 ) | ( n10837 & n21761 ) | ( n21760 & n21761 ) ;
  assign n21763 = n21759 & ~n21762 ;
  assign n21764 = n9475 & ~n10662 ;
  assign n21765 = n9021 & ~n10675 ;
  assign n21766 = n9024 & n10667 ;
  assign n21767 = n21765 | n21766 ;
  assign n21768 = n21764 | n21767 ;
  assign n21769 = n8970 | n21764 ;
  assign n21770 = n21767 | n21769 ;
  assign n21771 = ( n10850 & n21768 ) | ( n10850 & n21770 ) | ( n21768 & n21770 ) ;
  assign n21772 = x2 & n21770 ;
  assign n21773 = x2 & n21768 ;
  assign n21774 = ( n10850 & n21772 ) | ( n10850 & n21773 ) | ( n21772 & n21773 ) ;
  assign n21775 = x2 & ~n21774 ;
  assign n21776 = ( n21771 & ~n21774 ) | ( n21771 & n21775 ) | ( ~n21774 & n21775 ) ;
  assign n21777 = ( n21747 & n21763 ) | ( n21747 & n21776 ) | ( n21763 & n21776 ) ;
  assign n21778 = n9475 & n10654 ;
  assign n21779 = n9021 & n10667 ;
  assign n21780 = n9024 & ~n10662 ;
  assign n21781 = n21779 | n21780 ;
  assign n21782 = n21778 | n21781 ;
  assign n21783 = n8970 | n21778 ;
  assign n21784 = n21781 | n21783 ;
  assign n21785 = ( n10978 & n21782 ) | ( n10978 & n21784 ) | ( n21782 & n21784 ) ;
  assign n21786 = x2 & n21784 ;
  assign n21787 = x2 & n21782 ;
  assign n21788 = ( n10978 & n21786 ) | ( n10978 & n21787 ) | ( n21786 & n21787 ) ;
  assign n21789 = x2 & ~n21787 ;
  assign n21790 = x2 & ~n21786 ;
  assign n21791 = ( ~n10978 & n21789 ) | ( ~n10978 & n21790 ) | ( n21789 & n21790 ) ;
  assign n21792 = ( n21785 & ~n21788 ) | ( n21785 & n21791 ) | ( ~n21788 & n21791 ) ;
  assign n21793 = n21777 & n21792 ;
  assign n21794 = n21746 & n21793 ;
  assign n21795 = n21294 | n21297 ;
  assign n21796 = ~n21297 & n21299 ;
  assign n21797 = ( n21295 & n21795 ) | ( n21295 & ~n21796 ) | ( n21795 & ~n21796 ) ;
  assign n21798 = ~n21301 & n21797 ;
  assign n21799 = n21792 & n21798 ;
  assign n21800 = ( n21777 & n21798 ) | ( n21777 & n21799 ) | ( n21798 & n21799 ) ;
  assign n21801 = ( n21746 & n21794 ) | ( n21746 & n21800 ) | ( n21794 & n21800 ) ;
  assign n21802 = n21743 & n21801 ;
  assign n21803 = n21746 | n21793 ;
  assign n21804 = n9475 & n10325 ;
  assign n21805 = n9021 & ~n10662 ;
  assign n21806 = n9024 & n10654 ;
  assign n21807 = n21805 | n21806 ;
  assign n21808 = n21804 | n21807 ;
  assign n21809 = n8970 | n21808 ;
  assign n21810 = ( ~n10957 & n21808 ) | ( ~n10957 & n21809 ) | ( n21808 & n21809 ) ;
  assign n21811 = n21808 | n21809 ;
  assign n21812 = ( n10949 & n21810 ) | ( n10949 & n21811 ) | ( n21810 & n21811 ) ;
  assign n21813 = ~x2 & n21812 ;
  assign n21814 = x2 | n21812 ;
  assign n21815 = ( ~n21812 & n21813 ) | ( ~n21812 & n21814 ) | ( n21813 & n21814 ) ;
  assign n21816 = n21800 & n21815 ;
  assign n21817 = ( n21803 & n21815 ) | ( n21803 & n21816 ) | ( n21815 & n21816 ) ;
  assign n21818 = ( n21743 & n21802 ) | ( n21743 & n21817 ) | ( n21802 & n21817 ) ;
  assign n21819 = n21730 | n21818 ;
  assign n21820 = n21322 & ~n21333 ;
  assign n21821 = n21743 | n21801 ;
  assign n21822 = ( n21333 & n21817 ) | ( n21333 & n21820 ) | ( n21817 & n21820 ) ;
  assign n21823 = n21333 | n21820 ;
  assign n21824 = ( n21821 & n21822 ) | ( n21821 & n21823 ) | ( n21822 & n21823 ) ;
  assign n21825 = ( ~n21322 & n21820 ) | ( ~n21322 & n21824 ) | ( n21820 & n21824 ) ;
  assign n21826 = n21819 | n21825 ;
  assign n21827 = n9475 & n11363 ;
  assign n21828 = n9021 & n10325 ;
  assign n21829 = n9024 & n10649 ;
  assign n21830 = n21828 | n21829 ;
  assign n21831 = n21827 | n21830 ;
  assign n21832 = n8970 | n21831 ;
  assign n21833 = ( n12059 & n21831 ) | ( n12059 & n21832 ) | ( n21831 & n21832 ) ;
  assign n21834 = x2 & n21832 ;
  assign n21835 = x2 & n21831 ;
  assign n21836 = ( n12059 & n21834 ) | ( n12059 & n21835 ) | ( n21834 & n21835 ) ;
  assign n21837 = x2 & ~n21834 ;
  assign n21838 = x2 & ~n21835 ;
  assign n21839 = ( ~n12059 & n21837 ) | ( ~n12059 & n21838 ) | ( n21837 & n21838 ) ;
  assign n21840 = ( n21833 & ~n21836 ) | ( n21833 & n21839 ) | ( ~n21836 & n21839 ) ;
  assign n21841 = n21826 & n21840 ;
  assign n21842 = n9021 & n10649 ;
  assign n21843 = n9024 & n11363 ;
  assign n21844 = n21842 | n21843 ;
  assign n21845 = n9475 & ~n11663 ;
  assign n21846 = n8970 | n21845 ;
  assign n21847 = n21844 | n21846 ;
  assign n21848 = n21844 | n21845 ;
  assign n21849 = n12048 & ~n21848 ;
  assign n21850 = ( n11672 & ~n21848 ) | ( n11672 & n21849 ) | ( ~n21848 & n21849 ) ;
  assign n21851 = n21847 & ~n21850 ;
  assign n21852 = ( n12040 & n21847 ) | ( n12040 & n21851 ) | ( n21847 & n21851 ) ;
  assign n21853 = x2 & n21852 ;
  assign n21854 = x2 & ~n21852 ;
  assign n21855 = ( n21852 & ~n21853 ) | ( n21852 & n21854 ) | ( ~n21853 & n21854 ) ;
  assign n21856 = n21730 & n21818 ;
  assign n21857 = ( n21730 & n21825 ) | ( n21730 & n21856 ) | ( n21825 & n21856 ) ;
  assign n21858 = n21855 & n21857 ;
  assign n21859 = ( n21841 & n21855 ) | ( n21841 & n21858 ) | ( n21855 & n21858 ) ;
  assign n21861 = n9021 & n11363 ;
  assign n21862 = n9024 & ~n11663 ;
  assign n21863 = n21861 | n21862 ;
  assign n21860 = n9475 & n12010 ;
  assign n21865 = n8970 | n21860 ;
  assign n21866 = n21863 | n21865 ;
  assign n21864 = n21860 | n21863 ;
  assign n21867 = n21864 & n21866 ;
  assign n21868 = ( ~n12028 & n21866 ) | ( ~n12028 & n21867 ) | ( n21866 & n21867 ) ;
  assign n21869 = n21866 | n21867 ;
  assign n21870 = ( n12017 & n21868 ) | ( n12017 & n21869 ) | ( n21868 & n21869 ) ;
  assign n21871 = ~x2 & n21870 ;
  assign n21872 = x2 | n21870 ;
  assign n21873 = ( ~n21870 & n21871 ) | ( ~n21870 & n21872 ) | ( n21871 & n21872 ) ;
  assign n21874 = n21859 | n21873 ;
  assign n21875 = n21268 & ~n21339 ;
  assign n21876 = n21855 | n21857 ;
  assign n21877 = n21841 | n21876 ;
  assign n21878 = ( ~n21268 & n21339 ) | ( ~n21268 & n21875 ) | ( n21339 & n21875 ) ;
  assign n21879 = ( n21875 & n21877 ) | ( n21875 & n21878 ) | ( n21877 & n21878 ) ;
  assign n21880 = n21874 | n21879 ;
  assign n21881 = n21727 & n21880 ;
  assign n21883 = n9021 & ~n11663 ;
  assign n21884 = n9024 & n12010 ;
  assign n21885 = n21883 | n21884 ;
  assign n21882 = n9475 & ~n12616 ;
  assign n21887 = n8970 | n21882 ;
  assign n21888 = n21885 | n21887 ;
  assign n21886 = n21882 | n21885 ;
  assign n21889 = n21886 & n21888 ;
  assign n21890 = ( ~n12626 & n21888 ) | ( ~n12626 & n21889 ) | ( n21888 & n21889 ) ;
  assign n21891 = ~x2 & n21889 ;
  assign n21892 = ~x2 & n21888 ;
  assign n21893 = ( ~n12626 & n21891 ) | ( ~n12626 & n21892 ) | ( n21891 & n21892 ) ;
  assign n21894 = x2 | n21891 ;
  assign n21895 = x2 | n21892 ;
  assign n21896 = ( ~n12626 & n21894 ) | ( ~n12626 & n21895 ) | ( n21894 & n21895 ) ;
  assign n21897 = ( ~n21890 & n21893 ) | ( ~n21890 & n21896 ) | ( n21893 & n21896 ) ;
  assign n21898 = n21859 & n21873 ;
  assign n21899 = ( n21873 & n21879 ) | ( n21873 & n21898 ) | ( n21879 & n21898 ) ;
  assign n21900 = n21897 & n21899 ;
  assign n21901 = ( n21881 & n21897 ) | ( n21881 & n21900 ) | ( n21897 & n21900 ) ;
  assign n21902 = n21205 | n21347 ;
  assign n21903 = ~n21347 & n21902 ;
  assign n21904 = ( ~n21205 & n21902 ) | ( ~n21205 & n21903 ) | ( n21902 & n21903 ) ;
  assign n21905 = n21901 | n21904 ;
  assign n21906 = n21343 & ~n21345 ;
  assign n21907 = n21897 | n21899 ;
  assign n21908 = n21881 | n21907 ;
  assign n21909 = ( ~n21343 & n21345 ) | ( ~n21343 & n21906 ) | ( n21345 & n21906 ) ;
  assign n21910 = ( n21906 & n21908 ) | ( n21906 & n21909 ) | ( n21908 & n21909 ) ;
  assign n21911 = n21905 | n21910 ;
  assign n21912 = n9475 & n12936 ;
  assign n21913 = n9021 & n12010 ;
  assign n21914 = n9024 & ~n12616 ;
  assign n21915 = n21913 | n21914 ;
  assign n21916 = n21912 | n21915 ;
  assign n21917 = n8970 | n21912 ;
  assign n21918 = n21915 | n21917 ;
  assign n21919 = ( ~n13591 & n21916 ) | ( ~n13591 & n21918 ) | ( n21916 & n21918 ) ;
  assign n21920 = ~x2 & n21918 ;
  assign n21921 = ~x2 & n21916 ;
  assign n21922 = ( ~n13591 & n21920 ) | ( ~n13591 & n21921 ) | ( n21920 & n21921 ) ;
  assign n21923 = x2 | n21921 ;
  assign n21924 = x2 | n21920 ;
  assign n21925 = ( ~n13591 & n21923 ) | ( ~n13591 & n21924 ) | ( n21923 & n21924 ) ;
  assign n21926 = ( ~n21919 & n21922 ) | ( ~n21919 & n21925 ) | ( n21922 & n21925 ) ;
  assign n21927 = n21911 & n21926 ;
  assign n21928 = n21185 | n21349 ;
  assign n21929 = ~n21350 & n21928 ;
  assign n21930 = n21901 & n21904 ;
  assign n21931 = ( n21904 & n21910 ) | ( n21904 & n21930 ) | ( n21910 & n21930 ) ;
  assign n21932 = n21929 | n21931 ;
  assign n21933 = n21927 | n21932 ;
  assign n21934 = n9475 & n13235 ;
  assign n21935 = n9021 & ~n12616 ;
  assign n21936 = n9024 & n12936 ;
  assign n21937 = n21935 | n21936 ;
  assign n21938 = n21934 | n21937 ;
  assign n21939 = n8970 | n21934 ;
  assign n21940 = n21937 | n21939 ;
  assign n21941 = ( n13561 & n21938 ) | ( n13561 & n21940 ) | ( n21938 & n21940 ) ;
  assign n21942 = x2 & n21940 ;
  assign n21943 = x2 & n21938 ;
  assign n21944 = ( n13561 & n21942 ) | ( n13561 & n21943 ) | ( n21942 & n21943 ) ;
  assign n21945 = x2 & ~n21943 ;
  assign n21946 = x2 & ~n21942 ;
  assign n21947 = ( ~n13561 & n21945 ) | ( ~n13561 & n21946 ) | ( n21945 & n21946 ) ;
  assign n21948 = ( n21941 & ~n21944 ) | ( n21941 & n21947 ) | ( ~n21944 & n21947 ) ;
  assign n21949 = n21933 & n21948 ;
  assign n21950 = n21351 & n21353 ;
  assign n21951 = n21351 | n21353 ;
  assign n21952 = ~n21950 & n21951 ;
  assign n21953 = n21929 & n21931 ;
  assign n21954 = ( n21927 & n21929 ) | ( n21927 & n21953 ) | ( n21929 & n21953 ) ;
  assign n21955 = n21952 & n21954 ;
  assign n21956 = ( n21949 & n21952 ) | ( n21949 & n21955 ) | ( n21952 & n21955 ) ;
  assign n21957 = n21725 & n21956 ;
  assign n21958 = n21952 | n21954 ;
  assign n21959 = n21949 | n21958 ;
  assign n21960 = n9475 & n13522 ;
  assign n21961 = n9021 & n12936 ;
  assign n21962 = n9024 & n13235 ;
  assign n21963 = n21961 | n21962 ;
  assign n21964 = n21960 | n21963 ;
  assign n21965 = n8970 & n13537 ;
  assign n21966 = n8970 & n13539 ;
  assign n21967 = ( ~n13248 & n21965 ) | ( ~n13248 & n21966 ) | ( n21965 & n21966 ) ;
  assign n21968 = n21964 | n21967 ;
  assign n21969 = n8970 | n21964 ;
  assign n21970 = ( n13530 & n21968 ) | ( n13530 & n21969 ) | ( n21968 & n21969 ) ;
  assign n21971 = x2 & n21970 ;
  assign n21972 = n21970 & ~n21971 ;
  assign n21973 = x2 & ~n21971 ;
  assign n21974 = ( n21959 & n21972 ) | ( n21959 & n21973 ) | ( n21972 & n21973 ) ;
  assign n21975 = ( n21725 & n21957 ) | ( n21725 & n21974 ) | ( n21957 & n21974 ) ;
  assign n21976 = n21710 & n21975 ;
  assign n21977 = ~n21355 & n21357 ;
  assign n21978 = n21725 | n21956 ;
  assign n21979 = n21974 | n21978 ;
  assign n21980 = ( n21355 & ~n21357 ) | ( n21355 & n21977 ) | ( ~n21357 & n21977 ) ;
  assign n21981 = ( n21977 & n21979 ) | ( n21977 & n21980 ) | ( n21979 & n21980 ) ;
  assign n21982 = ( n21710 & n21976 ) | ( n21710 & n21981 ) | ( n21976 & n21981 ) ;
  assign n21984 = n9021 & n14607 ;
  assign n21985 = n9024 & n14329 ;
  assign n21986 = n21984 | n21985 ;
  assign n21983 = n9475 & n14591 ;
  assign n21988 = n8970 | n21983 ;
  assign n21989 = n21986 | n21988 ;
  assign n21987 = n21983 | n21986 ;
  assign n21990 = n21987 & n21989 ;
  assign n21991 = ( n14629 & n21989 ) | ( n14629 & n21990 ) | ( n21989 & n21990 ) ;
  assign n21992 = x2 & n21990 ;
  assign n21993 = x2 & n21989 ;
  assign n21994 = ( n14629 & n21992 ) | ( n14629 & n21993 ) | ( n21992 & n21993 ) ;
  assign n21995 = x2 & ~n21992 ;
  assign n21996 = x2 & ~n21993 ;
  assign n21997 = ( ~n14629 & n21995 ) | ( ~n14629 & n21996 ) | ( n21995 & n21996 ) ;
  assign n21998 = ( n21991 & ~n21994 ) | ( n21991 & n21997 ) | ( ~n21994 & n21997 ) ;
  assign n21999 = n21982 | n21998 ;
  assign n22000 = n21710 | n21975 ;
  assign n22001 = n21981 | n22000 ;
  assign n22002 = ~n21359 & n21360 ;
  assign n22003 = ( n21126 & ~n21359 ) | ( n21126 & n22002 ) | ( ~n21359 & n22002 ) ;
  assign n22004 = n21126 | n21360 ;
  assign n22005 = ( n21359 & n22003 ) | ( n21359 & ~n22004 ) | ( n22003 & ~n22004 ) ;
  assign n22006 = ( n22001 & n22003 ) | ( n22001 & n22005 ) | ( n22003 & n22005 ) ;
  assign n22007 = n21999 | n22006 ;
  assign n22008 = n21694 & n22007 ;
  assign n22009 = ( n21086 & n21087 ) | ( n21086 & ~n21367 ) | ( n21087 & ~n21367 ) ;
  assign n22010 = n21367 | n22009 ;
  assign n22011 = ~n21368 & n22010 ;
  assign n22012 = n21982 & n21998 ;
  assign n22013 = ( n21998 & n22006 ) | ( n21998 & n22012 ) | ( n22006 & n22012 ) ;
  assign n22014 = n22011 | n22013 ;
  assign n22015 = n22008 | n22014 ;
  assign n22016 = n9475 & n15434 ;
  assign n22017 = n9021 & n14329 ;
  assign n22018 = n9024 & n14591 ;
  assign n22019 = n22017 | n22018 ;
  assign n22020 = n22016 | n22019 ;
  assign n22021 = n8970 | n22016 ;
  assign n22022 = n22019 | n22021 ;
  assign n22023 = ( n15453 & n22020 ) | ( n15453 & n22022 ) | ( n22020 & n22022 ) ;
  assign n22024 = x2 & n22022 ;
  assign n22025 = x2 & n22020 ;
  assign n22026 = ( n15453 & n22024 ) | ( n15453 & n22025 ) | ( n22024 & n22025 ) ;
  assign n22027 = x2 & ~n22025 ;
  assign n22028 = x2 & ~n22024 ;
  assign n22029 = ( ~n15453 & n22027 ) | ( ~n15453 & n22028 ) | ( n22027 & n22028 ) ;
  assign n22030 = ( n22023 & ~n22026 ) | ( n22023 & n22029 ) | ( ~n22026 & n22029 ) ;
  assign n22031 = n22015 & n22030 ;
  assign n22032 = ( ~n21369 & n21370 ) | ( ~n21369 & n21371 ) | ( n21370 & n21371 ) ;
  assign n22033 = n21369 | n22032 ;
  assign n22034 = ~n21373 & n22033 ;
  assign n22035 = n22011 & n22013 ;
  assign n22036 = ( n22008 & n22011 ) | ( n22008 & n22035 ) | ( n22011 & n22035 ) ;
  assign n22037 = n22034 | n22036 ;
  assign n22038 = n22031 | n22037 ;
  assign n22039 = n9475 & ~n16085 ;
  assign n22040 = n9021 & n14591 ;
  assign n22041 = n9024 & n15434 ;
  assign n22042 = n22040 | n22041 ;
  assign n22043 = n22039 | n22042 ;
  assign n22044 = n8970 | n22039 ;
  assign n22045 = n22042 | n22044 ;
  assign n22046 = ( ~n16167 & n22043 ) | ( ~n16167 & n22045 ) | ( n22043 & n22045 ) ;
  assign n22047 = ~x2 & n22045 ;
  assign n22048 = ~x2 & n22043 ;
  assign n22049 = ( ~n16167 & n22047 ) | ( ~n16167 & n22048 ) | ( n22047 & n22048 ) ;
  assign n22050 = x2 | n22048 ;
  assign n22051 = x2 | n22047 ;
  assign n22052 = ( ~n16167 & n22050 ) | ( ~n16167 & n22051 ) | ( n22050 & n22051 ) ;
  assign n22053 = ( ~n22046 & n22049 ) | ( ~n22046 & n22052 ) | ( n22049 & n22052 ) ;
  assign n22054 = n22038 & n22053 ;
  assign n22055 = ( n21064 & n21065 ) | ( n21064 & n21373 ) | ( n21065 & n21373 ) ;
  assign n22056 = n21042 | n21064 ;
  assign n22057 = n21373 | n22056 ;
  assign n22058 = ~n22055 & n22057 ;
  assign n22059 = n22034 & n22036 ;
  assign n22060 = ( n22031 & n22034 ) | ( n22031 & n22059 ) | ( n22034 & n22059 ) ;
  assign n22061 = n22058 | n22060 ;
  assign n22062 = n22054 | n22061 ;
  assign n22063 = n9475 & n15886 ;
  assign n22064 = n9021 & n15434 ;
  assign n22065 = n9024 & ~n16085 ;
  assign n22066 = n22064 | n22065 ;
  assign n22067 = n22063 | n22066 ;
  assign n22068 = n8970 | n22063 ;
  assign n22069 = n22066 | n22068 ;
  assign n22070 = ( ~n16140 & n22067 ) | ( ~n16140 & n22069 ) | ( n22067 & n22069 ) ;
  assign n22071 = ~x2 & n22069 ;
  assign n22072 = ~x2 & n22067 ;
  assign n22073 = ( ~n16140 & n22071 ) | ( ~n16140 & n22072 ) | ( n22071 & n22072 ) ;
  assign n22074 = x2 | n22072 ;
  assign n22075 = x2 | n22071 ;
  assign n22076 = ( ~n16140 & n22074 ) | ( ~n16140 & n22075 ) | ( n22074 & n22075 ) ;
  assign n22077 = ( ~n22070 & n22073 ) | ( ~n22070 & n22076 ) | ( n22073 & n22076 ) ;
  assign n22078 = n22062 & n22077 ;
  assign n22079 = n9475 & ~n16069 ;
  assign n22080 = n9021 & ~n16085 ;
  assign n22081 = n9024 & n15886 ;
  assign n22082 = n22080 | n22081 ;
  assign n22083 = n22079 | n22082 ;
  assign n22084 = n8970 | n22083 ;
  assign n22085 = ( ~n16107 & n22083 ) | ( ~n16107 & n22084 ) | ( n22083 & n22084 ) ;
  assign n22086 = ~x2 & n22084 ;
  assign n22087 = ~x2 & n22083 ;
  assign n22088 = ( ~n16107 & n22086 ) | ( ~n16107 & n22087 ) | ( n22086 & n22087 ) ;
  assign n22089 = x2 | n22086 ;
  assign n22090 = x2 | n22087 ;
  assign n22091 = ( ~n16107 & n22089 ) | ( ~n16107 & n22090 ) | ( n22089 & n22090 ) ;
  assign n22092 = ( ~n22085 & n22088 ) | ( ~n22085 & n22091 ) | ( n22088 & n22091 ) ;
  assign n22093 = n22058 & n22060 ;
  assign n22094 = ( n22054 & n22058 ) | ( n22054 & n22093 ) | ( n22058 & n22093 ) ;
  assign n22095 = n22092 & n22094 ;
  assign n22096 = ( n22078 & n22092 ) | ( n22078 & n22095 ) | ( n22092 & n22095 ) ;
  assign n22097 = n21691 & n22096 ;
  assign n22098 = n21022 & ~n21375 ;
  assign n22099 = n22092 | n22094 ;
  assign n22100 = n22078 | n22099 ;
  assign n22101 = ( ~n21022 & n21375 ) | ( ~n21022 & n22098 ) | ( n21375 & n22098 ) ;
  assign n22102 = ( n22098 & n22100 ) | ( n22098 & n22101 ) | ( n22100 & n22101 ) ;
  assign n22103 = ( n21691 & n22097 ) | ( n21691 & n22102 ) | ( n22097 & n22102 ) ;
  assign n22104 = n21677 & n22103 ;
  assign n22105 = n21000 & ~n21377 ;
  assign n22106 = n21691 | n22096 ;
  assign n22107 = n22102 | n22106 ;
  assign n22108 = ( ~n21000 & n21377 ) | ( ~n21000 & n22105 ) | ( n21377 & n22105 ) ;
  assign n22109 = ( n22105 & n22107 ) | ( n22105 & n22108 ) | ( n22107 & n22108 ) ;
  assign n22110 = ( n21677 & n22104 ) | ( n21677 & n22109 ) | ( n22104 & n22109 ) ;
  assign n22111 = n20958 | n21383 ;
  assign n22112 = n20958 & ~n21383 ;
  assign n22113 = ( ~n20958 & n22111 ) | ( ~n20958 & n22112 ) | ( n22111 & n22112 ) ;
  assign n22114 = n22110 | n22113 ;
  assign n22115 = n21379 & ~n21381 ;
  assign n22116 = n21677 | n22103 ;
  assign n22117 = n22109 | n22116 ;
  assign n22118 = ( ~n21379 & n21381 ) | ( ~n21379 & n22115 ) | ( n21381 & n22115 ) ;
  assign n22119 = ( n22115 & n22117 ) | ( n22115 & n22118 ) | ( n22117 & n22118 ) ;
  assign n22120 = n22114 | n22119 ;
  assign n22121 = n9475 & ~n17092 ;
  assign n22122 = n9021 & n17111 ;
  assign n22123 = n9024 & n17100 ;
  assign n22124 = n22122 | n22123 ;
  assign n22125 = n22121 | n22124 ;
  assign n22126 = n8970 | n22121 ;
  assign n22127 = n22124 | n22126 ;
  assign n22128 = ( ~n17134 & n22125 ) | ( ~n17134 & n22127 ) | ( n22125 & n22127 ) ;
  assign n22129 = ~x2 & n22127 ;
  assign n22130 = ~x2 & n22125 ;
  assign n22131 = ( ~n17134 & n22129 ) | ( ~n17134 & n22130 ) | ( n22129 & n22130 ) ;
  assign n22132 = x2 | n22130 ;
  assign n22133 = x2 | n22129 ;
  assign n22134 = ( ~n17134 & n22132 ) | ( ~n17134 & n22133 ) | ( n22132 & n22133 ) ;
  assign n22135 = ( ~n22128 & n22131 ) | ( ~n22128 & n22134 ) | ( n22131 & n22134 ) ;
  assign n22136 = n22120 & n22135 ;
  assign n22137 = n22110 & n22113 ;
  assign n22138 = ( n22113 & n22119 ) | ( n22113 & n22137 ) | ( n22119 & n22137 ) ;
  assign n22139 = n20937 | n21385 ;
  assign n22140 = n20937 & ~n21385 ;
  assign n22141 = ( ~n20937 & n22139 ) | ( ~n20937 & n22140 ) | ( n22139 & n22140 ) ;
  assign n22142 = n22138 | n22141 ;
  assign n22143 = n22136 | n22142 ;
  assign n22144 = n9475 & n18037 ;
  assign n22145 = n9021 & n17100 ;
  assign n22146 = n9024 & ~n17092 ;
  assign n22147 = n22145 | n22146 ;
  assign n22148 = n22144 | n22147 ;
  assign n22149 = n8970 | n22144 ;
  assign n22150 = n22147 | n22149 ;
  assign n22151 = ( ~n18050 & n22148 ) | ( ~n18050 & n22150 ) | ( n22148 & n22150 ) ;
  assign n22152 = ~x2 & n22150 ;
  assign n22153 = ~x2 & n22148 ;
  assign n22154 = ( ~n18050 & n22152 ) | ( ~n18050 & n22153 ) | ( n22152 & n22153 ) ;
  assign n22155 = x2 | n22153 ;
  assign n22156 = x2 | n22152 ;
  assign n22157 = ( ~n18050 & n22155 ) | ( ~n18050 & n22156 ) | ( n22155 & n22156 ) ;
  assign n22158 = ( ~n22151 & n22154 ) | ( ~n22151 & n22157 ) | ( n22154 & n22157 ) ;
  assign n22159 = n22143 & n22158 ;
  assign n22160 = n21387 & n21389 ;
  assign n22161 = n21387 | n21389 ;
  assign n22162 = ~n22160 & n22161 ;
  assign n22163 = n22138 & n22141 ;
  assign n22164 = ( n22136 & n22141 ) | ( n22136 & n22163 ) | ( n22141 & n22163 ) ;
  assign n22165 = n22162 & n22164 ;
  assign n22166 = ( n22159 & n22162 ) | ( n22159 & n22165 ) | ( n22162 & n22165 ) ;
  assign n22167 = n21663 & n22166 ;
  assign n22168 = n22162 | n22164 ;
  assign n22169 = n22159 | n22168 ;
  assign n22170 = n8970 & ~n18675 ;
  assign n22171 = ( n8970 & n18672 ) | ( n8970 & n22170 ) | ( n18672 & n22170 ) ;
  assign n22172 = n9475 & ~n18585 ;
  assign n22173 = n9021 & ~n17092 ;
  assign n22174 = n9024 & n18037 ;
  assign n22175 = n22173 | n22174 ;
  assign n22176 = n22172 | n22175 ;
  assign n22177 = n22171 | n22176 ;
  assign n22178 = x2 & n22176 ;
  assign n22179 = ( x2 & n22171 ) | ( x2 & n22178 ) | ( n22171 & n22178 ) ;
  assign n22180 = n22177 & ~n22179 ;
  assign n22181 = x2 & ~n22179 ;
  assign n22182 = ( n22169 & n22180 ) | ( n22169 & n22181 ) | ( n22180 & n22181 ) ;
  assign n22183 = ( n21663 & n22167 ) | ( n21663 & n22182 ) | ( n22167 & n22182 ) ;
  assign n22184 = n21647 & n22183 ;
  assign n22185 = n20898 & ~n21391 ;
  assign n22186 = n21663 | n22166 ;
  assign n22187 = n22182 | n22186 ;
  assign n22188 = ( ~n20898 & n21391 ) | ( ~n20898 & n22185 ) | ( n21391 & n22185 ) ;
  assign n22189 = ( n22185 & n22187 ) | ( n22185 & n22188 ) | ( n22187 & n22188 ) ;
  assign n22190 = ( n21647 & n22184 ) | ( n21647 & n22189 ) | ( n22184 & n22189 ) ;
  assign n22192 = n9021 & n18410 ;
  assign n22193 = n9024 & n18576 ;
  assign n22194 = n22192 | n22193 ;
  assign n22191 = n9475 & n19352 ;
  assign n22196 = n8970 | n22191 ;
  assign n22197 = n22194 | n22196 ;
  assign n22195 = n22191 | n22194 ;
  assign n22198 = n22195 & n22197 ;
  assign n22199 = ( n19674 & n22197 ) | ( n19674 & n22198 ) | ( n22197 & n22198 ) ;
  assign n22200 = x2 & n22198 ;
  assign n22201 = x2 & n22197 ;
  assign n22202 = ( n19674 & n22200 ) | ( n19674 & n22201 ) | ( n22200 & n22201 ) ;
  assign n22203 = x2 & ~n22200 ;
  assign n22204 = x2 & ~n22201 ;
  assign n22205 = ( ~n19674 & n22203 ) | ( ~n19674 & n22204 ) | ( n22203 & n22204 ) ;
  assign n22206 = ( n22199 & ~n22202 ) | ( n22199 & n22205 ) | ( ~n22202 & n22205 ) ;
  assign n22207 = n22190 | n22206 ;
  assign n22208 = n20877 & ~n21393 ;
  assign n22209 = n21647 | n22183 ;
  assign n22210 = n22189 | n22209 ;
  assign n22211 = ( ~n20877 & n21393 ) | ( ~n20877 & n22208 ) | ( n21393 & n22208 ) ;
  assign n22212 = ( n22208 & n22210 ) | ( n22208 & n22211 ) | ( n22210 & n22211 ) ;
  assign n22213 = n22207 | n22212 ;
  assign n22214 = n21631 & n22213 ;
  assign n22215 = ( n20837 & n20838 ) | ( n20837 & ~n21399 ) | ( n20838 & ~n21399 ) ;
  assign n22216 = n21399 | n22215 ;
  assign n22217 = ~n21400 & n22216 ;
  assign n22218 = n22190 & n22206 ;
  assign n22219 = ( n22206 & n22212 ) | ( n22206 & n22218 ) | ( n22212 & n22218 ) ;
  assign n22220 = n22217 | n22219 ;
  assign n22221 = n22214 | n22220 ;
  assign n22222 = n9475 & n19494 ;
  assign n22223 = n9021 & n18576 ;
  assign n22224 = n9024 & n19352 ;
  assign n22225 = n22223 | n22224 ;
  assign n22226 = n22222 | n22225 ;
  assign n22227 = n8970 | n22222 ;
  assign n22228 = n22225 | n22227 ;
  assign n22229 = ( n20320 & n22226 ) | ( n20320 & n22228 ) | ( n22226 & n22228 ) ;
  assign n22230 = x2 & n22228 ;
  assign n22231 = x2 & n22226 ;
  assign n22232 = ( n20320 & n22230 ) | ( n20320 & n22231 ) | ( n22230 & n22231 ) ;
  assign n22233 = x2 & ~n22231 ;
  assign n22234 = x2 & ~n22230 ;
  assign n22235 = ( ~n20320 & n22233 ) | ( ~n20320 & n22234 ) | ( n22233 & n22234 ) ;
  assign n22236 = ( n22229 & ~n22232 ) | ( n22229 & n22235 ) | ( ~n22232 & n22235 ) ;
  assign n22237 = n22221 & n22236 ;
  assign n22238 = ( n20834 & n20835 ) | ( n20834 & n21400 ) | ( n20835 & n21400 ) ;
  assign n22239 = n20812 | n20834 ;
  assign n22240 = n21400 | n22239 ;
  assign n22241 = ~n22238 & n22240 ;
  assign n22242 = n22217 & n22219 ;
  assign n22243 = ( n22214 & n22217 ) | ( n22214 & n22242 ) | ( n22217 & n22242 ) ;
  assign n22244 = n22241 | n22243 ;
  assign n22245 = n22237 | n22244 ;
  assign n22246 = n9475 & n19631 ;
  assign n22247 = n9021 & n19352 ;
  assign n22248 = n9024 & n19494 ;
  assign n22249 = n22247 | n22248 ;
  assign n22250 = n22246 | n22249 ;
  assign n22251 = n8970 & n19652 ;
  assign n22252 = n8970 & n19655 ;
  assign n22253 = ( ~n18604 & n22251 ) | ( ~n18604 & n22252 ) | ( n22251 & n22252 ) ;
  assign n22254 = n22250 | n22253 ;
  assign n22255 = n8970 | n22250 ;
  assign n22256 = ( n19640 & n22254 ) | ( n19640 & n22255 ) | ( n22254 & n22255 ) ;
  assign n22257 = x2 & n22256 ;
  assign n22258 = n22256 & ~n22257 ;
  assign n22259 = x2 & ~n22257 ;
  assign n22260 = ( n22245 & n22258 ) | ( n22245 & n22259 ) | ( n22258 & n22259 ) ;
  assign n22261 = n22241 & n22243 ;
  assign n22262 = ( n22237 & n22241 ) | ( n22237 & n22261 ) | ( n22241 & n22261 ) ;
  assign n22263 = ~n21628 & n22262 ;
  assign n22264 = ( ~n21628 & n22260 ) | ( ~n21628 & n22263 ) | ( n22260 & n22263 ) ;
  assign n22265 = n20701 & ~n21410 ;
  assign n22266 = n21411 | n22265 ;
  assign n22267 = ( n21566 & ~n21569 ) | ( n21566 & n21572 ) | ( ~n21569 & n21572 ) ;
  assign n22268 = ( ~n20643 & n21579 ) | ( ~n20643 & n22267 ) | ( n21579 & n22267 ) ;
  assign n22269 = ( ~n20646 & n21579 ) | ( ~n20646 & n22267 ) | ( n21579 & n22267 ) ;
  assign n22270 = ( ~n18604 & n22268 ) | ( ~n18604 & n22269 ) | ( n22268 & n22269 ) ;
  assign n22271 = ~n21568 & n22270 ;
  assign n22273 = n9021 & n20609 ;
  assign n22274 = n9024 & ~n21563 ;
  assign n22275 = n22273 | n22274 ;
  assign n22272 = n9475 & ~n21517 ;
  assign n22277 = n8970 | n22272 ;
  assign n22278 = n22275 | n22277 ;
  assign n22276 = n22272 | n22275 ;
  assign n22279 = n22276 & n22278 ;
  assign n22280 = n21568 & ~n21579 ;
  assign n22281 = ( n20643 & n21575 ) | ( n20643 & n22280 ) | ( n21575 & n22280 ) ;
  assign n22282 = ( n20646 & n21575 ) | ( n20646 & n22280 ) | ( n21575 & n22280 ) ;
  assign n22283 = ( n18604 & n22281 ) | ( n18604 & n22282 ) | ( n22281 & n22282 ) ;
  assign n22284 = ( n22278 & n22279 ) | ( n22278 & ~n22283 ) | ( n22279 & ~n22283 ) ;
  assign n22285 = n22278 & n22279 ;
  assign n22286 = ( ~n22271 & n22284 ) | ( ~n22271 & n22285 ) | ( n22284 & n22285 ) ;
  assign n22287 = ~x2 & n22286 ;
  assign n22288 = x2 | n22286 ;
  assign n22289 = ( ~n22286 & n22287 ) | ( ~n22286 & n22288 ) | ( n22287 & n22288 ) ;
  assign n22290 = ~n22266 & n22289 ;
  assign n22291 = n22266 & ~n22289 ;
  assign n22292 = n22290 | n22291 ;
  assign n22293 = ~n20728 & n21408 ;
  assign n22294 = n20728 & ~n21408 ;
  assign n22295 = n22293 | n22294 ;
  assign n22296 = ( ~n20643 & n21566 ) | ( ~n20643 & n21578 ) | ( n21566 & n21578 ) ;
  assign n22297 = ( ~n20646 & n21566 ) | ( ~n20646 & n21578 ) | ( n21566 & n21578 ) ;
  assign n22298 = ( ~n18604 & n22296 ) | ( ~n18604 & n22297 ) | ( n22296 & n22297 ) ;
  assign n22299 = n21566 | n21571 ;
  assign n22300 = n21571 | n21578 ;
  assign n22301 = ( ~n20643 & n22299 ) | ( ~n20643 & n22300 ) | ( n22299 & n22300 ) ;
  assign n22302 = ( ~n20646 & n22299 ) | ( ~n20646 & n22300 ) | ( n22299 & n22300 ) ;
  assign n22303 = ( ~n18604 & n22301 ) | ( ~n18604 & n22302 ) | ( n22301 & n22302 ) ;
  assign n22304 = ~n22298 & n22303 ;
  assign n22305 = n9475 & ~n21563 ;
  assign n22306 = n9021 & ~n20618 ;
  assign n22307 = n9024 & n20609 ;
  assign n22308 = n22306 | n22307 ;
  assign n22309 = n22305 | n22308 ;
  assign n22310 = n21570 & ~n22309 ;
  assign n22311 = ( n22270 & n22309 ) | ( n22270 & ~n22310 ) | ( n22309 & ~n22310 ) ;
  assign n22312 = n22304 | n22311 ;
  assign n22313 = n8970 | n22305 ;
  assign n22314 = n22308 | n22313 ;
  assign n22315 = n22312 & n22314 ;
  assign n22316 = ~x2 & n22314 ;
  assign n22317 = n22312 & n22316 ;
  assign n22318 = x2 | n22316 ;
  assign n22319 = ( x2 & n22312 ) | ( x2 & n22318 ) | ( n22312 & n22318 ) ;
  assign n22320 = ( ~n22315 & n22317 ) | ( ~n22315 & n22319 ) | ( n22317 & n22319 ) ;
  assign n22321 = ~n22295 & n22320 ;
  assign n22322 = n22295 & ~n22320 ;
  assign n22323 = n22321 | n22322 ;
  assign n22324 = n20749 & n21406 ;
  assign n22325 = n20749 | n21406 ;
  assign n22326 = ~n22324 & n22325 ;
  assign n22328 = n9021 & ~n20630 ;
  assign n22329 = n9024 & ~n20618 ;
  assign n22330 = n22328 | n22329 ;
  assign n22327 = n9475 & n20609 ;
  assign n22332 = n8970 | n22327 ;
  assign n22333 = n22330 | n22332 ;
  assign n22331 = n22327 | n22330 ;
  assign n22334 = n22331 & n22333 ;
  assign n22335 = ( n20659 & n22333 ) | ( n20659 & n22334 ) | ( n22333 & n22334 ) ;
  assign n22336 = n22333 & n22334 ;
  assign n22337 = ( ~n20649 & n22335 ) | ( ~n20649 & n22336 ) | ( n22335 & n22336 ) ;
  assign n22338 = x2 & n22337 ;
  assign n22339 = x2 & ~n22337 ;
  assign n22340 = ( n22337 & ~n22338 ) | ( n22337 & n22339 ) | ( ~n22338 & n22339 ) ;
  assign n22341 = n22326 & n22340 ;
  assign n22342 = n22326 | n22340 ;
  assign n22343 = ~n22341 & n22342 ;
  assign n22344 = ~n20771 & n21404 ;
  assign n22345 = n20771 & ~n21404 ;
  assign n22346 = n22344 | n22345 ;
  assign n22347 = n9475 & ~n20618 ;
  assign n22348 = n9021 & n19631 ;
  assign n22349 = n9024 & ~n20630 ;
  assign n22350 = n22348 | n22349 ;
  assign n22351 = n22347 | n22350 ;
  assign n22352 = n20680 | n22351 ;
  assign n22353 = n8970 | n22347 ;
  assign n22354 = n22350 | n22353 ;
  assign n22355 = n20689 & n22354 ;
  assign n22356 = ( n22352 & n22354 ) | ( n22352 & n22355 ) | ( n22354 & n22355 ) ;
  assign n22357 = ~x2 & n22356 ;
  assign n22358 = x2 | n22356 ;
  assign n22359 = ( ~n22356 & n22357 ) | ( ~n22356 & n22358 ) | ( n22357 & n22358 ) ;
  assign n22360 = ~n22346 & n22359 ;
  assign n22361 = n22346 & ~n22359 ;
  assign n22362 = n22360 | n22361 ;
  assign n22363 = ~n22360 & n22362 ;
  assign n22364 = n22343 & ~n22363 ;
  assign n22365 = n22341 | n22364 ;
  assign n22366 = ~n22323 & n22365 ;
  assign n22367 = n22321 | n22366 ;
  assign n22368 = ~n22292 & n22367 ;
  assign n22369 = n21625 | n22360 ;
  assign n22370 = ( n22360 & ~n22362 ) | ( n22360 & n22369 ) | ( ~n22362 & n22369 ) ;
  assign n22371 = n22343 & n22370 ;
  assign n22372 = n22341 | n22371 ;
  assign n22373 = ~n22323 & n22372 ;
  assign n22374 = n22321 | n22373 ;
  assign n22375 = ~n22292 & n22374 ;
  assign n22376 = ( n22264 & n22368 ) | ( n22264 & n22375 ) | ( n22368 & n22375 ) ;
  assign n22377 = n21605 & n22290 ;
  assign n22378 = ( n21605 & n22376 ) | ( n21605 & n22377 ) | ( n22376 & n22377 ) ;
  assign n22379 = n21605 | n22290 ;
  assign n22380 = n22376 | n22379 ;
  assign n22381 = ~n22378 & n22380 ;
  assign n22382 = n22292 & ~n22367 ;
  assign n22383 = n22292 & ~n22374 ;
  assign n22384 = ( ~n22264 & n22382 ) | ( ~n22264 & n22383 ) | ( n22382 & n22383 ) ;
  assign n22385 = n22376 | n22384 ;
  assign n22386 = n22381 & ~n22385 ;
  assign n22387 = ~n22381 & n22385 ;
  assign n22388 = n22386 | n22387 ;
  assign n22389 = ( n22264 & n22364 ) | ( n22264 & n22371 ) | ( n22364 & n22371 ) ;
  assign n22390 = n22343 | n22370 ;
  assign n22391 = ~n22343 & n22363 ;
  assign n22392 = ( n22264 & n22390 ) | ( n22264 & ~n22391 ) | ( n22390 & ~n22391 ) ;
  assign n22393 = ~n22389 & n22392 ;
  assign n22394 = ( n22264 & n22366 ) | ( n22264 & n22373 ) | ( n22366 & n22373 ) ;
  assign n22395 = n22323 & ~n22365 ;
  assign n22396 = n22323 & ~n22372 ;
  assign n22397 = ( ~n22264 & n22395 ) | ( ~n22264 & n22396 ) | ( n22395 & n22396 ) ;
  assign n22398 = n22394 | n22397 ;
  assign n22399 = n22393 & ~n22398 ;
  assign n22400 = ~n22393 & n22398 ;
  assign n22401 = n22399 | n22400 ;
  assign n22402 = n21625 & ~n22362 ;
  assign n22403 = ( n22264 & ~n22362 ) | ( n22264 & n22402 ) | ( ~n22362 & n22402 ) ;
  assign n22404 = ~n21625 & n22362 ;
  assign n22405 = ~n22264 & n22404 ;
  assign n22406 = n22403 | n22405 ;
  assign n22407 = n21628 & ~n22262 ;
  assign n22408 = ~n22260 & n22407 ;
  assign n22409 = n22264 | n22408 ;
  assign n22410 = ~n22393 & n22409 ;
  assign n22411 = n22406 | n22410 ;
  assign n22412 = n22401 | n22411 ;
  assign n22413 = n22385 | n22398 ;
  assign n22414 = n22385 & n22398 ;
  assign n22415 = n22413 & ~n22414 ;
  assign n22416 = n22399 & n22415 ;
  assign n22417 = ( ~n22412 & n22415 ) | ( ~n22412 & n22416 ) | ( n22415 & n22416 ) ;
  assign n22418 = n22388 | n22413 ;
  assign n22419 = ( n22388 & ~n22417 ) | ( n22388 & n22418 ) | ( ~n22417 & n22418 ) ;
  assign n22420 = n22388 & n22413 ;
  assign n22421 = ~n22417 & n22420 ;
  assign n22422 = n22419 & ~n22421 ;
  assign n22423 = n1829 & n22381 ;
  assign n22424 = n1826 & ~n22398 ;
  assign n22425 = n1823 & ~n22385 ;
  assign n22426 = n22424 | n22425 ;
  assign n22427 = n22423 | n22426 ;
  assign n22428 = n1821 | n22427 ;
  assign n22429 = x29 & n22428 ;
  assign n22430 = x29 & n22427 ;
  assign n22431 = ( n22422 & n22429 ) | ( n22422 & n22430 ) | ( n22429 & n22430 ) ;
  assign n22432 = x29 | n22428 ;
  assign n22433 = x29 | n22427 ;
  assign n22434 = ( n22422 & n22432 ) | ( n22422 & n22433 ) | ( n22432 & n22433 ) ;
  assign n22435 = ~n22431 & n22434 ;
  assign n22436 = ~n22406 & n22409 ;
  assign n22437 = ~n22393 & n22436 ;
  assign n22438 = n22393 & ~n22436 ;
  assign n22439 = n22437 | n22438 ;
  assign n22440 = n1062 & n22439 ;
  assign n22441 = n1057 & n22393 ;
  assign n22442 = n1060 & ~n22409 ;
  assign n22443 = n1065 & ~n22406 ;
  assign n22444 = n22442 | n22443 ;
  assign n22445 = n22441 | n22444 ;
  assign n22446 = n22440 | n22445 ;
  assign n22447 = n1162 | n1186 ;
  assign n22448 = n159 | n511 ;
  assign n22449 = n263 | n22448 ;
  assign n22450 = n118 | n491 ;
  assign n22451 = n8052 | n22450 ;
  assign n22452 = n22449 | n22451 ;
  assign n22453 = n18475 | n22452 ;
  assign n22454 = n372 | n1637 ;
  assign n22455 = n16925 | n22454 ;
  assign n22456 = ( ~n1186 & n22453 ) | ( ~n1186 & n22455 ) | ( n22453 & n22455 ) ;
  assign n22457 = n22453 & n22455 ;
  assign n22458 = ( ~n1162 & n22456 ) | ( ~n1162 & n22457 ) | ( n22456 & n22457 ) ;
  assign n22459 = n22447 | n22458 ;
  assign n22460 = n1104 & ~n4287 ;
  assign n22461 = n1380 | n3467 ;
  assign n22462 = n22460 & ~n22461 ;
  assign n22463 = ~n2053 & n22462 ;
  assign n22464 = ~n22459 & n22463 ;
  assign n22465 = n176 | n594 ;
  assign n22466 = n226 | n527 ;
  assign n22467 = n22465 | n22466 ;
  assign n22468 = n381 | n22467 ;
  assign n22469 = n209 | n17724 ;
  assign n22470 = n17723 | n22469 ;
  assign n22471 = n22468 | n22470 ;
  assign n22472 = n22464 & ~n22471 ;
  assign n22473 = n22406 & ~n22409 ;
  assign n22474 = n22436 | n22473 ;
  assign n22475 = ( n1062 & n10826 ) | ( n1062 & ~n22409 ) | ( n10826 & ~n22409 ) ;
  assign n22476 = n17723 | n17724 ;
  assign n22477 = n926 & ~n8983 ;
  assign n22478 = ~n8990 & n22477 ;
  assign n22479 = ~n15914 & n22478 ;
  assign n22480 = n71 | n83 ;
  assign n22481 = n240 | n395 ;
  assign n22482 = n22480 | n22481 ;
  assign n22483 = n118 | n159 ;
  assign n22484 = n783 | n22483 ;
  assign n22485 = n22482 | n22484 ;
  assign n22486 = n22479 & ~n22485 ;
  assign n22487 = n1034 | n12387 ;
  assign n22488 = n952 | n966 ;
  assign n22489 = n22487 | n22488 ;
  assign n22490 = n2156 | n22489 ;
  assign n22491 = n22486 & ~n22490 ;
  assign n22492 = n1447 | n1742 ;
  assign n22493 = n264 | n2233 ;
  assign n22494 = n22492 | n22493 ;
  assign n22495 = n292 | n388 ;
  assign n22496 = n3425 | n22495 ;
  assign n22497 = n22494 | n22496 ;
  assign n22498 = n594 | n725 ;
  assign n22499 = n226 | n349 ;
  assign n22500 = n22498 | n22499 ;
  assign n22501 = n363 | n22500 ;
  assign n22502 = n22497 | n22501 ;
  assign n22503 = n478 | n2246 ;
  assign n22504 = n4253 | n22503 ;
  assign n22505 = n447 | n12269 ;
  assign n22506 = n141 | n237 ;
  assign n22507 = n203 | n312 ;
  assign n22508 = n22506 | n22507 ;
  assign n22509 = n22505 | n22508 ;
  assign n22510 = n22504 | n22509 ;
  assign n22511 = n22502 | n22510 ;
  assign n22512 = n22491 & ~n22511 ;
  assign n22513 = ~n22476 & n22512 ;
  assign n22514 = n1307 | n3430 ;
  assign n22515 = n550 | n748 ;
  assign n22516 = n22514 | n22515 ;
  assign n22517 = ~n153 & n15199 ;
  assign n22518 = ~n15199 & n22517 ;
  assign n22519 = ( n153 & n1005 ) | ( n153 & ~n15199 ) | ( n1005 & ~n15199 ) ;
  assign n22520 = n15199 | n22519 ;
  assign n22521 = ( n22516 & ~n22518 ) | ( n22516 & n22520 ) | ( ~n22518 & n22520 ) ;
  assign n22522 = n160 | n22521 ;
  assign n22523 = n305 | n491 ;
  assign n22524 = n22522 | n22523 ;
  assign n22525 = n22513 & ~n22524 ;
  assign n22526 = n1057 & ~n22525 ;
  assign n22527 = ~n22406 & n22526 ;
  assign n22528 = ( n22475 & ~n22525 ) | ( n22475 & n22527 ) | ( ~n22525 & n22527 ) ;
  assign n22529 = n1065 & ~n22409 ;
  assign n22530 = ( ~n22525 & n22527 ) | ( ~n22525 & n22529 ) | ( n22527 & n22529 ) ;
  assign n22531 = ( n22474 & n22528 ) | ( n22474 & n22530 ) | ( n22528 & n22530 ) ;
  assign n22532 = ~n22472 & n22531 ;
  assign n22533 = n22472 & ~n22531 ;
  assign n22534 = n22532 | n22533 ;
  assign n22535 = n22446 & ~n22534 ;
  assign n22536 = n22446 & ~n22535 ;
  assign n22537 = n22534 | n22535 ;
  assign n22538 = ~n22536 & n22537 ;
  assign n22539 = n22435 & ~n22538 ;
  assign n22540 = n22435 & ~n22539 ;
  assign n22541 = n22435 | n22538 ;
  assign n22542 = ~n22540 & n22541 ;
  assign n22543 = n22399 | n22415 ;
  assign n22544 = n22412 & ~n22543 ;
  assign n22545 = n22417 | n22544 ;
  assign n22546 = n1826 & n22393 ;
  assign n22547 = n1823 & ~n22398 ;
  assign n22548 = n22546 | n22547 ;
  assign n22549 = n1829 & ~n22385 ;
  assign n22550 = n1821 | n22549 ;
  assign n22551 = n22548 | n22550 ;
  assign n22552 = ~x29 & n22551 ;
  assign n22553 = n22548 | n22549 ;
  assign n22554 = ~x29 & n22553 ;
  assign n22555 = ( ~n22545 & n22552 ) | ( ~n22545 & n22554 ) | ( n22552 & n22554 ) ;
  assign n22556 = x29 & n22551 ;
  assign n22557 = x29 & ~n22556 ;
  assign n22558 = x29 & n22549 ;
  assign n22559 = ( x29 & n22548 ) | ( x29 & n22558 ) | ( n22548 & n22558 ) ;
  assign n22560 = x29 & ~n22559 ;
  assign n22561 = ( n22545 & n22557 ) | ( n22545 & n22560 ) | ( n22557 & n22560 ) ;
  assign n22562 = n22555 | n22561 ;
  assign n22563 = n1057 & ~n22406 ;
  assign n22564 = n22475 | n22563 ;
  assign n22565 = n22529 | n22563 ;
  assign n22566 = ( n22474 & n22564 ) | ( n22474 & n22565 ) | ( n22564 & n22565 ) ;
  assign n22567 = n22525 | n22566 ;
  assign n22568 = ~n22525 & n22566 ;
  assign n22569 = ( ~n22566 & n22567 ) | ( ~n22566 & n22568 ) | ( n22567 & n22568 ) ;
  assign n22570 = n22562 & ~n22569 ;
  assign n22571 = ~n22562 & n22569 ;
  assign n22572 = n22570 | n22571 ;
  assign n22573 = n2005 & ~n22409 ;
  assign n22574 = n1829 & n22393 ;
  assign n22575 = n1826 & ~n22409 ;
  assign n22576 = n1823 & ~n22406 ;
  assign n22577 = n22575 | n22576 ;
  assign n22578 = n22574 | n22577 ;
  assign n22579 = n22439 | n22578 ;
  assign n22580 = n1821 | n22574 ;
  assign n22581 = n22577 | n22580 ;
  assign n22582 = n22579 & n22581 ;
  assign n22583 = ~x29 & n22581 ;
  assign n22584 = n22579 & n22583 ;
  assign n22585 = x29 | n22584 ;
  assign n22586 = ( ~n22582 & n22584 ) | ( ~n22582 & n22585 ) | ( n22584 & n22585 ) ;
  assign n22587 = n1821 & n22474 ;
  assign n22588 = n1823 & ~n22409 ;
  assign n22589 = n1829 & ~n22406 ;
  assign n22590 = n22588 | n22589 ;
  assign n22591 = x29 | n22590 ;
  assign n22592 = n22587 | n22591 ;
  assign n22593 = ~x29 & n22592 ;
  assign n22594 = ( x29 & n11040 ) | ( x29 & n22409 ) | ( n11040 & n22409 ) ;
  assign n22595 = n22592 & n22594 ;
  assign n22596 = n22587 | n22590 ;
  assign n22597 = n22594 & ~n22596 ;
  assign n22598 = ( n22593 & n22595 ) | ( n22593 & n22597 ) | ( n22595 & n22597 ) ;
  assign n22599 = ~n22573 & n22598 ;
  assign n22600 = n22586 & n22599 ;
  assign n22601 = n22573 | n22600 ;
  assign n22602 = n1829 & ~n22398 ;
  assign n22603 = n1826 & ~n22406 ;
  assign n22604 = n1823 & n22393 ;
  assign n22605 = n22603 | n22604 ;
  assign n22606 = n22602 | n22605 ;
  assign n22607 = n22401 & n22411 ;
  assign n22608 = n22412 & ~n22607 ;
  assign n22609 = n1821 | n22602 ;
  assign n22610 = n22605 | n22609 ;
  assign n22611 = ( n22606 & n22608 ) | ( n22606 & n22610 ) | ( n22608 & n22610 ) ;
  assign n22612 = x29 & n22610 ;
  assign n22613 = x29 & n22606 ;
  assign n22614 = ( n22608 & n22612 ) | ( n22608 & n22613 ) | ( n22612 & n22613 ) ;
  assign n22615 = x29 & ~n22614 ;
  assign n22616 = ( n22611 & ~n22614 ) | ( n22611 & n22615 ) | ( ~n22614 & n22615 ) ;
  assign n22617 = n22600 & n22616 ;
  assign n22618 = n22586 & n22598 ;
  assign n22619 = n22616 & ~n22618 ;
  assign n22620 = ( n22601 & n22617 ) | ( n22601 & n22619 ) | ( n22617 & n22619 ) ;
  assign n22621 = n22573 & n22584 ;
  assign n22622 = n22573 & ~n22582 ;
  assign n22623 = ( n22585 & n22621 ) | ( n22585 & n22622 ) | ( n22621 & n22622 ) ;
  assign n22624 = n22598 & n22623 ;
  assign n22625 = ~n22572 & n22624 ;
  assign n22626 = ( ~n22572 & n22620 ) | ( ~n22572 & n22625 ) | ( n22620 & n22625 ) ;
  assign n22627 = n22570 | n22626 ;
  assign n22628 = n22542 & ~n22627 ;
  assign n22629 = ~n22542 & n22627 ;
  assign n22630 = n22628 | n22629 ;
  assign n22859 = n19663 | n20342 ;
  assign n22860 = ( n19663 & n19666 ) | ( n19663 & n22859 ) | ( n19666 & n22859 ) ;
  assign n22807 = n18067 | n18070 ;
  assign n22808 = ( n17658 & n18067 ) | ( n17658 & n22807 ) | ( n18067 & n22807 ) ;
  assign n22631 = n306 | n497 ;
  assign n22632 = n689 | n22631 ;
  assign n22633 = n1436 | n4180 ;
  assign n22634 = n18452 | n22633 ;
  assign n22635 = n17903 | n22634 ;
  assign n22636 = n18472 | n22635 ;
  assign n22637 = n1518 | n6813 ;
  assign n22638 = n1505 | n22637 ;
  assign n22639 = n1418 | n2188 ;
  assign n22640 = n1301 | n2809 ;
  assign n22641 = n22639 | n22640 ;
  assign n22642 = n10803 | n22641 ;
  assign n22643 = n450 | n574 ;
  assign n22644 = n510 | n22643 ;
  assign n22645 = n22642 | n22644 ;
  assign n22646 = n22638 | n22645 ;
  assign n22647 = n22636 | n22646 ;
  assign n22648 = n22632 | n22647 ;
  assign n22649 = n1057 & n11363 ;
  assign n22650 = n1065 & n10649 ;
  assign n22651 = n1060 & n10325 ;
  assign n22652 = n22650 | n22651 ;
  assign n22653 = n22649 | n22652 ;
  assign n22654 = n22648 & n22653 ;
  assign n22655 = n1062 | n22652 ;
  assign n22656 = n22648 & n22649 ;
  assign n22657 = ( n22648 & n22655 ) | ( n22648 & n22656 ) | ( n22655 & n22656 ) ;
  assign n22658 = ( n12059 & n22654 ) | ( n12059 & n22657 ) | ( n22654 & n22657 ) ;
  assign n22659 = n22649 | n22655 ;
  assign n22660 = ( n12059 & n22653 ) | ( n12059 & n22659 ) | ( n22653 & n22659 ) ;
  assign n22661 = ~n22658 & n22660 ;
  assign n22662 = n22648 & ~n22659 ;
  assign n22663 = n22648 & ~n22653 ;
  assign n22664 = ( ~n12059 & n22662 ) | ( ~n12059 & n22663 ) | ( n22662 & n22663 ) ;
  assign n22665 = n22661 | n22664 ;
  assign n22666 = n17741 | n17744 ;
  assign n22667 = ( n17741 & n17746 ) | ( n17741 & n22666 ) | ( n17746 & n22666 ) ;
  assign n22668 = n22665 & n22667 ;
  assign n22669 = n22665 | n22667 ;
  assign n22670 = ~n22668 & n22669 ;
  assign n22672 = n1826 & ~n11663 ;
  assign n22673 = n1823 & n12010 ;
  assign n22674 = n22672 | n22673 ;
  assign n22671 = n1829 & ~n12616 ;
  assign n22676 = n1821 | n22671 ;
  assign n22677 = n22674 | n22676 ;
  assign n22675 = n22671 | n22674 ;
  assign n22678 = n22675 & n22677 ;
  assign n22679 = ( ~n12626 & n22677 ) | ( ~n12626 & n22678 ) | ( n22677 & n22678 ) ;
  assign n22680 = ~x29 & n22678 ;
  assign n22681 = ~x29 & n22677 ;
  assign n22682 = ( ~n12626 & n22680 ) | ( ~n12626 & n22681 ) | ( n22680 & n22681 ) ;
  assign n22683 = x29 | n22680 ;
  assign n22684 = x29 | n22681 ;
  assign n22685 = ( ~n12626 & n22683 ) | ( ~n12626 & n22684 ) | ( n22683 & n22684 ) ;
  assign n22686 = ( ~n22679 & n22682 ) | ( ~n22679 & n22685 ) | ( n22682 & n22685 ) ;
  assign n22687 = n22670 & n22686 ;
  assign n22688 = n22670 | n22686 ;
  assign n22689 = ~n22687 & n22688 ;
  assign n22690 = n17765 & n22689 ;
  assign n22691 = ( n17770 & n22689 ) | ( n17770 & n22690 ) | ( n22689 & n22690 ) ;
  assign n22692 = n17765 | n22689 ;
  assign n22693 = n17770 | n22692 ;
  assign n22694 = ~n22691 & n22693 ;
  assign n22695 = n2312 & n12936 ;
  assign n22696 = n2308 & n13235 ;
  assign n22697 = n22695 | n22696 ;
  assign n22698 = n2315 & n13522 ;
  assign n22699 = n2306 | n22698 ;
  assign n22700 = n22697 | n22699 ;
  assign n22701 = n22697 | n22698 ;
  assign n22702 = n13537 | n22701 ;
  assign n22703 = n13539 | n22701 ;
  assign n22704 = ( ~n13248 & n22702 ) | ( ~n13248 & n22703 ) | ( n22702 & n22703 ) ;
  assign n22705 = n22700 & n22704 ;
  assign n22706 = ( n13530 & n22700 ) | ( n13530 & n22705 ) | ( n22700 & n22705 ) ;
  assign n22707 = ~x26 & n22706 ;
  assign n22708 = x26 | n22706 ;
  assign n22709 = ( ~n22706 & n22707 ) | ( ~n22706 & n22708 ) | ( n22707 & n22708 ) ;
  assign n22710 = n22694 & n22709 ;
  assign n22711 = n22694 & ~n22710 ;
  assign n22712 = ~n22694 & n22709 ;
  assign n22713 = n22711 | n22712 ;
  assign n22714 = n17790 | n17793 ;
  assign n22715 = ( n17790 & n17795 ) | ( n17790 & n22714 ) | ( n17795 & n22714 ) ;
  assign n22716 = n22713 & ~n22715 ;
  assign n22717 = ~n22713 & n22715 ;
  assign n22718 = n22716 | n22717 ;
  assign n22719 = n2932 & n14591 ;
  assign n22720 = n2925 & n14607 ;
  assign n22721 = n2928 & n14329 ;
  assign n22722 = n22720 | n22721 ;
  assign n22723 = n22719 | n22722 ;
  assign n22724 = n2936 | n22719 ;
  assign n22725 = n22722 | n22724 ;
  assign n22726 = ( n14629 & n22723 ) | ( n14629 & n22725 ) | ( n22723 & n22725 ) ;
  assign n22727 = x23 & n22725 ;
  assign n22728 = x23 & n22723 ;
  assign n22729 = ( n14629 & n22727 ) | ( n14629 & n22728 ) | ( n22727 & n22728 ) ;
  assign n22730 = x23 & ~n22728 ;
  assign n22731 = x23 & ~n22727 ;
  assign n22732 = ( ~n14629 & n22730 ) | ( ~n14629 & n22731 ) | ( n22730 & n22731 ) ;
  assign n22733 = ( n22726 & ~n22729 ) | ( n22726 & n22732 ) | ( ~n22729 & n22732 ) ;
  assign n22734 = n22718 & n22733 ;
  assign n22735 = n22718 | n22733 ;
  assign n22736 = ~n22734 & n22735 ;
  assign n22737 = n17814 | n17816 ;
  assign n22738 = ( n17814 & n17818 ) | ( n17814 & n22737 ) | ( n17818 & n22737 ) ;
  assign n22739 = n22736 & n22738 ;
  assign n22740 = n22736 | n22738 ;
  assign n22741 = ~n22739 & n22740 ;
  assign n22743 = n3544 & n15434 ;
  assign n22744 = n3541 & ~n16085 ;
  assign n22745 = n22743 | n22744 ;
  assign n22742 = n3547 & n15886 ;
  assign n22747 = n3537 | n22742 ;
  assign n22748 = n22745 | n22747 ;
  assign n22746 = n22742 | n22745 ;
  assign n22749 = n22746 & n22748 ;
  assign n22750 = ( ~n16140 & n22748 ) | ( ~n16140 & n22749 ) | ( n22748 & n22749 ) ;
  assign n22751 = ~x20 & n22749 ;
  assign n22752 = ~x20 & n22748 ;
  assign n22753 = ( ~n16140 & n22751 ) | ( ~n16140 & n22752 ) | ( n22751 & n22752 ) ;
  assign n22754 = x20 | n22751 ;
  assign n22755 = x20 | n22752 ;
  assign n22756 = ( ~n16140 & n22754 ) | ( ~n16140 & n22755 ) | ( n22754 & n22755 ) ;
  assign n22757 = ( ~n22750 & n22753 ) | ( ~n22750 & n22756 ) | ( n22753 & n22756 ) ;
  assign n22758 = n22741 & n22757 ;
  assign n22759 = n22741 & ~n22758 ;
  assign n22760 = ~n22741 & n22757 ;
  assign n22761 = n22759 | n22760 ;
  assign n22762 = n17838 | n17841 ;
  assign n22763 = ( n17838 & n17843 ) | ( n17838 & n22762 ) | ( n17843 & n22762 ) ;
  assign n22764 = n22761 & ~n22763 ;
  assign n22765 = ~n22761 & n22763 ;
  assign n22766 = n22764 | n22765 ;
  assign n22767 = n4471 & n17100 ;
  assign n22768 = n4466 & ~n16069 ;
  assign n22769 = n4468 & n17111 ;
  assign n22770 = n22768 | n22769 ;
  assign n22771 = n22767 | n22770 ;
  assign n22772 = n4475 & n17169 ;
  assign n22773 = ~n17129 & n22772 ;
  assign n22774 = n22771 | n22773 ;
  assign n22775 = n4475 | n22771 ;
  assign n22776 = ( n17161 & n22774 ) | ( n17161 & n22775 ) | ( n22774 & n22775 ) ;
  assign n22777 = x17 | n22776 ;
  assign n22778 = ~x17 & n22776 ;
  assign n22779 = ( ~n22776 & n22777 ) | ( ~n22776 & n22778 ) | ( n22777 & n22778 ) ;
  assign n22780 = n22766 & n22779 ;
  assign n22781 = n22766 | n22779 ;
  assign n22782 = ~n22780 & n22781 ;
  assign n22783 = n17860 & n22782 ;
  assign n22784 = ( n17864 & n22782 ) | ( n17864 & n22783 ) | ( n22782 & n22783 ) ;
  assign n22785 = n17860 | n22782 ;
  assign n22786 = n17864 | n22785 ;
  assign n22787 = ~n22784 & n22786 ;
  assign n22788 = n5234 & ~n18585 ;
  assign n22789 = n5237 & ~n17092 ;
  assign n22790 = n5231 & n18037 ;
  assign n22791 = n22789 | n22790 ;
  assign n22792 = n22788 | n22791 ;
  assign n22793 = n18675 & ~n22792 ;
  assign n22794 = ~n18672 & n22793 ;
  assign n22795 = n5227 | n22788 ;
  assign n22796 = n22791 | n22795 ;
  assign n22797 = ~n22794 & n22796 ;
  assign n22798 = x14 & n22796 ;
  assign n22799 = ~n22794 & n22798 ;
  assign n22800 = x14 & ~n22798 ;
  assign n22801 = ( x14 & n22794 ) | ( x14 & n22800 ) | ( n22794 & n22800 ) ;
  assign n22802 = ( n22797 & ~n22799 ) | ( n22797 & n22801 ) | ( ~n22799 & n22801 ) ;
  assign n22803 = n22787 & n22802 ;
  assign n22804 = n22787 & ~n22803 ;
  assign n22805 = ~n22787 & n22802 ;
  assign n22806 = n22804 | n22805 ;
  assign n22809 = n22806 & n22808 ;
  assign n22810 = n22808 & ~n22809 ;
  assign n22811 = n22806 & ~n22808 ;
  assign n22812 = n22810 | n22811 ;
  assign n22813 = n6122 & n19352 ;
  assign n22814 = n6125 & n18410 ;
  assign n22815 = n6119 & n18576 ;
  assign n22816 = n22814 | n22815 ;
  assign n22817 = n22813 | n22816 ;
  assign n22818 = n6115 | n22813 ;
  assign n22819 = n22816 | n22818 ;
  assign n22820 = ( n19674 & n22817 ) | ( n19674 & n22819 ) | ( n22817 & n22819 ) ;
  assign n22821 = x11 & n22819 ;
  assign n22822 = x11 & n22817 ;
  assign n22823 = ( n19674 & n22821 ) | ( n19674 & n22822 ) | ( n22821 & n22822 ) ;
  assign n22824 = x11 & ~n22822 ;
  assign n22825 = x11 & ~n22821 ;
  assign n22826 = ( ~n19674 & n22824 ) | ( ~n19674 & n22825 ) | ( n22824 & n22825 ) ;
  assign n22827 = ( n22820 & ~n22823 ) | ( n22820 & n22826 ) | ( ~n22823 & n22826 ) ;
  assign n22828 = n22811 & n22827 ;
  assign n22829 = ( n22810 & n22827 ) | ( n22810 & n22828 ) | ( n22827 & n22828 ) ;
  assign n22830 = n22812 & ~n22829 ;
  assign n22831 = ~n22811 & n22827 ;
  assign n22832 = ~n22810 & n22831 ;
  assign n22833 = n22830 | n22832 ;
  assign n22834 = n18629 | n19227 ;
  assign n22835 = ( n18629 & n18633 ) | ( n18629 & n22834 ) | ( n18633 & n22834 ) ;
  assign n22836 = n22833 & n22835 ;
  assign n22837 = n22833 | n22835 ;
  assign n22838 = ~n22836 & n22837 ;
  assign n22840 = n7074 & n19494 ;
  assign n22841 = n7068 & n19631 ;
  assign n22842 = n22840 | n22841 ;
  assign n22839 = n7079 & ~n20630 ;
  assign n22844 = n7078 | n22839 ;
  assign n22845 = n22842 | n22844 ;
  assign n22843 = n22839 | n22842 ;
  assign n22846 = n22843 & n22845 ;
  assign n22847 = ( ~n20709 & n22845 ) | ( ~n20709 & n22846 ) | ( n22845 & n22846 ) ;
  assign n22848 = ~x8 & n22846 ;
  assign n22849 = ~x8 & n22845 ;
  assign n22850 = ( ~n20709 & n22848 ) | ( ~n20709 & n22849 ) | ( n22848 & n22849 ) ;
  assign n22851 = x8 | n22848 ;
  assign n22852 = x8 | n22849 ;
  assign n22853 = ( ~n20709 & n22851 ) | ( ~n20709 & n22852 ) | ( n22851 & n22852 ) ;
  assign n22854 = ( ~n22847 & n22850 ) | ( ~n22847 & n22853 ) | ( n22850 & n22853 ) ;
  assign n22855 = n22838 & n22854 ;
  assign n22856 = n22838 & ~n22855 ;
  assign n22857 = ~n22838 & n22854 ;
  assign n22858 = n22856 | n22857 ;
  assign n22861 = n22858 & n22860 ;
  assign n22862 = n22860 & ~n22861 ;
  assign n22863 = n22858 & ~n22861 ;
  assign n22864 = n22862 | n22863 ;
  assign n22865 = n8122 & ~n21563 ;
  assign n22866 = n8115 & ~n20618 ;
  assign n22867 = n8118 & n20609 ;
  assign n22868 = n22866 | n22867 ;
  assign n22869 = n22865 | n22868 ;
  assign n22870 = n8125 & ~n21570 ;
  assign n22871 = n22270 & n22870 ;
  assign n22872 = ( n8125 & n22304 ) | ( n8125 & n22871 ) | ( n22304 & n22871 ) ;
  assign n22873 = n22869 | n22872 ;
  assign n22874 = x5 | n22869 ;
  assign n22875 = n22872 | n22874 ;
  assign n22876 = ~x5 & n22874 ;
  assign n22877 = ( ~x5 & n22872 ) | ( ~x5 & n22876 ) | ( n22872 & n22876 ) ;
  assign n22878 = ( ~n22873 & n22875 ) | ( ~n22873 & n22877 ) | ( n22875 & n22877 ) ;
  assign n22879 = n22864 & n22878 ;
  assign n22880 = n22864 & ~n22879 ;
  assign n22881 = ~n22864 & n22878 ;
  assign n22882 = n22880 | n22881 ;
  assign n22883 = n20669 | n21413 ;
  assign n22884 = n22882 & n22883 ;
  assign n22885 = n22855 | n22861 ;
  assign n22886 = n1829 & n12936 ;
  assign n22887 = n1826 & n12010 ;
  assign n22888 = n1823 & ~n12616 ;
  assign n22889 = n22887 | n22888 ;
  assign n22890 = n22886 | n22889 ;
  assign n22891 = n1821 | n22886 ;
  assign n22892 = n22889 | n22891 ;
  assign n22893 = ( ~n13591 & n22890 ) | ( ~n13591 & n22892 ) | ( n22890 & n22892 ) ;
  assign n22894 = ~x29 & n22892 ;
  assign n22895 = ~x29 & n22890 ;
  assign n22896 = ( ~n13591 & n22894 ) | ( ~n13591 & n22895 ) | ( n22894 & n22895 ) ;
  assign n22897 = x29 | n22895 ;
  assign n22898 = x29 | n22894 ;
  assign n22899 = ( ~n13591 & n22897 ) | ( ~n13591 & n22898 ) | ( n22897 & n22898 ) ;
  assign n22900 = ( ~n22893 & n22896 ) | ( ~n22893 & n22899 ) | ( n22896 & n22899 ) ;
  assign n22901 = n535 | n7929 ;
  assign n22902 = n2880 | n3465 ;
  assign n22903 = n22901 | n22902 ;
  assign n22904 = n805 | n22903 ;
  assign n22905 = n2861 | n22904 ;
  assign n22906 = n2147 | n22905 ;
  assign n22907 = n230 | n389 ;
  assign n22908 = n307 | n22907 ;
  assign n22909 = n10772 | n18447 ;
  assign n22910 = n22908 | n22909 ;
  assign n22911 = n2869 | n22910 ;
  assign n22912 = n96 | n343 ;
  assign n22913 = n4048 | n22912 ;
  assign n22914 = n513 | n1469 ;
  assign n22915 = n22913 | n22914 ;
  assign n22916 = n296 | n22915 ;
  assign n22917 = n1692 | n2146 ;
  assign n22918 = n209 | n654 ;
  assign n22919 = n213 | n22918 ;
  assign n22920 = n22917 | n22919 ;
  assign n22921 = n141 | n225 ;
  assign n22922 = n1723 | n22921 ;
  assign n22923 = n22920 | n22922 ;
  assign n22924 = n22916 | n22923 ;
  assign n22925 = n22911 | n22924 ;
  assign n22926 = n262 | n581 ;
  assign n22927 = n518 | n895 ;
  assign n22928 = n22926 | n22927 ;
  assign n22929 = n22925 | n22928 ;
  assign n22930 = n2809 | n14392 ;
  assign n22931 = n175 | n2696 ;
  assign n22932 = n205 | n22931 ;
  assign n22933 = n22930 | n22932 ;
  assign n22934 = n197 | n1114 ;
  assign n22935 = n245 | n22934 ;
  assign n22936 = n22933 | n22935 ;
  assign n22937 = n22929 | n22936 ;
  assign n22938 = n22906 | n22937 ;
  assign n22939 = n1057 & ~n11663 ;
  assign n22940 = n1065 & n11363 ;
  assign n22941 = n1060 & n10649 ;
  assign n22942 = n22940 | n22941 ;
  assign n22943 = n22939 | n22942 ;
  assign n22944 = n1062 & ~n12048 ;
  assign n22945 = ~n11672 & n22944 ;
  assign n22946 = n22943 | n22945 ;
  assign n22947 = n1062 | n22943 ;
  assign n22948 = ( n12040 & n22946 ) | ( n12040 & n22947 ) | ( n22946 & n22947 ) ;
  assign n22949 = ~n22938 & n22948 ;
  assign n22950 = n22938 & n22939 ;
  assign n22951 = ( n22938 & n22942 ) | ( n22938 & n22950 ) | ( n22942 & n22950 ) ;
  assign n22952 = ( n22938 & n22945 ) | ( n22938 & n22951 ) | ( n22945 & n22951 ) ;
  assign n22953 = ( n1062 & n22938 ) | ( n1062 & n22951 ) | ( n22938 & n22951 ) ;
  assign n22954 = ( n12040 & n22952 ) | ( n12040 & n22953 ) | ( n22952 & n22953 ) ;
  assign n22955 = ( n22938 & n22949 ) | ( n22938 & ~n22954 ) | ( n22949 & ~n22954 ) ;
  assign n22956 = n22658 | n22665 ;
  assign n22957 = ( n22658 & n22667 ) | ( n22658 & n22956 ) | ( n22667 & n22956 ) ;
  assign n22958 = ~n22955 & n22957 ;
  assign n22959 = n22900 & n22955 ;
  assign n22960 = ~n22957 & n22959 ;
  assign n22961 = ( n22900 & n22958 ) | ( n22900 & n22960 ) | ( n22958 & n22960 ) ;
  assign n22962 = n22900 | n22955 ;
  assign n22963 = ( n22900 & ~n22957 ) | ( n22900 & n22962 ) | ( ~n22957 & n22962 ) ;
  assign n22964 = n22958 | n22963 ;
  assign n22965 = ~n22961 & n22964 ;
  assign n22966 = n22687 & n22965 ;
  assign n22967 = ( n22691 & n22965 ) | ( n22691 & n22966 ) | ( n22965 & n22966 ) ;
  assign n22968 = n22687 | n22965 ;
  assign n22969 = n22691 | n22968 ;
  assign n22970 = ~n22967 & n22969 ;
  assign n22971 = n2312 & n13235 ;
  assign n22972 = n2308 & n13522 ;
  assign n22973 = n22971 | n22972 ;
  assign n22974 = n2315 & n14607 ;
  assign n22975 = n2306 | n22974 ;
  assign n22976 = n22973 | n22975 ;
  assign n22977 = n22973 | n22974 ;
  assign n22978 = n14696 | n22977 ;
  assign n22979 = n14698 | n22977 ;
  assign n22980 = ( ~n13248 & n22978 ) | ( ~n13248 & n22979 ) | ( n22978 & n22979 ) ;
  assign n22981 = n22976 & n22980 ;
  assign n22982 = ( n14687 & n22976 ) | ( n14687 & n22981 ) | ( n22976 & n22981 ) ;
  assign n22983 = ~x26 & n22982 ;
  assign n22984 = x26 | n22982 ;
  assign n22985 = ( ~n22982 & n22983 ) | ( ~n22982 & n22984 ) | ( n22983 & n22984 ) ;
  assign n22986 = n22970 & n22985 ;
  assign n22987 = n22970 & ~n22986 ;
  assign n22988 = ~n22970 & n22985 ;
  assign n22989 = n22987 | n22988 ;
  assign n22990 = n22710 | n22713 ;
  assign n22991 = ( n22710 & n22715 ) | ( n22710 & n22990 ) | ( n22715 & n22990 ) ;
  assign n22992 = n22989 & ~n22991 ;
  assign n22993 = ~n22989 & n22991 ;
  assign n22994 = n22992 | n22993 ;
  assign n22995 = n2932 & n15434 ;
  assign n22996 = n2925 & n14329 ;
  assign n22997 = n2928 & n14591 ;
  assign n22998 = n22996 | n22997 ;
  assign n22999 = n22995 | n22998 ;
  assign n23000 = n2936 | n22995 ;
  assign n23001 = n22998 | n23000 ;
  assign n23002 = ( n15453 & n22999 ) | ( n15453 & n23001 ) | ( n22999 & n23001 ) ;
  assign n23003 = x23 & n23001 ;
  assign n23004 = x23 & n22999 ;
  assign n23005 = ( n15453 & n23003 ) | ( n15453 & n23004 ) | ( n23003 & n23004 ) ;
  assign n23006 = x23 & ~n23004 ;
  assign n23007 = x23 & ~n23003 ;
  assign n23008 = ( ~n15453 & n23006 ) | ( ~n15453 & n23007 ) | ( n23006 & n23007 ) ;
  assign n23009 = ( n23002 & ~n23005 ) | ( n23002 & n23008 ) | ( ~n23005 & n23008 ) ;
  assign n23010 = n22994 & n23009 ;
  assign n23011 = n22994 | n23009 ;
  assign n23012 = ~n23010 & n23011 ;
  assign n23013 = n22734 | n22736 ;
  assign n23014 = ( n22734 & n22738 ) | ( n22734 & n23013 ) | ( n22738 & n23013 ) ;
  assign n23015 = n23012 & n23014 ;
  assign n23016 = n23012 | n23014 ;
  assign n23017 = ~n23015 & n23016 ;
  assign n23018 = n3547 & ~n16069 ;
  assign n23019 = n3544 & ~n16085 ;
  assign n23020 = n3541 & n15886 ;
  assign n23021 = n23019 | n23020 ;
  assign n23022 = n23018 | n23021 ;
  assign n23023 = n3537 | n23022 ;
  assign n23024 = ( ~n16107 & n23022 ) | ( ~n16107 & n23023 ) | ( n23022 & n23023 ) ;
  assign n23025 = ~x20 & n23023 ;
  assign n23026 = ~x20 & n23022 ;
  assign n23027 = ( ~n16107 & n23025 ) | ( ~n16107 & n23026 ) | ( n23025 & n23026 ) ;
  assign n23028 = x20 | n23025 ;
  assign n23029 = x20 | n23026 ;
  assign n23030 = ( ~n16107 & n23028 ) | ( ~n16107 & n23029 ) | ( n23028 & n23029 ) ;
  assign n23031 = ( ~n23024 & n23027 ) | ( ~n23024 & n23030 ) | ( n23027 & n23030 ) ;
  assign n23032 = n23017 & n23031 ;
  assign n23033 = n23017 & ~n23032 ;
  assign n23034 = ~n23017 & n23031 ;
  assign n23035 = n23033 | n23034 ;
  assign n23036 = n22758 | n22761 ;
  assign n23037 = ( n22758 & n22763 ) | ( n22758 & n23036 ) | ( n22763 & n23036 ) ;
  assign n23038 = n23035 & ~n23037 ;
  assign n23039 = ~n23035 & n23037 ;
  assign n23040 = n23038 | n23039 ;
  assign n23041 = n4471 & ~n17092 ;
  assign n23042 = n4466 & n17111 ;
  assign n23043 = n4468 & n17100 ;
  assign n23044 = n23042 | n23043 ;
  assign n23045 = n23041 | n23044 ;
  assign n23046 = n4475 | n23041 ;
  assign n23047 = n23044 | n23046 ;
  assign n23048 = ( ~n17134 & n23045 ) | ( ~n17134 & n23047 ) | ( n23045 & n23047 ) ;
  assign n23049 = ~x17 & n23047 ;
  assign n23050 = ~x17 & n23045 ;
  assign n23051 = ( ~n17134 & n23049 ) | ( ~n17134 & n23050 ) | ( n23049 & n23050 ) ;
  assign n23052 = x17 | n23050 ;
  assign n23053 = x17 | n23049 ;
  assign n23054 = ( ~n17134 & n23052 ) | ( ~n17134 & n23053 ) | ( n23052 & n23053 ) ;
  assign n23055 = ( ~n23048 & n23051 ) | ( ~n23048 & n23054 ) | ( n23051 & n23054 ) ;
  assign n23056 = n23040 & n23055 ;
  assign n23057 = n23040 | n23055 ;
  assign n23058 = ~n23056 & n23057 ;
  assign n23059 = n22780 & n23058 ;
  assign n23060 = ( n22784 & n23058 ) | ( n22784 & n23059 ) | ( n23058 & n23059 ) ;
  assign n23061 = n22780 | n23058 ;
  assign n23062 = n22784 | n23061 ;
  assign n23063 = ~n23060 & n23062 ;
  assign n23064 = n5234 & n18410 ;
  assign n23065 = n5237 & n18037 ;
  assign n23066 = n5231 & ~n18585 ;
  assign n23067 = n23065 | n23066 ;
  assign n23068 = n23064 | n23067 ;
  assign n23069 = n18586 & ~n23068 ;
  assign n23070 = ( n18609 & ~n23068 ) | ( n18609 & n23069 ) | ( ~n23068 & n23069 ) ;
  assign n23071 = ~n18650 & n23070 ;
  assign n23072 = n5227 | n23064 ;
  assign n23073 = n23067 | n23072 ;
  assign n23074 = ~n23071 & n23073 ;
  assign n23075 = x14 & n23073 ;
  assign n23076 = ~n23071 & n23075 ;
  assign n23077 = x14 & ~n23075 ;
  assign n23078 = ( x14 & n23071 ) | ( x14 & n23077 ) | ( n23071 & n23077 ) ;
  assign n23079 = ( n23074 & ~n23076 ) | ( n23074 & n23078 ) | ( ~n23076 & n23078 ) ;
  assign n23080 = n23063 & n23079 ;
  assign n23081 = n23063 & ~n23080 ;
  assign n23082 = ~n23063 & n23079 ;
  assign n23083 = n23081 | n23082 ;
  assign n23084 = n22803 | n22806 ;
  assign n23085 = ( n22803 & n22808 ) | ( n22803 & n23084 ) | ( n22808 & n23084 ) ;
  assign n23086 = n23083 & ~n23085 ;
  assign n23087 = ~n23083 & n23085 ;
  assign n23088 = n23086 | n23087 ;
  assign n23089 = n6122 & n19494 ;
  assign n23090 = n6125 & n18576 ;
  assign n23091 = n6119 & n19352 ;
  assign n23092 = n23090 | n23091 ;
  assign n23093 = n23089 | n23092 ;
  assign n23094 = n6115 | n23089 ;
  assign n23095 = n23092 | n23094 ;
  assign n23096 = ( n20320 & n23093 ) | ( n20320 & n23095 ) | ( n23093 & n23095 ) ;
  assign n23097 = x11 & n23095 ;
  assign n23098 = x11 & n23093 ;
  assign n23099 = ( n20320 & n23097 ) | ( n20320 & n23098 ) | ( n23097 & n23098 ) ;
  assign n23100 = x11 & ~n23098 ;
  assign n23101 = x11 & ~n23097 ;
  assign n23102 = ( ~n20320 & n23100 ) | ( ~n20320 & n23101 ) | ( n23100 & n23101 ) ;
  assign n23103 = ( n23096 & ~n23099 ) | ( n23096 & n23102 ) | ( ~n23099 & n23102 ) ;
  assign n23104 = n23088 & n23103 ;
  assign n23105 = n23088 | n23103 ;
  assign n23106 = ~n23104 & n23105 ;
  assign n23107 = n22829 & n23106 ;
  assign n23108 = ( n22836 & n23106 ) | ( n22836 & n23107 ) | ( n23106 & n23107 ) ;
  assign n23109 = n22829 | n23106 ;
  assign n23110 = n22836 | n23109 ;
  assign n23111 = ~n23108 & n23110 ;
  assign n23112 = n7079 & ~n20618 ;
  assign n23113 = n7074 & n19631 ;
  assign n23114 = n7068 & ~n20630 ;
  assign n23115 = n23113 | n23114 ;
  assign n23116 = n23112 | n23115 ;
  assign n23117 = n20680 | n23116 ;
  assign n23118 = n7078 | n23112 ;
  assign n23119 = n23115 | n23118 ;
  assign n23120 = n20689 & n23119 ;
  assign n23121 = ( n23117 & n23119 ) | ( n23117 & n23120 ) | ( n23119 & n23120 ) ;
  assign n23122 = ~x8 & n23121 ;
  assign n23123 = x8 | n23121 ;
  assign n23124 = ( ~n23121 & n23122 ) | ( ~n23121 & n23123 ) | ( n23122 & n23123 ) ;
  assign n23125 = n23111 & n23124 ;
  assign n23126 = n23111 & ~n23125 ;
  assign n23127 = ~n23111 & n23124 ;
  assign n23128 = n23126 | n23127 ;
  assign n23129 = ~n22885 & n23128 ;
  assign n23130 = n22885 & ~n23128 ;
  assign n23131 = n23129 | n23130 ;
  assign n23132 = n8122 & ~n21517 ;
  assign n23133 = n8115 & n20609 ;
  assign n23134 = n8118 & ~n21563 ;
  assign n23135 = n23133 | n23134 ;
  assign n23136 = n23132 | n23135 ;
  assign n23137 = n8125 | n23132 ;
  assign n23138 = n23135 | n23137 ;
  assign n23139 = ( ~n22283 & n23136 ) | ( ~n22283 & n23138 ) | ( n23136 & n23138 ) ;
  assign n23140 = n23136 & n23138 ;
  assign n23141 = ( ~n22271 & n23139 ) | ( ~n22271 & n23140 ) | ( n23139 & n23140 ) ;
  assign n23142 = ~x5 & n23141 ;
  assign n23143 = x5 | n23141 ;
  assign n23144 = ( ~n23141 & n23142 ) | ( ~n23141 & n23143 ) | ( n23142 & n23143 ) ;
  assign n23145 = n23131 & n23144 ;
  assign n23146 = n23131 | n23144 ;
  assign n23147 = ~n23145 & n23146 ;
  assign n23148 = n22879 & n23147 ;
  assign n23149 = ( n22884 & n23147 ) | ( n22884 & n23148 ) | ( n23147 & n23148 ) ;
  assign n23150 = n22879 | n23147 ;
  assign n23151 = n22884 | n23150 ;
  assign n23152 = ~n23149 & n23151 ;
  assign n23153 = ~n21537 & n21541 ;
  assign n23154 = ~n21538 & n23153 ;
  assign n23155 = ( n21537 & n21543 ) | ( n21537 & ~n23154 ) | ( n21543 & ~n23154 ) ;
  assign n23156 = ( n21537 & n21545 ) | ( n21537 & ~n23154 ) | ( n21545 & ~n23154 ) ;
  assign n23157 = ( n15882 & n23155 ) | ( n15882 & n23156 ) | ( n23155 & n23156 ) ;
  assign n23158 = n1260 | n2030 ;
  assign n23159 = n1081 | n23158 ;
  assign n23160 = n1156 | n19365 ;
  assign n23161 = n23159 | n23160 ;
  assign n23162 = n15058 | n23161 ;
  assign n23163 = n3292 | n23162 ;
  assign n23164 = n19386 | n23163 ;
  assign n23165 = n384 | n416 ;
  assign n23166 = n208 | n424 ;
  assign n23167 = n23165 | n23166 ;
  assign n23168 = n23164 | n23167 ;
  assign n23169 = n19394 | n19398 ;
  assign n23170 = n236 | n399 ;
  assign n23171 = n703 | n23170 ;
  assign n23172 = n75 | n23171 ;
  assign n23173 = n412 | n451 ;
  assign n23174 = n183 | n23173 ;
  assign n23175 = n79 | n306 ;
  assign n23176 = n277 | n23175 ;
  assign n23177 = n23174 | n23176 ;
  assign n23178 = n2787 | n23177 ;
  assign n23179 = ( ~n19398 & n23172 ) | ( ~n19398 & n23178 ) | ( n23172 & n23178 ) ;
  assign n23180 = n23172 & n23178 ;
  assign n23181 = ( ~n19394 & n23179 ) | ( ~n19394 & n23180 ) | ( n23179 & n23180 ) ;
  assign n23182 = n23169 | n23181 ;
  assign n23183 = n3371 | n3382 ;
  assign n23184 = n204 | n963 ;
  assign n23185 = n1663 | n23184 ;
  assign n23186 = n962 | n23185 ;
  assign n23187 = n364 | n2117 ;
  assign n23188 = n654 | n23187 ;
  assign n23189 = n23186 | n23188 ;
  assign n23190 = n23183 | n23189 ;
  assign n23191 = n23182 | n23190 ;
  assign n23192 = n23168 | n23191 ;
  assign n23193 = n1355 | n5860 ;
  assign n23194 = n2666 | n23193 ;
  assign n23195 = n763 | n821 ;
  assign n23196 = n153 | n23195 ;
  assign n23197 = n23194 | n23196 ;
  assign n23198 = n94 | n431 ;
  assign n23199 = n23197 | n23198 ;
  assign n23200 = n8973 | n8974 ;
  assign n23201 = n311 | n23200 ;
  assign n23202 = n23199 | n23201 ;
  assign n23203 = n434 | n23202 ;
  assign n23204 = n23192 | n23203 ;
  assign n23205 = n21531 & n23204 ;
  assign n23206 = n21531 | n23204 ;
  assign n23207 = ~n23205 & n23206 ;
  assign n23208 = ~n23154 & n23207 ;
  assign n23209 = n21534 & n23206 ;
  assign n23210 = ~n23205 & n23209 ;
  assign n23211 = n21536 & n23206 ;
  assign n23212 = ~n23205 & n23211 ;
  assign n23213 = ( ~n9072 & n23210 ) | ( ~n9072 & n23212 ) | ( n23210 & n23212 ) ;
  assign n23214 = ( n21543 & n23208 ) | ( n21543 & n23213 ) | ( n23208 & n23213 ) ;
  assign n23215 = ( n21545 & n23208 ) | ( n21545 & n23213 ) | ( n23208 & n23213 ) ;
  assign n23216 = ( n15882 & n23214 ) | ( n15882 & n23215 ) | ( n23214 & n23215 ) ;
  assign n23217 = n23157 & ~n23216 ;
  assign n23218 = n23206 & ~n23207 ;
  assign n23219 = ( n23154 & n23206 ) | ( n23154 & n23218 ) | ( n23206 & n23218 ) ;
  assign n23220 = n23206 & ~n23212 ;
  assign n23221 = n23206 & ~n23210 ;
  assign n23222 = ( n9072 & n23220 ) | ( n9072 & n23221 ) | ( n23220 & n23221 ) ;
  assign n23223 = ( ~n21543 & n23219 ) | ( ~n21543 & n23222 ) | ( n23219 & n23222 ) ;
  assign n23224 = ~n23205 & n23223 ;
  assign n23225 = ( ~n21545 & n23219 ) | ( ~n21545 & n23222 ) | ( n23219 & n23222 ) ;
  assign n23226 = ~n23205 & n23225 ;
  assign n23227 = ( ~n15882 & n23224 ) | ( ~n15882 & n23226 ) | ( n23224 & n23226 ) ;
  assign n23228 = n23217 | n23227 ;
  assign n23229 = n23204 & n23207 ;
  assign n23230 = ~n23154 & n23229 ;
  assign n23231 = n23204 & n23212 ;
  assign n23232 = n23204 & n23210 ;
  assign n23233 = ( ~n9072 & n23231 ) | ( ~n9072 & n23232 ) | ( n23231 & n23232 ) ;
  assign n23234 = ( n21543 & n23230 ) | ( n21543 & n23233 ) | ( n23230 & n23233 ) ;
  assign n23235 = ( n21545 & n23230 ) | ( n21545 & n23233 ) | ( n23230 & n23233 ) ;
  assign n23236 = ( n15882 & n23234 ) | ( n15882 & n23235 ) | ( n23234 & n23235 ) ;
  assign n23237 = ~n23204 & n23223 ;
  assign n23238 = ~n23204 & n23225 ;
  assign n23239 = ( ~n15882 & n23237 ) | ( ~n15882 & n23238 ) | ( n23237 & n23238 ) ;
  assign n23240 = n23236 | n23239 ;
  assign n23241 = n23228 & ~n23240 ;
  assign n23242 = ~n23228 & n23240 ;
  assign n23243 = n23241 | n23242 ;
  assign n23244 = ~n21551 & n23228 ;
  assign n23245 = n21551 & ~n23228 ;
  assign n23246 = n23244 | n23245 ;
  assign n23247 = n21552 & ~n23244 ;
  assign n23248 = ( ~n23244 & n23246 ) | ( ~n23244 & n23247 ) | ( n23246 & n23247 ) ;
  assign n23249 = n23243 | n23248 ;
  assign n23250 = ~n23244 & n23246 ;
  assign n23251 = n23243 | n23250 ;
  assign n23252 = ( ~n21554 & n23249 ) | ( ~n21554 & n23251 ) | ( n23249 & n23251 ) ;
  assign n23253 = n23249 | n23251 ;
  assign n23254 = ( n21584 & n23252 ) | ( n21584 & n23253 ) | ( n23252 & n23253 ) ;
  assign n23255 = n23248 | n23250 ;
  assign n23256 = n23243 & n23255 ;
  assign n23257 = ( ~n21554 & n23248 ) | ( ~n21554 & n23250 ) | ( n23248 & n23250 ) ;
  assign n23258 = n23243 & n23257 ;
  assign n23259 = ( n21584 & n23256 ) | ( n21584 & n23258 ) | ( n23256 & n23258 ) ;
  assign n23260 = n23254 & ~n23259 ;
  assign n23262 = n9021 & ~n21551 ;
  assign n23263 = n9024 & n23227 ;
  assign n23264 = ( n9024 & n23217 ) | ( n9024 & n23263 ) | ( n23217 & n23263 ) ;
  assign n23265 = n23262 | n23264 ;
  assign n23261 = n9475 & ~n23240 ;
  assign n23267 = n8970 | n23261 ;
  assign n23268 = n23265 | n23267 ;
  assign n23266 = n23261 | n23265 ;
  assign n23269 = n23266 & n23268 ;
  assign n23270 = ( n23260 & n23268 ) | ( n23260 & n23269 ) | ( n23268 & n23269 ) ;
  assign n23271 = x2 & n23269 ;
  assign n23272 = x2 & n23268 ;
  assign n23273 = ( n23260 & n23271 ) | ( n23260 & n23272 ) | ( n23271 & n23272 ) ;
  assign n23274 = x2 & ~n23271 ;
  assign n23275 = x2 & ~n23272 ;
  assign n23276 = ( ~n23260 & n23274 ) | ( ~n23260 & n23275 ) | ( n23274 & n23275 ) ;
  assign n23277 = ( n23270 & ~n23273 ) | ( n23270 & n23276 ) | ( ~n23273 & n23276 ) ;
  assign n23278 = n23152 & n23277 ;
  assign n23279 = n23152 | n23277 ;
  assign n23280 = ~n23278 & n23279 ;
  assign n23281 = n22882 | n22883 ;
  assign n23282 = ~n22884 & n23281 ;
  assign n23283 = n21552 & ~n21554 ;
  assign n23284 = ( n21552 & n21584 ) | ( n21552 & n23283 ) | ( n21584 & n23283 ) ;
  assign n23285 = n21552 | n23246 ;
  assign n23286 = ( ~n21554 & n23246 ) | ( ~n21554 & n23285 ) | ( n23246 & n23285 ) ;
  assign n23287 = n23246 | n23285 ;
  assign n23288 = ( n21584 & n23286 ) | ( n21584 & n23287 ) | ( n23286 & n23287 ) ;
  assign n23289 = ~n23284 & n23288 ;
  assign n23290 = n9021 & ~n21517 ;
  assign n23291 = n9024 & ~n21551 ;
  assign n23292 = n23290 | n23291 ;
  assign n23293 = n9475 & n23227 ;
  assign n23294 = ( n9475 & n23217 ) | ( n9475 & n23293 ) | ( n23217 & n23293 ) ;
  assign n23295 = n8970 | n23294 ;
  assign n23296 = n23292 | n23295 ;
  assign n23297 = n23292 | n23294 ;
  assign n23298 = ~n23245 & n23248 ;
  assign n23299 = ~n21554 & n23298 ;
  assign n23300 = n23297 | n23299 ;
  assign n23301 = n23297 | n23298 ;
  assign n23302 = ( n21584 & n23300 ) | ( n21584 & n23301 ) | ( n23300 & n23301 ) ;
  assign n23303 = n23296 & n23302 ;
  assign n23304 = ( n23289 & n23296 ) | ( n23289 & n23303 ) | ( n23296 & n23303 ) ;
  assign n23305 = ~x2 & n23304 ;
  assign n23306 = x2 | n23304 ;
  assign n23307 = ( ~n23304 & n23305 ) | ( ~n23304 & n23306 ) | ( n23305 & n23306 ) ;
  assign n23308 = n23282 & n23307 ;
  assign n23309 = n21603 | n22378 ;
  assign n23310 = n23282 | n23307 ;
  assign n23311 = ~n23308 & n23310 ;
  assign n23312 = n23308 | n23311 ;
  assign n23313 = ( n23308 & n23309 ) | ( n23308 & n23312 ) | ( n23309 & n23312 ) ;
  assign n23314 = n23280 & n23313 ;
  assign n23315 = n23280 | n23313 ;
  assign n23316 = ~n23314 & n23315 ;
  assign n23543 = n23125 | n23128 ;
  assign n23544 = ( n22885 & n23125 ) | ( n22885 & n23543 ) | ( n23125 & n23543 ) ;
  assign n23318 = n1826 & ~n12616 ;
  assign n23319 = n1823 & n12936 ;
  assign n23320 = n23318 | n23319 ;
  assign n23317 = n1829 & n13235 ;
  assign n23322 = n1821 | n23317 ;
  assign n23323 = n23320 | n23322 ;
  assign n23321 = n23317 | n23320 ;
  assign n23324 = n23321 & n23323 ;
  assign n23325 = ( n13561 & n23323 ) | ( n13561 & n23324 ) | ( n23323 & n23324 ) ;
  assign n23326 = x29 & n23324 ;
  assign n23327 = x29 & n23323 ;
  assign n23328 = ( n13561 & n23326 ) | ( n13561 & n23327 ) | ( n23326 & n23327 ) ;
  assign n23329 = x29 & ~n23326 ;
  assign n23330 = x29 & ~n23327 ;
  assign n23331 = ( ~n13561 & n23329 ) | ( ~n13561 & n23330 ) | ( n23329 & n23330 ) ;
  assign n23332 = ( n23325 & ~n23328 ) | ( n23325 & n23331 ) | ( ~n23328 & n23331 ) ;
  assign n23333 = n1057 & n12010 ;
  assign n23334 = n1065 & ~n11663 ;
  assign n23335 = n1060 & n11363 ;
  assign n23336 = n23334 | n23335 ;
  assign n23337 = n23333 | n23336 ;
  assign n23338 = n1062 | n23333 ;
  assign n23339 = n23336 | n23338 ;
  assign n23340 = ( ~n12028 & n23337 ) | ( ~n12028 & n23339 ) | ( n23337 & n23339 ) ;
  assign n23341 = n23337 | n23339 ;
  assign n23342 = ( n12017 & n23340 ) | ( n12017 & n23341 ) | ( n23340 & n23341 ) ;
  assign n23343 = n1473 | n18102 ;
  assign n23344 = n836 | n931 ;
  assign n23345 = n23343 | n23344 ;
  assign n23346 = n106 | n23345 ;
  assign n23347 = n11401 | n23346 ;
  assign n23348 = n20429 | n23347 ;
  assign n23349 = n2676 | n23348 ;
  assign n23350 = n5915 | n5941 ;
  assign n23351 = n23349 | n23350 ;
  assign n23352 = n1615 | n3995 ;
  assign n23353 = n364 | n638 ;
  assign n23354 = n297 | n23353 ;
  assign n23355 = n23352 | n23354 ;
  assign n23356 = n263 | n497 ;
  assign n23357 = n354 | n23356 ;
  assign n23358 = n23355 | n23357 ;
  assign n23359 = n23351 | n23358 ;
  assign n23360 = n23339 & n23359 ;
  assign n23361 = n23333 & n23359 ;
  assign n23362 = ( n23336 & n23359 ) | ( n23336 & n23361 ) | ( n23359 & n23361 ) ;
  assign n23363 = ( ~n12028 & n23360 ) | ( ~n12028 & n23362 ) | ( n23360 & n23362 ) ;
  assign n23364 = n23360 | n23362 ;
  assign n23365 = ( n12017 & n23363 ) | ( n12017 & n23364 ) | ( n23363 & n23364 ) ;
  assign n23366 = n23342 & ~n23365 ;
  assign n23367 = ~n23342 & n23359 ;
  assign n23368 = n23366 | n23367 ;
  assign n23369 = n22954 | n22955 ;
  assign n23370 = ( n22954 & n22957 ) | ( n22954 & n23369 ) | ( n22957 & n23369 ) ;
  assign n23371 = ~n23368 & n23370 ;
  assign n23372 = n23332 & n23368 ;
  assign n23373 = ~n23370 & n23372 ;
  assign n23374 = ( n23332 & n23371 ) | ( n23332 & n23373 ) | ( n23371 & n23373 ) ;
  assign n23375 = n23332 | n23368 ;
  assign n23376 = ( n23332 & ~n23370 ) | ( n23332 & n23375 ) | ( ~n23370 & n23375 ) ;
  assign n23377 = n23371 | n23376 ;
  assign n23378 = ~n23374 & n23377 ;
  assign n23379 = n22961 & n23378 ;
  assign n23380 = ( n22967 & n23378 ) | ( n22967 & n23379 ) | ( n23378 & n23379 ) ;
  assign n23381 = n22961 | n23378 ;
  assign n23382 = n22967 | n23381 ;
  assign n23383 = ~n23380 & n23382 ;
  assign n23385 = n2312 & n13522 ;
  assign n23386 = n2308 & n14607 ;
  assign n23387 = n23385 | n23386 ;
  assign n23384 = n2315 & n14329 ;
  assign n23389 = n2306 | n23384 ;
  assign n23390 = n23387 | n23389 ;
  assign n23388 = n23384 | n23387 ;
  assign n23391 = n23388 & n23390 ;
  assign n23392 = ( n14656 & n23390 ) | ( n14656 & n23391 ) | ( n23390 & n23391 ) ;
  assign n23393 = x26 & n23391 ;
  assign n23394 = x26 & n23390 ;
  assign n23395 = ( n14656 & n23393 ) | ( n14656 & n23394 ) | ( n23393 & n23394 ) ;
  assign n23396 = x26 & ~n23393 ;
  assign n23397 = x26 & ~n23394 ;
  assign n23398 = ( ~n14656 & n23396 ) | ( ~n14656 & n23397 ) | ( n23396 & n23397 ) ;
  assign n23399 = ( n23392 & ~n23395 ) | ( n23392 & n23398 ) | ( ~n23395 & n23398 ) ;
  assign n23400 = n23383 & n23399 ;
  assign n23401 = n23383 & ~n23400 ;
  assign n23402 = ~n23383 & n23399 ;
  assign n23403 = n23401 | n23402 ;
  assign n23404 = n22986 | n22989 ;
  assign n23405 = ( n22986 & n22991 ) | ( n22986 & n23404 ) | ( n22991 & n23404 ) ;
  assign n23406 = n23403 & ~n23405 ;
  assign n23407 = ~n23403 & n23405 ;
  assign n23408 = n23406 | n23407 ;
  assign n23409 = n2932 & ~n16085 ;
  assign n23410 = n2925 & n14591 ;
  assign n23411 = n2928 & n15434 ;
  assign n23412 = n23410 | n23411 ;
  assign n23413 = n23409 | n23412 ;
  assign n23414 = n2936 | n23409 ;
  assign n23415 = n23412 | n23414 ;
  assign n23416 = ( ~n16167 & n23413 ) | ( ~n16167 & n23415 ) | ( n23413 & n23415 ) ;
  assign n23417 = ~x23 & n23415 ;
  assign n23418 = ~x23 & n23413 ;
  assign n23419 = ( ~n16167 & n23417 ) | ( ~n16167 & n23418 ) | ( n23417 & n23418 ) ;
  assign n23420 = x23 | n23418 ;
  assign n23421 = x23 | n23417 ;
  assign n23422 = ( ~n16167 & n23420 ) | ( ~n16167 & n23421 ) | ( n23420 & n23421 ) ;
  assign n23423 = ( ~n23416 & n23419 ) | ( ~n23416 & n23422 ) | ( n23419 & n23422 ) ;
  assign n23424 = n23408 & n23423 ;
  assign n23425 = n23408 | n23423 ;
  assign n23426 = ~n23424 & n23425 ;
  assign n23427 = n23010 | n23012 ;
  assign n23428 = ( n23010 & n23014 ) | ( n23010 & n23427 ) | ( n23014 & n23427 ) ;
  assign n23429 = n23426 & n23428 ;
  assign n23430 = n23426 | n23428 ;
  assign n23431 = ~n23429 & n23430 ;
  assign n23432 = n3544 & n15886 ;
  assign n23433 = n3541 & ~n16069 ;
  assign n23434 = n23432 | n23433 ;
  assign n23435 = n3547 & n17111 ;
  assign n23436 = n3537 | n23435 ;
  assign n23437 = n23434 | n23436 ;
  assign n23438 = n23434 | n23435 ;
  assign n23439 = n17194 & ~n23438 ;
  assign n23440 = ( n17129 & ~n23438 ) | ( n17129 & n23439 ) | ( ~n23438 & n23439 ) ;
  assign n23441 = n23437 & ~n23440 ;
  assign n23442 = ( n17186 & n23437 ) | ( n17186 & n23441 ) | ( n23437 & n23441 ) ;
  assign n23443 = x20 & n23442 ;
  assign n23444 = x20 & ~n23442 ;
  assign n23445 = ( n23442 & ~n23443 ) | ( n23442 & n23444 ) | ( ~n23443 & n23444 ) ;
  assign n23446 = n23431 & n23445 ;
  assign n23447 = n23431 & ~n23446 ;
  assign n23448 = ~n23431 & n23445 ;
  assign n23449 = n23447 | n23448 ;
  assign n23450 = n23032 | n23035 ;
  assign n23451 = ( n23032 & n23037 ) | ( n23032 & n23450 ) | ( n23037 & n23450 ) ;
  assign n23452 = n23449 & ~n23451 ;
  assign n23453 = ~n23449 & n23451 ;
  assign n23454 = n23452 | n23453 ;
  assign n23455 = n4471 & n18037 ;
  assign n23456 = n4466 & n17100 ;
  assign n23457 = n4468 & ~n17092 ;
  assign n23458 = n23456 | n23457 ;
  assign n23459 = n23455 | n23458 ;
  assign n23460 = n4475 | n23455 ;
  assign n23461 = n23458 | n23460 ;
  assign n23462 = ( ~n18050 & n23459 ) | ( ~n18050 & n23461 ) | ( n23459 & n23461 ) ;
  assign n23463 = ~x17 & n23461 ;
  assign n23464 = ~x17 & n23459 ;
  assign n23465 = ( ~n18050 & n23463 ) | ( ~n18050 & n23464 ) | ( n23463 & n23464 ) ;
  assign n23466 = x17 | n23464 ;
  assign n23467 = x17 | n23463 ;
  assign n23468 = ( ~n18050 & n23466 ) | ( ~n18050 & n23467 ) | ( n23466 & n23467 ) ;
  assign n23469 = ( ~n23462 & n23465 ) | ( ~n23462 & n23468 ) | ( n23465 & n23468 ) ;
  assign n23470 = n23454 & n23469 ;
  assign n23471 = n23454 | n23469 ;
  assign n23472 = ~n23470 & n23471 ;
  assign n23473 = n23056 & n23472 ;
  assign n23474 = ( n23060 & n23472 ) | ( n23060 & n23473 ) | ( n23472 & n23473 ) ;
  assign n23475 = n23056 | n23472 ;
  assign n23476 = n23060 | n23475 ;
  assign n23477 = ~n23474 & n23476 ;
  assign n23479 = n5237 & ~n18585 ;
  assign n23480 = n5231 & n18410 ;
  assign n23481 = n23479 | n23480 ;
  assign n23478 = n5234 & n18576 ;
  assign n23483 = n5227 | n23478 ;
  assign n23484 = n23481 | n23483 ;
  assign n23482 = n23478 | n23481 ;
  assign n23485 = n23482 & n23484 ;
  assign n23486 = ( n18612 & n23484 ) | ( n18612 & n23485 ) | ( n23484 & n23485 ) ;
  assign n23487 = x14 & n23485 ;
  assign n23488 = x14 & n23484 ;
  assign n23489 = ( n18612 & n23487 ) | ( n18612 & n23488 ) | ( n23487 & n23488 ) ;
  assign n23490 = x14 & ~n23487 ;
  assign n23491 = x14 & ~n23488 ;
  assign n23492 = ( ~n18612 & n23490 ) | ( ~n18612 & n23491 ) | ( n23490 & n23491 ) ;
  assign n23493 = ( n23486 & ~n23489 ) | ( n23486 & n23492 ) | ( ~n23489 & n23492 ) ;
  assign n23494 = n23477 & n23493 ;
  assign n23495 = n23477 & ~n23494 ;
  assign n23496 = ~n23477 & n23493 ;
  assign n23497 = n23495 | n23496 ;
  assign n23498 = n23080 | n23083 ;
  assign n23499 = ( n23080 & n23085 ) | ( n23080 & n23498 ) | ( n23085 & n23498 ) ;
  assign n23500 = n23497 & ~n23499 ;
  assign n23501 = ~n23497 & n23499 ;
  assign n23502 = n23500 | n23501 ;
  assign n23503 = n6122 & n19631 ;
  assign n23504 = n6125 & n19352 ;
  assign n23505 = n6119 & n19494 ;
  assign n23506 = n23504 | n23505 ;
  assign n23507 = n23503 | n23506 ;
  assign n23508 = n6115 & n19652 ;
  assign n23509 = n6115 & n19655 ;
  assign n23510 = ( ~n18604 & n23508 ) | ( ~n18604 & n23509 ) | ( n23508 & n23509 ) ;
  assign n23511 = n23507 | n23510 ;
  assign n23512 = n6115 | n23507 ;
  assign n23513 = ( n19640 & n23511 ) | ( n19640 & n23512 ) | ( n23511 & n23512 ) ;
  assign n23514 = x11 | n23513 ;
  assign n23515 = ~x11 & n23513 ;
  assign n23516 = ( ~n23513 & n23514 ) | ( ~n23513 & n23515 ) | ( n23514 & n23515 ) ;
  assign n23517 = n23502 & n23516 ;
  assign n23518 = n23502 | n23516 ;
  assign n23519 = ~n23517 & n23518 ;
  assign n23520 = n23104 & n23519 ;
  assign n23521 = ( n23108 & n23519 ) | ( n23108 & n23520 ) | ( n23519 & n23520 ) ;
  assign n23522 = n23104 | n23519 ;
  assign n23523 = n23108 | n23522 ;
  assign n23524 = ~n23521 & n23523 ;
  assign n23526 = n7074 & ~n20630 ;
  assign n23527 = n7068 & ~n20618 ;
  assign n23528 = n23526 | n23527 ;
  assign n23525 = n7079 & n20609 ;
  assign n23530 = n7078 | n23525 ;
  assign n23531 = n23528 | n23530 ;
  assign n23529 = n23525 | n23528 ;
  assign n23532 = n23529 & n23531 ;
  assign n23533 = ( n20659 & n23531 ) | ( n20659 & n23532 ) | ( n23531 & n23532 ) ;
  assign n23534 = n23531 & n23532 ;
  assign n23535 = ( ~n20649 & n23533 ) | ( ~n20649 & n23534 ) | ( n23533 & n23534 ) ;
  assign n23536 = x8 & n23535 ;
  assign n23537 = x8 & ~n23535 ;
  assign n23538 = ( n23535 & ~n23536 ) | ( n23535 & n23537 ) | ( ~n23536 & n23537 ) ;
  assign n23539 = n23524 & n23538 ;
  assign n23540 = n23524 & ~n23539 ;
  assign n23541 = ~n23524 & n23538 ;
  assign n23542 = n23540 | n23541 ;
  assign n23545 = n23542 & n23544 ;
  assign n23546 = n23544 & ~n23545 ;
  assign n23547 = n23542 & ~n23544 ;
  assign n23548 = n23546 | n23547 ;
  assign n23549 = n8122 & ~n21551 ;
  assign n23550 = n8115 & ~n21563 ;
  assign n23551 = n8118 & ~n21517 ;
  assign n23552 = n23550 | n23551 ;
  assign n23553 = n23549 | n23552 ;
  assign n23554 = n8125 | n23549 ;
  assign n23555 = n23552 | n23554 ;
  assign n23556 = ( ~n21587 & n23553 ) | ( ~n21587 & n23555 ) | ( n23553 & n23555 ) ;
  assign n23557 = ~x5 & n23555 ;
  assign n23558 = ~x5 & n23553 ;
  assign n23559 = ( ~n21587 & n23557 ) | ( ~n21587 & n23558 ) | ( n23557 & n23558 ) ;
  assign n23560 = x5 | n23558 ;
  assign n23561 = x5 | n23557 ;
  assign n23562 = ( ~n21587 & n23560 ) | ( ~n21587 & n23561 ) | ( n23560 & n23561 ) ;
  assign n23563 = ( ~n23556 & n23559 ) | ( ~n23556 & n23562 ) | ( n23559 & n23562 ) ;
  assign n23564 = n23547 & n23563 ;
  assign n23565 = ( n23546 & n23563 ) | ( n23546 & n23564 ) | ( n23563 & n23564 ) ;
  assign n23566 = n23548 & ~n23565 ;
  assign n23567 = ~n23547 & n23563 ;
  assign n23568 = ~n23546 & n23567 ;
  assign n23569 = n23566 | n23568 ;
  assign n23570 = n23145 | n23149 ;
  assign n23571 = n23569 & n23570 ;
  assign n23572 = n23569 | n23570 ;
  assign n23573 = ~n23571 & n23572 ;
  assign n23574 = ~n23241 & n23243 ;
  assign n23575 = ( ~n23241 & n23248 ) | ( ~n23241 & n23574 ) | ( n23248 & n23574 ) ;
  assign n23576 = n23239 & ~n23575 ;
  assign n23577 = ( ~n23241 & n23250 ) | ( ~n23241 & n23574 ) | ( n23250 & n23574 ) ;
  assign n23578 = n23239 & ~n23577 ;
  assign n23579 = ( n21554 & n23576 ) | ( n21554 & n23578 ) | ( n23576 & n23578 ) ;
  assign n23580 = n23576 & n23578 ;
  assign n23581 = ( ~n21584 & n23579 ) | ( ~n21584 & n23580 ) | ( n23579 & n23580 ) ;
  assign n23582 = n23575 | n23577 ;
  assign n23583 = ~n23239 & n23582 ;
  assign n23584 = ( ~n21554 & n23575 ) | ( ~n21554 & n23577 ) | ( n23575 & n23577 ) ;
  assign n23585 = ~n23239 & n23584 ;
  assign n23586 = ( n21584 & n23583 ) | ( n21584 & n23585 ) | ( n23583 & n23585 ) ;
  assign n23587 = n23581 | n23586 ;
  assign n23588 = n9024 & ~n23240 ;
  assign n23589 = n9021 & n23227 ;
  assign n23590 = ( n9021 & n23217 ) | ( n9021 & n23589 ) | ( n23217 & n23589 ) ;
  assign n23591 = n23588 | n23590 ;
  assign n23592 = n9475 & ~n23234 ;
  assign n23593 = n9475 & ~n23235 ;
  assign n23594 = ( ~n15882 & n23592 ) | ( ~n15882 & n23593 ) | ( n23592 & n23593 ) ;
  assign n23596 = n8970 | n23594 ;
  assign n23597 = n23591 | n23596 ;
  assign n23595 = n23591 | n23594 ;
  assign n23598 = n23595 & n23597 ;
  assign n23599 = ( ~n23587 & n23597 ) | ( ~n23587 & n23598 ) | ( n23597 & n23598 ) ;
  assign n23600 = ~x2 & n23598 ;
  assign n23601 = ~x2 & n23597 ;
  assign n23602 = ( ~n23587 & n23600 ) | ( ~n23587 & n23601 ) | ( n23600 & n23601 ) ;
  assign n23603 = x2 | n23600 ;
  assign n23604 = x2 | n23601 ;
  assign n23605 = ( ~n23587 & n23603 ) | ( ~n23587 & n23604 ) | ( n23603 & n23604 ) ;
  assign n23606 = ( ~n23599 & n23602 ) | ( ~n23599 & n23605 ) | ( n23602 & n23605 ) ;
  assign n23607 = n23573 & n23606 ;
  assign n23608 = n23573 | n23606 ;
  assign n23609 = ~n23607 & n23608 ;
  assign n23610 = n23278 | n23280 ;
  assign n23611 = ( n23278 & n23313 ) | ( n23278 & n23610 ) | ( n23313 & n23610 ) ;
  assign n23612 = n23609 & n23611 ;
  assign n23613 = n23609 | n23611 ;
  assign n23614 = ~n23612 & n23613 ;
  assign n23615 = n23316 & n23614 ;
  assign n23616 = n23316 | n23614 ;
  assign n23617 = ~n23615 & n23616 ;
  assign n23618 = n23309 & n23311 ;
  assign n23619 = n23309 | n23311 ;
  assign n23620 = ~n23618 & n23619 ;
  assign n23621 = n23316 & n23620 ;
  assign n23622 = n22381 & n23620 ;
  assign n23623 = ~n22386 & n22419 ;
  assign n23624 = n22381 | n23620 ;
  assign n23625 = ~n23622 & n23624 ;
  assign n23626 = n23622 | n23625 ;
  assign n23627 = ( n23622 & ~n23623 ) | ( n23622 & n23626 ) | ( ~n23623 & n23626 ) ;
  assign n23628 = n23316 | n23620 ;
  assign n23629 = ~n23621 & n23628 ;
  assign n23630 = n23621 | n23629 ;
  assign n23631 = ( n23621 & n23627 ) | ( n23621 & n23630 ) | ( n23627 & n23630 ) ;
  assign n23632 = n23617 & n23631 ;
  assign n23633 = n23617 | n23631 ;
  assign n23634 = ~n23632 & n23633 ;
  assign n23635 = n2315 & n23614 ;
  assign n23636 = n2312 & n23620 ;
  assign n23637 = ( n2308 & n13089 ) | ( n2308 & n23620 ) | ( n13089 & n23620 ) ;
  assign n23638 = ( n23316 & n23636 ) | ( n23316 & n23637 ) | ( n23636 & n23637 ) ;
  assign n23640 = n2306 | n23638 ;
  assign n23641 = n23635 | n23640 ;
  assign n23639 = n23635 | n23638 ;
  assign n23642 = n23639 & n23641 ;
  assign n23643 = ( n23634 & n23641 ) | ( n23634 & n23642 ) | ( n23641 & n23642 ) ;
  assign n23644 = x26 & n23642 ;
  assign n23645 = x26 & n23641 ;
  assign n23646 = ( n23634 & n23644 ) | ( n23634 & n23645 ) | ( n23644 & n23645 ) ;
  assign n23647 = x26 & ~n23644 ;
  assign n23648 = x26 & ~n23645 ;
  assign n23649 = ( ~n23634 & n23647 ) | ( ~n23634 & n23648 ) | ( n23647 & n23648 ) ;
  assign n23650 = ( n23643 & ~n23646 ) | ( n23643 & n23649 ) | ( ~n23646 & n23649 ) ;
  assign n23651 = ~n22630 & n23650 ;
  assign n23652 = n22630 | n23651 ;
  assign n23653 = n22630 & n23650 ;
  assign n23654 = n23652 & ~n23653 ;
  assign n23655 = n22572 | n22626 ;
  assign n23659 = n23627 & n23629 ;
  assign n23660 = n23627 | n23629 ;
  assign n23661 = ~n23659 & n23660 ;
  assign n23662 = n2312 & n22381 ;
  assign n23663 = ( n2308 & n13089 ) | ( n2308 & n22381 ) | ( n13089 & n22381 ) ;
  assign n23664 = ( n23620 & n23662 ) | ( n23620 & n23663 ) | ( n23662 & n23663 ) ;
  assign n23665 = n2315 | n23663 ;
  assign n23666 = n2315 | n23662 ;
  assign n23667 = ( n23620 & n23665 ) | ( n23620 & n23666 ) | ( n23665 & n23666 ) ;
  assign n23668 = ( n23316 & n23664 ) | ( n23316 & n23667 ) | ( n23664 & n23667 ) ;
  assign n23669 = n2306 | n23668 ;
  assign n23670 = ( n23661 & n23668 ) | ( n23661 & n23669 ) | ( n23668 & n23669 ) ;
  assign n23671 = x26 & n23669 ;
  assign n23672 = x26 & n23668 ;
  assign n23673 = ( n23661 & n23671 ) | ( n23661 & n23672 ) | ( n23671 & n23672 ) ;
  assign n23674 = x26 & ~n23671 ;
  assign n23675 = x26 & ~n23672 ;
  assign n23676 = ( ~n23661 & n23674 ) | ( ~n23661 & n23675 ) | ( n23674 & n23675 ) ;
  assign n23677 = ( n23670 & ~n23673 ) | ( n23670 & n23676 ) | ( ~n23673 & n23676 ) ;
  assign n23656 = n22572 & n22624 ;
  assign n23657 = ( n22572 & n22620 ) | ( n22572 & n23656 ) | ( n22620 & n23656 ) ;
  assign n23678 = n23657 & n23677 ;
  assign n23679 = ( ~n23655 & n23677 ) | ( ~n23655 & n23678 ) | ( n23677 & n23678 ) ;
  assign n23658 = n23655 & ~n23657 ;
  assign n23680 = n23658 | n23679 ;
  assign n23681 = ~n23657 & n23677 ;
  assign n23682 = n23655 & n23681 ;
  assign n23683 = n23680 & ~n23682 ;
  assign n23684 = ~n23623 & n23625 ;
  assign n23685 = n23623 & ~n23625 ;
  assign n23686 = n23684 | n23685 ;
  assign n23687 = n2312 & ~n22385 ;
  assign n23688 = ( n2308 & n13089 ) | ( n2308 & ~n22385 ) | ( n13089 & ~n22385 ) ;
  assign n23689 = ( n22381 & n23687 ) | ( n22381 & n23688 ) | ( n23687 & n23688 ) ;
  assign n23690 = n2315 | n23689 ;
  assign n23691 = ( n23620 & n23689 ) | ( n23620 & n23690 ) | ( n23689 & n23690 ) ;
  assign n23692 = n2306 | n23691 ;
  assign n23693 = ~x26 & n23692 ;
  assign n23694 = ~x26 & n23691 ;
  assign n23695 = ( ~n23686 & n23693 ) | ( ~n23686 & n23694 ) | ( n23693 & n23694 ) ;
  assign n23696 = ( x26 & n12090 ) | ( x26 & n23691 ) | ( n12090 & n23691 ) ;
  assign n23697 = x26 & ~n23696 ;
  assign n23698 = x26 & n23691 ;
  assign n23699 = x26 & ~n23698 ;
  assign n23700 = ( n23686 & n23697 ) | ( n23686 & n23699 ) | ( n23697 & n23699 ) ;
  assign n23701 = n23695 | n23700 ;
  assign n23702 = n22600 | n22616 ;
  assign n23703 = ~n22616 & n22618 ;
  assign n23704 = ( n22601 & n23702 ) | ( n22601 & ~n23703 ) | ( n23702 & ~n23703 ) ;
  assign n23705 = ~n22620 & n23704 ;
  assign n23706 = n23701 & n23705 ;
  assign n23707 = n23701 | n23705 ;
  assign n23708 = ~n23706 & n23707 ;
  assign n23709 = n22586 | n22598 ;
  assign n23710 = ~n22618 & n23709 ;
  assign n23711 = n2315 & n22381 ;
  assign n23712 = n2312 & ~n22398 ;
  assign n23713 = n2308 & ~n22385 ;
  assign n23714 = n23712 | n23713 ;
  assign n23715 = n23711 | n23714 ;
  assign n23716 = n2306 | n23715 ;
  assign n23717 = x26 & n23716 ;
  assign n23718 = x26 & n23715 ;
  assign n23719 = ( n22422 & n23717 ) | ( n22422 & n23718 ) | ( n23717 & n23718 ) ;
  assign n23720 = x26 | n23716 ;
  assign n23721 = x26 | n23715 ;
  assign n23722 = ( n22422 & n23720 ) | ( n22422 & n23721 ) | ( n23720 & n23721 ) ;
  assign n23723 = ~n23719 & n23722 ;
  assign n23724 = n23710 & n23723 ;
  assign n23725 = ~n23710 & n23723 ;
  assign n23726 = ( n23710 & ~n23724 ) | ( n23710 & n23725 ) | ( ~n23724 & n23725 ) ;
  assign n23727 = n22592 | n22594 ;
  assign n23728 = ~n22594 & n22596 ;
  assign n23729 = ( n22593 & n23727 ) | ( n22593 & ~n23728 ) | ( n23727 & ~n23728 ) ;
  assign n23730 = ~n22598 & n23729 ;
  assign n23731 = n2315 & ~n22385 ;
  assign n23732 = n2312 & n22393 ;
  assign n23733 = n2308 & ~n22398 ;
  assign n23734 = n23732 | n23733 ;
  assign n23735 = n23731 | n23734 ;
  assign n23736 = n2306 | n23731 ;
  assign n23737 = n23734 | n23736 ;
  assign n23738 = ( ~n22545 & n23735 ) | ( ~n22545 & n23737 ) | ( n23735 & n23737 ) ;
  assign n23739 = ~x26 & n23737 ;
  assign n23740 = ~x26 & n23735 ;
  assign n23741 = ( ~n22545 & n23739 ) | ( ~n22545 & n23740 ) | ( n23739 & n23740 ) ;
  assign n23742 = x26 | n23740 ;
  assign n23743 = x26 | n23739 ;
  assign n23744 = ( ~n22545 & n23742 ) | ( ~n22545 & n23743 ) | ( n23742 & n23743 ) ;
  assign n23745 = ( ~n23738 & n23741 ) | ( ~n23738 & n23744 ) | ( n23741 & n23744 ) ;
  assign n23746 = n23730 & n23745 ;
  assign n23747 = n2306 & n22474 ;
  assign n23748 = n2308 & ~n22409 ;
  assign n23749 = n2315 & ~n22406 ;
  assign n23750 = n23748 | n23749 ;
  assign n23751 = x26 | n23750 ;
  assign n23752 = n23747 | n23751 ;
  assign n23753 = ~x26 & n23752 ;
  assign n23754 = ( x26 & n12161 ) | ( x26 & n22409 ) | ( n12161 & n22409 ) ;
  assign n23755 = n23752 & n23754 ;
  assign n23756 = n23747 | n23750 ;
  assign n23757 = n23754 & ~n23756 ;
  assign n23758 = ( n23753 & n23755 ) | ( n23753 & n23757 ) | ( n23755 & n23757 ) ;
  assign n23759 = n2315 & n22393 ;
  assign n23760 = n2312 & ~n22409 ;
  assign n23761 = n2308 & ~n22406 ;
  assign n23762 = n23760 | n23761 ;
  assign n23763 = n23759 | n23762 ;
  assign n23764 = n22439 | n23763 ;
  assign n23765 = n2306 | n23759 ;
  assign n23766 = n23762 | n23765 ;
  assign n23767 = ~x26 & n23766 ;
  assign n23768 = n23764 & n23767 ;
  assign n23769 = x26 | n23768 ;
  assign n23770 = n1820 & ~n22409 ;
  assign n23771 = n23768 & n23770 ;
  assign n23772 = n23764 & n23766 ;
  assign n23773 = n23770 & ~n23772 ;
  assign n23774 = ( n23769 & n23771 ) | ( n23769 & n23773 ) | ( n23771 & n23773 ) ;
  assign n23775 = n23758 & n23774 ;
  assign n23776 = ( n23768 & n23769 ) | ( n23768 & ~n23772 ) | ( n23769 & ~n23772 ) ;
  assign n23777 = n23758 | n23770 ;
  assign n23778 = ( n23770 & n23776 ) | ( n23770 & n23777 ) | ( n23776 & n23777 ) ;
  assign n23779 = ~n23775 & n23778 ;
  assign n23780 = n2312 & ~n22406 ;
  assign n23781 = n2308 & n22393 ;
  assign n23782 = n23780 | n23781 ;
  assign n23783 = n2315 & ~n22398 ;
  assign n23784 = n2306 | n23783 ;
  assign n23785 = n23782 | n23784 ;
  assign n23786 = x26 & n23785 ;
  assign n23787 = n23782 | n23783 ;
  assign n23788 = x26 & n23787 ;
  assign n23789 = ( n22608 & n23786 ) | ( n22608 & n23788 ) | ( n23786 & n23788 ) ;
  assign n23790 = x26 | n23785 ;
  assign n23791 = x26 | n23787 ;
  assign n23792 = ( n22608 & n23790 ) | ( n22608 & n23791 ) | ( n23790 & n23791 ) ;
  assign n23793 = ~n23789 & n23792 ;
  assign n23794 = n23775 | n23793 ;
  assign n23795 = ( n23775 & n23779 ) | ( n23775 & n23794 ) | ( n23779 & n23794 ) ;
  assign n23796 = n23730 | n23745 ;
  assign n23797 = ~n23746 & n23796 ;
  assign n23798 = n23746 | n23797 ;
  assign n23799 = ( n23746 & n23795 ) | ( n23746 & n23798 ) | ( n23795 & n23798 ) ;
  assign n23800 = n23726 & n23799 ;
  assign n23801 = n23724 | n23800 ;
  assign n23802 = n23708 & n23801 ;
  assign n23803 = n23706 | n23802 ;
  assign n23804 = ~n23683 & n23803 ;
  assign n23805 = n23679 | n23804 ;
  assign n23806 = ~n23654 & n23805 ;
  assign n23807 = n23651 | n23806 ;
  assign n23808 = n1826 & ~n22385 ;
  assign n23809 = ( n1823 & n13998 ) | ( n1823 & ~n22385 ) | ( n13998 & ~n22385 ) ;
  assign n23810 = ( n22381 & n23808 ) | ( n22381 & n23809 ) | ( n23808 & n23809 ) ;
  assign n23811 = n1829 | n23810 ;
  assign n23812 = ( n23620 & n23810 ) | ( n23620 & n23811 ) | ( n23810 & n23811 ) ;
  assign n23813 = n1821 | n23812 ;
  assign n23814 = ~x29 & n23813 ;
  assign n23815 = ~x29 & n23812 ;
  assign n23816 = ( ~n23686 & n23814 ) | ( ~n23686 & n23815 ) | ( n23814 & n23815 ) ;
  assign n23817 = ( x29 & n10963 ) | ( x29 & n23812 ) | ( n10963 & n23812 ) ;
  assign n23818 = x29 & ~n23817 ;
  assign n23819 = x29 & n23812 ;
  assign n23820 = x29 & ~n23819 ;
  assign n23821 = ( n23686 & n23818 ) | ( n23686 & n23820 ) | ( n23818 & n23820 ) ;
  assign n23822 = n23816 | n23821 ;
  assign n23823 = n22532 | n22535 ;
  assign n23824 = n12976 | n12977 ;
  assign n23825 = n5178 | n23824 ;
  assign n23826 = n236 | n461 ;
  assign n23827 = n1251 | n23826 ;
  assign n23828 = n2123 | n13310 ;
  assign n23829 = n2122 | n23828 ;
  assign n23830 = n23827 | n23829 ;
  assign n23831 = n110 | n13288 ;
  assign n23832 = n3461 | n23831 ;
  assign n23833 = n12997 | n23832 ;
  assign n23834 = n23830 | n23833 ;
  assign n23835 = n2115 | n23834 ;
  assign n23836 = n1723 | n5860 ;
  assign n23837 = n1301 | n5946 ;
  assign n23838 = n23836 | n23837 ;
  assign n23839 = n456 | n987 ;
  assign n23840 = n666 | n23839 ;
  assign n23841 = n23838 | n23840 ;
  assign n23842 = n349 | n566 ;
  assign n23843 = n23841 | n23842 ;
  assign n23844 = n23835 | n23843 ;
  assign n23845 = n23825 | n23844 ;
  assign n23846 = n1065 & n22393 ;
  assign n23847 = n1060 & ~n22406 ;
  assign n23848 = n23846 | n23847 ;
  assign n23849 = n1057 & ~n22398 ;
  assign n23850 = n1062 | n23849 ;
  assign n23851 = n23848 | n23850 ;
  assign n23852 = n23845 & n23851 ;
  assign n23853 = n23848 | n23849 ;
  assign n23854 = n23845 & n23853 ;
  assign n23855 = ( n22608 & n23852 ) | ( n22608 & n23854 ) | ( n23852 & n23854 ) ;
  assign n23856 = n23845 | n23851 ;
  assign n23857 = n23845 | n23853 ;
  assign n23858 = ( n22608 & n23856 ) | ( n22608 & n23857 ) | ( n23856 & n23857 ) ;
  assign n23859 = ~n23855 & n23858 ;
  assign n23860 = n23823 | n23859 ;
  assign n23861 = n23823 & ~n23859 ;
  assign n23862 = ( ~n23823 & n23860 ) | ( ~n23823 & n23861 ) | ( n23860 & n23861 ) ;
  assign n23863 = n23822 & n23862 ;
  assign n23864 = n23822 | n23862 ;
  assign n23865 = ~n23863 & n23864 ;
  assign n23866 = ~n22539 & n22542 ;
  assign n23867 = ( n22539 & n22627 ) | ( n22539 & ~n23866 ) | ( n22627 & ~n23866 ) ;
  assign n23868 = n23865 | n23867 ;
  assign n23869 = n23865 & n23867 ;
  assign n23870 = n23868 & ~n23869 ;
  assign n23871 = n1057 & ~n12616 ;
  assign n23872 = n1065 & n12010 ;
  assign n23873 = n1060 & ~n11663 ;
  assign n23874 = n23872 | n23873 ;
  assign n23875 = n23871 | n23874 ;
  assign n23876 = n1062 | n23871 ;
  assign n23877 = n23874 | n23876 ;
  assign n23878 = ( ~n12626 & n23875 ) | ( ~n12626 & n23877 ) | ( n23875 & n23877 ) ;
  assign n23879 = n269 | n497 ;
  assign n23880 = n623 | n23879 ;
  assign n23881 = n64 | n654 ;
  assign n23882 = n13826 | n23881 ;
  assign n23883 = n272 | n369 ;
  assign n23884 = n305 | n23883 ;
  assign n23885 = n23882 | n23884 ;
  assign n23886 = n5062 | n5066 ;
  assign n23887 = n954 | n17916 ;
  assign n23888 = n930 | n23887 ;
  assign n23889 = n1447 | n1667 ;
  assign n23890 = n23888 | n23889 ;
  assign n23891 = n5075 | n23890 ;
  assign n23892 = n23886 | n23891 ;
  assign n23893 = n23885 | n23892 ;
  assign n23894 = n283 | n1172 ;
  assign n23895 = n19366 | n23894 ;
  assign n23896 = n402 | n447 ;
  assign n23897 = n801 | n23896 ;
  assign n23898 = n23895 | n23897 ;
  assign n23899 = n357 | n758 ;
  assign n23900 = n442 | n23899 ;
  assign n23901 = n23898 | n23900 ;
  assign n23902 = n388 | n1251 ;
  assign n23903 = n321 | n23902 ;
  assign n23904 = n23901 | n23903 ;
  assign n23905 = n15215 | n23904 ;
  assign n23906 = n23893 | n23905 ;
  assign n23907 = n23880 | n23906 ;
  assign n23908 = n23877 & n23907 ;
  assign n23909 = n23871 & n23907 ;
  assign n23910 = ( n23874 & n23907 ) | ( n23874 & n23909 ) | ( n23907 & n23909 ) ;
  assign n23911 = ( ~n12626 & n23908 ) | ( ~n12626 & n23910 ) | ( n23908 & n23910 ) ;
  assign n23912 = n23878 & ~n23911 ;
  assign n23913 = ~n23877 & n23907 ;
  assign n23914 = ~n23875 & n23907 ;
  assign n23915 = ( n12626 & n23913 ) | ( n12626 & n23914 ) | ( n23913 & n23914 ) ;
  assign n23916 = n23912 | n23915 ;
  assign n23917 = n23365 | n23368 ;
  assign n23918 = n23916 & n23917 ;
  assign n23919 = n23365 & n23916 ;
  assign n23920 = ( n23370 & n23918 ) | ( n23370 & n23919 ) | ( n23918 & n23919 ) ;
  assign n23921 = n23916 | n23917 ;
  assign n23922 = n23365 | n23916 ;
  assign n23923 = ( n23370 & n23921 ) | ( n23370 & n23922 ) | ( n23921 & n23922 ) ;
  assign n23924 = ~n23920 & n23923 ;
  assign n23925 = n1826 & n12936 ;
  assign n23926 = n1823 & n13235 ;
  assign n23927 = n23925 | n23926 ;
  assign n23928 = n1829 & n13522 ;
  assign n23929 = n1821 | n23928 ;
  assign n23930 = n23927 | n23929 ;
  assign n23931 = n23927 | n23928 ;
  assign n23932 = n13537 | n23931 ;
  assign n23933 = n13539 | n23931 ;
  assign n23934 = ( ~n13248 & n23932 ) | ( ~n13248 & n23933 ) | ( n23932 & n23933 ) ;
  assign n23935 = n23930 & n23934 ;
  assign n23936 = ( n13530 & n23930 ) | ( n13530 & n23935 ) | ( n23930 & n23935 ) ;
  assign n23937 = ~x29 & n23936 ;
  assign n23938 = x29 | n23936 ;
  assign n23939 = ( ~n23936 & n23937 ) | ( ~n23936 & n23938 ) | ( n23937 & n23938 ) ;
  assign n23940 = n23924 & n23939 ;
  assign n23941 = n23924 | n23939 ;
  assign n23942 = ~n23940 & n23941 ;
  assign n23943 = n23374 & n23942 ;
  assign n23944 = ( n23380 & n23942 ) | ( n23380 & n23943 ) | ( n23942 & n23943 ) ;
  assign n23945 = n23374 | n23942 ;
  assign n23946 = n23380 | n23945 ;
  assign n23947 = ~n23944 & n23946 ;
  assign n23949 = n2312 & n14607 ;
  assign n23950 = n2308 & n14329 ;
  assign n23951 = n23949 | n23950 ;
  assign n23948 = n2315 & n14591 ;
  assign n23953 = n2306 | n23948 ;
  assign n23954 = n23951 | n23953 ;
  assign n23952 = n23948 | n23951 ;
  assign n23955 = n23952 & n23954 ;
  assign n23956 = ( n14629 & n23954 ) | ( n14629 & n23955 ) | ( n23954 & n23955 ) ;
  assign n23957 = x26 & n23955 ;
  assign n23958 = x26 & n23954 ;
  assign n23959 = ( n14629 & n23957 ) | ( n14629 & n23958 ) | ( n23957 & n23958 ) ;
  assign n23960 = x26 & ~n23957 ;
  assign n23961 = x26 & ~n23958 ;
  assign n23962 = ( ~n14629 & n23960 ) | ( ~n14629 & n23961 ) | ( n23960 & n23961 ) ;
  assign n23963 = ( n23956 & ~n23959 ) | ( n23956 & n23962 ) | ( ~n23959 & n23962 ) ;
  assign n23964 = n23947 & n23963 ;
  assign n23965 = n23947 | n23963 ;
  assign n23966 = ~n23964 & n23965 ;
  assign n23967 = n23400 | n23403 ;
  assign n23968 = ( n23400 & n23405 ) | ( n23400 & n23967 ) | ( n23405 & n23967 ) ;
  assign n23969 = n23966 & n23968 ;
  assign n23970 = n23966 | n23968 ;
  assign n23971 = ~n23969 & n23970 ;
  assign n23972 = n2932 & n15886 ;
  assign n23973 = n2925 & n15434 ;
  assign n23974 = n2928 & ~n16085 ;
  assign n23975 = n23973 | n23974 ;
  assign n23976 = n23972 | n23975 ;
  assign n23977 = n2936 | n23972 ;
  assign n23978 = n23975 | n23977 ;
  assign n23979 = ( ~n16140 & n23976 ) | ( ~n16140 & n23978 ) | ( n23976 & n23978 ) ;
  assign n23980 = ~x23 & n23978 ;
  assign n23981 = ~x23 & n23976 ;
  assign n23982 = ( ~n16140 & n23980 ) | ( ~n16140 & n23981 ) | ( n23980 & n23981 ) ;
  assign n23983 = x23 | n23981 ;
  assign n23984 = x23 | n23980 ;
  assign n23985 = ( ~n16140 & n23983 ) | ( ~n16140 & n23984 ) | ( n23983 & n23984 ) ;
  assign n23986 = ( ~n23979 & n23982 ) | ( ~n23979 & n23985 ) | ( n23982 & n23985 ) ;
  assign n23987 = n23971 & n23986 ;
  assign n23988 = ~n23971 & n23986 ;
  assign n23989 = ( n23971 & ~n23987 ) | ( n23971 & n23988 ) | ( ~n23987 & n23988 ) ;
  assign n23990 = n23424 | n23426 ;
  assign n23991 = ( n23424 & n23428 ) | ( n23424 & n23990 ) | ( n23428 & n23990 ) ;
  assign n23992 = n23989 & n23991 ;
  assign n23993 = n23989 | n23991 ;
  assign n23994 = ~n23992 & n23993 ;
  assign n23995 = n3544 & ~n16069 ;
  assign n23996 = n3541 & n17111 ;
  assign n23997 = n23995 | n23996 ;
  assign n23998 = n3547 & n17100 ;
  assign n23999 = n3537 | n23998 ;
  assign n24000 = n23997 | n23999 ;
  assign n24001 = n23997 | n23998 ;
  assign n24002 = n17169 | n24001 ;
  assign n24003 = ( ~n17129 & n24001 ) | ( ~n17129 & n24002 ) | ( n24001 & n24002 ) ;
  assign n24004 = n24000 & n24003 ;
  assign n24005 = ( n17161 & n24000 ) | ( n17161 & n24004 ) | ( n24000 & n24004 ) ;
  assign n24006 = ~x20 & n24005 ;
  assign n24007 = x20 | n24005 ;
  assign n24008 = ( ~n24005 & n24006 ) | ( ~n24005 & n24007 ) | ( n24006 & n24007 ) ;
  assign n24009 = n23994 & n24008 ;
  assign n24010 = n23994 | n24008 ;
  assign n24011 = ~n24009 & n24010 ;
  assign n24012 = n23446 | n23449 ;
  assign n24013 = ( n23446 & n23451 ) | ( n23446 & n24012 ) | ( n23451 & n24012 ) ;
  assign n24014 = n24011 & n24013 ;
  assign n24015 = n24011 | n24013 ;
  assign n24016 = ~n24014 & n24015 ;
  assign n24017 = n4471 & ~n18585 ;
  assign n24018 = n4466 & ~n17092 ;
  assign n24019 = n4468 & n18037 ;
  assign n24020 = n24018 | n24019 ;
  assign n24021 = n24017 | n24020 ;
  assign n24022 = n4475 & ~n18675 ;
  assign n24023 = ( n4475 & n18672 ) | ( n4475 & n24022 ) | ( n18672 & n24022 ) ;
  assign n24024 = n24021 | n24023 ;
  assign n24025 = x17 | n24021 ;
  assign n24026 = n24023 | n24025 ;
  assign n24027 = ~x17 & n24025 ;
  assign n24028 = ( ~x17 & n24023 ) | ( ~x17 & n24027 ) | ( n24023 & n24027 ) ;
  assign n24029 = ( ~n24024 & n24026 ) | ( ~n24024 & n24028 ) | ( n24026 & n24028 ) ;
  assign n24030 = n24016 & n24029 ;
  assign n24031 = ~n24016 & n24029 ;
  assign n24032 = ( n24016 & ~n24030 ) | ( n24016 & n24031 ) | ( ~n24030 & n24031 ) ;
  assign n24033 = n23470 & n24032 ;
  assign n24034 = ( n23474 & n24032 ) | ( n23474 & n24033 ) | ( n24032 & n24033 ) ;
  assign n24035 = n23470 | n24032 ;
  assign n24036 = n23474 | n24035 ;
  assign n24037 = ~n24034 & n24036 ;
  assign n24039 = n5237 & n18410 ;
  assign n24040 = n5231 & n18576 ;
  assign n24041 = n24039 | n24040 ;
  assign n24038 = n5234 & n19352 ;
  assign n24043 = n5227 | n24038 ;
  assign n24044 = n24041 | n24043 ;
  assign n24042 = n24038 | n24041 ;
  assign n24045 = n24042 & n24044 ;
  assign n24046 = ( n19674 & n24044 ) | ( n19674 & n24045 ) | ( n24044 & n24045 ) ;
  assign n24047 = x14 & n24045 ;
  assign n24048 = x14 & n24044 ;
  assign n24049 = ( n19674 & n24047 ) | ( n19674 & n24048 ) | ( n24047 & n24048 ) ;
  assign n24050 = x14 & ~n24047 ;
  assign n24051 = x14 & ~n24048 ;
  assign n24052 = ( ~n19674 & n24050 ) | ( ~n19674 & n24051 ) | ( n24050 & n24051 ) ;
  assign n24053 = ( n24046 & ~n24049 ) | ( n24046 & n24052 ) | ( ~n24049 & n24052 ) ;
  assign n24054 = n24037 & n24053 ;
  assign n24055 = n24037 | n24053 ;
  assign n24056 = ~n24054 & n24055 ;
  assign n24057 = n23494 | n23497 ;
  assign n24058 = ( n23494 & n23499 ) | ( n23494 & n24057 ) | ( n23499 & n24057 ) ;
  assign n24059 = n24056 & n24058 ;
  assign n24060 = n24056 | n24058 ;
  assign n24061 = ~n24059 & n24060 ;
  assign n24062 = n6122 & ~n20630 ;
  assign n24063 = n6125 & n19494 ;
  assign n24064 = n6119 & n19631 ;
  assign n24065 = n24063 | n24064 ;
  assign n24066 = n24062 | n24065 ;
  assign n24067 = n6115 | n24062 ;
  assign n24068 = n24065 | n24067 ;
  assign n24069 = ( ~n20709 & n24066 ) | ( ~n20709 & n24068 ) | ( n24066 & n24068 ) ;
  assign n24070 = ~x11 & n24068 ;
  assign n24071 = ~x11 & n24066 ;
  assign n24072 = ( ~n20709 & n24070 ) | ( ~n20709 & n24071 ) | ( n24070 & n24071 ) ;
  assign n24073 = x11 | n24071 ;
  assign n24074 = x11 | n24070 ;
  assign n24075 = ( ~n20709 & n24073 ) | ( ~n20709 & n24074 ) | ( n24073 & n24074 ) ;
  assign n24076 = ( ~n24069 & n24072 ) | ( ~n24069 & n24075 ) | ( n24072 & n24075 ) ;
  assign n24077 = n24061 & n24076 ;
  assign n24078 = ~n24061 & n24076 ;
  assign n24079 = ( n24061 & ~n24077 ) | ( n24061 & n24078 ) | ( ~n24077 & n24078 ) ;
  assign n24080 = n23517 & n24079 ;
  assign n24081 = ( n23521 & n24079 ) | ( n23521 & n24080 ) | ( n24079 & n24080 ) ;
  assign n24082 = n23517 | n24079 ;
  assign n24083 = n23521 | n24082 ;
  assign n24084 = ~n24081 & n24083 ;
  assign n24085 = n7079 & ~n21563 ;
  assign n24086 = n7074 & ~n20618 ;
  assign n24087 = n7068 & n20609 ;
  assign n24088 = n24086 | n24087 ;
  assign n24089 = n24085 | n24088 ;
  assign n24090 = n21570 & ~n24089 ;
  assign n24091 = ( n22270 & n24089 ) | ( n22270 & ~n24090 ) | ( n24089 & ~n24090 ) ;
  assign n24092 = n22304 | n24091 ;
  assign n24093 = n7078 | n24085 ;
  assign n24094 = n24088 | n24093 ;
  assign n24095 = n24092 & n24094 ;
  assign n24096 = ~x8 & n24094 ;
  assign n24097 = n24092 & n24096 ;
  assign n24098 = x8 | n24096 ;
  assign n24099 = ( x8 & n24092 ) | ( x8 & n24098 ) | ( n24092 & n24098 ) ;
  assign n24100 = ( ~n24095 & n24097 ) | ( ~n24095 & n24099 ) | ( n24097 & n24099 ) ;
  assign n24101 = n24084 & n24100 ;
  assign n24102 = n24084 | n24100 ;
  assign n24103 = ~n24101 & n24102 ;
  assign n24104 = n23539 & n24103 ;
  assign n24105 = ( n23545 & n24103 ) | ( n23545 & n24104 ) | ( n24103 & n24104 ) ;
  assign n24106 = n23539 | n24103 ;
  assign n24107 = n23545 | n24106 ;
  assign n24108 = ~n24105 & n24107 ;
  assign n24109 = n8115 & ~n21517 ;
  assign n24110 = n8118 & ~n21551 ;
  assign n24111 = n24109 | n24110 ;
  assign n24112 = n8122 & n23227 ;
  assign n24113 = ( n8122 & n23217 ) | ( n8122 & n24112 ) | ( n23217 & n24112 ) ;
  assign n24114 = n24111 | n24113 ;
  assign n24115 = n8125 & n23299 ;
  assign n24116 = n8125 & n23298 ;
  assign n24117 = ( n21584 & n24115 ) | ( n21584 & n24116 ) | ( n24115 & n24116 ) ;
  assign n24118 = n24114 | n24117 ;
  assign n24119 = n8125 | n24114 ;
  assign n24120 = ( n23289 & n24118 ) | ( n23289 & n24119 ) | ( n24118 & n24119 ) ;
  assign n24121 = x5 | n24120 ;
  assign n24122 = ~x5 & n24120 ;
  assign n24123 = ( ~n24120 & n24121 ) | ( ~n24120 & n24122 ) | ( n24121 & n24122 ) ;
  assign n24124 = n24108 & n24123 ;
  assign n24125 = n24108 & ~n24124 ;
  assign n24126 = x0 | n9024 ;
  assign n24127 = ( ~n8969 & n9024 ) | ( ~n8969 & n24126 ) | ( n9024 & n24126 ) ;
  assign n24128 = ~n23234 & n24127 ;
  assign n24129 = ~n23235 & n24127 ;
  assign n24130 = ( ~n15882 & n24128 ) | ( ~n15882 & n24129 ) | ( n24128 & n24129 ) ;
  assign n24131 = n9021 | n24128 ;
  assign n24132 = n9021 | n24129 ;
  assign n24133 = ( ~n15882 & n24131 ) | ( ~n15882 & n24132 ) | ( n24131 & n24132 ) ;
  assign n24134 = ( ~n23240 & n24130 ) | ( ~n23240 & n24133 ) | ( n24130 & n24133 ) ;
  assign n24135 = ~n23239 & n23240 ;
  assign n24136 = n8970 & ~n24135 ;
  assign n24137 = n8970 & ~n23240 ;
  assign n24138 = ( ~n23575 & n24136 ) | ( ~n23575 & n24137 ) | ( n24136 & n24137 ) ;
  assign n24139 = ( ~n23577 & n24136 ) | ( ~n23577 & n24137 ) | ( n24136 & n24137 ) ;
  assign n24140 = n24138 & n24139 ;
  assign n24141 = n24134 | n24140 ;
  assign n24142 = ( n21554 & n24138 ) | ( n21554 & n24139 ) | ( n24138 & n24139 ) ;
  assign n24143 = n24134 | n24142 ;
  assign n24144 = ( ~n21584 & n24141 ) | ( ~n21584 & n24143 ) | ( n24141 & n24143 ) ;
  assign n24145 = x2 & n24143 ;
  assign n24146 = x2 & n24141 ;
  assign n24147 = ( ~n21584 & n24145 ) | ( ~n21584 & n24146 ) | ( n24145 & n24146 ) ;
  assign n24148 = n24144 & ~n24147 ;
  assign n24149 = x2 & ~n24143 ;
  assign n24150 = x2 & ~n24141 ;
  assign n24151 = ( n21584 & n24149 ) | ( n21584 & n24150 ) | ( n24149 & n24150 ) ;
  assign n24152 = n24148 | n24151 ;
  assign n24153 = ~n24108 & n24123 ;
  assign n24154 = n24152 & n24153 ;
  assign n24155 = ( n24125 & n24152 ) | ( n24125 & n24154 ) | ( n24152 & n24154 ) ;
  assign n24156 = n24152 | n24153 ;
  assign n24157 = n24125 | n24156 ;
  assign n24158 = ~n24155 & n24157 ;
  assign n24159 = n23565 | n23569 ;
  assign n24160 = ( n23565 & n23570 ) | ( n23565 & n24159 ) | ( n23570 & n24159 ) ;
  assign n24161 = n24158 & n24160 ;
  assign n24162 = n24158 | n24160 ;
  assign n24163 = ~n24161 & n24162 ;
  assign n24164 = n23607 | n24163 ;
  assign n24165 = n23612 | n24164 ;
  assign n24166 = ( n23607 & n23612 ) | ( n23607 & n24163 ) | ( n23612 & n24163 ) ;
  assign n24167 = n24165 & ~n24166 ;
  assign n24168 = n23614 | n24167 ;
  assign n24169 = n23614 & n24167 ;
  assign n24170 = n23615 | n23617 ;
  assign n24171 = ( n23615 & n23631 ) | ( n23615 & n24170 ) | ( n23631 & n24170 ) ;
  assign n24172 = n24168 & ~n24169 ;
  assign n24173 = n24169 | n24172 ;
  assign n24174 = ( n24169 & n24171 ) | ( n24169 & n24173 ) | ( n24171 & n24173 ) ;
  assign n24175 = n24168 & ~n24174 ;
  assign n24176 = n2315 & n24167 ;
  assign n24177 = n2312 & n23316 ;
  assign n24178 = n2308 & n23614 ;
  assign n24179 = n24177 | n24178 ;
  assign n24180 = n24176 | n24179 ;
  assign n24181 = n2306 | n24180 ;
  assign n24182 = n24171 & ~n24172 ;
  assign n24183 = ( n24180 & n24181 ) | ( n24180 & n24182 ) | ( n24181 & n24182 ) ;
  assign n24184 = n24180 | n24181 ;
  assign n24185 = ( n24175 & n24183 ) | ( n24175 & n24184 ) | ( n24183 & n24184 ) ;
  assign n24186 = x26 & n24185 ;
  assign n24187 = x26 & ~n24185 ;
  assign n24188 = ( n24185 & ~n24186 ) | ( n24185 & n24187 ) | ( ~n24186 & n24187 ) ;
  assign n24189 = n23870 & n24188 ;
  assign n24190 = ~n23870 & n24188 ;
  assign n24191 = ( n23870 & ~n24189 ) | ( n23870 & n24190 ) | ( ~n24189 & n24190 ) ;
  assign n24192 = n23651 & n24191 ;
  assign n24193 = ( n23806 & n24191 ) | ( n23806 & n24192 ) | ( n24191 & n24192 ) ;
  assign n24194 = n23807 & ~n24193 ;
  assign n24195 = n24191 & ~n24193 ;
  assign n24196 = n24194 | n24195 ;
  assign n24197 = n8969 | n9020 ;
  assign n24198 = ~n23229 & n24197 ;
  assign n24199 = ( n23154 & n24197 ) | ( n23154 & n24198 ) | ( n24197 & n24198 ) ;
  assign n24200 = ~n23232 & n24197 ;
  assign n24201 = ~n23231 & n24197 ;
  assign n24202 = ( n9072 & n24200 ) | ( n9072 & n24201 ) | ( n24200 & n24201 ) ;
  assign n24203 = ( ~n21543 & n24199 ) | ( ~n21543 & n24202 ) | ( n24199 & n24202 ) ;
  assign n24204 = ( ~n21545 & n24199 ) | ( ~n21545 & n24202 ) | ( n24199 & n24202 ) ;
  assign n24205 = ( ~n15882 & n24203 ) | ( ~n15882 & n24204 ) | ( n24203 & n24204 ) ;
  assign n24206 = ~x2 & n24203 ;
  assign n24207 = ~x2 & n24204 ;
  assign n24208 = ( ~n15882 & n24206 ) | ( ~n15882 & n24207 ) | ( n24206 & n24207 ) ;
  assign n24209 = x2 | n24206 ;
  assign n24210 = x2 | n24207 ;
  assign n24211 = ( ~n15882 & n24209 ) | ( ~n15882 & n24210 ) | ( n24209 & n24210 ) ;
  assign n24212 = ( ~n24205 & n24208 ) | ( ~n24205 & n24211 ) | ( n24208 & n24211 ) ;
  assign n24213 = n10769 | n10774 ;
  assign n24214 = n926 & ~n2204 ;
  assign n24215 = ~n3305 & n24214 ;
  assign n24216 = ~n2873 & n24215 ;
  assign n24217 = ~n24213 & n24216 ;
  assign n24218 = n46 | n92 ;
  assign n24219 = n226 | n560 ;
  assign n24220 = n24218 | n24219 ;
  assign n24221 = n159 | n566 ;
  assign n24222 = n24220 | n24221 ;
  assign n24223 = n24217 & ~n24222 ;
  assign n24224 = n5923 | n6827 ;
  assign n24225 = n879 | n24224 ;
  assign n24226 = n649 | n24225 ;
  assign n24227 = n2179 | n24226 ;
  assign n24228 = n257 | n412 ;
  assign n24229 = n1663 | n3445 ;
  assign n24230 = n1307 | n24229 ;
  assign n24231 = n24228 | n24230 ;
  assign n24232 = n24227 | n24231 ;
  assign n24233 = n24223 & ~n24232 ;
  assign n24234 = ~n10727 & n24233 ;
  assign n24235 = n246 | n418 ;
  assign n24236 = n967 | n24235 ;
  assign n24237 = n456 | n775 ;
  assign n24238 = n643 | n24237 ;
  assign n24239 = n24236 | n24238 ;
  assign n24240 = n104 | n356 ;
  assign n24241 = n24239 | n24240 ;
  assign n24242 = n22929 | n24241 ;
  assign n24243 = n24234 & ~n24242 ;
  assign n24244 = n24212 & ~n24243 ;
  assign n24245 = n1057 & n12936 ;
  assign n24246 = n1060 & n12010 ;
  assign n24247 = n1065 & ~n12616 ;
  assign n24248 = n24246 | n24247 ;
  assign n24249 = n24245 | n24248 ;
  assign n24250 = ~n24212 & n24243 ;
  assign n24251 = n24244 | n24250 ;
  assign n24252 = n24249 & ~n24251 ;
  assign n24253 = n24244 | n24252 ;
  assign n24254 = n1062 | n24245 ;
  assign n24255 = n24248 | n24254 ;
  assign n24256 = ~n24251 & n24255 ;
  assign n24257 = n24244 | n24256 ;
  assign n24258 = ( ~n13591 & n24253 ) | ( ~n13591 & n24257 ) | ( n24253 & n24257 ) ;
  assign n24259 = n364 | n617 ;
  assign n24260 = n10727 | n24259 ;
  assign n24261 = n602 | n24260 ;
  assign n24262 = n728 | n1394 ;
  assign n24263 = n10853 | n24262 ;
  assign n24264 = n1232 | n5877 ;
  assign n24265 = n24263 | n24264 ;
  assign n24266 = n24261 | n24265 ;
  assign n24267 = n548 | n19377 ;
  assign n24268 = n24266 | n24267 ;
  assign n24269 = n1460 | n3467 ;
  assign n24270 = n24268 | n24269 ;
  assign n24271 = n630 | n13912 ;
  assign n24272 = n4369 | n24271 ;
  assign n24273 = n6926 | n24272 ;
  assign n24274 = n303 | n1114 ;
  assign n24275 = n250 | n254 ;
  assign n24276 = n24274 | n24275 ;
  assign n24277 = n245 | n24276 ;
  assign n24278 = n1631 | n3312 ;
  assign n24279 = n581 | n720 ;
  assign n24280 = n24278 | n24279 ;
  assign n24281 = n24277 | n24280 ;
  assign n24282 = n24273 | n24281 ;
  assign n24283 = n821 | n24282 ;
  assign n24284 = n966 | n22450 ;
  assign n24285 = n170 | n24284 ;
  assign n24286 = n23172 | n24285 ;
  assign n24287 = n341 | n929 ;
  assign n24288 = n24286 | n24287 ;
  assign n24289 = n2129 | n5907 ;
  assign n24290 = n24288 | n24289 ;
  assign n24291 = n24283 | n24290 ;
  assign n24292 = n24270 | n24291 ;
  assign n24293 = n235 | n711 ;
  assign n24294 = n4197 | n24293 ;
  assign n24295 = n2243 | n24294 ;
  assign n24296 = n5017 | n24295 ;
  assign n24297 = n282 | n15243 ;
  assign n24298 = n24296 | n24297 ;
  assign n24299 = n330 | n406 ;
  assign n24300 = n310 | n858 ;
  assign n24301 = n24299 | n24300 ;
  assign n24302 = n374 | n413 ;
  assign n24303 = n154 | n24302 ;
  assign n24304 = n24301 | n24303 ;
  assign n24305 = n24298 | n24304 ;
  assign n24306 = n24292 | n24305 ;
  assign n24307 = n24212 & n24306 ;
  assign n24308 = n24212 | n24306 ;
  assign n24309 = n24253 & n24308 ;
  assign n24310 = ~n24307 & n24309 ;
  assign n24311 = n24257 & n24308 ;
  assign n24312 = ~n24307 & n24311 ;
  assign n24313 = ( ~n13591 & n24310 ) | ( ~n13591 & n24312 ) | ( n24310 & n24312 ) ;
  assign n24314 = n24258 & ~n24313 ;
  assign n24315 = ~n24307 & n24308 ;
  assign n24316 = ~n24309 & n24315 ;
  assign n24317 = ~n24311 & n24315 ;
  assign n24318 = ( n13591 & n24316 ) | ( n13591 & n24317 ) | ( n24316 & n24317 ) ;
  assign n24319 = n24314 | n24318 ;
  assign n24320 = n1057 & n13235 ;
  assign n24321 = n1060 & ~n12616 ;
  assign n24322 = n1065 & n12936 ;
  assign n24323 = n24321 | n24322 ;
  assign n24324 = n24320 | n24323 ;
  assign n24325 = n1062 | n24320 ;
  assign n24326 = n24323 | n24325 ;
  assign n24327 = ( n13561 & n24324 ) | ( n13561 & n24326 ) | ( n24324 & n24326 ) ;
  assign n24328 = n24319 & n24327 ;
  assign n24329 = n24319 | n24327 ;
  assign n24330 = ~n24328 & n24329 ;
  assign n24331 = ( ~n13591 & n24249 ) | ( ~n13591 & n24255 ) | ( n24249 & n24255 ) ;
  assign n24332 = ( ~n13591 & n24252 ) | ( ~n13591 & n24256 ) | ( n24252 & n24256 ) ;
  assign n24333 = n24331 & ~n24332 ;
  assign n24334 = n24250 | n24257 ;
  assign n24335 = n24250 | n24253 ;
  assign n24336 = ( ~n13591 & n24334 ) | ( ~n13591 & n24335 ) | ( n24334 & n24335 ) ;
  assign n24337 = ~n24333 & n24336 ;
  assign n24338 = n23911 & ~n24336 ;
  assign n24339 = ( n23911 & n24333 ) | ( n23911 & n24338 ) | ( n24333 & n24338 ) ;
  assign n24340 = ( n23920 & ~n24337 ) | ( n23920 & n24339 ) | ( ~n24337 & n24339 ) ;
  assign n24341 = ~n23911 & n24336 ;
  assign n24342 = ~n24333 & n24341 ;
  assign n24343 = ~n23920 & n24342 ;
  assign n24344 = n24340 | n24343 ;
  assign n24345 = n1826 & n13235 ;
  assign n24346 = n1823 & n13522 ;
  assign n24347 = n24345 | n24346 ;
  assign n24348 = n1829 & n14607 ;
  assign n24349 = n1821 | n24348 ;
  assign n24350 = n24347 | n24349 ;
  assign n24351 = n24347 | n24348 ;
  assign n24352 = n14696 | n24351 ;
  assign n24353 = n14698 | n24351 ;
  assign n24354 = ( ~n13248 & n24352 ) | ( ~n13248 & n24353 ) | ( n24352 & n24353 ) ;
  assign n24355 = n24350 & n24354 ;
  assign n24356 = ( n14687 & n24350 ) | ( n14687 & n24355 ) | ( n24350 & n24355 ) ;
  assign n24357 = ~x29 & n24356 ;
  assign n24358 = x29 | n24356 ;
  assign n24359 = ( ~n24356 & n24357 ) | ( ~n24356 & n24358 ) | ( n24357 & n24358 ) ;
  assign n24360 = n24340 | n24359 ;
  assign n24361 = ( n24340 & ~n24344 ) | ( n24340 & n24360 ) | ( ~n24344 & n24360 ) ;
  assign n24362 = n24330 & n24361 ;
  assign n24363 = n24330 | n24361 ;
  assign n24364 = ~n24362 & n24363 ;
  assign n24365 = n1829 & n14329 ;
  assign n24366 = n1826 & n13522 ;
  assign n24367 = n1823 & n14607 ;
  assign n24368 = n24366 | n24367 ;
  assign n24369 = n24365 | n24368 ;
  assign n24370 = n1821 | n24365 ;
  assign n24371 = n24368 | n24370 ;
  assign n24372 = ( n14656 & n24369 ) | ( n14656 & n24371 ) | ( n24369 & n24371 ) ;
  assign n24373 = x29 & n24371 ;
  assign n24374 = x29 & n24369 ;
  assign n24375 = ( n14656 & n24373 ) | ( n14656 & n24374 ) | ( n24373 & n24374 ) ;
  assign n24376 = x29 & ~n24374 ;
  assign n24377 = x29 & ~n24373 ;
  assign n24378 = ( ~n14656 & n24376 ) | ( ~n14656 & n24377 ) | ( n24376 & n24377 ) ;
  assign n24379 = ( n24372 & ~n24375 ) | ( n24372 & n24378 ) | ( ~n24375 & n24378 ) ;
  assign n24380 = n24364 & n24379 ;
  assign n24381 = n24364 & ~n24380 ;
  assign n24382 = n2308 & n15434 ;
  assign n24383 = n2315 & ~n16085 ;
  assign n24384 = n2312 & n14591 ;
  assign n24385 = n24383 | n24384 ;
  assign n24386 = n24382 | n24385 ;
  assign n24387 = n2306 | n24382 ;
  assign n24388 = n24385 | n24387 ;
  assign n24389 = ( ~n16167 & n24386 ) | ( ~n16167 & n24388 ) | ( n24386 & n24388 ) ;
  assign n24390 = ~x26 & n24388 ;
  assign n24391 = ~x26 & n24386 ;
  assign n24392 = ( ~n16167 & n24390 ) | ( ~n16167 & n24391 ) | ( n24390 & n24391 ) ;
  assign n24393 = x26 | n24391 ;
  assign n24394 = x26 | n24390 ;
  assign n24395 = ( ~n16167 & n24393 ) | ( ~n16167 & n24394 ) | ( n24393 & n24394 ) ;
  assign n24396 = ( ~n24389 & n24392 ) | ( ~n24389 & n24395 ) | ( n24392 & n24395 ) ;
  assign n24397 = ~n24364 & n24379 ;
  assign n24398 = n24396 & n24397 ;
  assign n24399 = ( n24381 & n24396 ) | ( n24381 & n24398 ) | ( n24396 & n24398 ) ;
  assign n24400 = n24396 | n24397 ;
  assign n24401 = n24381 | n24400 ;
  assign n24402 = ~n24399 & n24401 ;
  assign n24403 = ~n24344 & n24359 ;
  assign n24404 = n24344 & ~n24359 ;
  assign n24405 = n24403 | n24404 ;
  assign n24406 = n23940 & ~n24405 ;
  assign n24407 = ( n23944 & ~n24405 ) | ( n23944 & n24406 ) | ( ~n24405 & n24406 ) ;
  assign n24408 = ~n23940 & n24405 ;
  assign n24409 = ~n23944 & n24408 ;
  assign n24410 = n24407 | n24409 ;
  assign n24411 = n2315 & n15434 ;
  assign n24412 = n2312 & n14329 ;
  assign n24413 = n2308 & n14591 ;
  assign n24414 = n24412 | n24413 ;
  assign n24415 = n24411 | n24414 ;
  assign n24416 = n2306 | n24411 ;
  assign n24417 = n24414 | n24416 ;
  assign n24418 = ( n15453 & n24415 ) | ( n15453 & n24417 ) | ( n24415 & n24417 ) ;
  assign n24419 = x26 & n24417 ;
  assign n24420 = x26 & n24415 ;
  assign n24421 = ( n15453 & n24419 ) | ( n15453 & n24420 ) | ( n24419 & n24420 ) ;
  assign n24422 = x26 & ~n24420 ;
  assign n24423 = x26 & ~n24419 ;
  assign n24424 = ( ~n15453 & n24422 ) | ( ~n15453 & n24423 ) | ( n24422 & n24423 ) ;
  assign n24425 = ( n24418 & ~n24421 ) | ( n24418 & n24424 ) | ( ~n24421 & n24424 ) ;
  assign n24426 = n24407 | n24425 ;
  assign n24427 = ( n24407 & ~n24410 ) | ( n24407 & n24426 ) | ( ~n24410 & n24426 ) ;
  assign n24428 = n24402 & n24427 ;
  assign n24429 = n24402 | n24427 ;
  assign n24430 = ~n24428 & n24429 ;
  assign n24431 = n2932 & n17111 ;
  assign n24432 = n2925 & n15886 ;
  assign n24433 = n2928 & ~n16069 ;
  assign n24434 = n24432 | n24433 ;
  assign n24435 = n24431 | n24434 ;
  assign n24436 = n2936 & ~n17194 ;
  assign n24437 = ~n17129 & n24436 ;
  assign n24438 = n24435 | n24437 ;
  assign n24439 = n2936 | n24435 ;
  assign n24440 = ( n17186 & n24438 ) | ( n17186 & n24439 ) | ( n24438 & n24439 ) ;
  assign n24441 = x23 | n24440 ;
  assign n24442 = ~x23 & n24440 ;
  assign n24443 = ( ~n24440 & n24441 ) | ( ~n24440 & n24442 ) | ( n24441 & n24442 ) ;
  assign n24444 = n24430 & ~n24443 ;
  assign n24445 = n24430 | n24443 ;
  assign n24446 = ( ~n24430 & n24444 ) | ( ~n24430 & n24445 ) | ( n24444 & n24445 ) ;
  assign n24447 = n24410 | n24425 ;
  assign n24448 = n24410 & ~n24425 ;
  assign n24449 = ( ~n24410 & n24447 ) | ( ~n24410 & n24448 ) | ( n24447 & n24448 ) ;
  assign n24450 = n23964 | n23966 ;
  assign n24451 = ~n24449 & n24450 ;
  assign n24452 = n23964 & ~n24449 ;
  assign n24453 = ( n23968 & n24451 ) | ( n23968 & n24452 ) | ( n24451 & n24452 ) ;
  assign n24454 = n24449 & ~n24450 ;
  assign n24455 = ~n23964 & n24449 ;
  assign n24456 = ( ~n23968 & n24454 ) | ( ~n23968 & n24455 ) | ( n24454 & n24455 ) ;
  assign n24457 = n24453 | n24456 ;
  assign n24458 = n2932 & ~n16069 ;
  assign n24459 = n2925 & ~n16085 ;
  assign n24460 = n2928 & n15886 ;
  assign n24461 = n24459 | n24460 ;
  assign n24462 = n24458 | n24461 ;
  assign n24463 = n2936 | n24462 ;
  assign n24464 = ( ~n16107 & n24462 ) | ( ~n16107 & n24463 ) | ( n24462 & n24463 ) ;
  assign n24465 = ~x23 & n24463 ;
  assign n24466 = ~x23 & n24462 ;
  assign n24467 = ( ~n16107 & n24465 ) | ( ~n16107 & n24466 ) | ( n24465 & n24466 ) ;
  assign n24468 = x23 | n24465 ;
  assign n24469 = x23 | n24466 ;
  assign n24470 = ( ~n16107 & n24468 ) | ( ~n16107 & n24469 ) | ( n24468 & n24469 ) ;
  assign n24471 = ( ~n24464 & n24467 ) | ( ~n24464 & n24470 ) | ( n24467 & n24470 ) ;
  assign n24472 = n24453 | n24471 ;
  assign n24473 = ( n24453 & ~n24457 ) | ( n24453 & n24472 ) | ( ~n24457 & n24472 ) ;
  assign n24474 = n24446 & n24473 ;
  assign n24475 = n24446 | n24473 ;
  assign n24476 = ~n24474 & n24475 ;
  assign n24477 = n3547 & n18037 ;
  assign n24478 = n3544 & n17100 ;
  assign n24479 = n3541 & ~n17092 ;
  assign n24480 = n24478 | n24479 ;
  assign n24481 = n24477 | n24480 ;
  assign n24482 = n3537 | n24477 ;
  assign n24483 = n24480 | n24482 ;
  assign n24484 = ( ~n18050 & n24481 ) | ( ~n18050 & n24483 ) | ( n24481 & n24483 ) ;
  assign n24485 = ~x20 & n24483 ;
  assign n24486 = ~x20 & n24481 ;
  assign n24487 = ( ~n18050 & n24485 ) | ( ~n18050 & n24486 ) | ( n24485 & n24486 ) ;
  assign n24488 = x20 | n24486 ;
  assign n24489 = x20 | n24485 ;
  assign n24490 = ( ~n18050 & n24488 ) | ( ~n18050 & n24489 ) | ( n24488 & n24489 ) ;
  assign n24491 = ( ~n24484 & n24487 ) | ( ~n24484 & n24490 ) | ( n24487 & n24490 ) ;
  assign n24492 = n24476 & ~n24491 ;
  assign n24493 = n24476 | n24491 ;
  assign n24494 = ( ~n24476 & n24492 ) | ( ~n24476 & n24493 ) | ( n24492 & n24493 ) ;
  assign n24495 = n24457 | n24471 ;
  assign n24496 = n24457 & ~n24471 ;
  assign n24497 = ( ~n24457 & n24495 ) | ( ~n24457 & n24496 ) | ( n24495 & n24496 ) ;
  assign n24498 = n23987 | n23989 ;
  assign n24499 = ( n23987 & n23991 ) | ( n23987 & n24498 ) | ( n23991 & n24498 ) ;
  assign n24500 = ~n24497 & n24499 ;
  assign n24501 = n24497 & ~n24499 ;
  assign n24502 = n24500 | n24501 ;
  assign n24503 = n3547 & ~n17092 ;
  assign n24504 = n3544 & n17111 ;
  assign n24505 = n3541 & n17100 ;
  assign n24506 = n24504 | n24505 ;
  assign n24507 = n24503 | n24506 ;
  assign n24508 = n3537 | n24503 ;
  assign n24509 = n24506 | n24508 ;
  assign n24510 = ( ~n17134 & n24507 ) | ( ~n17134 & n24509 ) | ( n24507 & n24509 ) ;
  assign n24511 = ~x20 & n24509 ;
  assign n24512 = ~x20 & n24507 ;
  assign n24513 = ( ~n17134 & n24511 ) | ( ~n17134 & n24512 ) | ( n24511 & n24512 ) ;
  assign n24514 = x20 | n24512 ;
  assign n24515 = x20 | n24511 ;
  assign n24516 = ( ~n17134 & n24514 ) | ( ~n17134 & n24515 ) | ( n24514 & n24515 ) ;
  assign n24517 = ( ~n24510 & n24513 ) | ( ~n24510 & n24516 ) | ( n24513 & n24516 ) ;
  assign n24518 = n24500 | n24517 ;
  assign n24519 = ( n24500 & ~n24502 ) | ( n24500 & n24518 ) | ( ~n24502 & n24518 ) ;
  assign n24520 = n24494 & n24519 ;
  assign n24521 = n24494 | n24519 ;
  assign n24522 = ~n24520 & n24521 ;
  assign n24523 = n4471 & n18576 ;
  assign n24524 = n4466 & ~n18585 ;
  assign n24525 = n4468 & n18410 ;
  assign n24526 = n24524 | n24525 ;
  assign n24527 = n24523 | n24526 ;
  assign n24528 = n4475 | n24523 ;
  assign n24529 = n24526 | n24528 ;
  assign n24530 = ( n18612 & n24527 ) | ( n18612 & n24529 ) | ( n24527 & n24529 ) ;
  assign n24531 = x17 & n24529 ;
  assign n24532 = x17 & n24527 ;
  assign n24533 = ( n18612 & n24531 ) | ( n18612 & n24532 ) | ( n24531 & n24532 ) ;
  assign n24534 = x17 & ~n24532 ;
  assign n24535 = x17 & ~n24531 ;
  assign n24536 = ( ~n18612 & n24534 ) | ( ~n18612 & n24535 ) | ( n24534 & n24535 ) ;
  assign n24537 = ( n24530 & ~n24533 ) | ( n24530 & n24536 ) | ( ~n24533 & n24536 ) ;
  assign n24538 = n24522 & ~n24537 ;
  assign n24539 = n24522 | n24537 ;
  assign n24540 = ( ~n24522 & n24538 ) | ( ~n24522 & n24539 ) | ( n24538 & n24539 ) ;
  assign n24541 = n24502 | n24517 ;
  assign n24542 = n24502 & ~n24517 ;
  assign n24543 = ( ~n24502 & n24541 ) | ( ~n24502 & n24542 ) | ( n24541 & n24542 ) ;
  assign n24544 = n24009 | n24011 ;
  assign n24545 = ~n24543 & n24544 ;
  assign n24546 = n24009 & ~n24543 ;
  assign n24547 = ( n24013 & n24545 ) | ( n24013 & n24546 ) | ( n24545 & n24546 ) ;
  assign n24548 = n24543 & ~n24544 ;
  assign n24549 = ~n24009 & n24543 ;
  assign n24550 = ( ~n24013 & n24548 ) | ( ~n24013 & n24549 ) | ( n24548 & n24549 ) ;
  assign n24551 = n24547 | n24550 ;
  assign n24552 = n4471 & n18410 ;
  assign n24553 = n4466 & n18037 ;
  assign n24554 = n4468 & ~n18585 ;
  assign n24555 = n24553 | n24554 ;
  assign n24556 = n24552 | n24555 ;
  assign n24557 = n4475 & ~n18586 ;
  assign n24558 = ~n18609 & n24557 ;
  assign n24559 = ( n4475 & n18650 ) | ( n4475 & n24558 ) | ( n18650 & n24558 ) ;
  assign n24560 = n24556 | n24559 ;
  assign n24561 = x17 | n24556 ;
  assign n24562 = n24559 | n24561 ;
  assign n24563 = ~x17 & n24561 ;
  assign n24564 = ( ~x17 & n24559 ) | ( ~x17 & n24563 ) | ( n24559 & n24563 ) ;
  assign n24565 = ( ~n24560 & n24562 ) | ( ~n24560 & n24564 ) | ( n24562 & n24564 ) ;
  assign n24566 = n24547 | n24565 ;
  assign n24567 = ( n24547 & ~n24551 ) | ( n24547 & n24566 ) | ( ~n24551 & n24566 ) ;
  assign n24568 = n24540 & n24567 ;
  assign n24569 = n24540 | n24567 ;
  assign n24570 = ~n24568 & n24569 ;
  assign n24571 = n5234 & n19631 ;
  assign n24572 = n5237 & n19352 ;
  assign n24573 = n5231 & n19494 ;
  assign n24574 = n24572 | n24573 ;
  assign n24575 = n24571 | n24574 ;
  assign n24576 = n5227 & n19652 ;
  assign n24577 = n5227 & n19655 ;
  assign n24578 = ( ~n18604 & n24576 ) | ( ~n18604 & n24577 ) | ( n24576 & n24577 ) ;
  assign n24579 = n24575 | n24578 ;
  assign n24580 = n5227 | n24575 ;
  assign n24581 = ( n19640 & n24579 ) | ( n19640 & n24580 ) | ( n24579 & n24580 ) ;
  assign n24582 = x14 | n24581 ;
  assign n24583 = ~x14 & n24581 ;
  assign n24584 = ( ~n24581 & n24582 ) | ( ~n24581 & n24583 ) | ( n24582 & n24583 ) ;
  assign n24585 = n24570 & ~n24584 ;
  assign n24586 = n24570 | n24584 ;
  assign n24587 = ( ~n24570 & n24585 ) | ( ~n24570 & n24586 ) | ( n24585 & n24586 ) ;
  assign n24588 = n24551 | n24565 ;
  assign n24589 = n24551 & ~n24565 ;
  assign n24590 = ( ~n24551 & n24588 ) | ( ~n24551 & n24589 ) | ( n24588 & n24589 ) ;
  assign n24591 = n24030 & ~n24590 ;
  assign n24592 = ( n24034 & ~n24590 ) | ( n24034 & n24591 ) | ( ~n24590 & n24591 ) ;
  assign n24593 = ~n24030 & n24590 ;
  assign n24594 = ~n24034 & n24593 ;
  assign n24595 = n24592 | n24594 ;
  assign n24596 = n5234 & n19494 ;
  assign n24597 = n5237 & n18576 ;
  assign n24598 = n5231 & n19352 ;
  assign n24599 = n24597 | n24598 ;
  assign n24600 = n24596 | n24599 ;
  assign n24601 = n5227 | n24596 ;
  assign n24602 = n24599 | n24601 ;
  assign n24603 = ( n20320 & n24600 ) | ( n20320 & n24602 ) | ( n24600 & n24602 ) ;
  assign n24604 = x14 & n24602 ;
  assign n24605 = x14 & n24600 ;
  assign n24606 = ( n20320 & n24604 ) | ( n20320 & n24605 ) | ( n24604 & n24605 ) ;
  assign n24607 = x14 & ~n24605 ;
  assign n24608 = x14 & ~n24604 ;
  assign n24609 = ( ~n20320 & n24607 ) | ( ~n20320 & n24608 ) | ( n24607 & n24608 ) ;
  assign n24610 = ( n24603 & ~n24606 ) | ( n24603 & n24609 ) | ( ~n24606 & n24609 ) ;
  assign n24611 = n24592 | n24610 ;
  assign n24612 = ( n24592 & ~n24595 ) | ( n24592 & n24611 ) | ( ~n24595 & n24611 ) ;
  assign n24613 = n24587 & n24612 ;
  assign n24614 = n24587 | n24612 ;
  assign n24615 = ~n24613 & n24614 ;
  assign n24616 = n6122 & n20609 ;
  assign n24617 = n6125 & ~n20630 ;
  assign n24618 = n6119 & ~n20618 ;
  assign n24619 = n24617 | n24618 ;
  assign n24620 = n24616 | n24619 ;
  assign n24621 = n6115 | n24616 ;
  assign n24622 = n24619 | n24621 ;
  assign n24623 = ( n20659 & n24620 ) | ( n20659 & n24622 ) | ( n24620 & n24622 ) ;
  assign n24624 = n24620 & n24622 ;
  assign n24625 = ( ~n20649 & n24623 ) | ( ~n20649 & n24624 ) | ( n24623 & n24624 ) ;
  assign n24626 = x11 & n24625 ;
  assign n24627 = x11 & ~n24625 ;
  assign n24628 = ( n24625 & ~n24626 ) | ( n24625 & n24627 ) | ( ~n24626 & n24627 ) ;
  assign n24629 = n24615 & ~n24628 ;
  assign n24630 = n24615 | n24628 ;
  assign n24631 = ( ~n24615 & n24629 ) | ( ~n24615 & n24630 ) | ( n24629 & n24630 ) ;
  assign n24632 = n24595 | n24610 ;
  assign n24633 = n24595 & ~n24610 ;
  assign n24634 = ( ~n24595 & n24632 ) | ( ~n24595 & n24633 ) | ( n24632 & n24633 ) ;
  assign n24635 = n24054 | n24056 ;
  assign n24636 = ~n24634 & n24635 ;
  assign n24637 = n24054 & ~n24634 ;
  assign n24638 = ( n24058 & n24636 ) | ( n24058 & n24637 ) | ( n24636 & n24637 ) ;
  assign n24639 = n24634 & ~n24635 ;
  assign n24640 = ~n24054 & n24634 ;
  assign n24641 = ( ~n24058 & n24639 ) | ( ~n24058 & n24640 ) | ( n24639 & n24640 ) ;
  assign n24642 = n24638 | n24641 ;
  assign n24643 = n6115 & n20680 ;
  assign n24644 = n6122 & ~n20618 ;
  assign n24645 = n6125 & n19631 ;
  assign n24646 = n6119 & ~n20630 ;
  assign n24647 = n24645 | n24646 ;
  assign n24648 = n24644 | n24647 ;
  assign n24649 = n20689 | n24648 ;
  assign n24650 = n6115 | n24648 ;
  assign n24651 = ( n24643 & n24649 ) | ( n24643 & n24650 ) | ( n24649 & n24650 ) ;
  assign n24652 = x11 | n24651 ;
  assign n24653 = ~x11 & n24651 ;
  assign n24654 = ( ~n24651 & n24652 ) | ( ~n24651 & n24653 ) | ( n24652 & n24653 ) ;
  assign n24655 = n24638 | n24654 ;
  assign n24656 = ( n24638 & ~n24642 ) | ( n24638 & n24655 ) | ( ~n24642 & n24655 ) ;
  assign n24657 = n24631 & n24656 ;
  assign n24658 = n24631 | n24656 ;
  assign n24659 = ~n24657 & n24658 ;
  assign n24660 = n7079 & ~n21551 ;
  assign n24661 = n7074 & ~n21563 ;
  assign n24662 = n7068 & ~n21517 ;
  assign n24663 = n24661 | n24662 ;
  assign n24664 = n24660 | n24663 ;
  assign n24665 = n7078 | n24660 ;
  assign n24666 = n24663 | n24665 ;
  assign n24667 = ( ~n21587 & n24664 ) | ( ~n21587 & n24666 ) | ( n24664 & n24666 ) ;
  assign n24668 = ~x8 & n24666 ;
  assign n24669 = ~x8 & n24664 ;
  assign n24670 = ( ~n21587 & n24668 ) | ( ~n21587 & n24669 ) | ( n24668 & n24669 ) ;
  assign n24671 = x8 | n24669 ;
  assign n24672 = x8 | n24668 ;
  assign n24673 = ( ~n21587 & n24671 ) | ( ~n21587 & n24672 ) | ( n24671 & n24672 ) ;
  assign n24674 = ( ~n24667 & n24670 ) | ( ~n24667 & n24673 ) | ( n24670 & n24673 ) ;
  assign n24675 = n24659 & ~n24674 ;
  assign n24676 = n24659 | n24674 ;
  assign n24677 = ( ~n24659 & n24675 ) | ( ~n24659 & n24676 ) | ( n24675 & n24676 ) ;
  assign n24678 = n24642 | n24654 ;
  assign n24679 = n24642 & ~n24654 ;
  assign n24680 = ( ~n24642 & n24678 ) | ( ~n24642 & n24679 ) | ( n24678 & n24679 ) ;
  assign n24681 = n24077 & ~n24680 ;
  assign n24682 = ( n24081 & ~n24680 ) | ( n24081 & n24681 ) | ( ~n24680 & n24681 ) ;
  assign n24683 = ~n24077 & n24680 ;
  assign n24684 = ~n24081 & n24683 ;
  assign n24685 = n24682 | n24684 ;
  assign n24686 = n7079 & ~n21517 ;
  assign n24687 = n7074 & n20609 ;
  assign n24688 = n7068 & ~n21563 ;
  assign n24689 = n24687 | n24688 ;
  assign n24690 = n24686 | n24689 ;
  assign n24691 = n7078 | n24686 ;
  assign n24692 = n24689 | n24691 ;
  assign n24693 = ( ~n22283 & n24690 ) | ( ~n22283 & n24692 ) | ( n24690 & n24692 ) ;
  assign n24694 = n24690 & n24692 ;
  assign n24695 = ( ~n22271 & n24693 ) | ( ~n22271 & n24694 ) | ( n24693 & n24694 ) ;
  assign n24696 = ~x8 & n24695 ;
  assign n24697 = x8 | n24695 ;
  assign n24698 = ( ~n24695 & n24696 ) | ( ~n24695 & n24697 ) | ( n24696 & n24697 ) ;
  assign n24699 = n24682 | n24698 ;
  assign n24700 = ( n24682 & ~n24685 ) | ( n24682 & n24699 ) | ( ~n24685 & n24699 ) ;
  assign n24701 = n24677 & n24700 ;
  assign n24702 = n24677 | n24700 ;
  assign n24703 = ~n24701 & n24702 ;
  assign n24704 = n8118 & ~n23240 ;
  assign n24705 = n8115 & n23227 ;
  assign n24706 = ( n8115 & n23217 ) | ( n8115 & n24705 ) | ( n23217 & n24705 ) ;
  assign n24707 = n24704 | n24706 ;
  assign n24708 = n8122 & ~n23234 ;
  assign n24709 = n8122 & ~n23235 ;
  assign n24710 = ( ~n15882 & n24708 ) | ( ~n15882 & n24709 ) | ( n24708 & n24709 ) ;
  assign n24711 = n24707 | n24710 ;
  assign n24712 = n8125 | n24710 ;
  assign n24713 = n24707 | n24712 ;
  assign n24714 = ( ~n23587 & n24711 ) | ( ~n23587 & n24713 ) | ( n24711 & n24713 ) ;
  assign n24715 = ~x5 & n24713 ;
  assign n24716 = ~x5 & n24711 ;
  assign n24717 = ( ~n23587 & n24715 ) | ( ~n23587 & n24716 ) | ( n24715 & n24716 ) ;
  assign n24718 = x5 | n24716 ;
  assign n24719 = x5 | n24715 ;
  assign n24720 = ( ~n23587 & n24718 ) | ( ~n23587 & n24719 ) | ( n24718 & n24719 ) ;
  assign n24721 = ( ~n24714 & n24717 ) | ( ~n24714 & n24720 ) | ( n24717 & n24720 ) ;
  assign n24722 = n24703 & ~n24721 ;
  assign n24723 = n24703 | n24721 ;
  assign n24724 = ( ~n24703 & n24722 ) | ( ~n24703 & n24723 ) | ( n24722 & n24723 ) ;
  assign n24725 = n24685 | n24698 ;
  assign n24726 = n24685 & ~n24698 ;
  assign n24727 = ( ~n24685 & n24725 ) | ( ~n24685 & n24726 ) | ( n24725 & n24726 ) ;
  assign n24728 = n24101 | n24104 ;
  assign n24729 = n24101 | n24103 ;
  assign n24730 = ( n23545 & n24728 ) | ( n23545 & n24729 ) | ( n24728 & n24729 ) ;
  assign n24731 = ~n24727 & n24730 ;
  assign n24732 = n24727 & ~n24730 ;
  assign n24733 = n24731 | n24732 ;
  assign n24734 = n8122 & ~n23240 ;
  assign n24735 = n8115 & ~n21551 ;
  assign n24736 = n8118 & n23227 ;
  assign n24737 = ( n8118 & n23217 ) | ( n8118 & n24736 ) | ( n23217 & n24736 ) ;
  assign n24738 = n24735 | n24737 ;
  assign n24739 = n24734 | n24738 ;
  assign n24740 = n8125 | n24734 ;
  assign n24741 = n24738 | n24740 ;
  assign n24742 = ( n23260 & n24739 ) | ( n23260 & n24741 ) | ( n24739 & n24741 ) ;
  assign n24743 = x5 & n24741 ;
  assign n24744 = x5 & n24739 ;
  assign n24745 = ( n23260 & n24743 ) | ( n23260 & n24744 ) | ( n24743 & n24744 ) ;
  assign n24746 = x5 & ~n24744 ;
  assign n24747 = x5 & ~n24743 ;
  assign n24748 = ( ~n23260 & n24746 ) | ( ~n23260 & n24747 ) | ( n24746 & n24747 ) ;
  assign n24749 = ( n24742 & ~n24745 ) | ( n24742 & n24748 ) | ( ~n24745 & n24748 ) ;
  assign n24750 = n24731 | n24749 ;
  assign n24751 = ( n24731 & ~n24733 ) | ( n24731 & n24750 ) | ( ~n24733 & n24750 ) ;
  assign n24752 = n24724 & n24751 ;
  assign n24753 = n24724 | n24751 ;
  assign n24754 = ~n24752 & n24753 ;
  assign n24755 = n24124 | n24155 ;
  assign n24756 = n24733 | n24749 ;
  assign n24757 = n24733 & ~n24749 ;
  assign n24758 = ( ~n24733 & n24756 ) | ( ~n24733 & n24757 ) | ( n24756 & n24757 ) ;
  assign n24759 = n24755 & ~n24758 ;
  assign n24760 = ~n24755 & n24758 ;
  assign n24761 = n24759 | n24760 ;
  assign n24762 = n24161 & ~n24761 ;
  assign n24763 = ( n24163 & ~n24761 ) | ( n24163 & n24762 ) | ( ~n24761 & n24762 ) ;
  assign n24764 = ( n23607 & ~n24761 ) | ( n23607 & n24762 ) | ( ~n24761 & n24762 ) ;
  assign n24765 = ( n23612 & n24763 ) | ( n23612 & n24764 ) | ( n24763 & n24764 ) ;
  assign n24766 = n24754 & n24759 ;
  assign n24767 = ( n24754 & n24765 ) | ( n24754 & n24766 ) | ( n24765 & n24766 ) ;
  assign n24768 = n24754 | n24759 ;
  assign n24769 = n24765 | n24768 ;
  assign n24770 = ~n24767 & n24769 ;
  assign n24771 = n8118 | n8122 ;
  assign n24772 = ~n23234 & n24771 ;
  assign n24773 = n8115 | n24772 ;
  assign n24774 = ~n23235 & n24771 ;
  assign n24775 = n8115 | n24774 ;
  assign n24776 = ( ~n15882 & n24773 ) | ( ~n15882 & n24775 ) | ( n24773 & n24775 ) ;
  assign n24777 = n8125 | n24776 ;
  assign n24778 = ( ~n15882 & n24772 ) | ( ~n15882 & n24774 ) | ( n24772 & n24774 ) ;
  assign n24779 = n8125 | n24778 ;
  assign n24780 = ( ~n23240 & n24777 ) | ( ~n23240 & n24779 ) | ( n24777 & n24779 ) ;
  assign n24781 = ( ~n23240 & n24776 ) | ( ~n23240 & n24778 ) | ( n24776 & n24778 ) ;
  assign n24782 = n24135 & ~n24781 ;
  assign n24783 = n23240 & ~n24781 ;
  assign n24784 = ( n23575 & n24782 ) | ( n23575 & n24783 ) | ( n24782 & n24783 ) ;
  assign n24785 = ( n23577 & n24782 ) | ( n23577 & n24783 ) | ( n24782 & n24783 ) ;
  assign n24786 = ( ~n21554 & n24784 ) | ( ~n21554 & n24785 ) | ( n24784 & n24785 ) ;
  assign n24787 = n24780 & ~n24786 ;
  assign n24788 = x5 & ~n24787 ;
  assign n24789 = n24784 | n24785 ;
  assign n24790 = n24780 & ~n24789 ;
  assign n24791 = x5 & ~n24790 ;
  assign n24792 = ( n21584 & n24788 ) | ( n21584 & n24791 ) | ( n24788 & n24791 ) ;
  assign n24793 = ~x5 & n24787 ;
  assign n24794 = ~x5 & n24790 ;
  assign n24795 = ( ~n21584 & n24793 ) | ( ~n21584 & n24794 ) | ( n24793 & n24794 ) ;
  assign n24796 = n24792 | n24795 ;
  assign n24797 = n24657 | n24674 ;
  assign n24798 = ( n24657 & n24659 ) | ( n24657 & n24797 ) | ( n24659 & n24797 ) ;
  assign n24799 = n24796 & n24798 ;
  assign n24800 = n24796 | n24798 ;
  assign n24801 = ~n24799 & n24800 ;
  assign n24802 = n24380 | n24399 ;
  assign n24803 = n514 | n895 ;
  assign n24804 = n104 | n348 ;
  assign n24805 = n24803 | n24804 ;
  assign n24806 = n324 | n24805 ;
  assign n24807 = n483 | n554 ;
  assign n24808 = n704 | n24807 ;
  assign n24809 = n2614 | n24808 ;
  assign n24810 = n18244 | n24809 ;
  assign n24811 = n7837 | n24810 ;
  assign n24812 = n11744 | n24811 ;
  assign n24813 = n138 | n550 ;
  assign n24814 = n638 | n24813 ;
  assign n24815 = n978 | n24814 ;
  assign n24816 = n223 | n370 ;
  assign n24817 = n143 & ~n24816 ;
  assign n24818 = ~n24815 & n24817 ;
  assign n24819 = ~n24812 & n24818 ;
  assign n24820 = ~n18243 & n24819 ;
  assign n24821 = ~n24806 & n24820 ;
  assign n24822 = n24307 | n24309 ;
  assign n24823 = n24307 | n24311 ;
  assign n24824 = ( ~n13591 & n24822 ) | ( ~n13591 & n24823 ) | ( n24822 & n24823 ) ;
  assign n24825 = ( n24212 & n24821 ) | ( n24212 & ~n24824 ) | ( n24821 & ~n24824 ) ;
  assign n24826 = ( ~n24212 & n24824 ) | ( ~n24212 & n24825 ) | ( n24824 & n24825 ) ;
  assign n24827 = ( ~n24821 & n24825 ) | ( ~n24821 & n24826 ) | ( n24825 & n24826 ) ;
  assign n24828 = n1057 & n13522 ;
  assign n24829 = n1060 & n12936 ;
  assign n24830 = n1065 & n13235 ;
  assign n24831 = n24829 | n24830 ;
  assign n24832 = n24828 | n24831 ;
  assign n24833 = n1062 & n13537 ;
  assign n24834 = n1062 & n13539 ;
  assign n24835 = ( ~n13248 & n24833 ) | ( ~n13248 & n24834 ) | ( n24833 & n24834 ) ;
  assign n24836 = n24832 | n24835 ;
  assign n24837 = n1062 | n24832 ;
  assign n24838 = ( n13530 & n24836 ) | ( n13530 & n24837 ) | ( n24836 & n24837 ) ;
  assign n24839 = ~n24825 & n24838 ;
  assign n24840 = n24821 & n24838 ;
  assign n24841 = ( ~n24826 & n24839 ) | ( ~n24826 & n24840 ) | ( n24839 & n24840 ) ;
  assign n24842 = n24827 | n24841 ;
  assign n24843 = n24825 & n24838 ;
  assign n24844 = ~n24821 & n24838 ;
  assign n24845 = ( n24826 & n24843 ) | ( n24826 & n24844 ) | ( n24843 & n24844 ) ;
  assign n24846 = n24842 & ~n24845 ;
  assign n24847 = n24328 | n24330 ;
  assign n24848 = ~n24846 & n24847 ;
  assign n24849 = n24328 & ~n24846 ;
  assign n24850 = ( n24361 & n24848 ) | ( n24361 & n24849 ) | ( n24848 & n24849 ) ;
  assign n24851 = n24846 & ~n24847 ;
  assign n24852 = ~n24328 & n24846 ;
  assign n24853 = ( ~n24361 & n24851 ) | ( ~n24361 & n24852 ) | ( n24851 & n24852 ) ;
  assign n24854 = n24850 | n24853 ;
  assign n24855 = n1829 & n14591 ;
  assign n24856 = n1826 & n14607 ;
  assign n24857 = n1823 & n14329 ;
  assign n24858 = n24856 | n24857 ;
  assign n24859 = n24855 | n24858 ;
  assign n24860 = n1821 | n24855 ;
  assign n24861 = n24858 | n24860 ;
  assign n24862 = ( n14629 & n24859 ) | ( n14629 & n24861 ) | ( n24859 & n24861 ) ;
  assign n24863 = x29 & n24861 ;
  assign n24864 = x29 & n24859 ;
  assign n24865 = ( n14629 & n24863 ) | ( n14629 & n24864 ) | ( n24863 & n24864 ) ;
  assign n24866 = x29 & ~n24864 ;
  assign n24867 = x29 & ~n24863 ;
  assign n24868 = ( ~n14629 & n24866 ) | ( ~n14629 & n24867 ) | ( n24866 & n24867 ) ;
  assign n24869 = ( n24862 & ~n24865 ) | ( n24862 & n24868 ) | ( ~n24865 & n24868 ) ;
  assign n24870 = ~n24854 & n24869 ;
  assign n24871 = n24854 | n24870 ;
  assign n24872 = n2312 & n15434 ;
  assign n24873 = n2308 & ~n16085 ;
  assign n24874 = n2315 & n15886 ;
  assign n24875 = n24873 | n24874 ;
  assign n24876 = n24872 | n24875 ;
  assign n24877 = n2306 | n24872 ;
  assign n24878 = n24875 | n24877 ;
  assign n24879 = ( ~n16140 & n24876 ) | ( ~n16140 & n24878 ) | ( n24876 & n24878 ) ;
  assign n24880 = ~x26 & n24878 ;
  assign n24881 = ~x26 & n24876 ;
  assign n24882 = ( ~n16140 & n24880 ) | ( ~n16140 & n24881 ) | ( n24880 & n24881 ) ;
  assign n24883 = x26 | n24881 ;
  assign n24884 = x26 | n24880 ;
  assign n24885 = ( ~n16140 & n24883 ) | ( ~n16140 & n24884 ) | ( n24883 & n24884 ) ;
  assign n24886 = ( ~n24879 & n24882 ) | ( ~n24879 & n24885 ) | ( n24882 & n24885 ) ;
  assign n24887 = n24854 & n24869 ;
  assign n24888 = n24886 & n24887 ;
  assign n24889 = ( ~n24871 & n24886 ) | ( ~n24871 & n24888 ) | ( n24886 & n24888 ) ;
  assign n24890 = n24886 | n24887 ;
  assign n24891 = n24871 & ~n24890 ;
  assign n24892 = n24889 | n24891 ;
  assign n24893 = n24802 & ~n24892 ;
  assign n24894 = ~n24802 & n24892 ;
  assign n24895 = n24893 | n24894 ;
  assign n24896 = n2932 & n17100 ;
  assign n24897 = n2925 & ~n16069 ;
  assign n24898 = n2928 & n17111 ;
  assign n24899 = n24897 | n24898 ;
  assign n24900 = n24896 | n24899 ;
  assign n24901 = n2936 & n17169 ;
  assign n24902 = ~n17129 & n24901 ;
  assign n24903 = n24900 | n24902 ;
  assign n24904 = n2936 | n24900 ;
  assign n24905 = ( n17161 & n24903 ) | ( n17161 & n24904 ) | ( n24903 & n24904 ) ;
  assign n24906 = x23 | n24905 ;
  assign n24907 = ~x23 & n24905 ;
  assign n24908 = ( ~n24905 & n24906 ) | ( ~n24905 & n24907 ) | ( n24906 & n24907 ) ;
  assign n24909 = ~n24895 & n24908 ;
  assign n24910 = n24895 | n24909 ;
  assign n24912 = n24428 | n24443 ;
  assign n24913 = ( n24428 & n24430 ) | ( n24428 & n24912 ) | ( n24430 & n24912 ) ;
  assign n24911 = n24895 & n24908 ;
  assign n24914 = n24911 & n24913 ;
  assign n24915 = ( ~n24910 & n24913 ) | ( ~n24910 & n24914 ) | ( n24913 & n24914 ) ;
  assign n24916 = n24911 | n24913 ;
  assign n24917 = n24910 & ~n24916 ;
  assign n24918 = n24915 | n24917 ;
  assign n24919 = n3547 & ~n18585 ;
  assign n24920 = n3544 & ~n17092 ;
  assign n24921 = n3541 & n18037 ;
  assign n24922 = n24920 | n24921 ;
  assign n24923 = n24919 | n24922 ;
  assign n24924 = n3537 & ~n18675 ;
  assign n24925 = ( n3537 & n18672 ) | ( n3537 & n24924 ) | ( n18672 & n24924 ) ;
  assign n24926 = n24923 | n24925 ;
  assign n24927 = x20 | n24923 ;
  assign n24928 = n24925 | n24927 ;
  assign n24929 = ~x20 & n24927 ;
  assign n24930 = ( ~x20 & n24925 ) | ( ~x20 & n24929 ) | ( n24925 & n24929 ) ;
  assign n24931 = ( ~n24926 & n24928 ) | ( ~n24926 & n24930 ) | ( n24928 & n24930 ) ;
  assign n24932 = n24918 | n24931 ;
  assign n24933 = n24918 & ~n24931 ;
  assign n24934 = ( ~n24918 & n24932 ) | ( ~n24918 & n24933 ) | ( n24932 & n24933 ) ;
  assign n24935 = n24474 | n24491 ;
  assign n24936 = ( n24474 & n24476 ) | ( n24474 & n24935 ) | ( n24476 & n24935 ) ;
  assign n24937 = ~n24934 & n24936 ;
  assign n24938 = n24934 & ~n24936 ;
  assign n24939 = n24937 | n24938 ;
  assign n24940 = n4471 & n19352 ;
  assign n24941 = n4466 & n18410 ;
  assign n24942 = n4468 & n18576 ;
  assign n24943 = n24941 | n24942 ;
  assign n24944 = n24940 | n24943 ;
  assign n24945 = n4475 | n24940 ;
  assign n24946 = n24943 | n24945 ;
  assign n24947 = ( n19674 & n24944 ) | ( n19674 & n24946 ) | ( n24944 & n24946 ) ;
  assign n24948 = x17 & n24946 ;
  assign n24949 = x17 & n24944 ;
  assign n24950 = ( n19674 & n24948 ) | ( n19674 & n24949 ) | ( n24948 & n24949 ) ;
  assign n24951 = x17 & ~n24949 ;
  assign n24952 = x17 & ~n24948 ;
  assign n24953 = ( ~n19674 & n24951 ) | ( ~n19674 & n24952 ) | ( n24951 & n24952 ) ;
  assign n24954 = ( n24947 & ~n24950 ) | ( n24947 & n24953 ) | ( ~n24950 & n24953 ) ;
  assign n24955 = n24939 | n24954 ;
  assign n24956 = n24939 & ~n24954 ;
  assign n24957 = ( ~n24939 & n24955 ) | ( ~n24939 & n24956 ) | ( n24955 & n24956 ) ;
  assign n24958 = n24520 | n24537 ;
  assign n24959 = ( n24520 & n24522 ) | ( n24520 & n24958 ) | ( n24522 & n24958 ) ;
  assign n24960 = ~n24957 & n24959 ;
  assign n24961 = n24957 & ~n24959 ;
  assign n24962 = n24960 | n24961 ;
  assign n24963 = n5234 & ~n20630 ;
  assign n24964 = n5237 & n19494 ;
  assign n24965 = n5231 & n19631 ;
  assign n24966 = n24964 | n24965 ;
  assign n24967 = n24963 | n24966 ;
  assign n24968 = n5227 | n24963 ;
  assign n24969 = n24966 | n24968 ;
  assign n24970 = ( ~n20709 & n24967 ) | ( ~n20709 & n24969 ) | ( n24967 & n24969 ) ;
  assign n24971 = ~x14 & n24969 ;
  assign n24972 = ~x14 & n24967 ;
  assign n24973 = ( ~n20709 & n24971 ) | ( ~n20709 & n24972 ) | ( n24971 & n24972 ) ;
  assign n24974 = x14 | n24972 ;
  assign n24975 = x14 | n24971 ;
  assign n24976 = ( ~n20709 & n24974 ) | ( ~n20709 & n24975 ) | ( n24974 & n24975 ) ;
  assign n24977 = ( ~n24970 & n24973 ) | ( ~n24970 & n24976 ) | ( n24973 & n24976 ) ;
  assign n24978 = n24962 | n24977 ;
  assign n24979 = n24962 & ~n24977 ;
  assign n24980 = ( ~n24962 & n24978 ) | ( ~n24962 & n24979 ) | ( n24978 & n24979 ) ;
  assign n24981 = n24568 | n24584 ;
  assign n24982 = ( n24568 & n24570 ) | ( n24568 & n24981 ) | ( n24570 & n24981 ) ;
  assign n24983 = ~n24980 & n24982 ;
  assign n24984 = n24980 & ~n24982 ;
  assign n24985 = n24983 | n24984 ;
  assign n24986 = n6122 & ~n21563 ;
  assign n24987 = n6125 & ~n20618 ;
  assign n24988 = n6119 & n20609 ;
  assign n24989 = n24987 | n24988 ;
  assign n24990 = n24986 | n24989 ;
  assign n24991 = n6115 & ~n21570 ;
  assign n24992 = n22270 & n24991 ;
  assign n24993 = ( n6115 & n22304 ) | ( n6115 & n24992 ) | ( n22304 & n24992 ) ;
  assign n24994 = n24990 | n24993 ;
  assign n24995 = x11 | n24990 ;
  assign n24996 = n24993 | n24995 ;
  assign n24997 = ~x11 & n24995 ;
  assign n24998 = ( ~x11 & n24993 ) | ( ~x11 & n24997 ) | ( n24993 & n24997 ) ;
  assign n24999 = ( ~n24994 & n24996 ) | ( ~n24994 & n24998 ) | ( n24996 & n24998 ) ;
  assign n25000 = n24985 | n24999 ;
  assign n25001 = n24985 & ~n24999 ;
  assign n25002 = ( ~n24985 & n25000 ) | ( ~n24985 & n25001 ) | ( n25000 & n25001 ) ;
  assign n25003 = n24613 | n24628 ;
  assign n25004 = ( n24613 & n24615 ) | ( n24613 & n25003 ) | ( n24615 & n25003 ) ;
  assign n25005 = ~n25002 & n25004 ;
  assign n25006 = n25002 & ~n25004 ;
  assign n25007 = n25005 | n25006 ;
  assign n25008 = n7074 & ~n21517 ;
  assign n25009 = n7068 & ~n21551 ;
  assign n25010 = n25008 | n25009 ;
  assign n25011 = n7079 & n23227 ;
  assign n25012 = ( n7079 & n23217 ) | ( n7079 & n25011 ) | ( n23217 & n25011 ) ;
  assign n25013 = n25010 | n25012 ;
  assign n25014 = n7078 & n23299 ;
  assign n25015 = n7078 & n23298 ;
  assign n25016 = ( n21584 & n25014 ) | ( n21584 & n25015 ) | ( n25014 & n25015 ) ;
  assign n25017 = n25013 | n25016 ;
  assign n25018 = n7078 | n25013 ;
  assign n25019 = ( n23289 & n25017 ) | ( n23289 & n25018 ) | ( n25017 & n25018 ) ;
  assign n25020 = x8 | n25019 ;
  assign n25021 = ~x8 & n25019 ;
  assign n25022 = ( ~n25019 & n25020 ) | ( ~n25019 & n25021 ) | ( n25020 & n25021 ) ;
  assign n25023 = n25007 | n25022 ;
  assign n25024 = n25007 & ~n25022 ;
  assign n25025 = ( ~n25007 & n25023 ) | ( ~n25007 & n25024 ) | ( n25023 & n25024 ) ;
  assign n25026 = n24801 & ~n25025 ;
  assign n25027 = n24801 | n25025 ;
  assign n25028 = ( ~n24801 & n25026 ) | ( ~n24801 & n25027 ) | ( n25026 & n25027 ) ;
  assign n25029 = n24701 | n24721 ;
  assign n25030 = ( n24701 & n24703 ) | ( n24701 & n25029 ) | ( n24703 & n25029 ) ;
  assign n25031 = ~n25028 & n25030 ;
  assign n25032 = n25028 & ~n25030 ;
  assign n25033 = n25031 | n25032 ;
  assign n25034 = n24724 & ~n25033 ;
  assign n25035 = n24751 & n25034 ;
  assign n25036 = ( n24754 & ~n25033 ) | ( n24754 & n25035 ) | ( ~n25033 & n25035 ) ;
  assign n25037 = ( n24759 & n25035 ) | ( n24759 & n25036 ) | ( n25035 & n25036 ) ;
  assign n25038 = n25035 | n25036 ;
  assign n25039 = ( n24765 & n25037 ) | ( n24765 & n25038 ) | ( n25037 & n25038 ) ;
  assign n25040 = n24752 | n24754 ;
  assign n25041 = n24752 | n25040 ;
  assign n25042 = n25033 & ~n25041 ;
  assign n25043 = ( n24752 & n24759 ) | ( n24752 & n25040 ) | ( n24759 & n25040 ) ;
  assign n25044 = n25033 & ~n25043 ;
  assign n25045 = ( ~n24765 & n25042 ) | ( ~n24765 & n25044 ) | ( n25042 & n25044 ) ;
  assign n25046 = n25039 | n25045 ;
  assign n25047 = n24770 & ~n25046 ;
  assign n25048 = ~n24770 & n25046 ;
  assign n25049 = n25047 | n25048 ;
  assign n25050 = ~n24161 & n24761 ;
  assign n25051 = ~n24163 & n25050 ;
  assign n25052 = ~n23607 & n25050 ;
  assign n25053 = ( ~n23612 & n25051 ) | ( ~n23612 & n25052 ) | ( n25051 & n25052 ) ;
  assign n25054 = n24765 | n25053 ;
  assign n25055 = n24770 & ~n25054 ;
  assign n25056 = ~n24770 & n25054 ;
  assign n25057 = n25055 | n25056 ;
  assign n25058 = n24167 & ~n25054 ;
  assign n25059 = ~n24167 & n25054 ;
  assign n25060 = n25058 | n25059 ;
  assign n25061 = ~n25058 & n25060 ;
  assign n25062 = n25057 | n25061 ;
  assign n25063 = ~n25057 & n25058 ;
  assign n25064 = ( n24174 & ~n25062 ) | ( n24174 & n25063 ) | ( ~n25062 & n25063 ) ;
  assign n25065 = ~n25049 & n25055 ;
  assign n25066 = ( ~n25049 & n25064 ) | ( ~n25049 & n25065 ) | ( n25064 & n25065 ) ;
  assign n25067 = n25049 & ~n25055 ;
  assign n25068 = ~n25064 & n25067 ;
  assign n25069 = n25066 | n25068 ;
  assign n25070 = n2932 & ~n25046 ;
  assign n25071 = n2925 & ~n25054 ;
  assign n25072 = n2928 & n24770 ;
  assign n25073 = n25071 | n25072 ;
  assign n25074 = n25070 | n25073 ;
  assign n25075 = n2936 | n25070 ;
  assign n25076 = n25073 | n25075 ;
  assign n25077 = ( ~n25069 & n25074 ) | ( ~n25069 & n25076 ) | ( n25074 & n25076 ) ;
  assign n25078 = ~x23 & n25076 ;
  assign n25079 = ~x23 & n25074 ;
  assign n25080 = ( ~n25069 & n25078 ) | ( ~n25069 & n25079 ) | ( n25078 & n25079 ) ;
  assign n25081 = x23 | n25079 ;
  assign n25082 = x23 | n25078 ;
  assign n25083 = ( ~n25069 & n25081 ) | ( ~n25069 & n25082 ) | ( n25081 & n25082 ) ;
  assign n25084 = ( ~n25077 & n25080 ) | ( ~n25077 & n25083 ) | ( n25080 & n25083 ) ;
  assign n25085 = n24196 & n25084 ;
  assign n25086 = n24196 & ~n25085 ;
  assign n25087 = ~n24196 & n25084 ;
  assign n25088 = n25086 | n25087 ;
  assign n25089 = n23805 & ~n23806 ;
  assign n25090 = n23654 | n23806 ;
  assign n25091 = ~n25089 & n25090 ;
  assign n25092 = n25057 & n25061 ;
  assign n25093 = n25057 & ~n25058 ;
  assign n25094 = ( ~n24174 & n25092 ) | ( ~n24174 & n25093 ) | ( n25092 & n25093 ) ;
  assign n25095 = n25064 | n25094 ;
  assign n25096 = n2932 & n24770 ;
  assign n25097 = n2925 & n24167 ;
  assign n25098 = n2928 & ~n25054 ;
  assign n25099 = n25097 | n25098 ;
  assign n25100 = n25096 | n25099 ;
  assign n25101 = n2936 | n25100 ;
  assign n25102 = ( ~n25095 & n25100 ) | ( ~n25095 & n25101 ) | ( n25100 & n25101 ) ;
  assign n25103 = ~x23 & n25101 ;
  assign n25104 = ~x23 & n25100 ;
  assign n25105 = ( ~n25095 & n25103 ) | ( ~n25095 & n25104 ) | ( n25103 & n25104 ) ;
  assign n25106 = x23 | n25103 ;
  assign n25107 = x23 | n25104 ;
  assign n25108 = ( ~n25095 & n25106 ) | ( ~n25095 & n25107 ) | ( n25106 & n25107 ) ;
  assign n25109 = ( ~n25102 & n25105 ) | ( ~n25102 & n25108 ) | ( n25105 & n25108 ) ;
  assign n25110 = ~n25091 & n25109 ;
  assign n25111 = n25091 | n25110 ;
  assign n25112 = n23683 & n23803 ;
  assign n25113 = n23683 | n23803 ;
  assign n25114 = ~n25112 & n25113 ;
  assign n25115 = n2932 & ~n25054 ;
  assign n25116 = n2925 & n23614 ;
  assign n25117 = n2928 & n24167 ;
  assign n25118 = n25116 | n25117 ;
  assign n25119 = n25115 | n25118 ;
  assign n25120 = n24174 & ~n25060 ;
  assign n25121 = ~n24174 & n25060 ;
  assign n25122 = n25120 | n25121 ;
  assign n25123 = n2936 | n25115 ;
  assign n25124 = n25118 | n25123 ;
  assign n25125 = ( n25119 & ~n25122 ) | ( n25119 & n25124 ) | ( ~n25122 & n25124 ) ;
  assign n25126 = ~x23 & n25124 ;
  assign n25127 = ~x23 & n25119 ;
  assign n25128 = ( ~n25122 & n25126 ) | ( ~n25122 & n25127 ) | ( n25126 & n25127 ) ;
  assign n25129 = x23 | n25127 ;
  assign n25130 = x23 | n25126 ;
  assign n25131 = ( ~n25122 & n25129 ) | ( ~n25122 & n25130 ) | ( n25129 & n25130 ) ;
  assign n25132 = ( ~n25125 & n25128 ) | ( ~n25125 & n25131 ) | ( n25128 & n25131 ) ;
  assign n25133 = ~n25114 & n25132 ;
  assign n25134 = n25114 & ~n25132 ;
  assign n25135 = n25133 | n25134 ;
  assign n25136 = n23708 | n23801 ;
  assign n25137 = ~n23802 & n25136 ;
  assign n25138 = n2932 & n24167 ;
  assign n25139 = n2925 & n23316 ;
  assign n25140 = n2928 & n23614 ;
  assign n25141 = n25139 | n25140 ;
  assign n25142 = n25138 | n25141 ;
  assign n25143 = n2936 | n25142 ;
  assign n25144 = ( n24182 & n25142 ) | ( n24182 & n25143 ) | ( n25142 & n25143 ) ;
  assign n25145 = n25142 | n25143 ;
  assign n25146 = ( n24175 & n25144 ) | ( n24175 & n25145 ) | ( n25144 & n25145 ) ;
  assign n25147 = x23 & n25146 ;
  assign n25148 = x23 & ~n25146 ;
  assign n25149 = ( n25146 & ~n25147 ) | ( n25146 & n25148 ) | ( ~n25147 & n25148 ) ;
  assign n25150 = n25137 & n25149 ;
  assign n25151 = n23726 | n23799 ;
  assign n25152 = ~n23800 & n25151 ;
  assign n25153 = n2932 & n23614 ;
  assign n25154 = n2925 & n23620 ;
  assign n25155 = ( n2928 & n11882 ) | ( n2928 & n23620 ) | ( n11882 & n23620 ) ;
  assign n25156 = ( n23316 & n25154 ) | ( n23316 & n25155 ) | ( n25154 & n25155 ) ;
  assign n25158 = n2936 | n25156 ;
  assign n25159 = n25153 | n25158 ;
  assign n25157 = n25153 | n25156 ;
  assign n25160 = n25157 & n25159 ;
  assign n25161 = ( n23634 & n25159 ) | ( n23634 & n25160 ) | ( n25159 & n25160 ) ;
  assign n25162 = x23 & n25160 ;
  assign n25163 = x23 & n25159 ;
  assign n25164 = ( n23634 & n25162 ) | ( n23634 & n25163 ) | ( n25162 & n25163 ) ;
  assign n25165 = x23 & ~n25162 ;
  assign n25166 = x23 & ~n25163 ;
  assign n25167 = ( ~n23634 & n25165 ) | ( ~n23634 & n25166 ) | ( n25165 & n25166 ) ;
  assign n25168 = ( n25161 & ~n25164 ) | ( n25161 & n25167 ) | ( ~n25164 & n25167 ) ;
  assign n25169 = n25152 & n25168 ;
  assign n25170 = n25152 & ~n25169 ;
  assign n25171 = ~n25152 & n25168 ;
  assign n25172 = n25170 | n25171 ;
  assign n25173 = n23779 & n23793 ;
  assign n25174 = n23779 & ~n25173 ;
  assign n25175 = n2925 & ~n22385 ;
  assign n25176 = ( n2928 & n11882 ) | ( n2928 & ~n22385 ) | ( n11882 & ~n22385 ) ;
  assign n25177 = ( n22381 & n25175 ) | ( n22381 & n25176 ) | ( n25175 & n25176 ) ;
  assign n25178 = n2932 | n25177 ;
  assign n25179 = ( n23620 & n25177 ) | ( n23620 & n25178 ) | ( n25177 & n25178 ) ;
  assign n25180 = n2936 | n25179 ;
  assign n25181 = ( ~n23686 & n25179 ) | ( ~n23686 & n25180 ) | ( n25179 & n25180 ) ;
  assign n25182 = ~x23 & n25180 ;
  assign n25183 = ~x23 & n25179 ;
  assign n25184 = ( ~n23686 & n25182 ) | ( ~n23686 & n25183 ) | ( n25182 & n25183 ) ;
  assign n25185 = x23 | n25182 ;
  assign n25186 = x23 | n25183 ;
  assign n25187 = ( ~n23686 & n25185 ) | ( ~n23686 & n25186 ) | ( n25185 & n25186 ) ;
  assign n25188 = ( ~n25181 & n25184 ) | ( ~n25181 & n25187 ) | ( n25184 & n25187 ) ;
  assign n25189 = ~n23779 & n23793 ;
  assign n25190 = n25188 & n25189 ;
  assign n25191 = ( n25174 & n25188 ) | ( n25174 & n25190 ) | ( n25188 & n25190 ) ;
  assign n25192 = n25188 | n25189 ;
  assign n25193 = n25174 | n25192 ;
  assign n25194 = ~n25191 & n25193 ;
  assign n25195 = n23758 & n23776 ;
  assign n25196 = n23758 | n23776 ;
  assign n25197 = ~n25195 & n25196 ;
  assign n25198 = n2932 & n22381 ;
  assign n25199 = n2925 & ~n22398 ;
  assign n25200 = n2928 & ~n22385 ;
  assign n25201 = n25199 | n25200 ;
  assign n25202 = n25198 | n25201 ;
  assign n25203 = n2936 | n25202 ;
  assign n25204 = x23 & n25203 ;
  assign n25205 = x23 & n25202 ;
  assign n25206 = ( n22422 & n25204 ) | ( n22422 & n25205 ) | ( n25204 & n25205 ) ;
  assign n25207 = x23 | n25203 ;
  assign n25208 = x23 | n25202 ;
  assign n25209 = ( n22422 & n25207 ) | ( n22422 & n25208 ) | ( n25207 & n25208 ) ;
  assign n25210 = ~n25206 & n25209 ;
  assign n25211 = n25197 & n25210 ;
  assign n25212 = ~n25197 & n25210 ;
  assign n25213 = ( n25197 & ~n25211 ) | ( n25197 & n25212 ) | ( ~n25211 & n25212 ) ;
  assign n25214 = n23752 | n23754 ;
  assign n25215 = ~n23754 & n23756 ;
  assign n25216 = ( n23753 & n25214 ) | ( n23753 & ~n25215 ) | ( n25214 & ~n25215 ) ;
  assign n25217 = ~n23758 & n25216 ;
  assign n25218 = n2932 & ~n22385 ;
  assign n25219 = n2925 & n22393 ;
  assign n25220 = n2928 & ~n22398 ;
  assign n25221 = n25219 | n25220 ;
  assign n25222 = n25218 | n25221 ;
  assign n25223 = n2936 | n25218 ;
  assign n25224 = n25221 | n25223 ;
  assign n25225 = ( ~n22545 & n25222 ) | ( ~n22545 & n25224 ) | ( n25222 & n25224 ) ;
  assign n25226 = ~x23 & n25224 ;
  assign n25227 = ~x23 & n25222 ;
  assign n25228 = ( ~n22545 & n25226 ) | ( ~n22545 & n25227 ) | ( n25226 & n25227 ) ;
  assign n25229 = x23 | n25227 ;
  assign n25230 = x23 | n25226 ;
  assign n25231 = ( ~n22545 & n25229 ) | ( ~n22545 & n25230 ) | ( n25229 & n25230 ) ;
  assign n25232 = ( ~n25225 & n25228 ) | ( ~n25225 & n25231 ) | ( n25228 & n25231 ) ;
  assign n25233 = n25217 & n25232 ;
  assign n25234 = n2936 & n22474 ;
  assign n25235 = n2928 & ~n22409 ;
  assign n25236 = n2932 & ~n22406 ;
  assign n25237 = n25235 | n25236 ;
  assign n25238 = x23 | n25237 ;
  assign n25239 = n25234 | n25238 ;
  assign n25240 = ~x23 & n25239 ;
  assign n25241 = ( x23 & n13753 ) | ( x23 & n22409 ) | ( n13753 & n22409 ) ;
  assign n25242 = n25239 & n25241 ;
  assign n25243 = n25234 | n25237 ;
  assign n25244 = n25241 & ~n25243 ;
  assign n25245 = ( n25240 & n25242 ) | ( n25240 & n25244 ) | ( n25242 & n25244 ) ;
  assign n25246 = n2932 & n22393 ;
  assign n25247 = n2925 & ~n22409 ;
  assign n25248 = n2928 & ~n22406 ;
  assign n25249 = n25247 | n25248 ;
  assign n25250 = n25246 | n25249 ;
  assign n25251 = n22439 | n25250 ;
  assign n25252 = n2936 | n25246 ;
  assign n25253 = n25249 | n25252 ;
  assign n25254 = ~x23 & n25253 ;
  assign n25255 = n25251 & n25254 ;
  assign n25256 = x23 | n25255 ;
  assign n25257 = n2302 & ~n22409 ;
  assign n25258 = n25255 & n25257 ;
  assign n25259 = n25251 & n25253 ;
  assign n25260 = n25257 & ~n25259 ;
  assign n25261 = ( n25256 & n25258 ) | ( n25256 & n25260 ) | ( n25258 & n25260 ) ;
  assign n25262 = n25245 & n25261 ;
  assign n25263 = ( n25255 & n25256 ) | ( n25255 & ~n25259 ) | ( n25256 & ~n25259 ) ;
  assign n25264 = n25245 | n25257 ;
  assign n25265 = ( n25257 & n25263 ) | ( n25257 & n25264 ) | ( n25263 & n25264 ) ;
  assign n25266 = ~n25262 & n25265 ;
  assign n25267 = n2925 & ~n22406 ;
  assign n25268 = n2928 & n22393 ;
  assign n25269 = n25267 | n25268 ;
  assign n25270 = n2932 & ~n22398 ;
  assign n25271 = n2936 | n25270 ;
  assign n25272 = n25269 | n25271 ;
  assign n25273 = x23 & n25272 ;
  assign n25274 = n25269 | n25270 ;
  assign n25275 = x23 & n25274 ;
  assign n25276 = ( n22608 & n25273 ) | ( n22608 & n25275 ) | ( n25273 & n25275 ) ;
  assign n25277 = x23 | n25272 ;
  assign n25278 = x23 | n25274 ;
  assign n25279 = ( n22608 & n25277 ) | ( n22608 & n25278 ) | ( n25277 & n25278 ) ;
  assign n25280 = ~n25276 & n25279 ;
  assign n25281 = n25262 | n25280 ;
  assign n25282 = ( n25262 & n25266 ) | ( n25262 & n25281 ) | ( n25266 & n25281 ) ;
  assign n25283 = n25217 | n25232 ;
  assign n25284 = ~n25233 & n25283 ;
  assign n25285 = n25233 | n25284 ;
  assign n25286 = ( n25233 & n25282 ) | ( n25233 & n25285 ) | ( n25282 & n25285 ) ;
  assign n25287 = n25213 & n25286 ;
  assign n25288 = n25211 | n25287 ;
  assign n25289 = n25194 & n25288 ;
  assign n25290 = n25191 | n25289 ;
  assign n25291 = n2925 & n22381 ;
  assign n25292 = ( n2928 & n11882 ) | ( n2928 & n22381 ) | ( n11882 & n22381 ) ;
  assign n25293 = ( n23620 & n25291 ) | ( n23620 & n25292 ) | ( n25291 & n25292 ) ;
  assign n25294 = n2932 | n25292 ;
  assign n25295 = n2932 | n25291 ;
  assign n25296 = ( n23620 & n25294 ) | ( n23620 & n25295 ) | ( n25294 & n25295 ) ;
  assign n25297 = ( n23316 & n25293 ) | ( n23316 & n25296 ) | ( n25293 & n25296 ) ;
  assign n25298 = n2936 | n25297 ;
  assign n25299 = ~x23 & n25298 ;
  assign n25300 = ~x23 & n25297 ;
  assign n25301 = ( n23661 & n25299 ) | ( n23661 & n25300 ) | ( n25299 & n25300 ) ;
  assign n25302 = ( x23 & n13713 ) | ( x23 & n25297 ) | ( n13713 & n25297 ) ;
  assign n25303 = x23 & ~n25302 ;
  assign n25304 = x23 & n25297 ;
  assign n25305 = x23 & ~n25304 ;
  assign n25306 = ( ~n23661 & n25303 ) | ( ~n23661 & n25305 ) | ( n25303 & n25305 ) ;
  assign n25307 = n25301 | n25306 ;
  assign n25308 = n23795 & n23797 ;
  assign n25309 = n23795 | n23797 ;
  assign n25310 = ~n25308 & n25309 ;
  assign n25311 = n25307 & n25310 ;
  assign n25312 = n25307 | n25310 ;
  assign n25313 = ~n25311 & n25312 ;
  assign n25314 = n25311 | n25313 ;
  assign n25315 = ( n25290 & n25311 ) | ( n25290 & n25314 ) | ( n25311 & n25314 ) ;
  assign n25316 = n25172 & n25315 ;
  assign n25317 = n25169 | n25316 ;
  assign n25318 = n25137 | n25149 ;
  assign n25319 = ~n25150 & n25318 ;
  assign n25320 = n25150 | n25319 ;
  assign n25321 = ( n25150 & n25317 ) | ( n25150 & n25320 ) | ( n25317 & n25320 ) ;
  assign n25322 = ~n25135 & n25321 ;
  assign n25323 = n25133 | n25322 ;
  assign n25324 = n25091 & n25109 ;
  assign n25325 = n25323 & n25324 ;
  assign n25326 = ( ~n25111 & n25323 ) | ( ~n25111 & n25325 ) | ( n25323 & n25325 ) ;
  assign n25327 = n25110 | n25326 ;
  assign n25328 = n25088 & n25327 ;
  assign n25329 = n24189 | n24193 ;
  assign n25330 = n1826 & n22381 ;
  assign n25331 = ( n1823 & n13998 ) | ( n1823 & n22381 ) | ( n13998 & n22381 ) ;
  assign n25332 = ( n23620 & n25330 ) | ( n23620 & n25331 ) | ( n25330 & n25331 ) ;
  assign n25333 = n1829 | n25331 ;
  assign n25334 = n1829 | n25330 ;
  assign n25335 = ( n23620 & n25333 ) | ( n23620 & n25334 ) | ( n25333 & n25334 ) ;
  assign n25336 = ( n23316 & n25332 ) | ( n23316 & n25335 ) | ( n25332 & n25335 ) ;
  assign n25337 = n1821 | n25336 ;
  assign n25338 = ~x29 & n25337 ;
  assign n25339 = ~x29 & n25336 ;
  assign n25340 = ( n23661 & n25338 ) | ( n23661 & n25339 ) | ( n25338 & n25339 ) ;
  assign n25341 = ( x29 & n10963 ) | ( x29 & n25336 ) | ( n10963 & n25336 ) ;
  assign n25342 = x29 & ~n25341 ;
  assign n25343 = x29 & n25336 ;
  assign n25344 = x29 & ~n25343 ;
  assign n25345 = ( ~n23661 & n25342 ) | ( ~n23661 & n25344 ) | ( n25342 & n25344 ) ;
  assign n25346 = n25340 | n25345 ;
  assign n25347 = n1057 & ~n22385 ;
  assign n25348 = n1065 & ~n22398 ;
  assign n25349 = n1060 & n22393 ;
  assign n25350 = n25348 | n25349 ;
  assign n25351 = n25347 | n25350 ;
  assign n25352 = n1062 | n25347 ;
  assign n25353 = n25350 | n25352 ;
  assign n25354 = ( ~n22545 & n25351 ) | ( ~n22545 & n25353 ) | ( n25351 & n25353 ) ;
  assign n25355 = n1270 | n1364 ;
  assign n25356 = n12683 | n25355 ;
  assign n25357 = n950 | n5069 ;
  assign n25358 = n7882 | n15196 ;
  assign n25359 = n606 | n779 ;
  assign n25360 = n6932 | n25359 ;
  assign n25361 = n25358 | n25360 ;
  assign n25362 = n67 | n503 ;
  assign n25363 = n4197 | n25362 ;
  assign n25364 = n257 | n25363 ;
  assign n25365 = n886 | n18439 ;
  assign n25366 = n25364 | n25365 ;
  assign n25367 = n25361 | n25366 ;
  assign n25368 = ( n25356 & n25357 ) | ( n25356 & ~n25367 ) | ( n25357 & ~n25367 ) ;
  assign n25369 = n648 | n938 ;
  assign n25370 = n479 | n638 ;
  assign n25371 = n25369 | n25370 ;
  assign n25372 = n321 | n858 ;
  assign n25373 = n395 | n25372 ;
  assign n25374 = n25371 | n25373 ;
  assign n25375 = n501 | n25374 ;
  assign n25376 = n857 | n980 ;
  assign n25377 = n9111 | n25376 ;
  assign n25378 = n263 | n402 ;
  assign n25379 = n112 | n246 ;
  assign n25380 = n128 | n171 ;
  assign n25381 = n25379 | n25380 ;
  assign n25382 = n25378 | n25381 ;
  assign n25383 = n25377 | n25382 ;
  assign n25384 = n25375 | n25383 ;
  assign n25385 = n25367 | n25384 ;
  assign n25386 = n25368 | n25385 ;
  assign n25387 = n654 | n979 ;
  assign n25388 = n25386 | n25387 ;
  assign n25389 = n15046 & ~n25388 ;
  assign n25390 = n123 | n288 ;
  assign n25391 = n160 | n566 ;
  assign n25392 = n25390 | n25391 ;
  assign n25393 = n25389 & ~n25392 ;
  assign n25394 = n25353 & ~n25393 ;
  assign n25395 = n25347 & ~n25393 ;
  assign n25396 = ( n25350 & ~n25393 ) | ( n25350 & n25395 ) | ( ~n25393 & n25395 ) ;
  assign n25397 = ( ~n22545 & n25394 ) | ( ~n22545 & n25396 ) | ( n25394 & n25396 ) ;
  assign n25398 = n25354 & ~n25397 ;
  assign n25399 = n25353 | n25393 ;
  assign n25400 = n25351 | n25393 ;
  assign n25401 = ( ~n22545 & n25399 ) | ( ~n22545 & n25400 ) | ( n25399 & n25400 ) ;
  assign n25402 = ~n25398 & n25401 ;
  assign n25403 = n23855 | n23859 ;
  assign n25404 = ( n23823 & n23855 ) | ( n23823 & n25403 ) | ( n23855 & n25403 ) ;
  assign n25405 = n25402 & n25404 ;
  assign n25406 = n25402 | n25404 ;
  assign n25407 = ~n25405 & n25406 ;
  assign n25408 = n25346 & ~n25407 ;
  assign n25409 = ~n25346 & n25407 ;
  assign n25410 = n25408 | n25409 ;
  assign n25411 = n23863 | n23865 ;
  assign n25412 = ( n23863 & n23867 ) | ( n23863 & n25411 ) | ( n23867 & n25411 ) ;
  assign n25413 = n25410 & ~n25412 ;
  assign n25414 = ~n25410 & n25412 ;
  assign n25415 = n25413 | n25414 ;
  assign n25416 = n2315 & ~n25054 ;
  assign n25417 = n2312 & n23614 ;
  assign n25418 = n2308 & n24167 ;
  assign n25419 = n25417 | n25418 ;
  assign n25420 = n25416 | n25419 ;
  assign n25421 = n2306 | n25416 ;
  assign n25422 = n25419 | n25421 ;
  assign n25423 = ( ~n25122 & n25420 ) | ( ~n25122 & n25422 ) | ( n25420 & n25422 ) ;
  assign n25424 = ~x26 & n25422 ;
  assign n25425 = ~x26 & n25420 ;
  assign n25426 = ( ~n25122 & n25424 ) | ( ~n25122 & n25425 ) | ( n25424 & n25425 ) ;
  assign n25427 = x26 | n25425 ;
  assign n25428 = x26 | n25424 ;
  assign n25429 = ( ~n25122 & n25427 ) | ( ~n25122 & n25428 ) | ( n25427 & n25428 ) ;
  assign n25430 = ( ~n25423 & n25426 ) | ( ~n25423 & n25429 ) | ( n25426 & n25429 ) ;
  assign n25431 = ~n25415 & n25430 ;
  assign n25432 = n25415 | n25431 ;
  assign n25433 = n25415 & n25430 ;
  assign n25434 = n25432 & ~n25433 ;
  assign n25435 = n25329 | n25434 ;
  assign n25436 = n25329 & n25434 ;
  assign n25437 = n25435 & ~n25436 ;
  assign n25438 = ~n25047 & n25049 ;
  assign n25439 = ( n25047 & n25055 ) | ( n25047 & ~n25438 ) | ( n25055 & ~n25438 ) ;
  assign n25440 = ~n25047 & n25438 ;
  assign n25441 = ( n25064 & n25439 ) | ( n25064 & ~n25440 ) | ( n25439 & ~n25440 ) ;
  assign n25458 = n25005 | n25022 ;
  assign n25459 = ( n25005 & ~n25007 ) | ( n25005 & n25458 ) | ( ~n25007 & n25458 ) ;
  assign n25442 = n7079 & ~n23240 ;
  assign n25443 = n7074 & ~n21551 ;
  assign n25444 = n7068 & n23227 ;
  assign n25445 = ( n7068 & n23217 ) | ( n7068 & n25444 ) | ( n23217 & n25444 ) ;
  assign n25446 = n25443 | n25445 ;
  assign n25447 = n25442 | n25446 ;
  assign n25448 = n7078 | n25442 ;
  assign n25449 = n25446 | n25448 ;
  assign n25450 = ( n23260 & n25447 ) | ( n23260 & n25449 ) | ( n25447 & n25449 ) ;
  assign n25451 = x8 & n25449 ;
  assign n25452 = x8 & n25447 ;
  assign n25453 = ( n23260 & n25451 ) | ( n23260 & n25452 ) | ( n25451 & n25452 ) ;
  assign n25454 = x8 & ~n25452 ;
  assign n25455 = x8 & ~n25451 ;
  assign n25456 = ( ~n23260 & n25454 ) | ( ~n23260 & n25455 ) | ( n25454 & n25455 ) ;
  assign n25457 = ( n25450 & ~n25453 ) | ( n25450 & n25456 ) | ( ~n25453 & n25456 ) ;
  assign n25460 = n25457 & n25459 ;
  assign n25461 = n25459 & ~n25460 ;
  assign n25462 = n24870 | n24889 ;
  assign n25510 = n24212 & ~n24821 ;
  assign n25511 = ~n24212 & n24821 ;
  assign n25512 = n25510 | n25511 ;
  assign n25513 = ~n25510 & n25512 ;
  assign n25514 = n24307 & ~n25511 ;
  assign n25515 = n25510 | n25514 ;
  assign n25516 = ( n24309 & ~n25513 ) | ( n24309 & n25515 ) | ( ~n25513 & n25515 ) ;
  assign n25517 = ( n24311 & ~n25513 ) | ( n24311 & n25515 ) | ( ~n25513 & n25515 ) ;
  assign n25518 = ( ~n13591 & n25516 ) | ( ~n13591 & n25517 ) | ( n25516 & n25517 ) ;
  assign n25463 = n8115 | n24771 ;
  assign n25464 = n8125 | n25463 ;
  assign n25465 = ~n23229 & n25464 ;
  assign n25466 = ( n23154 & n25464 ) | ( n23154 & n25465 ) | ( n25464 & n25465 ) ;
  assign n25467 = ~n23232 & n25464 ;
  assign n25468 = ~n23231 & n25464 ;
  assign n25469 = ( n9072 & n25467 ) | ( n9072 & n25468 ) | ( n25467 & n25468 ) ;
  assign n25470 = ( ~n21543 & n25466 ) | ( ~n21543 & n25469 ) | ( n25466 & n25469 ) ;
  assign n25471 = ~x5 & n25470 ;
  assign n25472 = ( ~n21545 & n25466 ) | ( ~n21545 & n25469 ) | ( n25466 & n25469 ) ;
  assign n25473 = ~x5 & n25472 ;
  assign n25474 = ( ~n15882 & n25471 ) | ( ~n15882 & n25473 ) | ( n25471 & n25473 ) ;
  assign n25475 = x5 & ~n25470 ;
  assign n25476 = x5 & ~n25472 ;
  assign n25477 = ( n15882 & n25475 ) | ( n15882 & n25476 ) | ( n25475 & n25476 ) ;
  assign n25478 = n25474 | n25477 ;
  assign n25479 = n24270 | n24283 ;
  assign n25480 = n290 | n10851 ;
  assign n25481 = n10366 | n25480 ;
  assign n25482 = n1263 | n25481 ;
  assign n25483 = n573 | n869 ;
  assign n25484 = n4186 | n25483 ;
  assign n25485 = n85 | n460 ;
  assign n25486 = n370 | n775 ;
  assign n25487 = n25485 | n25486 ;
  assign n25488 = n237 | n696 ;
  assign n25489 = n143 & ~n309 ;
  assign n25490 = ~n25488 & n25489 ;
  assign n25491 = ~n25487 & n25490 ;
  assign n25492 = ~n25484 & n25491 ;
  assign n25493 = ~n18441 & n25492 ;
  assign n25494 = ~n25482 & n25493 ;
  assign n25495 = ~n341 & n25494 ;
  assign n25496 = n1287 | n3986 ;
  assign n25497 = n258 | n11076 ;
  assign n25498 = n25496 | n25497 ;
  assign n25499 = n450 | n456 ;
  assign n25500 = n518 | n25499 ;
  assign n25501 = n25498 | n25500 ;
  assign n25502 = n25495 & ~n25501 ;
  assign n25503 = ~n25479 & n25502 ;
  assign n25504 = ~n24212 & n25503 ;
  assign n25505 = n24212 & ~n25503 ;
  assign n25506 = n25504 | n25505 ;
  assign n25507 = n25478 | n25506 ;
  assign n25508 = ~n25506 & n25507 ;
  assign n25509 = ( ~n25478 & n25507 ) | ( ~n25478 & n25508 ) | ( n25507 & n25508 ) ;
  assign n25519 = n25509 & ~n25518 ;
  assign n25520 = n25509 & n25518 ;
  assign n25521 = ( n25518 & n25519 ) | ( n25518 & ~n25520 ) | ( n25519 & ~n25520 ) ;
  assign n25522 = n1057 & n14607 ;
  assign n25523 = n1060 & n13235 ;
  assign n25524 = n1065 & n13522 ;
  assign n25525 = n25523 | n25524 ;
  assign n25526 = n25522 | n25525 ;
  assign n25527 = n1062 & n14696 ;
  assign n25528 = n1062 & n14698 ;
  assign n25529 = ( ~n13248 & n25527 ) | ( ~n13248 & n25528 ) | ( n25527 & n25528 ) ;
  assign n25530 = n25526 | n25529 ;
  assign n25531 = n1062 | n25526 ;
  assign n25532 = ( n14687 & n25530 ) | ( n14687 & n25531 ) | ( n25530 & n25531 ) ;
  assign n25533 = ~n25521 & n25532 ;
  assign n25534 = n25521 & ~n25532 ;
  assign n25535 = n25533 | n25534 ;
  assign n25536 = n24841 & ~n25535 ;
  assign n25537 = ( n24849 & ~n25535 ) | ( n24849 & n25536 ) | ( ~n25535 & n25536 ) ;
  assign n25538 = ( n24848 & ~n25535 ) | ( n24848 & n25536 ) | ( ~n25535 & n25536 ) ;
  assign n25539 = ( n24361 & n25537 ) | ( n24361 & n25538 ) | ( n25537 & n25538 ) ;
  assign n25540 = ~n24841 & n25535 ;
  assign n25541 = ~n24849 & n25540 ;
  assign n25542 = ~n24848 & n25540 ;
  assign n25543 = ( ~n24361 & n25541 ) | ( ~n24361 & n25542 ) | ( n25541 & n25542 ) ;
  assign n25544 = n25539 | n25543 ;
  assign n25545 = n1829 & n15434 ;
  assign n25546 = n1826 & n14329 ;
  assign n25547 = n1823 & n14591 ;
  assign n25548 = n25546 | n25547 ;
  assign n25549 = n25545 | n25548 ;
  assign n25550 = n1821 | n25545 ;
  assign n25551 = n25548 | n25550 ;
  assign n25552 = ( n15453 & n25549 ) | ( n15453 & n25551 ) | ( n25549 & n25551 ) ;
  assign n25553 = x29 & n25551 ;
  assign n25554 = x29 & n25549 ;
  assign n25555 = ( n15453 & n25553 ) | ( n15453 & n25554 ) | ( n25553 & n25554 ) ;
  assign n25556 = x29 & ~n25554 ;
  assign n25557 = x29 & ~n25553 ;
  assign n25558 = ( ~n15453 & n25556 ) | ( ~n15453 & n25557 ) | ( n25556 & n25557 ) ;
  assign n25559 = ( n25552 & ~n25555 ) | ( n25552 & n25558 ) | ( ~n25555 & n25558 ) ;
  assign n25560 = ~n25544 & n25559 ;
  assign n25561 = n25544 | n25560 ;
  assign n25562 = n2315 & ~n16069 ;
  assign n25563 = n2312 & ~n16085 ;
  assign n25564 = n2308 & n15886 ;
  assign n25565 = n25563 | n25564 ;
  assign n25566 = n25562 | n25565 ;
  assign n25567 = n2306 | n25566 ;
  assign n25568 = ( ~n16107 & n25566 ) | ( ~n16107 & n25567 ) | ( n25566 & n25567 ) ;
  assign n25569 = ~x26 & n25567 ;
  assign n25570 = ~x26 & n25566 ;
  assign n25571 = ( ~n16107 & n25569 ) | ( ~n16107 & n25570 ) | ( n25569 & n25570 ) ;
  assign n25572 = x26 | n25569 ;
  assign n25573 = x26 | n25570 ;
  assign n25574 = ( ~n16107 & n25572 ) | ( ~n16107 & n25573 ) | ( n25572 & n25573 ) ;
  assign n25575 = ( ~n25568 & n25571 ) | ( ~n25568 & n25574 ) | ( n25571 & n25574 ) ;
  assign n25576 = n25544 & n25559 ;
  assign n25577 = n25575 & n25576 ;
  assign n25578 = ( ~n25561 & n25575 ) | ( ~n25561 & n25577 ) | ( n25575 & n25577 ) ;
  assign n25579 = n25575 | n25576 ;
  assign n25580 = n25561 & ~n25579 ;
  assign n25581 = n25578 | n25580 ;
  assign n25582 = n25462 & ~n25581 ;
  assign n25583 = ~n25462 & n25581 ;
  assign n25584 = n25582 | n25583 ;
  assign n25585 = n2932 & ~n17092 ;
  assign n25586 = n2925 & n17111 ;
  assign n25587 = n2928 & n17100 ;
  assign n25588 = n25586 | n25587 ;
  assign n25589 = n25585 | n25588 ;
  assign n25590 = n2936 | n25585 ;
  assign n25591 = n25588 | n25590 ;
  assign n25592 = ( ~n17134 & n25589 ) | ( ~n17134 & n25591 ) | ( n25589 & n25591 ) ;
  assign n25593 = ~x23 & n25591 ;
  assign n25594 = ~x23 & n25589 ;
  assign n25595 = ( ~n17134 & n25593 ) | ( ~n17134 & n25594 ) | ( n25593 & n25594 ) ;
  assign n25596 = x23 | n25594 ;
  assign n25597 = x23 | n25593 ;
  assign n25598 = ( ~n17134 & n25596 ) | ( ~n17134 & n25597 ) | ( n25596 & n25597 ) ;
  assign n25599 = ( ~n25592 & n25595 ) | ( ~n25592 & n25598 ) | ( n25595 & n25598 ) ;
  assign n25600 = ~n25584 & n25599 ;
  assign n25601 = n25584 | n25600 ;
  assign n25603 = n24893 | n24908 ;
  assign n25604 = ( n24893 & ~n24895 ) | ( n24893 & n25603 ) | ( ~n24895 & n25603 ) ;
  assign n25602 = n25584 & n25599 ;
  assign n25605 = n25602 & n25604 ;
  assign n25606 = ( ~n25601 & n25604 ) | ( ~n25601 & n25605 ) | ( n25604 & n25605 ) ;
  assign n25607 = n25602 | n25604 ;
  assign n25608 = n25601 & ~n25607 ;
  assign n25609 = n25606 | n25608 ;
  assign n25610 = n3547 & n18410 ;
  assign n25611 = n3544 & n18037 ;
  assign n25612 = n3541 & ~n18585 ;
  assign n25613 = n25611 | n25612 ;
  assign n25614 = n25610 | n25613 ;
  assign n25615 = n3537 & ~n18586 ;
  assign n25616 = ~n18609 & n25615 ;
  assign n25617 = ( n3537 & n18650 ) | ( n3537 & n25616 ) | ( n18650 & n25616 ) ;
  assign n25618 = n25614 | n25617 ;
  assign n25619 = x20 | n25614 ;
  assign n25620 = n25617 | n25619 ;
  assign n25621 = ~x20 & n25619 ;
  assign n25622 = ( ~x20 & n25617 ) | ( ~x20 & n25621 ) | ( n25617 & n25621 ) ;
  assign n25623 = ( ~n25618 & n25620 ) | ( ~n25618 & n25622 ) | ( n25620 & n25622 ) ;
  assign n25624 = ~n25609 & n25623 ;
  assign n25625 = n25609 | n25624 ;
  assign n25627 = n24915 | n24931 ;
  assign n25628 = ( n24915 & ~n24918 ) | ( n24915 & n25627 ) | ( ~n24918 & n25627 ) ;
  assign n25626 = n25609 & n25623 ;
  assign n25629 = n25626 & n25628 ;
  assign n25630 = ( ~n25625 & n25628 ) | ( ~n25625 & n25629 ) | ( n25628 & n25629 ) ;
  assign n25631 = n25626 | n25628 ;
  assign n25632 = n25625 & ~n25631 ;
  assign n25633 = n25630 | n25632 ;
  assign n25634 = n4471 & n19494 ;
  assign n25635 = n4466 & n18576 ;
  assign n25636 = n4468 & n19352 ;
  assign n25637 = n25635 | n25636 ;
  assign n25638 = n25634 | n25637 ;
  assign n25639 = n4475 | n25634 ;
  assign n25640 = n25637 | n25639 ;
  assign n25641 = ( n20320 & n25638 ) | ( n20320 & n25640 ) | ( n25638 & n25640 ) ;
  assign n25642 = x17 & n25640 ;
  assign n25643 = x17 & n25638 ;
  assign n25644 = ( n20320 & n25642 ) | ( n20320 & n25643 ) | ( n25642 & n25643 ) ;
  assign n25645 = x17 & ~n25643 ;
  assign n25646 = x17 & ~n25642 ;
  assign n25647 = ( ~n20320 & n25645 ) | ( ~n20320 & n25646 ) | ( n25645 & n25646 ) ;
  assign n25648 = ( n25641 & ~n25644 ) | ( n25641 & n25647 ) | ( ~n25644 & n25647 ) ;
  assign n25649 = ~n25633 & n25648 ;
  assign n25650 = n25633 | n25649 ;
  assign n25652 = n24937 | n24954 ;
  assign n25653 = ( n24937 & ~n24939 ) | ( n24937 & n25652 ) | ( ~n24939 & n25652 ) ;
  assign n25651 = n25633 & n25648 ;
  assign n25654 = n25651 & n25653 ;
  assign n25655 = ( ~n25650 & n25653 ) | ( ~n25650 & n25654 ) | ( n25653 & n25654 ) ;
  assign n25656 = n25651 | n25653 ;
  assign n25657 = n25650 & ~n25656 ;
  assign n25658 = n25655 | n25657 ;
  assign n25659 = n5227 & n20680 ;
  assign n25660 = n5234 & ~n20618 ;
  assign n25661 = n5237 & n19631 ;
  assign n25662 = n5231 & ~n20630 ;
  assign n25663 = n25661 | n25662 ;
  assign n25664 = n25660 | n25663 ;
  assign n25665 = n20689 | n25664 ;
  assign n25666 = n5227 | n25664 ;
  assign n25667 = ( n25659 & n25665 ) | ( n25659 & n25666 ) | ( n25665 & n25666 ) ;
  assign n25668 = x14 | n25667 ;
  assign n25669 = ~x14 & n25667 ;
  assign n25670 = ( ~n25667 & n25668 ) | ( ~n25667 & n25669 ) | ( n25668 & n25669 ) ;
  assign n25671 = ~n25658 & n25670 ;
  assign n25672 = n25658 | n25671 ;
  assign n25673 = n25658 & n25670 ;
  assign n25674 = n25672 & ~n25673 ;
  assign n25675 = n24960 | n24977 ;
  assign n25676 = ( n24960 & ~n24962 ) | ( n24960 & n25675 ) | ( ~n24962 & n25675 ) ;
  assign n25677 = ~n25674 & n25676 ;
  assign n25678 = n25674 & ~n25676 ;
  assign n25679 = n25677 | n25678 ;
  assign n25680 = n6122 & ~n21517 ;
  assign n25681 = n6125 & n20609 ;
  assign n25682 = n6119 & ~n21563 ;
  assign n25683 = n25681 | n25682 ;
  assign n25684 = n25680 | n25683 ;
  assign n25685 = n6115 | n25680 ;
  assign n25686 = n25683 | n25685 ;
  assign n25687 = ( ~n22283 & n25684 ) | ( ~n22283 & n25686 ) | ( n25684 & n25686 ) ;
  assign n25688 = n25684 & n25686 ;
  assign n25689 = ( ~n22271 & n25687 ) | ( ~n22271 & n25688 ) | ( n25687 & n25688 ) ;
  assign n25690 = ~x11 & n25689 ;
  assign n25691 = x11 | n25689 ;
  assign n25692 = ( ~n25689 & n25690 ) | ( ~n25689 & n25691 ) | ( n25690 & n25691 ) ;
  assign n25693 = ~n25679 & n25692 ;
  assign n25694 = n25679 | n25693 ;
  assign n25695 = n25679 & n25692 ;
  assign n25696 = n25694 & ~n25695 ;
  assign n25697 = n24983 | n24999 ;
  assign n25698 = ( n24983 & ~n24985 ) | ( n24983 & n25697 ) | ( ~n24985 & n25697 ) ;
  assign n25699 = ~n25696 & n25698 ;
  assign n25700 = n25696 & ~n25698 ;
  assign n25701 = n25699 | n25700 ;
  assign n25702 = n25457 & ~n25701 ;
  assign n25703 = ~n25459 & n25702 ;
  assign n25704 = ( n25461 & ~n25701 ) | ( n25461 & n25703 ) | ( ~n25701 & n25703 ) ;
  assign n25705 = ~n25457 & n25701 ;
  assign n25706 = ( n25459 & n25701 ) | ( n25459 & n25705 ) | ( n25701 & n25705 ) ;
  assign n25707 = ~n25461 & n25706 ;
  assign n25708 = n25704 | n25707 ;
  assign n25709 = ~n24799 & n25025 ;
  assign n25710 = ( n24799 & n24801 ) | ( n24799 & ~n25709 ) | ( n24801 & ~n25709 ) ;
  assign n25711 = ~n25708 & n25710 ;
  assign n25712 = n25708 & ~n25710 ;
  assign n25713 = n25711 | n25712 ;
  assign n25714 = n25031 | n25035 ;
  assign n25715 = ~n25031 & n25033 ;
  assign n25716 = ( n24754 & n25714 ) | ( n24754 & ~n25715 ) | ( n25714 & ~n25715 ) ;
  assign n25717 = ~n25713 & n25716 ;
  assign n25718 = n25031 & ~n25713 ;
  assign n25719 = ( n25035 & ~n25713 ) | ( n25035 & n25718 ) | ( ~n25713 & n25718 ) ;
  assign n25720 = ( n24759 & n25717 ) | ( n24759 & n25719 ) | ( n25717 & n25719 ) ;
  assign n25721 = n25717 | n25719 ;
  assign n25722 = ( n24765 & n25720 ) | ( n24765 & n25721 ) | ( n25720 & n25721 ) ;
  assign n25723 = n25714 | n25716 ;
  assign n25724 = n25713 & ~n25723 ;
  assign n25725 = ( n24759 & n25714 ) | ( n24759 & n25716 ) | ( n25714 & n25716 ) ;
  assign n25726 = n25713 & ~n25725 ;
  assign n25727 = ( ~n24765 & n25724 ) | ( ~n24765 & n25726 ) | ( n25724 & n25726 ) ;
  assign n25728 = n25722 | n25727 ;
  assign n25729 = n25046 | n25728 ;
  assign n25730 = n25046 & n25728 ;
  assign n25731 = n25729 & ~n25730 ;
  assign n25732 = n25441 & n25731 ;
  assign n25733 = ( n25047 & n25066 ) | ( n25047 & ~n25732 ) | ( n25066 & ~n25732 ) ;
  assign n25734 = n2932 & ~n25728 ;
  assign n25735 = n2925 & n24770 ;
  assign n25736 = n2928 & ~n25046 ;
  assign n25737 = n25735 | n25736 ;
  assign n25738 = n25734 | n25737 ;
  assign n25739 = n25729 & n25730 ;
  assign n25740 = ~n25730 & n25739 ;
  assign n25741 = n2936 & n25740 ;
  assign n25742 = n2936 & n25731 ;
  assign n25743 = ( ~n25441 & n25741 ) | ( ~n25441 & n25742 ) | ( n25741 & n25742 ) ;
  assign n25744 = n25738 | n25743 ;
  assign n25745 = n2936 | n25738 ;
  assign n25746 = ( n25733 & n25744 ) | ( n25733 & n25745 ) | ( n25744 & n25745 ) ;
  assign n25747 = x23 | n25746 ;
  assign n25748 = ~x23 & n25746 ;
  assign n25749 = ( ~n25746 & n25747 ) | ( ~n25746 & n25748 ) | ( n25747 & n25748 ) ;
  assign n25750 = ~n25437 & n25749 ;
  assign n25751 = n25437 & ~n25749 ;
  assign n25752 = n25750 | n25751 ;
  assign n25753 = ~n25085 & n25752 ;
  assign n25754 = ~n25328 & n25753 ;
  assign n25755 = n25085 & ~n25752 ;
  assign n25756 = ( n25328 & ~n25752 ) | ( n25328 & n25755 ) | ( ~n25752 & n25755 ) ;
  assign n25757 = n25754 | n25756 ;
  assign n25758 = n25693 | n25699 ;
  assign n25759 = n25624 | n25630 ;
  assign n25760 = n25600 | n25606 ;
  assign n25761 = ( n24212 & n25478 ) | ( n24212 & n25503 ) | ( n25478 & n25503 ) ;
  assign n25762 = n1775 | n1780 ;
  assign n25763 = n391 | n6031 ;
  assign n25764 = n1776 | n6976 ;
  assign n25765 = n25763 | n25764 ;
  assign n25766 = n16775 | n25765 ;
  assign n25767 = n2630 | n5901 ;
  assign n25768 = n1467 | n1673 ;
  assign n25769 = n25767 | n25768 ;
  assign n25770 = n510 | n801 ;
  assign n25771 = n623 | n25770 ;
  assign n25772 = n1404 | n4046 ;
  assign n25773 = n1592 | n25772 ;
  assign n25774 = n25771 | n25773 ;
  assign n25775 = n25769 | n25774 ;
  assign n25776 = n25766 | n25775 ;
  assign n25777 = n25762 | n25776 ;
  assign n25778 = n104 | n134 ;
  assign n25779 = n1035 | n25778 ;
  assign n25780 = n157 | n25779 ;
  assign n25781 = n1282 | n4369 ;
  assign n25782 = n67 | n25781 ;
  assign n25783 = n25780 | n25782 ;
  assign n25784 = n160 | n247 ;
  assign n25785 = n306 | n527 ;
  assign n25786 = n25784 | n25785 ;
  assign n25787 = n437 | n25786 ;
  assign n25788 = n25783 | n25787 ;
  assign n25789 = n304 | n2051 ;
  assign n25790 = n17671 | n25789 ;
  assign n25791 = n189 | n775 ;
  assign n25792 = n250 | n501 ;
  assign n25793 = n25791 | n25792 ;
  assign n25794 = n758 | n25793 ;
  assign n25795 = n25790 | n25794 ;
  assign n25796 = n661 | n25795 ;
  assign n25797 = n25788 | n25796 ;
  assign n25798 = n12280 | n25797 ;
  assign n25799 = n274 | n442 ;
  assign n25800 = n483 | n550 ;
  assign n25801 = n25799 | n25800 ;
  assign n25802 = n163 | n886 ;
  assign n25803 = n25801 | n25802 ;
  assign n25804 = n25798 | n25803 ;
  assign n25805 = n25777 | n25804 ;
  assign n25806 = n25761 | n25805 ;
  assign n25807 = n25761 & n25805 ;
  assign n25808 = n25806 & ~n25807 ;
  assign n25809 = n1065 & n14607 ;
  assign n25810 = n1060 & n13522 ;
  assign n25811 = n25809 | n25810 ;
  assign n25812 = n1057 & n14329 ;
  assign n25813 = n1062 | n25812 ;
  assign n25814 = n25811 | n25813 ;
  assign n25815 = n25808 & n25814 ;
  assign n25816 = n25811 | n25812 ;
  assign n25817 = n25808 & n25816 ;
  assign n25818 = ( n14656 & n25815 ) | ( n14656 & n25817 ) | ( n25815 & n25817 ) ;
  assign n25819 = n25808 | n25814 ;
  assign n25820 = n25808 | n25816 ;
  assign n25821 = ( n14656 & n25819 ) | ( n14656 & n25820 ) | ( n25819 & n25820 ) ;
  assign n25822 = ~n25818 & n25821 ;
  assign n25823 = ~n25509 & n25518 ;
  assign n25824 = n25532 | n25823 ;
  assign n25825 = ( ~n25521 & n25823 ) | ( ~n25521 & n25824 ) | ( n25823 & n25824 ) ;
  assign n25826 = n25822 & n25825 ;
  assign n25827 = n25822 | n25825 ;
  assign n25828 = ~n25826 & n25827 ;
  assign n25830 = n1826 & n14591 ;
  assign n25831 = n1823 & n15434 ;
  assign n25832 = n25830 | n25831 ;
  assign n25829 = n1829 & ~n16085 ;
  assign n25834 = n1821 | n25829 ;
  assign n25835 = n25832 | n25834 ;
  assign n25833 = n25829 | n25832 ;
  assign n25836 = n25833 & n25835 ;
  assign n25837 = ( ~n16167 & n25835 ) | ( ~n16167 & n25836 ) | ( n25835 & n25836 ) ;
  assign n25838 = ~x29 & n25836 ;
  assign n25839 = ~x29 & n25835 ;
  assign n25840 = ( ~n16167 & n25838 ) | ( ~n16167 & n25839 ) | ( n25838 & n25839 ) ;
  assign n25841 = x29 | n25838 ;
  assign n25842 = x29 | n25839 ;
  assign n25843 = ( ~n16167 & n25841 ) | ( ~n16167 & n25842 ) | ( n25841 & n25842 ) ;
  assign n25844 = ( ~n25837 & n25840 ) | ( ~n25837 & n25843 ) | ( n25840 & n25843 ) ;
  assign n25845 = n25828 & n25844 ;
  assign n25846 = n25828 | n25844 ;
  assign n25847 = ~n25845 & n25846 ;
  assign n25848 = n25539 | n25559 ;
  assign n25849 = ( n25539 & ~n25544 ) | ( n25539 & n25848 ) | ( ~n25544 & n25848 ) ;
  assign n25850 = n25847 & n25849 ;
  assign n25851 = n25847 | n25849 ;
  assign n25852 = ~n25850 & n25851 ;
  assign n25853 = n2315 & n17111 ;
  assign n25854 = n2312 & n15886 ;
  assign n25855 = n2308 & ~n16069 ;
  assign n25856 = n25854 | n25855 ;
  assign n25857 = n25853 | n25856 ;
  assign n25858 = n2306 & ~n17194 ;
  assign n25859 = ~n17129 & n25858 ;
  assign n25860 = n25857 | n25859 ;
  assign n25861 = n2306 | n25857 ;
  assign n25862 = ( n17186 & n25860 ) | ( n17186 & n25861 ) | ( n25860 & n25861 ) ;
  assign n25863 = x26 | n25862 ;
  assign n25864 = ~x26 & n25862 ;
  assign n25865 = ( ~n25862 & n25863 ) | ( ~n25862 & n25864 ) | ( n25863 & n25864 ) ;
  assign n25866 = n25852 & ~n25865 ;
  assign n25867 = n25852 | n25865 ;
  assign n25868 = ( ~n25852 & n25866 ) | ( ~n25852 & n25867 ) | ( n25866 & n25867 ) ;
  assign n25869 = n25578 | n25582 ;
  assign n25870 = n25868 & n25869 ;
  assign n25871 = n25868 | n25869 ;
  assign n25872 = ~n25870 & n25871 ;
  assign n25873 = n2932 & n18037 ;
  assign n25874 = n2925 & n17100 ;
  assign n25875 = n2928 & ~n17092 ;
  assign n25876 = n25874 | n25875 ;
  assign n25877 = n25873 | n25876 ;
  assign n25878 = n2936 | n25873 ;
  assign n25879 = n25876 | n25878 ;
  assign n25880 = ( ~n18050 & n25877 ) | ( ~n18050 & n25879 ) | ( n25877 & n25879 ) ;
  assign n25881 = ~x23 & n25879 ;
  assign n25882 = ~x23 & n25877 ;
  assign n25883 = ( ~n18050 & n25881 ) | ( ~n18050 & n25882 ) | ( n25881 & n25882 ) ;
  assign n25884 = x23 | n25882 ;
  assign n25885 = x23 | n25881 ;
  assign n25886 = ( ~n18050 & n25884 ) | ( ~n18050 & n25885 ) | ( n25884 & n25885 ) ;
  assign n25887 = ( ~n25880 & n25883 ) | ( ~n25880 & n25886 ) | ( n25883 & n25886 ) ;
  assign n25888 = n25872 & ~n25887 ;
  assign n25889 = n25872 | n25887 ;
  assign n25890 = ( ~n25872 & n25888 ) | ( ~n25872 & n25889 ) | ( n25888 & n25889 ) ;
  assign n25891 = n25760 & n25890 ;
  assign n25892 = n25760 | n25890 ;
  assign n25893 = ~n25891 & n25892 ;
  assign n25894 = n3547 & n18576 ;
  assign n25895 = n3544 & ~n18585 ;
  assign n25896 = n3541 & n18410 ;
  assign n25897 = n25895 | n25896 ;
  assign n25898 = n25894 | n25897 ;
  assign n25899 = n3537 | n25894 ;
  assign n25900 = n25897 | n25899 ;
  assign n25901 = ( n18612 & n25898 ) | ( n18612 & n25900 ) | ( n25898 & n25900 ) ;
  assign n25902 = x20 & n25900 ;
  assign n25903 = x20 & n25898 ;
  assign n25904 = ( n18612 & n25902 ) | ( n18612 & n25903 ) | ( n25902 & n25903 ) ;
  assign n25905 = x20 & ~n25903 ;
  assign n25906 = x20 & ~n25902 ;
  assign n25907 = ( ~n18612 & n25905 ) | ( ~n18612 & n25906 ) | ( n25905 & n25906 ) ;
  assign n25908 = ( n25901 & ~n25904 ) | ( n25901 & n25907 ) | ( ~n25904 & n25907 ) ;
  assign n25909 = n25893 & ~n25908 ;
  assign n25910 = n25893 | n25908 ;
  assign n25911 = ( ~n25893 & n25909 ) | ( ~n25893 & n25910 ) | ( n25909 & n25910 ) ;
  assign n25912 = n25759 & n25911 ;
  assign n25913 = n25759 | n25911 ;
  assign n25914 = ~n25912 & n25913 ;
  assign n25915 = n4471 & n19631 ;
  assign n25916 = n4466 & n19352 ;
  assign n25917 = n4468 & n19494 ;
  assign n25918 = n25916 | n25917 ;
  assign n25919 = n25915 | n25918 ;
  assign n25920 = n4475 & n19652 ;
  assign n25921 = n4475 & n19655 ;
  assign n25922 = ( ~n18604 & n25920 ) | ( ~n18604 & n25921 ) | ( n25920 & n25921 ) ;
  assign n25923 = n25919 | n25922 ;
  assign n25924 = n4475 | n25919 ;
  assign n25925 = ( n19640 & n25923 ) | ( n19640 & n25924 ) | ( n25923 & n25924 ) ;
  assign n25926 = x17 | n25925 ;
  assign n25927 = ~x17 & n25925 ;
  assign n25928 = ( ~n25925 & n25926 ) | ( ~n25925 & n25927 ) | ( n25926 & n25927 ) ;
  assign n25929 = n25914 & n25928 ;
  assign n25930 = n25914 & ~n25929 ;
  assign n25931 = n25649 | n25655 ;
  assign n25932 = ~n25914 & n25928 ;
  assign n25933 = n25931 & n25932 ;
  assign n25934 = ( n25930 & n25931 ) | ( n25930 & n25933 ) | ( n25931 & n25933 ) ;
  assign n25935 = n25931 | n25932 ;
  assign n25936 = n25930 | n25935 ;
  assign n25937 = ~n25934 & n25936 ;
  assign n25938 = n5234 & n20609 ;
  assign n25939 = n5237 & ~n20630 ;
  assign n25940 = n5231 & ~n20618 ;
  assign n25941 = n25939 | n25940 ;
  assign n25942 = n25938 | n25941 ;
  assign n25943 = n5227 | n25938 ;
  assign n25944 = n25941 | n25943 ;
  assign n25945 = ( n20659 & n25942 ) | ( n20659 & n25944 ) | ( n25942 & n25944 ) ;
  assign n25946 = n25942 & n25944 ;
  assign n25947 = ( ~n20649 & n25945 ) | ( ~n20649 & n25946 ) | ( n25945 & n25946 ) ;
  assign n25948 = x14 & n25947 ;
  assign n25949 = x14 & ~n25947 ;
  assign n25950 = ( n25947 & ~n25948 ) | ( n25947 & n25949 ) | ( ~n25948 & n25949 ) ;
  assign n25951 = n25937 & n25950 ;
  assign n25952 = n25937 & ~n25951 ;
  assign n25953 = n25671 | n25677 ;
  assign n25954 = ~n25937 & n25950 ;
  assign n25955 = n25953 & n25954 ;
  assign n25956 = ( n25952 & n25953 ) | ( n25952 & n25955 ) | ( n25953 & n25955 ) ;
  assign n25957 = n25953 | n25954 ;
  assign n25958 = n25952 | n25957 ;
  assign n25959 = ~n25956 & n25958 ;
  assign n25960 = n6122 & ~n21551 ;
  assign n25961 = n6125 & ~n21563 ;
  assign n25962 = n6119 & ~n21517 ;
  assign n25963 = n25961 | n25962 ;
  assign n25964 = n25960 | n25963 ;
  assign n25965 = n6115 | n25960 ;
  assign n25966 = n25963 | n25965 ;
  assign n25967 = ( ~n21587 & n25964 ) | ( ~n21587 & n25966 ) | ( n25964 & n25966 ) ;
  assign n25968 = ~x11 & n25966 ;
  assign n25969 = ~x11 & n25964 ;
  assign n25970 = ( ~n21587 & n25968 ) | ( ~n21587 & n25969 ) | ( n25968 & n25969 ) ;
  assign n25971 = x11 | n25969 ;
  assign n25972 = x11 | n25968 ;
  assign n25973 = ( ~n21587 & n25971 ) | ( ~n21587 & n25972 ) | ( n25971 & n25972 ) ;
  assign n25974 = ( ~n25967 & n25970 ) | ( ~n25967 & n25973 ) | ( n25970 & n25973 ) ;
  assign n25975 = n25959 & ~n25974 ;
  assign n25976 = n25959 | n25974 ;
  assign n25977 = ( ~n25959 & n25975 ) | ( ~n25959 & n25976 ) | ( n25975 & n25976 ) ;
  assign n25978 = n25758 & n25977 ;
  assign n25979 = n25758 | n25977 ;
  assign n25980 = ~n25978 & n25979 ;
  assign n25981 = n7068 & ~n23240 ;
  assign n25982 = n7074 & n23227 ;
  assign n25983 = ( n7074 & n23217 ) | ( n7074 & n25982 ) | ( n23217 & n25982 ) ;
  assign n25984 = n25981 | n25983 ;
  assign n25985 = n7079 & ~n23234 ;
  assign n25986 = n7079 & ~n23235 ;
  assign n25987 = ( ~n15882 & n25985 ) | ( ~n15882 & n25986 ) | ( n25985 & n25986 ) ;
  assign n25988 = n25984 | n25987 ;
  assign n25989 = n7078 | n25987 ;
  assign n25990 = n25984 | n25989 ;
  assign n25991 = ( ~n23587 & n25988 ) | ( ~n23587 & n25990 ) | ( n25988 & n25990 ) ;
  assign n25992 = ~x8 & n25990 ;
  assign n25993 = ~x8 & n25988 ;
  assign n25994 = ( ~n23587 & n25992 ) | ( ~n23587 & n25993 ) | ( n25992 & n25993 ) ;
  assign n25995 = x8 | n25993 ;
  assign n25996 = x8 | n25992 ;
  assign n25997 = ( ~n23587 & n25995 ) | ( ~n23587 & n25996 ) | ( n25995 & n25996 ) ;
  assign n25998 = ( ~n25991 & n25994 ) | ( ~n25991 & n25997 ) | ( n25994 & n25997 ) ;
  assign n25999 = n25980 & ~n25998 ;
  assign n26000 = n25980 | n25998 ;
  assign n26001 = ( ~n25980 & n25999 ) | ( ~n25980 & n26000 ) | ( n25999 & n26000 ) ;
  assign n26002 = n25460 & n26001 ;
  assign n26003 = ( n25704 & n26001 ) | ( n25704 & n26002 ) | ( n26001 & n26002 ) ;
  assign n26004 = n25460 | n25703 ;
  assign n26005 = ~n25460 & n25701 ;
  assign n26006 = ( n25461 & n26004 ) | ( n25461 & ~n26005 ) | ( n26004 & ~n26005 ) ;
  assign n26007 = ~n26001 & n26006 ;
  assign n26008 = ( n26001 & ~n26003 ) | ( n26001 & n26007 ) | ( ~n26003 & n26007 ) ;
  assign n26009 = n25711 | n25720 ;
  assign n26010 = n26008 & n26009 ;
  assign n26011 = n25711 | n25721 ;
  assign n26012 = n26008 & n26011 ;
  assign n26013 = ( n24765 & n26010 ) | ( n24765 & n26012 ) | ( n26010 & n26012 ) ;
  assign n26014 = n26008 | n26009 ;
  assign n26015 = n26008 | n26011 ;
  assign n26016 = ( n24765 & n26014 ) | ( n24765 & n26015 ) | ( n26014 & n26015 ) ;
  assign n26017 = ~n26013 & n26016 ;
  assign n26018 = n7068 | n7079 ;
  assign n26019 = ~n23234 & n26018 ;
  assign n26020 = n7074 | n26019 ;
  assign n26021 = ~n23235 & n26018 ;
  assign n26022 = n7074 | n26021 ;
  assign n26023 = ( ~n15882 & n26020 ) | ( ~n15882 & n26022 ) | ( n26020 & n26022 ) ;
  assign n26024 = n7078 | n26023 ;
  assign n26025 = ( ~n15882 & n26019 ) | ( ~n15882 & n26021 ) | ( n26019 & n26021 ) ;
  assign n26026 = n7078 | n26025 ;
  assign n26027 = ( ~n23240 & n26024 ) | ( ~n23240 & n26026 ) | ( n26024 & n26026 ) ;
  assign n26028 = ( ~n23240 & n26023 ) | ( ~n23240 & n26025 ) | ( n26023 & n26025 ) ;
  assign n26029 = n24135 & ~n26028 ;
  assign n26030 = n23240 & ~n26028 ;
  assign n26031 = ( n23575 & n26029 ) | ( n23575 & n26030 ) | ( n26029 & n26030 ) ;
  assign n26032 = ( n23577 & n26029 ) | ( n23577 & n26030 ) | ( n26029 & n26030 ) ;
  assign n26033 = ( ~n21554 & n26031 ) | ( ~n21554 & n26032 ) | ( n26031 & n26032 ) ;
  assign n26034 = n26027 & ~n26033 ;
  assign n26035 = x8 & ~n26034 ;
  assign n26036 = n26031 | n26032 ;
  assign n26037 = n26027 & ~n26036 ;
  assign n26038 = x8 & ~n26037 ;
  assign n26039 = ( n21584 & n26035 ) | ( n21584 & n26038 ) | ( n26035 & n26038 ) ;
  assign n26040 = ~x8 & n26034 ;
  assign n26041 = ~x8 & n26037 ;
  assign n26042 = ( ~n21584 & n26040 ) | ( ~n21584 & n26041 ) | ( n26040 & n26041 ) ;
  assign n26043 = n26039 | n26042 ;
  assign n26044 = n25956 | n25974 ;
  assign n26045 = ( n25956 & n25959 ) | ( n25956 & n26044 ) | ( n25959 & n26044 ) ;
  assign n26046 = n26043 & n26045 ;
  assign n26047 = n26043 | n26045 ;
  assign n26048 = ~n26046 & n26047 ;
  assign n26049 = n25806 & ~n25817 ;
  assign n26050 = n25806 & ~n25815 ;
  assign n26051 = ( ~n14656 & n26049 ) | ( ~n14656 & n26050 ) | ( n26049 & n26050 ) ;
  assign n26052 = n3984 | n12377 ;
  assign n26053 = n413 | n648 ;
  assign n26054 = n1355 | n26053 ;
  assign n26055 = n1221 | n26054 ;
  assign n26056 = n26052 | n26055 ;
  assign n26057 = n2182 | n26056 ;
  assign n26058 = n1014 | n6910 ;
  assign n26059 = n26057 | n26058 ;
  assign n26060 = n2171 & ~n26059 ;
  assign n26061 = n796 | n5946 ;
  assign n26062 = n2108 | n26061 ;
  assign n26063 = n26060 & ~n26062 ;
  assign n26064 = n281 | n2756 ;
  assign n26065 = n2765 | n26064 ;
  assign n26066 = n2751 | n26065 ;
  assign n26067 = n588 | n26066 ;
  assign n26068 = n175 | n1172 ;
  assign n26069 = n85 | n623 ;
  assign n26070 = n26068 | n26069 ;
  assign n26071 = n280 | n26070 ;
  assign n26072 = n26067 | n26071 ;
  assign n26073 = n26063 & ~n26072 ;
  assign n26074 = n25805 | n26073 ;
  assign n26075 = n25805 & n26073 ;
  assign n26076 = n26074 & ~n26075 ;
  assign n26077 = ~n26050 & n26076 ;
  assign n26078 = ~n26049 & n26076 ;
  assign n26079 = ( n14656 & n26077 ) | ( n14656 & n26078 ) | ( n26077 & n26078 ) ;
  assign n26080 = n26051 | n26079 ;
  assign n26081 = n1057 & n14591 ;
  assign n26082 = n1060 & n14607 ;
  assign n26083 = n1065 & n14329 ;
  assign n26084 = n26082 | n26083 ;
  assign n26085 = n26081 | n26084 ;
  assign n26086 = n1062 | n26081 ;
  assign n26087 = n26084 | n26086 ;
  assign n26088 = ( n14629 & n26085 ) | ( n14629 & n26087 ) | ( n26085 & n26087 ) ;
  assign n26089 = n26050 & n26076 ;
  assign n26090 = n26049 & n26076 ;
  assign n26091 = ( ~n14656 & n26089 ) | ( ~n14656 & n26090 ) | ( n26089 & n26090 ) ;
  assign n26092 = n26088 & n26091 ;
  assign n26093 = ( ~n26080 & n26088 ) | ( ~n26080 & n26092 ) | ( n26088 & n26092 ) ;
  assign n26094 = n26088 | n26091 ;
  assign n26095 = n26080 & ~n26094 ;
  assign n26096 = n26093 | n26095 ;
  assign n26097 = n25826 | n25844 ;
  assign n26098 = ( n25826 & n25828 ) | ( n25826 & n26097 ) | ( n25828 & n26097 ) ;
  assign n26099 = ~n26096 & n26098 ;
  assign n26100 = n26096 & ~n26098 ;
  assign n26101 = n26099 | n26100 ;
  assign n26102 = n1829 & n15886 ;
  assign n26103 = n1826 & n15434 ;
  assign n26104 = n1823 & ~n16085 ;
  assign n26105 = n26103 | n26104 ;
  assign n26106 = n26102 | n26105 ;
  assign n26107 = n1821 | n26102 ;
  assign n26108 = n26105 | n26107 ;
  assign n26109 = ( ~n16140 & n26106 ) | ( ~n16140 & n26108 ) | ( n26106 & n26108 ) ;
  assign n26110 = ~x29 & n26108 ;
  assign n26111 = ~x29 & n26106 ;
  assign n26112 = ( ~n16140 & n26110 ) | ( ~n16140 & n26111 ) | ( n26110 & n26111 ) ;
  assign n26113 = x29 | n26111 ;
  assign n26114 = x29 | n26110 ;
  assign n26115 = ( ~n16140 & n26113 ) | ( ~n16140 & n26114 ) | ( n26113 & n26114 ) ;
  assign n26116 = ( ~n26109 & n26112 ) | ( ~n26109 & n26115 ) | ( n26112 & n26115 ) ;
  assign n26117 = ~n26101 & n26116 ;
  assign n26118 = n26101 | n26117 ;
  assign n26119 = n2315 & n17100 ;
  assign n26120 = n2312 & ~n16069 ;
  assign n26121 = n2308 & n17111 ;
  assign n26122 = n26120 | n26121 ;
  assign n26123 = n26119 | n26122 ;
  assign n26124 = n2306 & n17169 ;
  assign n26125 = ~n17129 & n26124 ;
  assign n26126 = n26123 | n26125 ;
  assign n26127 = n2306 | n26123 ;
  assign n26128 = ( n17161 & n26126 ) | ( n17161 & n26127 ) | ( n26126 & n26127 ) ;
  assign n26129 = x26 | n26128 ;
  assign n26130 = ~x26 & n26128 ;
  assign n26131 = ( ~n26128 & n26129 ) | ( ~n26128 & n26130 ) | ( n26129 & n26130 ) ;
  assign n26132 = n26101 & n26116 ;
  assign n26133 = n26131 & n26132 ;
  assign n26134 = ( ~n26118 & n26131 ) | ( ~n26118 & n26133 ) | ( n26131 & n26133 ) ;
  assign n26135 = n26131 | n26132 ;
  assign n26136 = n26118 & ~n26135 ;
  assign n26137 = n26134 | n26136 ;
  assign n26138 = n25850 | n25865 ;
  assign n26139 = ( n25850 & n25852 ) | ( n25850 & n26138 ) | ( n25852 & n26138 ) ;
  assign n26140 = ~n26137 & n26139 ;
  assign n26141 = n26137 & ~n26139 ;
  assign n26142 = n26140 | n26141 ;
  assign n26143 = n2932 & ~n18585 ;
  assign n26144 = n2925 & ~n17092 ;
  assign n26145 = n2928 & n18037 ;
  assign n26146 = n26144 | n26145 ;
  assign n26147 = n26143 | n26146 ;
  assign n26148 = n2936 & ~n18675 ;
  assign n26149 = ( n2936 & n18672 ) | ( n2936 & n26148 ) | ( n18672 & n26148 ) ;
  assign n26150 = n26147 | n26149 ;
  assign n26151 = x23 | n26147 ;
  assign n26152 = n26149 | n26151 ;
  assign n26153 = ~x23 & n26151 ;
  assign n26154 = ( ~x23 & n26149 ) | ( ~x23 & n26153 ) | ( n26149 & n26153 ) ;
  assign n26155 = ( ~n26150 & n26152 ) | ( ~n26150 & n26154 ) | ( n26152 & n26154 ) ;
  assign n26156 = n26142 | n26155 ;
  assign n26157 = n26142 & ~n26155 ;
  assign n26158 = ( ~n26142 & n26156 ) | ( ~n26142 & n26157 ) | ( n26156 & n26157 ) ;
  assign n26159 = n25870 | n25887 ;
  assign n26160 = ( n25870 & n25872 ) | ( n25870 & n26159 ) | ( n25872 & n26159 ) ;
  assign n26161 = ~n26158 & n26160 ;
  assign n26162 = n26158 & ~n26160 ;
  assign n26163 = n26161 | n26162 ;
  assign n26164 = n3547 & n19352 ;
  assign n26165 = n3544 & n18410 ;
  assign n26166 = n3541 & n18576 ;
  assign n26167 = n26165 | n26166 ;
  assign n26168 = n26164 | n26167 ;
  assign n26169 = n3537 | n26164 ;
  assign n26170 = n26167 | n26169 ;
  assign n26171 = ( n19674 & n26168 ) | ( n19674 & n26170 ) | ( n26168 & n26170 ) ;
  assign n26172 = x20 & n26170 ;
  assign n26173 = x20 & n26168 ;
  assign n26174 = ( n19674 & n26172 ) | ( n19674 & n26173 ) | ( n26172 & n26173 ) ;
  assign n26175 = x20 & ~n26173 ;
  assign n26176 = x20 & ~n26172 ;
  assign n26177 = ( ~n19674 & n26175 ) | ( ~n19674 & n26176 ) | ( n26175 & n26176 ) ;
  assign n26178 = ( n26171 & ~n26174 ) | ( n26171 & n26177 ) | ( ~n26174 & n26177 ) ;
  assign n26179 = n26163 | n26178 ;
  assign n26180 = n26163 & ~n26178 ;
  assign n26181 = ( ~n26163 & n26179 ) | ( ~n26163 & n26180 ) | ( n26179 & n26180 ) ;
  assign n26182 = n25891 | n25908 ;
  assign n26183 = ( n25891 & n25893 ) | ( n25891 & n26182 ) | ( n25893 & n26182 ) ;
  assign n26184 = ~n26181 & n26183 ;
  assign n26185 = n26181 & ~n26183 ;
  assign n26186 = n26184 | n26185 ;
  assign n26187 = n4471 & ~n20630 ;
  assign n26188 = n4466 & n19494 ;
  assign n26189 = n4468 & n19631 ;
  assign n26190 = n26188 | n26189 ;
  assign n26191 = n26187 | n26190 ;
  assign n26192 = n4475 | n26187 ;
  assign n26193 = n26190 | n26192 ;
  assign n26194 = ( ~n20709 & n26191 ) | ( ~n20709 & n26193 ) | ( n26191 & n26193 ) ;
  assign n26195 = ~x17 & n26193 ;
  assign n26196 = ~x17 & n26191 ;
  assign n26197 = ( ~n20709 & n26195 ) | ( ~n20709 & n26196 ) | ( n26195 & n26196 ) ;
  assign n26198 = x17 | n26196 ;
  assign n26199 = x17 | n26195 ;
  assign n26200 = ( ~n20709 & n26198 ) | ( ~n20709 & n26199 ) | ( n26198 & n26199 ) ;
  assign n26201 = ( ~n26194 & n26197 ) | ( ~n26194 & n26200 ) | ( n26197 & n26200 ) ;
  assign n26202 = n26186 | n26201 ;
  assign n26203 = n26186 & ~n26201 ;
  assign n26204 = ( ~n26186 & n26202 ) | ( ~n26186 & n26203 ) | ( n26202 & n26203 ) ;
  assign n26205 = n25912 | n25928 ;
  assign n26206 = ( n25912 & n25914 ) | ( n25912 & n26205 ) | ( n25914 & n26205 ) ;
  assign n26207 = ~n26204 & n26206 ;
  assign n26208 = n26204 & ~n26206 ;
  assign n26209 = n26207 | n26208 ;
  assign n26210 = n5234 & ~n21563 ;
  assign n26211 = n5237 & ~n20618 ;
  assign n26212 = n5231 & n20609 ;
  assign n26213 = n26211 | n26212 ;
  assign n26214 = n26210 | n26213 ;
  assign n26215 = n5227 & ~n21570 ;
  assign n26216 = n22270 & n26215 ;
  assign n26217 = ( n5227 & n22304 ) | ( n5227 & n26216 ) | ( n22304 & n26216 ) ;
  assign n26218 = n26214 | n26217 ;
  assign n26219 = x14 | n26214 ;
  assign n26220 = n26217 | n26219 ;
  assign n26221 = ~x14 & n26219 ;
  assign n26222 = ( ~x14 & n26217 ) | ( ~x14 & n26221 ) | ( n26217 & n26221 ) ;
  assign n26223 = ( ~n26218 & n26220 ) | ( ~n26218 & n26222 ) | ( n26220 & n26222 ) ;
  assign n26224 = n26209 | n26223 ;
  assign n26225 = n26209 & ~n26223 ;
  assign n26226 = ( ~n26209 & n26224 ) | ( ~n26209 & n26225 ) | ( n26224 & n26225 ) ;
  assign n26227 = n25934 | n25950 ;
  assign n26228 = ( n25934 & n25937 ) | ( n25934 & n26227 ) | ( n25937 & n26227 ) ;
  assign n26229 = ~n26226 & n26228 ;
  assign n26230 = n26226 & ~n26228 ;
  assign n26231 = n26229 | n26230 ;
  assign n26232 = n6125 & ~n21517 ;
  assign n26233 = n6119 & ~n21551 ;
  assign n26234 = n26232 | n26233 ;
  assign n26235 = n6122 & n23227 ;
  assign n26236 = ( n6122 & n23217 ) | ( n6122 & n26235 ) | ( n23217 & n26235 ) ;
  assign n26237 = n26234 | n26236 ;
  assign n26238 = n6115 & n23299 ;
  assign n26239 = n6115 & n23298 ;
  assign n26240 = ( n21584 & n26238 ) | ( n21584 & n26239 ) | ( n26238 & n26239 ) ;
  assign n26241 = n26237 | n26240 ;
  assign n26242 = n6115 | n26237 ;
  assign n26243 = ( n23289 & n26241 ) | ( n23289 & n26242 ) | ( n26241 & n26242 ) ;
  assign n26244 = x11 | n26243 ;
  assign n26245 = ~x11 & n26243 ;
  assign n26246 = ( ~n26243 & n26244 ) | ( ~n26243 & n26245 ) | ( n26244 & n26245 ) ;
  assign n26247 = n26231 | n26246 ;
  assign n26248 = n26231 & ~n26246 ;
  assign n26249 = ( ~n26231 & n26247 ) | ( ~n26231 & n26248 ) | ( n26247 & n26248 ) ;
  assign n26250 = n26048 & ~n26249 ;
  assign n26251 = n26048 & ~n26250 ;
  assign n26252 = n26048 | n26249 ;
  assign n26253 = ~n26251 & n26252 ;
  assign n26254 = n25978 | n25998 ;
  assign n26255 = ( n25978 & n25980 ) | ( n25978 & n26254 ) | ( n25980 & n26254 ) ;
  assign n26256 = ~n26253 & n26255 ;
  assign n26257 = n26253 & ~n26255 ;
  assign n26258 = n26256 | n26257 ;
  assign n26259 = n26003 | n26008 ;
  assign n26260 = ( n26003 & n26009 ) | ( n26003 & n26259 ) | ( n26009 & n26259 ) ;
  assign n26261 = ( n26003 & n26011 ) | ( n26003 & n26259 ) | ( n26011 & n26259 ) ;
  assign n26262 = ( n24765 & n26260 ) | ( n24765 & n26261 ) | ( n26260 & n26261 ) ;
  assign n26263 = n26258 & ~n26262 ;
  assign n26264 = n26002 & ~n26258 ;
  assign n26265 = n26001 & ~n26258 ;
  assign n26266 = ( n25704 & n26264 ) | ( n25704 & n26265 ) | ( n26264 & n26265 ) ;
  assign n26267 = ( n26008 & ~n26258 ) | ( n26008 & n26266 ) | ( ~n26258 & n26266 ) ;
  assign n26268 = ( n26009 & n26266 ) | ( n26009 & n26267 ) | ( n26266 & n26267 ) ;
  assign n26269 = ( n26011 & n26266 ) | ( n26011 & n26267 ) | ( n26266 & n26267 ) ;
  assign n26270 = ( n24765 & n26268 ) | ( n24765 & n26269 ) | ( n26268 & n26269 ) ;
  assign n26271 = n26263 | n26270 ;
  assign n26272 = n26017 & ~n26271 ;
  assign n26273 = n128 | n1763 ;
  assign n26274 = n2615 | n26273 ;
  assign n26275 = n5068 | n13293 ;
  assign n26276 = n26274 | n26275 ;
  assign n26277 = n1469 | n26276 ;
  assign n26278 = n468 | n15027 ;
  assign n26279 = n15025 & ~n26278 ;
  assign n26280 = ~n26277 & n26279 ;
  assign n26281 = ~n19540 & n26280 ;
  assign n26282 = n4380 | n4388 ;
  assign n26283 = n26281 & ~n26282 ;
  assign n26284 = n277 | n1114 ;
  assign n26285 = n189 | n297 ;
  assign n26286 = n160 | n202 ;
  assign n26287 = n26285 | n26286 ;
  assign n26288 = n383 | n1172 ;
  assign n26289 = n280 | n26288 ;
  assign n26290 = n26287 | n26289 ;
  assign n26291 = n445 | n2050 ;
  assign n26292 = n588 | n26291 ;
  assign n26293 = n26290 | n26292 ;
  assign n26294 = n193 | n667 ;
  assign n26295 = n616 | n26294 ;
  assign n26296 = n26293 | n26295 ;
  assign n26297 = n26284 | n26296 ;
  assign n26298 = n26283 & ~n26297 ;
  assign n26299 = n25805 & ~n26298 ;
  assign n26300 = ~n25805 & n26298 ;
  assign n26301 = n26299 | n26300 ;
  assign n26302 = n7074 | n26018 ;
  assign n26303 = n7078 | n26302 ;
  assign n26304 = ~n23229 & n26303 ;
  assign n26305 = ( n23154 & n26303 ) | ( n23154 & n26304 ) | ( n26303 & n26304 ) ;
  assign n26306 = ~n23232 & n26303 ;
  assign n26307 = ~n23231 & n26303 ;
  assign n26308 = ( n9072 & n26306 ) | ( n9072 & n26307 ) | ( n26306 & n26307 ) ;
  assign n26309 = ( ~n21543 & n26305 ) | ( ~n21543 & n26308 ) | ( n26305 & n26308 ) ;
  assign n26310 = ( ~n21545 & n26305 ) | ( ~n21545 & n26308 ) | ( n26305 & n26308 ) ;
  assign n26311 = ( ~n15882 & n26309 ) | ( ~n15882 & n26310 ) | ( n26309 & n26310 ) ;
  assign n26312 = ~x8 & n26309 ;
  assign n26313 = ~x8 & n26310 ;
  assign n26314 = ( ~n15882 & n26312 ) | ( ~n15882 & n26313 ) | ( n26312 & n26313 ) ;
  assign n26315 = x8 | n26312 ;
  assign n26316 = x8 | n26313 ;
  assign n26317 = ( ~n15882 & n26315 ) | ( ~n15882 & n26316 ) | ( n26315 & n26316 ) ;
  assign n26318 = ( ~n26311 & n26314 ) | ( ~n26311 & n26317 ) | ( n26314 & n26317 ) ;
  assign n26319 = n26301 | n26318 ;
  assign n26320 = n26301 & n26318 ;
  assign n26321 = n26319 & ~n26320 ;
  assign n26322 = ( ~n26074 & n26078 ) | ( ~n26074 & n26321 ) | ( n26078 & n26321 ) ;
  assign n26323 = ( ~n26074 & n26077 ) | ( ~n26074 & n26321 ) | ( n26077 & n26321 ) ;
  assign n26324 = ( n14656 & n26322 ) | ( n14656 & n26323 ) | ( n26322 & n26323 ) ;
  assign n26325 = n26074 & ~n26076 ;
  assign n26326 = ( n26049 & n26074 ) | ( n26049 & n26325 ) | ( n26074 & n26325 ) ;
  assign n26327 = ~n26321 & n26326 ;
  assign n26328 = ( n26050 & n26074 ) | ( n26050 & n26325 ) | ( n26074 & n26325 ) ;
  assign n26329 = ~n26321 & n26328 ;
  assign n26330 = ( ~n14656 & n26327 ) | ( ~n14656 & n26329 ) | ( n26327 & n26329 ) ;
  assign n26331 = n26324 | n26330 ;
  assign n26332 = n1057 & n15434 ;
  assign n26333 = n1060 & n14329 ;
  assign n26334 = n1065 & n14591 ;
  assign n26335 = n26333 | n26334 ;
  assign n26336 = n26332 | n26335 ;
  assign n26337 = n1062 | n26332 ;
  assign n26338 = n26335 | n26337 ;
  assign n26339 = ( n15453 & n26336 ) | ( n15453 & n26338 ) | ( n26336 & n26338 ) ;
  assign n26340 = n26331 & n26339 ;
  assign n26341 = n26331 | n26339 ;
  assign n26342 = ~n26340 & n26341 ;
  assign n26343 = n1829 & ~n16069 ;
  assign n26344 = n1826 & ~n16085 ;
  assign n26345 = n1823 & n15886 ;
  assign n26346 = n26344 | n26345 ;
  assign n26347 = n26343 | n26346 ;
  assign n26348 = n1821 | n26347 ;
  assign n26349 = ( ~n16107 & n26347 ) | ( ~n16107 & n26348 ) | ( n26347 & n26348 ) ;
  assign n26350 = ~x29 & n26348 ;
  assign n26351 = ~x29 & n26347 ;
  assign n26352 = ( ~n16107 & n26350 ) | ( ~n16107 & n26351 ) | ( n26350 & n26351 ) ;
  assign n26353 = x29 | n26350 ;
  assign n26354 = x29 | n26351 ;
  assign n26355 = ( ~n16107 & n26353 ) | ( ~n16107 & n26354 ) | ( n26353 & n26354 ) ;
  assign n26356 = ( ~n26349 & n26352 ) | ( ~n26349 & n26355 ) | ( n26352 & n26355 ) ;
  assign n26357 = ~n26342 & n26356 ;
  assign n26358 = n26342 & ~n26356 ;
  assign n26359 = n26357 | n26358 ;
  assign n26360 = ~n26093 & n26096 ;
  assign n26361 = ( n26093 & n26098 ) | ( n26093 & ~n26360 ) | ( n26098 & ~n26360 ) ;
  assign n26362 = ~n26359 & n26361 ;
  assign n26363 = n26359 & ~n26361 ;
  assign n26364 = n26362 | n26363 ;
  assign n26365 = n2315 & ~n17092 ;
  assign n26366 = n2312 & n17111 ;
  assign n26367 = n2308 & n17100 ;
  assign n26368 = n26366 | n26367 ;
  assign n26369 = n26365 | n26368 ;
  assign n26370 = n2306 | n26365 ;
  assign n26371 = n26368 | n26370 ;
  assign n26372 = ( ~n17134 & n26369 ) | ( ~n17134 & n26371 ) | ( n26369 & n26371 ) ;
  assign n26373 = ~x26 & n26371 ;
  assign n26374 = ~x26 & n26369 ;
  assign n26375 = ( ~n17134 & n26373 ) | ( ~n17134 & n26374 ) | ( n26373 & n26374 ) ;
  assign n26376 = x26 | n26374 ;
  assign n26377 = x26 | n26373 ;
  assign n26378 = ( ~n17134 & n26376 ) | ( ~n17134 & n26377 ) | ( n26376 & n26377 ) ;
  assign n26379 = ( ~n26372 & n26375 ) | ( ~n26372 & n26378 ) | ( n26375 & n26378 ) ;
  assign n26380 = ~n26364 & n26379 ;
  assign n26381 = n26364 | n26380 ;
  assign n26382 = n26364 & n26379 ;
  assign n26383 = n26381 & ~n26382 ;
  assign n26384 = n26117 | n26134 ;
  assign n26385 = ~n26383 & n26384 ;
  assign n26386 = n26383 & ~n26384 ;
  assign n26387 = n26385 | n26386 ;
  assign n26388 = n2932 & n18410 ;
  assign n26389 = n2925 & n18037 ;
  assign n26390 = n2928 & ~n18585 ;
  assign n26391 = n26389 | n26390 ;
  assign n26392 = n26388 | n26391 ;
  assign n26393 = n2936 & ~n18586 ;
  assign n26394 = ~n18609 & n26393 ;
  assign n26395 = ( n2936 & n18650 ) | ( n2936 & n26394 ) | ( n18650 & n26394 ) ;
  assign n26396 = n26392 | n26395 ;
  assign n26397 = x23 | n26392 ;
  assign n26398 = n26395 | n26397 ;
  assign n26399 = ~x23 & n26397 ;
  assign n26400 = ( ~x23 & n26395 ) | ( ~x23 & n26399 ) | ( n26395 & n26399 ) ;
  assign n26401 = ( ~n26396 & n26398 ) | ( ~n26396 & n26400 ) | ( n26398 & n26400 ) ;
  assign n26402 = ~n26387 & n26401 ;
  assign n26403 = n26387 | n26402 ;
  assign n26405 = n26140 | n26155 ;
  assign n26406 = ( n26140 & ~n26142 ) | ( n26140 & n26405 ) | ( ~n26142 & n26405 ) ;
  assign n26404 = n26387 & n26401 ;
  assign n26407 = n26404 & n26406 ;
  assign n26408 = ( ~n26403 & n26406 ) | ( ~n26403 & n26407 ) | ( n26406 & n26407 ) ;
  assign n26409 = n26403 & ~n26404 ;
  assign n26410 = ~n26406 & n26409 ;
  assign n26411 = n26408 | n26410 ;
  assign n26412 = n3547 & n19494 ;
  assign n26413 = n3544 & n18576 ;
  assign n26414 = n3541 & n19352 ;
  assign n26415 = n26413 | n26414 ;
  assign n26416 = n26412 | n26415 ;
  assign n26417 = n3537 | n26412 ;
  assign n26418 = n26415 | n26417 ;
  assign n26419 = ( n20320 & n26416 ) | ( n20320 & n26418 ) | ( n26416 & n26418 ) ;
  assign n26420 = x20 & n26418 ;
  assign n26421 = x20 & n26416 ;
  assign n26422 = ( n20320 & n26420 ) | ( n20320 & n26421 ) | ( n26420 & n26421 ) ;
  assign n26423 = x20 & ~n26421 ;
  assign n26424 = x20 & ~n26420 ;
  assign n26425 = ( ~n20320 & n26423 ) | ( ~n20320 & n26424 ) | ( n26423 & n26424 ) ;
  assign n26426 = ( n26419 & ~n26422 ) | ( n26419 & n26425 ) | ( ~n26422 & n26425 ) ;
  assign n26427 = ~n26410 & n26426 ;
  assign n26428 = ~n26408 & n26427 ;
  assign n26429 = n26411 | n26428 ;
  assign n26430 = n26410 & n26426 ;
  assign n26431 = ( n26408 & n26426 ) | ( n26408 & n26430 ) | ( n26426 & n26430 ) ;
  assign n26432 = n26429 & ~n26431 ;
  assign n26433 = n26161 | n26178 ;
  assign n26434 = ( n26161 & ~n26163 ) | ( n26161 & n26433 ) | ( ~n26163 & n26433 ) ;
  assign n26435 = ~n26432 & n26434 ;
  assign n26436 = n26432 & ~n26434 ;
  assign n26437 = n26435 | n26436 ;
  assign n26438 = n4475 & n20680 ;
  assign n26439 = n4471 & ~n20618 ;
  assign n26440 = n4466 & n19631 ;
  assign n26441 = n4468 & ~n20630 ;
  assign n26442 = n26440 | n26441 ;
  assign n26443 = n26439 | n26442 ;
  assign n26444 = n20689 | n26443 ;
  assign n26445 = n4475 | n26443 ;
  assign n26446 = ( n26438 & n26444 ) | ( n26438 & n26445 ) | ( n26444 & n26445 ) ;
  assign n26447 = x17 | n26446 ;
  assign n26448 = ~x17 & n26446 ;
  assign n26449 = ( ~n26446 & n26447 ) | ( ~n26446 & n26448 ) | ( n26447 & n26448 ) ;
  assign n26450 = ~n26437 & n26449 ;
  assign n26451 = n26437 | n26450 ;
  assign n26452 = n26437 & n26449 ;
  assign n26453 = n26451 & ~n26452 ;
  assign n26454 = n26184 | n26201 ;
  assign n26455 = ( n26184 & ~n26186 ) | ( n26184 & n26454 ) | ( ~n26186 & n26454 ) ;
  assign n26456 = ~n26453 & n26455 ;
  assign n26457 = n26453 & ~n26455 ;
  assign n26458 = n26456 | n26457 ;
  assign n26459 = n5234 & ~n21517 ;
  assign n26460 = n5237 & n20609 ;
  assign n26461 = n5231 & ~n21563 ;
  assign n26462 = n26460 | n26461 ;
  assign n26463 = n26459 | n26462 ;
  assign n26464 = n5227 | n26459 ;
  assign n26465 = n26462 | n26464 ;
  assign n26466 = ( ~n22283 & n26463 ) | ( ~n22283 & n26465 ) | ( n26463 & n26465 ) ;
  assign n26467 = n26463 & n26465 ;
  assign n26468 = ( ~n22271 & n26466 ) | ( ~n22271 & n26467 ) | ( n26466 & n26467 ) ;
  assign n26469 = ~x14 & n26468 ;
  assign n26470 = x14 | n26468 ;
  assign n26471 = ( ~n26468 & n26469 ) | ( ~n26468 & n26470 ) | ( n26469 & n26470 ) ;
  assign n26472 = ~n26458 & n26471 ;
  assign n26473 = n26458 | n26472 ;
  assign n26474 = n26207 | n26223 ;
  assign n26475 = ( n26207 & ~n26209 ) | ( n26207 & n26474 ) | ( ~n26209 & n26474 ) ;
  assign n26476 = n26458 & n26471 ;
  assign n26477 = n26475 & n26476 ;
  assign n26478 = ( ~n26473 & n26475 ) | ( ~n26473 & n26477 ) | ( n26475 & n26477 ) ;
  assign n26479 = n26475 | n26476 ;
  assign n26480 = n26473 & ~n26479 ;
  assign n26481 = n26478 | n26480 ;
  assign n26498 = n26229 | n26246 ;
  assign n26499 = ( n26229 & ~n26231 ) | ( n26229 & n26498 ) | ( ~n26231 & n26498 ) ;
  assign n26482 = n6122 & ~n23240 ;
  assign n26483 = n6125 & ~n21551 ;
  assign n26484 = n6119 & n23227 ;
  assign n26485 = ( n6119 & n23217 ) | ( n6119 & n26484 ) | ( n23217 & n26484 ) ;
  assign n26486 = n26483 | n26485 ;
  assign n26487 = n26482 | n26486 ;
  assign n26488 = n6115 | n26482 ;
  assign n26489 = n26486 | n26488 ;
  assign n26490 = ( n23260 & n26487 ) | ( n23260 & n26489 ) | ( n26487 & n26489 ) ;
  assign n26491 = x11 & n26489 ;
  assign n26492 = x11 & n26487 ;
  assign n26493 = ( n23260 & n26491 ) | ( n23260 & n26492 ) | ( n26491 & n26492 ) ;
  assign n26494 = x11 & ~n26492 ;
  assign n26495 = x11 & ~n26491 ;
  assign n26496 = ( ~n23260 & n26494 ) | ( ~n23260 & n26495 ) | ( n26494 & n26495 ) ;
  assign n26497 = ( n26490 & ~n26493 ) | ( n26490 & n26496 ) | ( ~n26493 & n26496 ) ;
  assign n26500 = n26497 & n26499 ;
  assign n26501 = n26499 & ~n26500 ;
  assign n26502 = ~n26481 & n26497 ;
  assign n26503 = ~n26499 & n26502 ;
  assign n26504 = ( ~n26481 & n26501 ) | ( ~n26481 & n26503 ) | ( n26501 & n26503 ) ;
  assign n26505 = n26481 & ~n26497 ;
  assign n26506 = ( n26481 & n26499 ) | ( n26481 & n26505 ) | ( n26499 & n26505 ) ;
  assign n26507 = ~n26501 & n26506 ;
  assign n26508 = n26504 | n26507 ;
  assign n26509 = ~n26046 & n26249 ;
  assign n26510 = ( n26046 & n26048 ) | ( n26046 & ~n26509 ) | ( n26048 & ~n26509 ) ;
  assign n26511 = ~n26508 & n26510 ;
  assign n26512 = n26508 & ~n26510 ;
  assign n26513 = n26511 | n26512 ;
  assign n26514 = n26256 | n26266 ;
  assign n26515 = ~n26256 & n26258 ;
  assign n26516 = ( n26008 & n26514 ) | ( n26008 & ~n26515 ) | ( n26514 & ~n26515 ) ;
  assign n26517 = ( n26009 & n26514 ) | ( n26009 & n26516 ) | ( n26514 & n26516 ) ;
  assign n26518 = ( n26011 & n26514 ) | ( n26011 & n26516 ) | ( n26514 & n26516 ) ;
  assign n26519 = ( n24765 & n26517 ) | ( n24765 & n26518 ) | ( n26517 & n26518 ) ;
  assign n26520 = n26513 & ~n26519 ;
  assign n26521 = ~n26513 & n26516 ;
  assign n26522 = n26256 & ~n26513 ;
  assign n26523 = ( n26266 & ~n26513 ) | ( n26266 & n26522 ) | ( ~n26513 & n26522 ) ;
  assign n26524 = ( n26009 & n26521 ) | ( n26009 & n26523 ) | ( n26521 & n26523 ) ;
  assign n26525 = ( n26011 & n26521 ) | ( n26011 & n26523 ) | ( n26521 & n26523 ) ;
  assign n26526 = ( n24765 & n26524 ) | ( n24765 & n26525 ) | ( n26524 & n26525 ) ;
  assign n26527 = n26520 | n26526 ;
  assign n26528 = n26271 | n26527 ;
  assign n26529 = n26271 & n26527 ;
  assign n26530 = n26272 & ~n26529 ;
  assign n26531 = ( n25728 & n25739 ) | ( n25728 & ~n26017 ) | ( n25739 & ~n26017 ) ;
  assign n26532 = ~n26017 & n26271 ;
  assign n26533 = n26272 | n26532 ;
  assign n26534 = ( n26529 & ~n26530 ) | ( n26529 & n26533 ) | ( ~n26530 & n26533 ) ;
  assign n26535 = ( ~n26530 & n26531 ) | ( ~n26530 & n26534 ) | ( n26531 & n26534 ) ;
  assign n26536 = ( n25728 & n25729 ) | ( n25728 & ~n26017 ) | ( n25729 & ~n26017 ) ;
  assign n26537 = ( ~n26530 & n26534 ) | ( ~n26530 & n26536 ) | ( n26534 & n26536 ) ;
  assign n26538 = ( ~n25441 & n26535 ) | ( ~n25441 & n26537 ) | ( n26535 & n26537 ) ;
  assign n26539 = n26528 & ~n26538 ;
  assign n26540 = n26531 | n26533 ;
  assign n26541 = n26533 | n26536 ;
  assign n26542 = ( ~n25441 & n26540 ) | ( ~n25441 & n26541 ) | ( n26540 & n26541 ) ;
  assign n26543 = ( ~n26272 & n26539 ) | ( ~n26272 & n26542 ) | ( n26539 & n26542 ) ;
  assign n26544 = n3544 & n26017 ;
  assign n26545 = n3541 & ~n26270 ;
  assign n26546 = ~n26263 & n26545 ;
  assign n26547 = n26544 | n26546 ;
  assign n26548 = n3547 & ~n26526 ;
  assign n26549 = ~n26520 & n26548 ;
  assign n26551 = n3537 | n26549 ;
  assign n26552 = n26547 | n26551 ;
  assign n26550 = n26547 | n26549 ;
  assign n26553 = n26550 & n26552 ;
  assign n26554 = ( n26271 & n26527 ) | ( n26271 & n26528 ) | ( n26527 & n26528 ) ;
  assign n26555 = ( n26529 & ~n26538 ) | ( n26529 & n26554 ) | ( ~n26538 & n26554 ) ;
  assign n26556 = ( n26552 & n26553 ) | ( n26552 & ~n26555 ) | ( n26553 & ~n26555 ) ;
  assign n26557 = ( n26528 & n26552 ) | ( n26528 & n26553 ) | ( n26552 & n26553 ) ;
  assign n26558 = ( ~n26543 & n26556 ) | ( ~n26543 & n26557 ) | ( n26556 & n26557 ) ;
  assign n26559 = ~x20 & n26558 ;
  assign n26560 = x20 | n26558 ;
  assign n26561 = ( ~n26558 & n26559 ) | ( ~n26558 & n26560 ) | ( n26559 & n26560 ) ;
  assign n26562 = ~n25757 & n26561 ;
  assign n26563 = n25757 | n26562 ;
  assign n26564 = n25757 & n26561 ;
  assign n26565 = n26563 & ~n26564 ;
  assign n26566 = n25088 | n25327 ;
  assign n26567 = ~n25328 & n26566 ;
  assign n26568 = n26531 & n26533 ;
  assign n26569 = n26533 & n26536 ;
  assign n26570 = ( ~n25441 & n26568 ) | ( ~n25441 & n26569 ) | ( n26568 & n26569 ) ;
  assign n26571 = n26542 & ~n26570 ;
  assign n26572 = n3544 & ~n25728 ;
  assign n26573 = n3541 & n26017 ;
  assign n26574 = n26572 | n26573 ;
  assign n26575 = n3547 & ~n26270 ;
  assign n26576 = ~n26263 & n26575 ;
  assign n26578 = n3537 | n26576 ;
  assign n26579 = n26574 | n26578 ;
  assign n26577 = n26574 | n26576 ;
  assign n26580 = n26577 & n26579 ;
  assign n26581 = ( n26571 & n26579 ) | ( n26571 & n26580 ) | ( n26579 & n26580 ) ;
  assign n26582 = x20 & n26580 ;
  assign n26583 = x20 & n26579 ;
  assign n26584 = ( n26571 & n26582 ) | ( n26571 & n26583 ) | ( n26582 & n26583 ) ;
  assign n26585 = x20 & ~n26582 ;
  assign n26586 = x20 & ~n26583 ;
  assign n26587 = ( ~n26571 & n26585 ) | ( ~n26571 & n26586 ) | ( n26585 & n26586 ) ;
  assign n26588 = ( n26581 & ~n26584 ) | ( n26581 & n26587 ) | ( ~n26584 & n26587 ) ;
  assign n26589 = n26567 & n26588 ;
  assign n26590 = n26567 & ~n26589 ;
  assign n26591 = ~n26567 & n26588 ;
  assign n26592 = n26590 | n26591 ;
  assign n26593 = n25323 | n25324 ;
  assign n26594 = n25111 & ~n26593 ;
  assign n26595 = n25326 | n26594 ;
  assign n26596 = ( ~n25441 & n25729 ) | ( ~n25441 & n25739 ) | ( n25729 & n25739 ) ;
  assign n26597 = ~n25728 & n26017 ;
  assign n26598 = n25728 & ~n26017 ;
  assign n26599 = n25729 | n26598 ;
  assign n26600 = n26597 | n26599 ;
  assign n26601 = n26597 | n26598 ;
  assign n26602 = ( n25730 & n26600 ) | ( n25730 & n26601 ) | ( n26600 & n26601 ) ;
  assign n26603 = n26600 | n26601 ;
  assign n26604 = ( ~n25441 & n26602 ) | ( ~n25441 & n26603 ) | ( n26602 & n26603 ) ;
  assign n26605 = ~n26596 & n26604 ;
  assign n26606 = n3547 & n26017 ;
  assign n26607 = n3544 & ~n25046 ;
  assign n26608 = n3541 & ~n25728 ;
  assign n26609 = n26607 | n26608 ;
  assign n26610 = n26606 | n26609 ;
  assign n26611 = n26531 & ~n26598 ;
  assign n26612 = n26536 & ~n26598 ;
  assign n26613 = ( ~n25441 & n26611 ) | ( ~n25441 & n26612 ) | ( n26611 & n26612 ) ;
  assign n26614 = n3537 | n26606 ;
  assign n26615 = n26609 | n26614 ;
  assign n26616 = ( n26610 & n26613 ) | ( n26610 & n26615 ) | ( n26613 & n26615 ) ;
  assign n26617 = n26610 | n26615 ;
  assign n26618 = ( n26605 & n26616 ) | ( n26605 & n26617 ) | ( n26616 & n26617 ) ;
  assign n26619 = x20 & n26618 ;
  assign n26620 = x20 & ~n26618 ;
  assign n26621 = ( n26618 & ~n26619 ) | ( n26618 & n26620 ) | ( ~n26619 & n26620 ) ;
  assign n26622 = ~n26595 & n26621 ;
  assign n26623 = n26595 | n26622 ;
  assign n26624 = n26595 & n26621 ;
  assign n26625 = n26623 & ~n26624 ;
  assign n26626 = n25135 & ~n25321 ;
  assign n26627 = n25322 | n26626 ;
  assign n26628 = n3544 & n24770 ;
  assign n26629 = n3541 & ~n25046 ;
  assign n26630 = n26628 | n26629 ;
  assign n26631 = n3547 & ~n25728 ;
  assign n26632 = n3537 | n26631 ;
  assign n26633 = n26630 | n26632 ;
  assign n26634 = n26630 | n26631 ;
  assign n26635 = n25740 | n26634 ;
  assign n26636 = n25731 | n26634 ;
  assign n26637 = ( ~n25441 & n26635 ) | ( ~n25441 & n26636 ) | ( n26635 & n26636 ) ;
  assign n26638 = n26633 & n26637 ;
  assign n26639 = ( n25733 & n26633 ) | ( n25733 & n26638 ) | ( n26633 & n26638 ) ;
  assign n26640 = ~x20 & n26639 ;
  assign n26641 = x20 | n26639 ;
  assign n26642 = ( ~n26639 & n26640 ) | ( ~n26639 & n26641 ) | ( n26640 & n26641 ) ;
  assign n26643 = ~n26627 & n26642 ;
  assign n26644 = n26627 | n26643 ;
  assign n26645 = n26627 & n26642 ;
  assign n26646 = n26644 & ~n26645 ;
  assign n26647 = n25317 & n25319 ;
  assign n26648 = n25317 | n25319 ;
  assign n26649 = ~n26647 & n26648 ;
  assign n26650 = n3547 & ~n25046 ;
  assign n26651 = n3544 & ~n25054 ;
  assign n26652 = n3541 & n24770 ;
  assign n26653 = n26651 | n26652 ;
  assign n26654 = n26650 | n26653 ;
  assign n26655 = n3537 | n26650 ;
  assign n26656 = n26653 | n26655 ;
  assign n26657 = ( ~n25069 & n26654 ) | ( ~n25069 & n26656 ) | ( n26654 & n26656 ) ;
  assign n26658 = ~x20 & n26656 ;
  assign n26659 = ~x20 & n26654 ;
  assign n26660 = ( ~n25069 & n26658 ) | ( ~n25069 & n26659 ) | ( n26658 & n26659 ) ;
  assign n26661 = x20 | n26659 ;
  assign n26662 = x20 | n26658 ;
  assign n26663 = ( ~n25069 & n26661 ) | ( ~n25069 & n26662 ) | ( n26661 & n26662 ) ;
  assign n26664 = ( ~n26657 & n26660 ) | ( ~n26657 & n26663 ) | ( n26660 & n26663 ) ;
  assign n26665 = n26649 & n26664 ;
  assign n26666 = n25315 & ~n25316 ;
  assign n26667 = n25172 & ~n25316 ;
  assign n26668 = n26666 | n26667 ;
  assign n26669 = n3547 & n24770 ;
  assign n26670 = n3544 & n24167 ;
  assign n26671 = n3541 & ~n25054 ;
  assign n26672 = n26670 | n26671 ;
  assign n26673 = n26669 | n26672 ;
  assign n26674 = n3537 | n26673 ;
  assign n26675 = ( ~n25095 & n26673 ) | ( ~n25095 & n26674 ) | ( n26673 & n26674 ) ;
  assign n26676 = ~x20 & n26674 ;
  assign n26677 = ~x20 & n26673 ;
  assign n26678 = ( ~n25095 & n26676 ) | ( ~n25095 & n26677 ) | ( n26676 & n26677 ) ;
  assign n26679 = x20 | n26676 ;
  assign n26680 = x20 | n26677 ;
  assign n26681 = ( ~n25095 & n26679 ) | ( ~n25095 & n26680 ) | ( n26679 & n26680 ) ;
  assign n26682 = ( ~n26675 & n26678 ) | ( ~n26675 & n26681 ) | ( n26678 & n26681 ) ;
  assign n26683 = n26668 & n26682 ;
  assign n26684 = n26668 & ~n26683 ;
  assign n26685 = ~n26668 & n26682 ;
  assign n26686 = n26684 | n26685 ;
  assign n26687 = n25194 | n25288 ;
  assign n26688 = ~n25289 & n26687 ;
  assign n26689 = n3547 & n24167 ;
  assign n26690 = n3544 & n23316 ;
  assign n26691 = n3541 & n23614 ;
  assign n26692 = n26690 | n26691 ;
  assign n26693 = n26689 | n26692 ;
  assign n26694 = n3537 | n26693 ;
  assign n26695 = ( n24182 & n26693 ) | ( n24182 & n26694 ) | ( n26693 & n26694 ) ;
  assign n26696 = n26693 | n26694 ;
  assign n26697 = ( n24175 & n26695 ) | ( n24175 & n26696 ) | ( n26695 & n26696 ) ;
  assign n26698 = x20 & n26697 ;
  assign n26699 = x20 & ~n26697 ;
  assign n26700 = ( n26697 & ~n26698 ) | ( n26697 & n26699 ) | ( ~n26698 & n26699 ) ;
  assign n26701 = n26688 & n26700 ;
  assign n26702 = n25290 & n25313 ;
  assign n26703 = n25290 | n25313 ;
  assign n26704 = ~n26702 & n26703 ;
  assign n26705 = n3547 & ~n25054 ;
  assign n26706 = n3544 & n23614 ;
  assign n26707 = n3541 & n24167 ;
  assign n26708 = n26706 | n26707 ;
  assign n26709 = n26705 | n26708 ;
  assign n26710 = n3537 | n26705 ;
  assign n26711 = n26708 | n26710 ;
  assign n26712 = ( ~n25122 & n26709 ) | ( ~n25122 & n26711 ) | ( n26709 & n26711 ) ;
  assign n26713 = ~x20 & n26711 ;
  assign n26714 = ~x20 & n26709 ;
  assign n26715 = ( ~n25122 & n26713 ) | ( ~n25122 & n26714 ) | ( n26713 & n26714 ) ;
  assign n26716 = x20 | n26714 ;
  assign n26717 = x20 | n26713 ;
  assign n26718 = ( ~n25122 & n26716 ) | ( ~n25122 & n26717 ) | ( n26716 & n26717 ) ;
  assign n26719 = ( ~n26712 & n26715 ) | ( ~n26712 & n26718 ) | ( n26715 & n26718 ) ;
  assign n26720 = n26704 & n26719 ;
  assign n26721 = n26704 | n26719 ;
  assign n26722 = ~n26720 & n26721 ;
  assign n26723 = n26701 & n26722 ;
  assign n26724 = n26720 | n26722 ;
  assign n26725 = n25213 | n25286 ;
  assign n26726 = ~n25287 & n26725 ;
  assign n26727 = n3547 & n23614 ;
  assign n26728 = n3544 & n23620 ;
  assign n26729 = ( n3541 & n10490 ) | ( n3541 & n23620 ) | ( n10490 & n23620 ) ;
  assign n26730 = ( n23316 & n26728 ) | ( n23316 & n26729 ) | ( n26728 & n26729 ) ;
  assign n26732 = n3537 | n26730 ;
  assign n26733 = n26727 | n26732 ;
  assign n26731 = n26727 | n26730 ;
  assign n26734 = n26731 & n26733 ;
  assign n26735 = ( n23634 & n26733 ) | ( n23634 & n26734 ) | ( n26733 & n26734 ) ;
  assign n26736 = x20 & n26734 ;
  assign n26737 = x20 & n26733 ;
  assign n26738 = ( n23634 & n26736 ) | ( n23634 & n26737 ) | ( n26736 & n26737 ) ;
  assign n26739 = x20 & ~n26736 ;
  assign n26740 = x20 & ~n26737 ;
  assign n26741 = ( ~n23634 & n26739 ) | ( ~n23634 & n26740 ) | ( n26739 & n26740 ) ;
  assign n26742 = ( n26735 & ~n26738 ) | ( n26735 & n26741 ) | ( ~n26738 & n26741 ) ;
  assign n26743 = n26726 & n26742 ;
  assign n26744 = n26726 & ~n26743 ;
  assign n26745 = ~n26726 & n26742 ;
  assign n26746 = n26744 | n26745 ;
  assign n26747 = n25266 & n25280 ;
  assign n26748 = n25266 & ~n26747 ;
  assign n26749 = n3544 & ~n22385 ;
  assign n26750 = ( n3541 & n10490 ) | ( n3541 & ~n22385 ) | ( n10490 & ~n22385 ) ;
  assign n26751 = ( n22381 & n26749 ) | ( n22381 & n26750 ) | ( n26749 & n26750 ) ;
  assign n26752 = n3547 | n26751 ;
  assign n26753 = ( n23620 & n26751 ) | ( n23620 & n26752 ) | ( n26751 & n26752 ) ;
  assign n26754 = n3537 | n26753 ;
  assign n26755 = ( ~n23686 & n26753 ) | ( ~n23686 & n26754 ) | ( n26753 & n26754 ) ;
  assign n26756 = ~x20 & n26754 ;
  assign n26757 = ~x20 & n26753 ;
  assign n26758 = ( ~n23686 & n26756 ) | ( ~n23686 & n26757 ) | ( n26756 & n26757 ) ;
  assign n26759 = x20 | n26756 ;
  assign n26760 = x20 | n26757 ;
  assign n26761 = ( ~n23686 & n26759 ) | ( ~n23686 & n26760 ) | ( n26759 & n26760 ) ;
  assign n26762 = ( ~n26755 & n26758 ) | ( ~n26755 & n26761 ) | ( n26758 & n26761 ) ;
  assign n26763 = ~n25266 & n25280 ;
  assign n26764 = n26762 & n26763 ;
  assign n26765 = ( n26748 & n26762 ) | ( n26748 & n26764 ) | ( n26762 & n26764 ) ;
  assign n26766 = n26762 | n26763 ;
  assign n26767 = n26748 | n26766 ;
  assign n26768 = ~n26765 & n26767 ;
  assign n26769 = n25245 & n25263 ;
  assign n26770 = n25245 | n25263 ;
  assign n26771 = ~n26769 & n26770 ;
  assign n26772 = n3547 & n22381 ;
  assign n26773 = n3544 & ~n22398 ;
  assign n26774 = n3541 & ~n22385 ;
  assign n26775 = n26773 | n26774 ;
  assign n26776 = n26772 | n26775 ;
  assign n26777 = n3537 | n26776 ;
  assign n26778 = x20 & n26777 ;
  assign n26779 = x20 & n26776 ;
  assign n26780 = ( n22422 & n26778 ) | ( n22422 & n26779 ) | ( n26778 & n26779 ) ;
  assign n26781 = x20 | n26777 ;
  assign n26782 = x20 | n26776 ;
  assign n26783 = ( n22422 & n26781 ) | ( n22422 & n26782 ) | ( n26781 & n26782 ) ;
  assign n26784 = ~n26780 & n26783 ;
  assign n26785 = n26771 & n26784 ;
  assign n26786 = ~n26771 & n26784 ;
  assign n26787 = ( n26771 & ~n26785 ) | ( n26771 & n26786 ) | ( ~n26785 & n26786 ) ;
  assign n26788 = n25239 | n25241 ;
  assign n26789 = ~n25241 & n25243 ;
  assign n26790 = ( n25240 & n26788 ) | ( n25240 & ~n26789 ) | ( n26788 & ~n26789 ) ;
  assign n26791 = ~n25245 & n26790 ;
  assign n26792 = n3547 & ~n22385 ;
  assign n26793 = n3544 & n22393 ;
  assign n26794 = n3541 & ~n22398 ;
  assign n26795 = n26793 | n26794 ;
  assign n26796 = n26792 | n26795 ;
  assign n26797 = n3537 | n26792 ;
  assign n26798 = n26795 | n26797 ;
  assign n26799 = ( ~n22545 & n26796 ) | ( ~n22545 & n26798 ) | ( n26796 & n26798 ) ;
  assign n26800 = ~x20 & n26798 ;
  assign n26801 = ~x20 & n26796 ;
  assign n26802 = ( ~n22545 & n26800 ) | ( ~n22545 & n26801 ) | ( n26800 & n26801 ) ;
  assign n26803 = x20 | n26801 ;
  assign n26804 = x20 | n26800 ;
  assign n26805 = ( ~n22545 & n26803 ) | ( ~n22545 & n26804 ) | ( n26803 & n26804 ) ;
  assign n26806 = ( ~n26799 & n26802 ) | ( ~n26799 & n26805 ) | ( n26802 & n26805 ) ;
  assign n26807 = n26791 & n26806 ;
  assign n26808 = n3537 & n22474 ;
  assign n26809 = n3541 & ~n22409 ;
  assign n26810 = n3547 & ~n22406 ;
  assign n26811 = n26809 | n26810 ;
  assign n26812 = x20 | n26811 ;
  assign n26813 = n26808 | n26812 ;
  assign n26814 = ~x20 & n26813 ;
  assign n26815 = ( x20 & n14923 ) | ( x20 & n22409 ) | ( n14923 & n22409 ) ;
  assign n26816 = n26813 & n26815 ;
  assign n26817 = n26808 | n26811 ;
  assign n26818 = n26815 & ~n26817 ;
  assign n26819 = ( n26814 & n26816 ) | ( n26814 & n26818 ) | ( n26816 & n26818 ) ;
  assign n26820 = n3547 & n22393 ;
  assign n26821 = n3544 & ~n22409 ;
  assign n26822 = n3541 & ~n22406 ;
  assign n26823 = n26821 | n26822 ;
  assign n26824 = n26820 | n26823 ;
  assign n26825 = n22439 | n26824 ;
  assign n26826 = n3537 | n26820 ;
  assign n26827 = n26823 | n26826 ;
  assign n26828 = ~x20 & n26827 ;
  assign n26829 = n26825 & n26828 ;
  assign n26830 = x20 | n26829 ;
  assign n26831 = n2920 & ~n22409 ;
  assign n26832 = n26829 & n26831 ;
  assign n26833 = n26825 & n26827 ;
  assign n26834 = n26831 & ~n26833 ;
  assign n26835 = ( n26830 & n26832 ) | ( n26830 & n26834 ) | ( n26832 & n26834 ) ;
  assign n26836 = n26819 & n26835 ;
  assign n26837 = ( n26829 & n26830 ) | ( n26829 & ~n26833 ) | ( n26830 & ~n26833 ) ;
  assign n26838 = n26819 | n26831 ;
  assign n26839 = ( n26831 & n26837 ) | ( n26831 & n26838 ) | ( n26837 & n26838 ) ;
  assign n26840 = ~n26836 & n26839 ;
  assign n26841 = n3544 & ~n22406 ;
  assign n26842 = n3541 & n22393 ;
  assign n26843 = n26841 | n26842 ;
  assign n26844 = n3547 & ~n22398 ;
  assign n26845 = n3537 | n26844 ;
  assign n26846 = n26843 | n26845 ;
  assign n26847 = x20 & n26846 ;
  assign n26848 = n26843 | n26844 ;
  assign n26849 = x20 & n26848 ;
  assign n26850 = ( n22608 & n26847 ) | ( n22608 & n26849 ) | ( n26847 & n26849 ) ;
  assign n26851 = x20 | n26846 ;
  assign n26852 = x20 | n26848 ;
  assign n26853 = ( n22608 & n26851 ) | ( n22608 & n26852 ) | ( n26851 & n26852 ) ;
  assign n26854 = ~n26850 & n26853 ;
  assign n26855 = n26836 | n26854 ;
  assign n26856 = ( n26836 & n26840 ) | ( n26836 & n26855 ) | ( n26840 & n26855 ) ;
  assign n26857 = n26791 | n26806 ;
  assign n26858 = ~n26807 & n26857 ;
  assign n26859 = n26807 | n26858 ;
  assign n26860 = ( n26807 & n26856 ) | ( n26807 & n26859 ) | ( n26856 & n26859 ) ;
  assign n26861 = n26787 & n26860 ;
  assign n26862 = n26785 | n26861 ;
  assign n26863 = n26768 & n26862 ;
  assign n26864 = n26765 | n26863 ;
  assign n26865 = n3544 & n22381 ;
  assign n26866 = ( n3541 & n10490 ) | ( n3541 & n22381 ) | ( n10490 & n22381 ) ;
  assign n26867 = ( n23620 & n26865 ) | ( n23620 & n26866 ) | ( n26865 & n26866 ) ;
  assign n26868 = n3547 | n26866 ;
  assign n26869 = n3547 | n26865 ;
  assign n26870 = ( n23620 & n26868 ) | ( n23620 & n26869 ) | ( n26868 & n26869 ) ;
  assign n26871 = ( n23316 & n26867 ) | ( n23316 & n26870 ) | ( n26867 & n26870 ) ;
  assign n26872 = n3537 | n26871 ;
  assign n26873 = ~x20 & n26872 ;
  assign n26874 = ~x20 & n26871 ;
  assign n26875 = ( n23661 & n26873 ) | ( n23661 & n26874 ) | ( n26873 & n26874 ) ;
  assign n26876 = ( x20 & n14883 ) | ( x20 & n26871 ) | ( n14883 & n26871 ) ;
  assign n26877 = x20 & ~n26876 ;
  assign n26878 = x20 & n26871 ;
  assign n26879 = x20 & ~n26878 ;
  assign n26880 = ( ~n23661 & n26877 ) | ( ~n23661 & n26879 ) | ( n26877 & n26879 ) ;
  assign n26881 = n26875 | n26880 ;
  assign n26882 = n25282 & n25284 ;
  assign n26883 = n25282 | n25284 ;
  assign n26884 = ~n26882 & n26883 ;
  assign n26885 = n26881 & n26884 ;
  assign n26886 = n26881 | n26884 ;
  assign n26887 = ~n26885 & n26886 ;
  assign n26888 = n26885 | n26887 ;
  assign n26889 = ( n26864 & n26885 ) | ( n26864 & n26888 ) | ( n26885 & n26888 ) ;
  assign n26890 = n26746 & n26889 ;
  assign n26891 = n26743 | n26890 ;
  assign n26892 = ~n26688 & n26700 ;
  assign n26893 = ( n26688 & ~n26701 ) | ( n26688 & n26892 ) | ( ~n26701 & n26892 ) ;
  assign n26894 = n26891 & n26893 ;
  assign n26895 = n26720 | n26894 ;
  assign n26896 = ( n26723 & n26724 ) | ( n26723 & n26895 ) | ( n26724 & n26895 ) ;
  assign n26897 = n26683 | n26896 ;
  assign n26898 = ( n26683 & n26686 ) | ( n26683 & n26897 ) | ( n26686 & n26897 ) ;
  assign n26899 = ~n26649 & n26664 ;
  assign n26900 = ( n26649 & ~n26665 ) | ( n26649 & n26899 ) | ( ~n26665 & n26899 ) ;
  assign n26901 = n26665 | n26900 ;
  assign n26902 = ( n26665 & n26898 ) | ( n26665 & n26901 ) | ( n26898 & n26901 ) ;
  assign n26903 = ~n26646 & n26902 ;
  assign n26904 = n26643 | n26903 ;
  assign n26905 = n26622 | n26904 ;
  assign n26906 = ( n26622 & ~n26625 ) | ( n26622 & n26905 ) | ( ~n26625 & n26905 ) ;
  assign n26907 = n26589 | n26906 ;
  assign n26908 = ( n26589 & n26592 ) | ( n26589 & n26907 ) | ( n26592 & n26907 ) ;
  assign n26909 = n26565 | n26908 ;
  assign n26910 = n26565 & n26908 ;
  assign n26911 = n26909 & ~n26910 ;
  assign n27111 = n26500 | n26503 ;
  assign n27112 = n26481 & ~n26500 ;
  assign n27113 = ( n26501 & n27111 ) | ( n26501 & ~n27112 ) | ( n27111 & ~n27112 ) ;
  assign n26912 = n2064 | n20382 ;
  assign n26913 = n1463 | n26912 ;
  assign n26914 = n407 | n23885 ;
  assign n26915 = ( ~n1025 & n26913 ) | ( ~n1025 & n26914 ) | ( n26913 & n26914 ) ;
  assign n26916 = n26913 & n26914 ;
  assign n26917 = ( ~n1022 & n26915 ) | ( ~n1022 & n26916 ) | ( n26915 & n26916 ) ;
  assign n26918 = n1026 | n26917 ;
  assign n26919 = ~n10356 & n25492 ;
  assign n26920 = n575 | n3425 ;
  assign n26921 = n209 | n821 ;
  assign n26922 = n26920 | n26921 ;
  assign n26923 = n175 | n14391 ;
  assign n26924 = n295 | n26923 ;
  assign n26925 = n26922 | n26924 ;
  assign n26926 = n196 | n468 ;
  assign n26927 = n26925 | n26926 ;
  assign n26928 = n26919 & ~n26927 ;
  assign n26929 = ~n26918 & n26928 ;
  assign n26930 = ~n675 & n26929 ;
  assign n26931 = ( n26299 & ~n26301 ) | ( n26299 & n26930 ) | ( ~n26301 & n26930 ) ;
  assign n26932 = n26299 & n26930 ;
  assign n26933 = ( ~n26318 & n26931 ) | ( ~n26318 & n26932 ) | ( n26931 & n26932 ) ;
  assign n26934 = ~n26299 & n26301 ;
  assign n26935 = ~n26930 & n26934 ;
  assign n26936 = n26299 | n26930 ;
  assign n26937 = ( n26318 & n26935 ) | ( n26318 & ~n26936 ) | ( n26935 & ~n26936 ) ;
  assign n26938 = n26933 | n26937 ;
  assign n26939 = n1057 & ~n16085 ;
  assign n26940 = n1065 & n15434 ;
  assign n26941 = n1060 & n14591 ;
  assign n26942 = n26940 | n26941 ;
  assign n26943 = n26939 | n26942 ;
  assign n26944 = ~n26938 & n26943 ;
  assign n26945 = n1062 | n26939 ;
  assign n26946 = n26942 | n26945 ;
  assign n26947 = ~n26938 & n26946 ;
  assign n26948 = ( ~n16167 & n26944 ) | ( ~n16167 & n26947 ) | ( n26944 & n26947 ) ;
  assign n26949 = n26938 & ~n26946 ;
  assign n26950 = n26938 & ~n26943 ;
  assign n26951 = ( n16167 & n26949 ) | ( n16167 & n26950 ) | ( n26949 & n26950 ) ;
  assign n26952 = n26948 | n26951 ;
  assign n26953 = ~n26331 & n26339 ;
  assign n26954 = n26324 | n26953 ;
  assign n26955 = ~n26952 & n26954 ;
  assign n26956 = n26952 & ~n26954 ;
  assign n26957 = n26955 | n26956 ;
  assign n26958 = n1826 & n15886 ;
  assign n26959 = n1823 & ~n16069 ;
  assign n26960 = n26958 | n26959 ;
  assign n26961 = n1829 & n17111 ;
  assign n26962 = n1821 | n26961 ;
  assign n26963 = n26960 | n26962 ;
  assign n26964 = n26960 | n26961 ;
  assign n26965 = n17194 & ~n26964 ;
  assign n26966 = ( n17129 & ~n26964 ) | ( n17129 & n26965 ) | ( ~n26964 & n26965 ) ;
  assign n26967 = n26963 & ~n26966 ;
  assign n26968 = ( n17186 & n26963 ) | ( n17186 & n26967 ) | ( n26963 & n26967 ) ;
  assign n26969 = x29 & n26968 ;
  assign n26970 = x29 & ~n26968 ;
  assign n26971 = ( n26968 & ~n26969 ) | ( n26968 & n26970 ) | ( ~n26969 & n26970 ) ;
  assign n26972 = ~n26957 & n26971 ;
  assign n26973 = n26957 & ~n26971 ;
  assign n26974 = n26972 | n26973 ;
  assign n26975 = n26357 & ~n26974 ;
  assign n26976 = ( n26362 & ~n26974 ) | ( n26362 & n26975 ) | ( ~n26974 & n26975 ) ;
  assign n26977 = ~n26357 & n26974 ;
  assign n26978 = ~n26362 & n26977 ;
  assign n26979 = n26976 | n26978 ;
  assign n26980 = n2315 & n18037 ;
  assign n26981 = n2312 & n17100 ;
  assign n26982 = n2308 & ~n17092 ;
  assign n26983 = n26981 | n26982 ;
  assign n26984 = n26980 | n26983 ;
  assign n26985 = n2306 | n26980 ;
  assign n26986 = n26983 | n26985 ;
  assign n26987 = ( ~n18050 & n26984 ) | ( ~n18050 & n26986 ) | ( n26984 & n26986 ) ;
  assign n26988 = ~x26 & n26986 ;
  assign n26989 = ~x26 & n26984 ;
  assign n26990 = ( ~n18050 & n26988 ) | ( ~n18050 & n26989 ) | ( n26988 & n26989 ) ;
  assign n26991 = x26 | n26989 ;
  assign n26992 = x26 | n26988 ;
  assign n26993 = ( ~n18050 & n26991 ) | ( ~n18050 & n26992 ) | ( n26991 & n26992 ) ;
  assign n26994 = ( ~n26987 & n26990 ) | ( ~n26987 & n26993 ) | ( n26990 & n26993 ) ;
  assign n26995 = n26979 | n26994 ;
  assign n26996 = n26979 & ~n26994 ;
  assign n26997 = ( ~n26979 & n26995 ) | ( ~n26979 & n26996 ) | ( n26995 & n26996 ) ;
  assign n26998 = n26380 | n26385 ;
  assign n26999 = ~n26997 & n26998 ;
  assign n27000 = n26997 & ~n26998 ;
  assign n27001 = n26999 | n27000 ;
  assign n27002 = n2932 & n18576 ;
  assign n27003 = n2925 & ~n18585 ;
  assign n27004 = n2928 & n18410 ;
  assign n27005 = n27003 | n27004 ;
  assign n27006 = n27002 | n27005 ;
  assign n27007 = n2936 | n27002 ;
  assign n27008 = n27005 | n27007 ;
  assign n27009 = ( n18612 & n27006 ) | ( n18612 & n27008 ) | ( n27006 & n27008 ) ;
  assign n27010 = x23 & n27008 ;
  assign n27011 = x23 & n27006 ;
  assign n27012 = ( n18612 & n27010 ) | ( n18612 & n27011 ) | ( n27010 & n27011 ) ;
  assign n27013 = x23 & ~n27011 ;
  assign n27014 = x23 & ~n27010 ;
  assign n27015 = ( ~n18612 & n27013 ) | ( ~n18612 & n27014 ) | ( n27013 & n27014 ) ;
  assign n27016 = ( n27009 & ~n27012 ) | ( n27009 & n27015 ) | ( ~n27012 & n27015 ) ;
  assign n27017 = n27001 | n27016 ;
  assign n27018 = n27001 & ~n27016 ;
  assign n27019 = ( ~n27001 & n27017 ) | ( ~n27001 & n27018 ) | ( n27017 & n27018 ) ;
  assign n27020 = n26402 | n26406 ;
  assign n27021 = ~n26402 & n26403 ;
  assign n27022 = ( n26407 & n27020 ) | ( n26407 & ~n27021 ) | ( n27020 & ~n27021 ) ;
  assign n27023 = ~n27019 & n27022 ;
  assign n27024 = n27019 & ~n27022 ;
  assign n27025 = n27023 | n27024 ;
  assign n27026 = n3547 & n19631 ;
  assign n27027 = n3544 & n19352 ;
  assign n27028 = n3541 & n19494 ;
  assign n27029 = n27027 | n27028 ;
  assign n27030 = n27026 | n27029 ;
  assign n27031 = n3537 & n19652 ;
  assign n27032 = n3537 & n19655 ;
  assign n27033 = ( ~n18604 & n27031 ) | ( ~n18604 & n27032 ) | ( n27031 & n27032 ) ;
  assign n27034 = n27030 | n27033 ;
  assign n27035 = n3537 | n27030 ;
  assign n27036 = ( n19640 & n27034 ) | ( n19640 & n27035 ) | ( n27034 & n27035 ) ;
  assign n27037 = x20 | n27036 ;
  assign n27038 = ~x20 & n27036 ;
  assign n27039 = ( ~n27036 & n27037 ) | ( ~n27036 & n27038 ) | ( n27037 & n27038 ) ;
  assign n27040 = n27025 | n27039 ;
  assign n27041 = n27025 & ~n27039 ;
  assign n27042 = ( ~n27025 & n27040 ) | ( ~n27025 & n27041 ) | ( n27040 & n27041 ) ;
  assign n27043 = n26428 | n26435 ;
  assign n27044 = ~n27042 & n27043 ;
  assign n27045 = n27042 & ~n27043 ;
  assign n27046 = n27044 | n27045 ;
  assign n27047 = n4471 & n20609 ;
  assign n27048 = n4466 & ~n20630 ;
  assign n27049 = n4468 & ~n20618 ;
  assign n27050 = n27048 | n27049 ;
  assign n27051 = n27047 | n27050 ;
  assign n27052 = n4475 | n27047 ;
  assign n27053 = n27050 | n27052 ;
  assign n27054 = ( n20659 & n27051 ) | ( n20659 & n27053 ) | ( n27051 & n27053 ) ;
  assign n27055 = n27051 & n27053 ;
  assign n27056 = ( ~n20649 & n27054 ) | ( ~n20649 & n27055 ) | ( n27054 & n27055 ) ;
  assign n27057 = x17 & n27056 ;
  assign n27058 = x17 & ~n27056 ;
  assign n27059 = ( n27056 & ~n27057 ) | ( n27056 & n27058 ) | ( ~n27057 & n27058 ) ;
  assign n27060 = n27046 | n27059 ;
  assign n27061 = n27046 & ~n27059 ;
  assign n27062 = ( ~n27046 & n27060 ) | ( ~n27046 & n27061 ) | ( n27060 & n27061 ) ;
  assign n27063 = n26450 | n26455 ;
  assign n27064 = ( n26450 & ~n26453 ) | ( n26450 & n27063 ) | ( ~n26453 & n27063 ) ;
  assign n27065 = ~n27062 & n27064 ;
  assign n27066 = n27062 & ~n27064 ;
  assign n27067 = n27065 | n27066 ;
  assign n27068 = n5234 & ~n21551 ;
  assign n27069 = n5237 & ~n21563 ;
  assign n27070 = n5231 & ~n21517 ;
  assign n27071 = n27069 | n27070 ;
  assign n27072 = n27068 | n27071 ;
  assign n27073 = n5227 | n27068 ;
  assign n27074 = n27071 | n27073 ;
  assign n27075 = ( ~n21587 & n27072 ) | ( ~n21587 & n27074 ) | ( n27072 & n27074 ) ;
  assign n27076 = ~x14 & n27074 ;
  assign n27077 = ~x14 & n27072 ;
  assign n27078 = ( ~n21587 & n27076 ) | ( ~n21587 & n27077 ) | ( n27076 & n27077 ) ;
  assign n27079 = x14 | n27077 ;
  assign n27080 = x14 | n27076 ;
  assign n27081 = ( ~n21587 & n27079 ) | ( ~n21587 & n27080 ) | ( n27079 & n27080 ) ;
  assign n27082 = ( ~n27075 & n27078 ) | ( ~n27075 & n27081 ) | ( n27078 & n27081 ) ;
  assign n27083 = n27067 | n27082 ;
  assign n27084 = n27067 & ~n27082 ;
  assign n27085 = ( ~n27067 & n27083 ) | ( ~n27067 & n27084 ) | ( n27083 & n27084 ) ;
  assign n27086 = n26472 | n26478 ;
  assign n27087 = ~n27085 & n27086 ;
  assign n27088 = n27085 & ~n27086 ;
  assign n27089 = n27087 | n27088 ;
  assign n27090 = n6119 & ~n23240 ;
  assign n27091 = n6125 & n23227 ;
  assign n27092 = ( n6125 & n23217 ) | ( n6125 & n27091 ) | ( n23217 & n27091 ) ;
  assign n27093 = n27090 | n27092 ;
  assign n27094 = n6122 & ~n23234 ;
  assign n27095 = n6122 & ~n23235 ;
  assign n27096 = ( ~n15882 & n27094 ) | ( ~n15882 & n27095 ) | ( n27094 & n27095 ) ;
  assign n27097 = n27093 | n27096 ;
  assign n27098 = n6115 | n27096 ;
  assign n27099 = n27093 | n27098 ;
  assign n27100 = ( ~n23587 & n27097 ) | ( ~n23587 & n27099 ) | ( n27097 & n27099 ) ;
  assign n27101 = ~x11 & n27099 ;
  assign n27102 = ~x11 & n27097 ;
  assign n27103 = ( ~n23587 & n27101 ) | ( ~n23587 & n27102 ) | ( n27101 & n27102 ) ;
  assign n27104 = x11 | n27102 ;
  assign n27105 = x11 | n27101 ;
  assign n27106 = ( ~n23587 & n27104 ) | ( ~n23587 & n27105 ) | ( n27104 & n27105 ) ;
  assign n27107 = ( ~n27100 & n27103 ) | ( ~n27100 & n27106 ) | ( n27103 & n27106 ) ;
  assign n27108 = n27089 | n27107 ;
  assign n27109 = n27089 & ~n27107 ;
  assign n27110 = ( ~n27089 & n27108 ) | ( ~n27089 & n27109 ) | ( n27108 & n27109 ) ;
  assign n27114 = ~n27110 & n27113 ;
  assign n27115 = n27113 & ~n27114 ;
  assign n27116 = n27110 | n27113 ;
  assign n27117 = ~n27115 & n27116 ;
  assign n27118 = ~n26511 & n26513 ;
  assign n27119 = ( n26511 & n26516 ) | ( n26511 & ~n27118 ) | ( n26516 & ~n27118 ) ;
  assign n27120 = n26511 | n26522 ;
  assign n27121 = ( n26266 & ~n27118 ) | ( n26266 & n27120 ) | ( ~n27118 & n27120 ) ;
  assign n27122 = ( n26009 & n27119 ) | ( n26009 & n27121 ) | ( n27119 & n27121 ) ;
  assign n27123 = ( n26011 & n27119 ) | ( n26011 & n27121 ) | ( n27119 & n27121 ) ;
  assign n27124 = ( n24765 & n27122 ) | ( n24765 & n27123 ) | ( n27122 & n27123 ) ;
  assign n27125 = n27117 & ~n27124 ;
  assign n27126 = n27117 | n27118 ;
  assign n27127 = n26511 & ~n27117 ;
  assign n27128 = ( n26516 & ~n27126 ) | ( n26516 & n27127 ) | ( ~n27126 & n27127 ) ;
  assign n27129 = ~n27117 & n27120 ;
  assign n27130 = ( n26266 & ~n27126 ) | ( n26266 & n27129 ) | ( ~n27126 & n27129 ) ;
  assign n27131 = ( n26009 & n27128 ) | ( n26009 & n27130 ) | ( n27128 & n27130 ) ;
  assign n27132 = ( n26011 & n27128 ) | ( n26011 & n27130 ) | ( n27128 & n27130 ) ;
  assign n27133 = ( n24765 & n27131 ) | ( n24765 & n27132 ) | ( n27131 & n27132 ) ;
  assign n27134 = n4466 & ~n27133 ;
  assign n27135 = ~n27125 & n27134 ;
  assign n27136 = n6119 | n6122 ;
  assign n27137 = ~n23234 & n27136 ;
  assign n27138 = n6125 | n27137 ;
  assign n27139 = ~n23235 & n27136 ;
  assign n27140 = n6125 | n27139 ;
  assign n27141 = ( ~n15882 & n27138 ) | ( ~n15882 & n27140 ) | ( n27138 & n27140 ) ;
  assign n27142 = n6115 | n27141 ;
  assign n27143 = ( ~n15882 & n27137 ) | ( ~n15882 & n27139 ) | ( n27137 & n27139 ) ;
  assign n27144 = n6115 | n27143 ;
  assign n27145 = ( ~n23240 & n27142 ) | ( ~n23240 & n27144 ) | ( n27142 & n27144 ) ;
  assign n27146 = ( ~n23240 & n27141 ) | ( ~n23240 & n27143 ) | ( n27141 & n27143 ) ;
  assign n27147 = n24135 & ~n27146 ;
  assign n27148 = n23240 & ~n27146 ;
  assign n27149 = ( n23575 & n27147 ) | ( n23575 & n27148 ) | ( n27147 & n27148 ) ;
  assign n27150 = ( n23577 & n27147 ) | ( n23577 & n27148 ) | ( n27147 & n27148 ) ;
  assign n27151 = ( ~n21554 & n27149 ) | ( ~n21554 & n27150 ) | ( n27149 & n27150 ) ;
  assign n27152 = n27145 & ~n27151 ;
  assign n27153 = x11 & ~n27152 ;
  assign n27154 = n27149 | n27150 ;
  assign n27155 = n27145 & ~n27154 ;
  assign n27156 = x11 & ~n27155 ;
  assign n27157 = ( n21584 & n27153 ) | ( n21584 & n27156 ) | ( n27153 & n27156 ) ;
  assign n27158 = ~x11 & n27152 ;
  assign n27159 = ~x11 & n27155 ;
  assign n27160 = ( ~n21584 & n27158 ) | ( ~n21584 & n27159 ) | ( n27158 & n27159 ) ;
  assign n27161 = n27157 | n27160 ;
  assign n27162 = n27065 | n27082 ;
  assign n27163 = ( n27065 & ~n27067 ) | ( n27065 & n27162 ) | ( ~n27067 & n27162 ) ;
  assign n27164 = n27161 & n27163 ;
  assign n27165 = n27161 | n27163 ;
  assign n27166 = ~n27164 & n27165 ;
  assign n27167 = n26933 | n26944 ;
  assign n27168 = n26933 | n26947 ;
  assign n27169 = ( ~n16167 & n27167 ) | ( ~n16167 & n27168 ) | ( n27167 & n27168 ) ;
  assign n27170 = n5058 | n7927 ;
  assign n27171 = n3447 | n27170 ;
  assign n27172 = n1771 | n27171 ;
  assign n27173 = n10754 | n27172 ;
  assign n27174 = n10730 | n27173 ;
  assign n27175 = n10724 & ~n27174 ;
  assign n27176 = n679 | n1001 ;
  assign n27177 = n442 | n602 ;
  assign n27178 = n27176 | n27177 ;
  assign n27179 = n64 | n258 ;
  assign n27180 = n725 | n27179 ;
  assign n27181 = n623 | n27180 ;
  assign n27182 = n27178 | n27181 ;
  assign n27183 = n75 | n27182 ;
  assign n27184 = n12266 | n12270 ;
  assign n27185 = n12263 | n27184 ;
  assign n27186 = n4293 | n27185 ;
  assign n27187 = n15584 | n27186 ;
  assign n27188 = n27183 | n27187 ;
  assign n27189 = n27175 & ~n27188 ;
  assign n27190 = n675 & n27189 ;
  assign n27191 = ( ~n26929 & n27189 ) | ( ~n26929 & n27190 ) | ( n27189 & n27190 ) ;
  assign n27192 = n675 | n27189 ;
  assign n27193 = n26929 & ~n27192 ;
  assign n27194 = n26933 & ~n27193 ;
  assign n27195 = ~n27191 & n27194 ;
  assign n27196 = n27191 | n27193 ;
  assign n27197 = ( n26944 & n27195 ) | ( n26944 & ~n27196 ) | ( n27195 & ~n27196 ) ;
  assign n27198 = ( n26947 & n27195 ) | ( n26947 & ~n27196 ) | ( n27195 & ~n27196 ) ;
  assign n27199 = ( ~n16167 & n27197 ) | ( ~n16167 & n27198 ) | ( n27197 & n27198 ) ;
  assign n27200 = n27169 & ~n27199 ;
  assign n27201 = n1057 & n15886 ;
  assign n27202 = n1060 & n15434 ;
  assign n27203 = n1065 & ~n16085 ;
  assign n27204 = n27202 | n27203 ;
  assign n27205 = n27201 | n27204 ;
  assign n27206 = n1062 | n27201 ;
  assign n27207 = n27204 | n27206 ;
  assign n27208 = ( ~n16140 & n27205 ) | ( ~n16140 & n27207 ) | ( n27205 & n27207 ) ;
  assign n27209 = n27193 | n27198 ;
  assign n27210 = n27191 | n27209 ;
  assign n27211 = n27193 | n27197 ;
  assign n27212 = n27191 | n27211 ;
  assign n27213 = ( ~n16167 & n27210 ) | ( ~n16167 & n27212 ) | ( n27210 & n27212 ) ;
  assign n27214 = n27208 & ~n27213 ;
  assign n27215 = ( n27200 & n27208 ) | ( n27200 & n27214 ) | ( n27208 & n27214 ) ;
  assign n27216 = ~n27208 & n27213 ;
  assign n27217 = ~n27200 & n27216 ;
  assign n27218 = n27215 | n27217 ;
  assign n27219 = n1826 & ~n16069 ;
  assign n27220 = n1823 & n17111 ;
  assign n27221 = n27219 | n27220 ;
  assign n27222 = n1829 & n17100 ;
  assign n27223 = n1821 | n27222 ;
  assign n27224 = n27221 | n27223 ;
  assign n27225 = n27221 | n27222 ;
  assign n27226 = n17169 | n27225 ;
  assign n27227 = ( ~n17129 & n27225 ) | ( ~n17129 & n27226 ) | ( n27225 & n27226 ) ;
  assign n27228 = n27224 & n27227 ;
  assign n27229 = ( n17161 & n27224 ) | ( n17161 & n27228 ) | ( n27224 & n27228 ) ;
  assign n27230 = ~x29 & n27229 ;
  assign n27231 = x29 | n27229 ;
  assign n27232 = ( ~n27229 & n27230 ) | ( ~n27229 & n27231 ) | ( n27230 & n27231 ) ;
  assign n27233 = ~n27218 & n27232 ;
  assign n27234 = n27218 & ~n27232 ;
  assign n27235 = n27233 | n27234 ;
  assign n27236 = n26955 | n26971 ;
  assign n27237 = ( n26955 & ~n26957 ) | ( n26955 & n27236 ) | ( ~n26957 & n27236 ) ;
  assign n27238 = ~n27235 & n27237 ;
  assign n27239 = n27235 & ~n27237 ;
  assign n27240 = n27238 | n27239 ;
  assign n27241 = n2315 & ~n18585 ;
  assign n27242 = n2312 & ~n17092 ;
  assign n27243 = n2308 & n18037 ;
  assign n27244 = n27242 | n27243 ;
  assign n27245 = n27241 | n27244 ;
  assign n27246 = n2306 & ~n18675 ;
  assign n27247 = ( n2306 & n18672 ) | ( n2306 & n27246 ) | ( n18672 & n27246 ) ;
  assign n27248 = n27245 | n27247 ;
  assign n27249 = x26 | n27245 ;
  assign n27250 = n27247 | n27249 ;
  assign n27251 = ~x26 & n27249 ;
  assign n27252 = ( ~x26 & n27247 ) | ( ~x26 & n27251 ) | ( n27247 & n27251 ) ;
  assign n27253 = ( ~n27248 & n27250 ) | ( ~n27248 & n27252 ) | ( n27250 & n27252 ) ;
  assign n27254 = n27240 | n27253 ;
  assign n27255 = n27240 & ~n27253 ;
  assign n27256 = ( ~n27240 & n27254 ) | ( ~n27240 & n27255 ) | ( n27254 & n27255 ) ;
  assign n27257 = n26976 | n26994 ;
  assign n27258 = ( n26976 & ~n26979 ) | ( n26976 & n27257 ) | ( ~n26979 & n27257 ) ;
  assign n27259 = ~n27256 & n27258 ;
  assign n27260 = n27256 & ~n27258 ;
  assign n27261 = n27259 | n27260 ;
  assign n27262 = n2932 & n19352 ;
  assign n27263 = n2925 & n18410 ;
  assign n27264 = n2928 & n18576 ;
  assign n27265 = n27263 | n27264 ;
  assign n27266 = n27262 | n27265 ;
  assign n27267 = n2936 | n27262 ;
  assign n27268 = n27265 | n27267 ;
  assign n27269 = ( n19674 & n27266 ) | ( n19674 & n27268 ) | ( n27266 & n27268 ) ;
  assign n27270 = x23 & n27268 ;
  assign n27271 = x23 & n27266 ;
  assign n27272 = ( n19674 & n27270 ) | ( n19674 & n27271 ) | ( n27270 & n27271 ) ;
  assign n27273 = x23 & ~n27271 ;
  assign n27274 = x23 & ~n27270 ;
  assign n27275 = ( ~n19674 & n27273 ) | ( ~n19674 & n27274 ) | ( n27273 & n27274 ) ;
  assign n27276 = ( n27269 & ~n27272 ) | ( n27269 & n27275 ) | ( ~n27272 & n27275 ) ;
  assign n27277 = n27261 | n27276 ;
  assign n27278 = n27261 & ~n27276 ;
  assign n27279 = ( ~n27261 & n27277 ) | ( ~n27261 & n27278 ) | ( n27277 & n27278 ) ;
  assign n27280 = n26999 | n27016 ;
  assign n27281 = ( n26999 & ~n27001 ) | ( n26999 & n27280 ) | ( ~n27001 & n27280 ) ;
  assign n27282 = ~n27279 & n27281 ;
  assign n27283 = n27279 & ~n27281 ;
  assign n27284 = n27282 | n27283 ;
  assign n27285 = n3547 & ~n20630 ;
  assign n27286 = n3544 & n19494 ;
  assign n27287 = n3541 & n19631 ;
  assign n27288 = n27286 | n27287 ;
  assign n27289 = n27285 | n27288 ;
  assign n27290 = n3537 | n27285 ;
  assign n27291 = n27288 | n27290 ;
  assign n27292 = ( ~n20709 & n27289 ) | ( ~n20709 & n27291 ) | ( n27289 & n27291 ) ;
  assign n27293 = ~x20 & n27291 ;
  assign n27294 = ~x20 & n27289 ;
  assign n27295 = ( ~n20709 & n27293 ) | ( ~n20709 & n27294 ) | ( n27293 & n27294 ) ;
  assign n27296 = x20 | n27294 ;
  assign n27297 = x20 | n27293 ;
  assign n27298 = ( ~n20709 & n27296 ) | ( ~n20709 & n27297 ) | ( n27296 & n27297 ) ;
  assign n27299 = ( ~n27292 & n27295 ) | ( ~n27292 & n27298 ) | ( n27295 & n27298 ) ;
  assign n27300 = n27284 | n27299 ;
  assign n27301 = n27284 & ~n27299 ;
  assign n27302 = ( ~n27284 & n27300 ) | ( ~n27284 & n27301 ) | ( n27300 & n27301 ) ;
  assign n27303 = n27023 | n27039 ;
  assign n27304 = ( n27023 & ~n27025 ) | ( n27023 & n27303 ) | ( ~n27025 & n27303 ) ;
  assign n27305 = ~n27302 & n27304 ;
  assign n27306 = n27302 & ~n27304 ;
  assign n27307 = n27305 | n27306 ;
  assign n27308 = n4471 & ~n21563 ;
  assign n27309 = n4466 & ~n20618 ;
  assign n27310 = n4468 & n20609 ;
  assign n27311 = n27309 | n27310 ;
  assign n27312 = n27308 | n27311 ;
  assign n27313 = n4475 & ~n21570 ;
  assign n27314 = n22270 & n27313 ;
  assign n27315 = ( n4475 & n22304 ) | ( n4475 & n27314 ) | ( n22304 & n27314 ) ;
  assign n27316 = n27312 | n27315 ;
  assign n27317 = x17 | n27312 ;
  assign n27318 = n27315 | n27317 ;
  assign n27319 = ~x17 & n27317 ;
  assign n27320 = ( ~x17 & n27315 ) | ( ~x17 & n27319 ) | ( n27315 & n27319 ) ;
  assign n27321 = ( ~n27316 & n27318 ) | ( ~n27316 & n27320 ) | ( n27318 & n27320 ) ;
  assign n27322 = n27307 | n27321 ;
  assign n27323 = n27307 & ~n27321 ;
  assign n27324 = ( ~n27307 & n27322 ) | ( ~n27307 & n27323 ) | ( n27322 & n27323 ) ;
  assign n27325 = n27044 | n27059 ;
  assign n27326 = ( n27044 & ~n27046 ) | ( n27044 & n27325 ) | ( ~n27046 & n27325 ) ;
  assign n27327 = ~n27324 & n27326 ;
  assign n27328 = n27324 & ~n27326 ;
  assign n27329 = n27327 | n27328 ;
  assign n27330 = n5237 & ~n21517 ;
  assign n27331 = n5231 & ~n21551 ;
  assign n27332 = n27330 | n27331 ;
  assign n27333 = n5234 & n23227 ;
  assign n27334 = ( n5234 & n23217 ) | ( n5234 & n27333 ) | ( n23217 & n27333 ) ;
  assign n27335 = n27332 | n27334 ;
  assign n27336 = n5227 & n23299 ;
  assign n27337 = n5227 & n23298 ;
  assign n27338 = ( n21584 & n27336 ) | ( n21584 & n27337 ) | ( n27336 & n27337 ) ;
  assign n27339 = n27335 | n27338 ;
  assign n27340 = n5227 | n27335 ;
  assign n27341 = ( n23289 & n27339 ) | ( n23289 & n27340 ) | ( n27339 & n27340 ) ;
  assign n27342 = x14 | n27341 ;
  assign n27343 = ~x14 & n27341 ;
  assign n27344 = ( ~n27341 & n27342 ) | ( ~n27341 & n27343 ) | ( n27342 & n27343 ) ;
  assign n27345 = n27329 | n27344 ;
  assign n27346 = n27329 & ~n27344 ;
  assign n27347 = ( ~n27329 & n27345 ) | ( ~n27329 & n27346 ) | ( n27345 & n27346 ) ;
  assign n27348 = n27166 & ~n27347 ;
  assign n27349 = n27166 | n27347 ;
  assign n27350 = ( ~n27166 & n27348 ) | ( ~n27166 & n27349 ) | ( n27348 & n27349 ) ;
  assign n27351 = n27087 | n27107 ;
  assign n27352 = ( n27087 & ~n27089 ) | ( n27087 & n27351 ) | ( ~n27089 & n27351 ) ;
  assign n27353 = ~n27350 & n27352 ;
  assign n27354 = n27350 & ~n27352 ;
  assign n27355 = n27353 | n27354 ;
  assign n27356 = n27114 | n27130 ;
  assign n27357 = ~n27114 & n27126 ;
  assign n27358 = n27114 | n27127 ;
  assign n27359 = ( n26516 & ~n27357 ) | ( n26516 & n27358 ) | ( ~n27357 & n27358 ) ;
  assign n27360 = ( n26009 & n27356 ) | ( n26009 & n27359 ) | ( n27356 & n27359 ) ;
  assign n27361 = ( n26011 & n27356 ) | ( n26011 & n27359 ) | ( n27356 & n27359 ) ;
  assign n27362 = ( n24765 & n27360 ) | ( n24765 & n27361 ) | ( n27360 & n27361 ) ;
  assign n27363 = n27355 & ~n27362 ;
  assign n27364 = n27355 | n27357 ;
  assign n27365 = ~n27355 & n27358 ;
  assign n27366 = ( n26516 & ~n27364 ) | ( n26516 & n27365 ) | ( ~n27364 & n27365 ) ;
  assign n27367 = n27114 & ~n27355 ;
  assign n27368 = ( n27130 & ~n27355 ) | ( n27130 & n27367 ) | ( ~n27355 & n27367 ) ;
  assign n27369 = ( n26009 & n27366 ) | ( n26009 & n27368 ) | ( n27366 & n27368 ) ;
  assign n27370 = ( n26011 & n27366 ) | ( n26011 & n27368 ) | ( n27366 & n27368 ) ;
  assign n27371 = ( n24765 & n27369 ) | ( n24765 & n27370 ) | ( n27369 & n27370 ) ;
  assign n27372 = n4468 & ~n27371 ;
  assign n27373 = ~n27363 & n27372 ;
  assign n27374 = n27135 | n27373 ;
  assign n27375 = n27215 | n27233 ;
  assign n27376 = ( ~n16167 & n27209 ) | ( ~n16167 & n27211 ) | ( n27209 & n27211 ) ;
  assign n27377 = n1135 | n5158 ;
  assign n27378 = n795 | n2256 ;
  assign n27379 = n27377 | n27378 ;
  assign n27380 = n12702 | n27379 ;
  assign n27381 = n3999 | n4352 ;
  assign n27382 = n27380 | n27381 ;
  assign n27383 = n6868 & ~n6992 ;
  assign n27384 = ~n27382 & n27383 ;
  assign n27385 = n257 | n1693 ;
  assign n27386 = n4305 | n27385 ;
  assign n27387 = n514 | n886 ;
  assign n27388 = n663 | n27387 ;
  assign n27389 = n14392 | n27388 ;
  assign n27390 = n27386 | n27389 ;
  assign n27391 = n581 | n841 ;
  assign n27392 = n193 | n27391 ;
  assign n27393 = n27390 | n27392 ;
  assign n27394 = n131 | n27393 ;
  assign n27395 = n27384 & ~n27394 ;
  assign n27396 = n26930 | n27395 ;
  assign n27397 = n26930 & n27395 ;
  assign n27398 = n27396 & ~n27397 ;
  assign n27399 = n6125 | n27136 ;
  assign n27400 = n6115 | n27399 ;
  assign n27401 = ~n23229 & n27400 ;
  assign n27402 = ( n23154 & n27400 ) | ( n23154 & n27401 ) | ( n27400 & n27401 ) ;
  assign n27403 = ~n23232 & n27400 ;
  assign n27404 = ~n23231 & n27400 ;
  assign n27405 = ( n9072 & n27403 ) | ( n9072 & n27404 ) | ( n27403 & n27404 ) ;
  assign n27406 = ( ~n21543 & n27402 ) | ( ~n21543 & n27405 ) | ( n27402 & n27405 ) ;
  assign n27407 = ( ~n21545 & n27402 ) | ( ~n21545 & n27405 ) | ( n27402 & n27405 ) ;
  assign n27408 = ( ~n15882 & n27406 ) | ( ~n15882 & n27407 ) | ( n27406 & n27407 ) ;
  assign n27409 = ~x11 & n27406 ;
  assign n27410 = ~x11 & n27407 ;
  assign n27411 = ( ~n15882 & n27409 ) | ( ~n15882 & n27410 ) | ( n27409 & n27410 ) ;
  assign n27412 = x11 | n27409 ;
  assign n27413 = x11 | n27410 ;
  assign n27414 = ( ~n15882 & n27412 ) | ( ~n15882 & n27413 ) | ( n27412 & n27413 ) ;
  assign n27415 = ( ~n27408 & n27411 ) | ( ~n27408 & n27414 ) | ( n27411 & n27414 ) ;
  assign n27416 = n27398 & ~n27415 ;
  assign n27417 = ~n27398 & n27415 ;
  assign n27418 = n27416 | n27417 ;
  assign n27419 = n1057 & ~n16069 ;
  assign n27420 = n1060 & ~n16085 ;
  assign n27421 = n1065 & n15886 ;
  assign n27422 = n27420 | n27421 ;
  assign n27423 = n27419 | n27422 ;
  assign n27424 = n1062 | n27423 ;
  assign n27425 = ~n27418 & n27424 ;
  assign n27426 = ~n27418 & n27423 ;
  assign n27427 = ( ~n16107 & n27425 ) | ( ~n16107 & n27426 ) | ( n27425 & n27426 ) ;
  assign n27428 = ( ~n16107 & n27423 ) | ( ~n16107 & n27424 ) | ( n27423 & n27424 ) ;
  assign n27429 = ~n27427 & n27428 ;
  assign n27430 = n27418 | n27424 ;
  assign n27431 = n27418 | n27423 ;
  assign n27432 = ( ~n16107 & n27430 ) | ( ~n16107 & n27431 ) | ( n27430 & n27431 ) ;
  assign n27433 = n27376 & ~n27432 ;
  assign n27434 = ( n27376 & n27429 ) | ( n27376 & n27433 ) | ( n27429 & n27433 ) ;
  assign n27435 = ~n27376 & n27432 ;
  assign n27436 = ~n27429 & n27435 ;
  assign n27437 = n27434 | n27436 ;
  assign n27438 = n27215 & ~n27437 ;
  assign n27439 = ( n27233 & ~n27437 ) | ( n27233 & n27438 ) | ( ~n27437 & n27438 ) ;
  assign n27440 = n27375 & ~n27439 ;
  assign n27441 = n1829 & ~n17092 ;
  assign n27442 = n1826 & n17111 ;
  assign n27443 = n1823 & n17100 ;
  assign n27444 = n27442 | n27443 ;
  assign n27445 = n27441 | n27444 ;
  assign n27446 = n1821 | n27441 ;
  assign n27447 = n27444 | n27446 ;
  assign n27448 = ( ~n17134 & n27445 ) | ( ~n17134 & n27447 ) | ( n27445 & n27447 ) ;
  assign n27449 = ~x29 & n27447 ;
  assign n27450 = ~x29 & n27445 ;
  assign n27451 = ( ~n17134 & n27449 ) | ( ~n17134 & n27450 ) | ( n27449 & n27450 ) ;
  assign n27452 = x29 | n27450 ;
  assign n27453 = x29 | n27449 ;
  assign n27454 = ( ~n17134 & n27452 ) | ( ~n17134 & n27453 ) | ( n27452 & n27453 ) ;
  assign n27455 = ( ~n27448 & n27451 ) | ( ~n27448 & n27454 ) | ( n27451 & n27454 ) ;
  assign n27456 = n27215 | n27437 ;
  assign n27457 = n27233 | n27456 ;
  assign n27458 = n27455 & ~n27457 ;
  assign n27459 = ( n27440 & n27455 ) | ( n27440 & n27458 ) | ( n27455 & n27458 ) ;
  assign n27460 = ~n27455 & n27457 ;
  assign n27461 = ~n27440 & n27460 ;
  assign n27462 = n27459 | n27461 ;
  assign n27463 = n2315 & n18410 ;
  assign n27464 = n2312 & n18037 ;
  assign n27465 = n2308 & ~n18585 ;
  assign n27466 = n27464 | n27465 ;
  assign n27467 = n27463 | n27466 ;
  assign n27468 = n2306 & ~n18586 ;
  assign n27469 = ~n18609 & n27468 ;
  assign n27470 = ( n2306 & n18650 ) | ( n2306 & n27469 ) | ( n18650 & n27469 ) ;
  assign n27471 = n27467 | n27470 ;
  assign n27472 = x26 | n27467 ;
  assign n27473 = n27470 | n27472 ;
  assign n27474 = ~x26 & n27472 ;
  assign n27475 = ( ~x26 & n27470 ) | ( ~x26 & n27474 ) | ( n27470 & n27474 ) ;
  assign n27476 = ( ~n27471 & n27473 ) | ( ~n27471 & n27475 ) | ( n27473 & n27475 ) ;
  assign n27477 = ~n27462 & n27476 ;
  assign n27478 = n27462 | n27477 ;
  assign n27480 = n27238 | n27253 ;
  assign n27481 = ( n27238 & ~n27240 ) | ( n27238 & n27480 ) | ( ~n27240 & n27480 ) ;
  assign n27479 = n27462 & n27476 ;
  assign n27482 = n27479 & n27481 ;
  assign n27483 = ( ~n27478 & n27481 ) | ( ~n27478 & n27482 ) | ( n27481 & n27482 ) ;
  assign n27484 = n27479 | n27481 ;
  assign n27485 = n27478 & ~n27484 ;
  assign n27486 = n27483 | n27485 ;
  assign n27487 = n2932 & n19494 ;
  assign n27488 = n2925 & n18576 ;
  assign n27489 = n2928 & n19352 ;
  assign n27490 = n27488 | n27489 ;
  assign n27491 = n27487 | n27490 ;
  assign n27492 = n2936 | n27487 ;
  assign n27493 = n27490 | n27492 ;
  assign n27494 = ( n20320 & n27491 ) | ( n20320 & n27493 ) | ( n27491 & n27493 ) ;
  assign n27495 = x23 & n27493 ;
  assign n27496 = x23 & n27491 ;
  assign n27497 = ( n20320 & n27495 ) | ( n20320 & n27496 ) | ( n27495 & n27496 ) ;
  assign n27498 = x23 & ~n27496 ;
  assign n27499 = x23 & ~n27495 ;
  assign n27500 = ( ~n20320 & n27498 ) | ( ~n20320 & n27499 ) | ( n27498 & n27499 ) ;
  assign n27501 = ( n27494 & ~n27497 ) | ( n27494 & n27500 ) | ( ~n27497 & n27500 ) ;
  assign n27502 = ~n27486 & n27501 ;
  assign n27503 = n27486 | n27502 ;
  assign n27505 = n27259 | n27276 ;
  assign n27506 = ( n27259 & ~n27261 ) | ( n27259 & n27505 ) | ( ~n27261 & n27505 ) ;
  assign n27504 = n27486 & n27501 ;
  assign n27507 = n27504 & n27506 ;
  assign n27508 = ( ~n27503 & n27506 ) | ( ~n27503 & n27507 ) | ( n27506 & n27507 ) ;
  assign n27509 = n27504 | n27506 ;
  assign n27510 = n27503 & ~n27509 ;
  assign n27511 = n27508 | n27510 ;
  assign n27512 = n3537 & n20680 ;
  assign n27513 = n3547 & ~n20618 ;
  assign n27514 = n3544 & n19631 ;
  assign n27515 = n3541 & ~n20630 ;
  assign n27516 = n27514 | n27515 ;
  assign n27517 = n27513 | n27516 ;
  assign n27518 = n20689 | n27517 ;
  assign n27519 = n3537 | n27517 ;
  assign n27520 = ( n27512 & n27518 ) | ( n27512 & n27519 ) | ( n27518 & n27519 ) ;
  assign n27521 = x20 | n27520 ;
  assign n27522 = ~x20 & n27520 ;
  assign n27523 = ( ~n27520 & n27521 ) | ( ~n27520 & n27522 ) | ( n27521 & n27522 ) ;
  assign n27524 = ~n27511 & n27523 ;
  assign n27525 = n27511 | n27524 ;
  assign n27527 = n27282 | n27299 ;
  assign n27528 = ( n27282 & ~n27284 ) | ( n27282 & n27527 ) | ( ~n27284 & n27527 ) ;
  assign n27526 = n27511 & n27523 ;
  assign n27529 = n27526 & n27528 ;
  assign n27530 = ( ~n27525 & n27528 ) | ( ~n27525 & n27529 ) | ( n27528 & n27529 ) ;
  assign n27531 = n27526 | n27528 ;
  assign n27532 = n27525 & ~n27531 ;
  assign n27533 = n27530 | n27532 ;
  assign n27534 = n4471 & ~n21517 ;
  assign n27535 = n4466 & n20609 ;
  assign n27536 = n4468 & ~n21563 ;
  assign n27537 = n27535 | n27536 ;
  assign n27538 = n27534 | n27537 ;
  assign n27539 = n4475 | n27534 ;
  assign n27540 = n27537 | n27539 ;
  assign n27541 = ( ~n22283 & n27538 ) | ( ~n22283 & n27540 ) | ( n27538 & n27540 ) ;
  assign n27542 = n27538 & n27540 ;
  assign n27543 = ( ~n22271 & n27541 ) | ( ~n22271 & n27542 ) | ( n27541 & n27542 ) ;
  assign n27544 = ~x17 & n27543 ;
  assign n27545 = x17 | n27543 ;
  assign n27546 = ( ~n27543 & n27544 ) | ( ~n27543 & n27545 ) | ( n27544 & n27545 ) ;
  assign n27547 = ~n27533 & n27546 ;
  assign n27548 = n27533 | n27547 ;
  assign n27549 = n27533 & n27546 ;
  assign n27550 = n27548 & ~n27549 ;
  assign n27551 = n27305 | n27321 ;
  assign n27552 = ( n27305 & ~n27307 ) | ( n27305 & n27551 ) | ( ~n27307 & n27551 ) ;
  assign n27553 = ~n27550 & n27552 ;
  assign n27554 = n27550 & ~n27552 ;
  assign n27555 = n27553 | n27554 ;
  assign n27572 = n27327 | n27344 ;
  assign n27573 = ( n27327 & ~n27329 ) | ( n27327 & n27572 ) | ( ~n27329 & n27572 ) ;
  assign n27556 = n5234 & ~n23240 ;
  assign n27557 = n5237 & ~n21551 ;
  assign n27558 = n5231 & n23227 ;
  assign n27559 = ( n5231 & n23217 ) | ( n5231 & n27558 ) | ( n23217 & n27558 ) ;
  assign n27560 = n27557 | n27559 ;
  assign n27561 = n27556 | n27560 ;
  assign n27562 = n5227 | n27556 ;
  assign n27563 = n27560 | n27562 ;
  assign n27564 = ( n23260 & n27561 ) | ( n23260 & n27563 ) | ( n27561 & n27563 ) ;
  assign n27565 = x14 & n27563 ;
  assign n27566 = x14 & n27561 ;
  assign n27567 = ( n23260 & n27565 ) | ( n23260 & n27566 ) | ( n27565 & n27566 ) ;
  assign n27568 = x14 & ~n27566 ;
  assign n27569 = x14 & ~n27565 ;
  assign n27570 = ( ~n23260 & n27568 ) | ( ~n23260 & n27569 ) | ( n27568 & n27569 ) ;
  assign n27571 = ( n27564 & ~n27567 ) | ( n27564 & n27570 ) | ( ~n27567 & n27570 ) ;
  assign n27574 = n27571 & n27573 ;
  assign n27575 = n27573 & ~n27574 ;
  assign n27576 = ~n27555 & n27571 ;
  assign n27577 = ~n27573 & n27576 ;
  assign n27578 = ( ~n27555 & n27575 ) | ( ~n27555 & n27577 ) | ( n27575 & n27577 ) ;
  assign n27579 = n27555 & ~n27571 ;
  assign n27580 = ( n27555 & n27573 ) | ( n27555 & n27579 ) | ( n27573 & n27579 ) ;
  assign n27581 = ~n27575 & n27580 ;
  assign n27582 = n27578 | n27581 ;
  assign n27583 = ~n27164 & n27347 ;
  assign n27584 = ( n27164 & n27166 ) | ( n27164 & ~n27583 ) | ( n27166 & ~n27583 ) ;
  assign n27585 = ~n27582 & n27584 ;
  assign n27586 = n27582 & ~n27584 ;
  assign n27587 = n27585 | n27586 ;
  assign n27588 = ~n27353 & n27364 ;
  assign n27589 = n27353 | n27365 ;
  assign n27590 = ( n26516 & ~n27588 ) | ( n26516 & n27589 ) | ( ~n27588 & n27589 ) ;
  assign n27591 = n27353 | n27367 ;
  assign n27592 = ~n27353 & n27355 ;
  assign n27593 = ( n27130 & n27591 ) | ( n27130 & ~n27592 ) | ( n27591 & ~n27592 ) ;
  assign n27594 = ( n26009 & n27590 ) | ( n26009 & n27593 ) | ( n27590 & n27593 ) ;
  assign n27595 = ( n26011 & n27590 ) | ( n26011 & n27593 ) | ( n27590 & n27593 ) ;
  assign n27596 = ( n24765 & n27594 ) | ( n24765 & n27595 ) | ( n27594 & n27595 ) ;
  assign n27597 = n27587 & ~n27596 ;
  assign n27598 = n27587 | n27588 ;
  assign n27599 = ~n27587 & n27589 ;
  assign n27600 = ( n26516 & ~n27598 ) | ( n26516 & n27599 ) | ( ~n27598 & n27599 ) ;
  assign n27601 = ~n27587 & n27591 ;
  assign n27602 = n27587 | n27592 ;
  assign n27603 = ( n27130 & n27601 ) | ( n27130 & ~n27602 ) | ( n27601 & ~n27602 ) ;
  assign n27604 = ( n26009 & n27600 ) | ( n26009 & n27603 ) | ( n27600 & n27603 ) ;
  assign n27605 = ( n26011 & n27600 ) | ( n26011 & n27603 ) | ( n27600 & n27603 ) ;
  assign n27606 = ( n24765 & n27604 ) | ( n24765 & n27605 ) | ( n27604 & n27605 ) ;
  assign n27607 = n4471 & ~n27606 ;
  assign n27608 = ~n27597 & n27607 ;
  assign n27609 = n27374 | n27608 ;
  assign n27610 = n27125 | n27133 ;
  assign n27611 = n27363 | n27371 ;
  assign n27612 = n27610 | n27611 ;
  assign n27613 = n27610 & n27611 ;
  assign n27614 = n27612 & ~n27613 ;
  assign n27615 = n26527 | n27610 ;
  assign n27616 = n26527 & n27610 ;
  assign n27617 = n27615 & ~n27616 ;
  assign n27618 = n26528 & n27615 ;
  assign n27619 = ( n27615 & ~n27617 ) | ( n27615 & n27618 ) | ( ~n27617 & n27618 ) ;
  assign n27620 = n27614 & ~n27619 ;
  assign n27621 = n27615 & ~n27617 ;
  assign n27622 = n27614 & ~n27621 ;
  assign n27623 = ( n26528 & n27620 ) | ( n26528 & n27622 ) | ( n27620 & n27622 ) ;
  assign n27624 = n27620 & n27622 ;
  assign n27625 = ( ~n26538 & n27623 ) | ( ~n26538 & n27624 ) | ( n27623 & n27624 ) ;
  assign n27626 = n27597 | n27606 ;
  assign n27627 = n27611 | n27626 ;
  assign n27628 = n27611 & n27626 ;
  assign n27629 = n27627 & ~n27628 ;
  assign n27630 = n27612 & n27629 ;
  assign n27631 = n4475 & n27630 ;
  assign n27632 = ~n27625 & n27631 ;
  assign n27633 = n27612 | n27629 ;
  assign n27634 = ( ~n27625 & n27629 ) | ( ~n27625 & n27633 ) | ( n27629 & n27633 ) ;
  assign n27635 = ( n4475 & n27632 ) | ( n4475 & ~n27634 ) | ( n27632 & ~n27634 ) ;
  assign n27636 = n27609 | n27635 ;
  assign n27637 = x17 | n27609 ;
  assign n27638 = n27635 | n27637 ;
  assign n27639 = ~x17 & n27637 ;
  assign n27640 = ( ~x17 & n27635 ) | ( ~x17 & n27639 ) | ( n27635 & n27639 ) ;
  assign n27641 = ( ~n27636 & n27638 ) | ( ~n27636 & n27640 ) | ( n27638 & n27640 ) ;
  assign n27642 = ~n26911 & n27641 ;
  assign n27643 = n26911 & ~n27641 ;
  assign n27644 = n27642 | n27643 ;
  assign n27645 = n26592 & n26906 ;
  assign n27646 = n26592 & ~n27645 ;
  assign n27649 = n27619 | n27621 ;
  assign n27650 = ~n27614 & n27649 ;
  assign n27651 = ( ~n26528 & n27619 ) | ( ~n26528 & n27621 ) | ( n27619 & n27621 ) ;
  assign n27652 = ~n27614 & n27651 ;
  assign n27653 = ( n26538 & n27650 ) | ( n26538 & n27652 ) | ( n27650 & n27652 ) ;
  assign n27654 = n27625 | n27653 ;
  assign n27655 = n4466 & ~n26526 ;
  assign n27656 = ~n26520 & n27655 ;
  assign n27657 = n4468 & ~n27133 ;
  assign n27658 = ~n27125 & n27657 ;
  assign n27659 = n27656 | n27658 ;
  assign n27660 = n4471 & ~n27371 ;
  assign n27661 = ~n27363 & n27660 ;
  assign n27662 = n27659 | n27661 ;
  assign n27663 = n4475 | n27661 ;
  assign n27664 = n27659 | n27663 ;
  assign n27665 = ( ~n27654 & n27662 ) | ( ~n27654 & n27664 ) | ( n27662 & n27664 ) ;
  assign n27666 = ~x17 & n27664 ;
  assign n27667 = ~x17 & n27662 ;
  assign n27668 = ( ~n27654 & n27666 ) | ( ~n27654 & n27667 ) | ( n27666 & n27667 ) ;
  assign n27669 = x17 | n27667 ;
  assign n27670 = x17 | n27666 ;
  assign n27671 = ( ~n27654 & n27669 ) | ( ~n27654 & n27670 ) | ( n27669 & n27670 ) ;
  assign n27672 = ( ~n27665 & n27668 ) | ( ~n27665 & n27671 ) | ( n27668 & n27671 ) ;
  assign n27647 = ~n26592 & n26906 ;
  assign n27673 = n27647 & n27672 ;
  assign n27674 = ( n27646 & n27672 ) | ( n27646 & n27673 ) | ( n27672 & n27673 ) ;
  assign n27648 = n27646 | n27647 ;
  assign n27675 = n27648 & ~n27674 ;
  assign n27676 = ~n27647 & n27672 ;
  assign n27677 = ~n27646 & n27676 ;
  assign n27678 = n27675 | n27677 ;
  assign n27679 = ~n26625 & n26904 ;
  assign n27680 = n26625 | n27679 ;
  assign n27683 = n4466 & ~n26270 ;
  assign n27684 = ~n26263 & n27683 ;
  assign n27685 = n4468 & ~n26526 ;
  assign n27686 = ~n26520 & n27685 ;
  assign n27687 = n27684 | n27686 ;
  assign n27688 = n4471 & ~n27133 ;
  assign n27689 = ~n27125 & n27688 ;
  assign n27690 = n27687 | n27689 ;
  assign n27691 = n26528 & n26538 ;
  assign n27692 = ~n26528 & n27617 ;
  assign n27693 = ( n26528 & n27617 ) | ( n26528 & n27692 ) | ( n27617 & n27692 ) ;
  assign n27694 = n27617 & n27692 ;
  assign n27695 = ( ~n26538 & n27693 ) | ( ~n26538 & n27694 ) | ( n27693 & n27694 ) ;
  assign n27696 = n27691 | n27695 ;
  assign n27697 = ~n27616 & n27619 ;
  assign n27698 = ~n26528 & n27697 ;
  assign n27699 = ( n26538 & n27697 ) | ( n26538 & n27698 ) | ( n27697 & n27698 ) ;
  assign n27700 = n4475 & n27699 ;
  assign n27701 = ( n4475 & ~n27696 ) | ( n4475 & n27700 ) | ( ~n27696 & n27700 ) ;
  assign n27702 = n27690 | n27701 ;
  assign n27703 = x17 | n27690 ;
  assign n27704 = n27701 | n27703 ;
  assign n27705 = ~x17 & n27703 ;
  assign n27706 = ( ~x17 & n27701 ) | ( ~x17 & n27705 ) | ( n27701 & n27705 ) ;
  assign n27707 = ( ~n27702 & n27704 ) | ( ~n27702 & n27706 ) | ( n27704 & n27706 ) ;
  assign n27681 = n26625 & n26904 ;
  assign n27708 = n27681 & n27707 ;
  assign n27709 = ( ~n27680 & n27707 ) | ( ~n27680 & n27708 ) | ( n27707 & n27708 ) ;
  assign n27682 = n27680 & ~n27681 ;
  assign n27710 = n27682 | n27709 ;
  assign n27711 = ~n27681 & n27707 ;
  assign n27712 = n27680 & n27711 ;
  assign n27713 = n27710 & ~n27712 ;
  assign n27714 = n26902 & ~n26903 ;
  assign n27715 = n26646 | n26903 ;
  assign n27716 = ~n27714 & n27715 ;
  assign n27717 = n4466 & n26017 ;
  assign n27718 = n4468 & ~n26270 ;
  assign n27719 = ~n26263 & n27718 ;
  assign n27720 = n27717 | n27719 ;
  assign n27721 = n4471 & ~n26526 ;
  assign n27722 = ~n26520 & n27721 ;
  assign n27723 = n27720 | n27722 ;
  assign n27724 = n4475 | n27722 ;
  assign n27725 = n27720 | n27724 ;
  assign n27726 = ( ~n26555 & n27723 ) | ( ~n26555 & n27725 ) | ( n27723 & n27725 ) ;
  assign n27727 = ( n26528 & n27723 ) | ( n26528 & n27725 ) | ( n27723 & n27725 ) ;
  assign n27728 = ( ~n26543 & n27726 ) | ( ~n26543 & n27727 ) | ( n27726 & n27727 ) ;
  assign n27729 = ~x17 & n27728 ;
  assign n27730 = x17 | n27728 ;
  assign n27731 = ( ~n27728 & n27729 ) | ( ~n27728 & n27730 ) | ( n27729 & n27730 ) ;
  assign n27732 = n27716 & n27731 ;
  assign n27733 = n26898 & n26900 ;
  assign n27734 = n26898 | n26900 ;
  assign n27735 = ~n27733 & n27734 ;
  assign n27736 = n4466 & ~n25728 ;
  assign n27737 = n4468 & n26017 ;
  assign n27738 = n27736 | n27737 ;
  assign n27739 = n4471 & ~n26270 ;
  assign n27740 = ~n26263 & n27739 ;
  assign n27742 = n4475 | n27740 ;
  assign n27743 = n27738 | n27742 ;
  assign n27741 = n27738 | n27740 ;
  assign n27744 = n27741 & n27743 ;
  assign n27745 = ( n26571 & n27743 ) | ( n26571 & n27744 ) | ( n27743 & n27744 ) ;
  assign n27746 = x17 & n27744 ;
  assign n27747 = x17 & n27743 ;
  assign n27748 = ( n26571 & n27746 ) | ( n26571 & n27747 ) | ( n27746 & n27747 ) ;
  assign n27749 = x17 & ~n27746 ;
  assign n27750 = x17 & ~n27747 ;
  assign n27751 = ( ~n26571 & n27749 ) | ( ~n26571 & n27750 ) | ( n27749 & n27750 ) ;
  assign n27752 = ( n27745 & ~n27748 ) | ( n27745 & n27751 ) | ( ~n27748 & n27751 ) ;
  assign n27753 = n27735 & n27752 ;
  assign n27754 = n26686 & n26896 ;
  assign n27755 = n26686 | n26896 ;
  assign n27756 = ~n27754 & n27755 ;
  assign n27757 = n4471 & n26017 ;
  assign n27758 = n4466 & ~n25046 ;
  assign n27759 = n4468 & ~n25728 ;
  assign n27760 = n27758 | n27759 ;
  assign n27761 = n27757 | n27760 ;
  assign n27762 = n4475 | n27757 ;
  assign n27763 = n27760 | n27762 ;
  assign n27764 = ( n26613 & n27761 ) | ( n26613 & n27763 ) | ( n27761 & n27763 ) ;
  assign n27765 = n27761 | n27763 ;
  assign n27766 = ( n26605 & n27764 ) | ( n26605 & n27765 ) | ( n27764 & n27765 ) ;
  assign n27767 = x17 & n27766 ;
  assign n27768 = x17 & ~n27766 ;
  assign n27769 = ( n27766 & ~n27767 ) | ( n27766 & n27768 ) | ( ~n27767 & n27768 ) ;
  assign n27770 = n27756 & n27769 ;
  assign n27771 = n27756 & ~n27770 ;
  assign n27772 = ~n27756 & n27769 ;
  assign n27773 = n27771 | n27772 ;
  assign n27774 = ( n26722 & n26723 ) | ( n26722 & n26894 ) | ( n26723 & n26894 ) ;
  assign n27775 = n26701 | n26722 ;
  assign n27776 = n26894 | n27775 ;
  assign n27777 = ~n27774 & n27776 ;
  assign n27778 = n4471 & ~n25728 ;
  assign n27779 = n4466 & n24770 ;
  assign n27780 = n4468 & ~n25046 ;
  assign n27781 = n27779 | n27780 ;
  assign n27782 = n27778 | n27781 ;
  assign n27783 = n4475 & n25740 ;
  assign n27784 = n4475 & n25731 ;
  assign n27785 = ( ~n25441 & n27783 ) | ( ~n25441 & n27784 ) | ( n27783 & n27784 ) ;
  assign n27786 = n27782 | n27785 ;
  assign n27787 = n4475 | n27782 ;
  assign n27788 = ( n25733 & n27786 ) | ( n25733 & n27787 ) | ( n27786 & n27787 ) ;
  assign n27789 = x17 | n27788 ;
  assign n27790 = ~x17 & n27788 ;
  assign n27791 = ( ~n27788 & n27789 ) | ( ~n27788 & n27790 ) | ( n27789 & n27790 ) ;
  assign n27792 = n27777 & n27791 ;
  assign n27793 = n26891 & ~n26894 ;
  assign n27796 = n4471 & ~n25046 ;
  assign n27797 = n4466 & ~n25054 ;
  assign n27798 = n4468 & n24770 ;
  assign n27799 = n27797 | n27798 ;
  assign n27800 = n27796 | n27799 ;
  assign n27801 = n4475 | n27796 ;
  assign n27802 = n27799 | n27801 ;
  assign n27803 = ( ~n25069 & n27800 ) | ( ~n25069 & n27802 ) | ( n27800 & n27802 ) ;
  assign n27804 = ~x17 & n27802 ;
  assign n27805 = ~x17 & n27800 ;
  assign n27806 = ( ~n25069 & n27804 ) | ( ~n25069 & n27805 ) | ( n27804 & n27805 ) ;
  assign n27807 = x17 | n27805 ;
  assign n27808 = x17 | n27804 ;
  assign n27809 = ( ~n25069 & n27807 ) | ( ~n25069 & n27808 ) | ( n27807 & n27808 ) ;
  assign n27810 = ( ~n27803 & n27806 ) | ( ~n27803 & n27809 ) | ( n27806 & n27809 ) ;
  assign n27794 = ~n26891 & n26893 ;
  assign n27811 = n27794 & n27810 ;
  assign n27812 = ( n27793 & n27810 ) | ( n27793 & n27811 ) | ( n27810 & n27811 ) ;
  assign n27795 = n27793 | n27794 ;
  assign n27813 = n27795 & ~n27812 ;
  assign n27814 = ~n27794 & n27810 ;
  assign n27815 = ~n27793 & n27814 ;
  assign n27816 = n27813 | n27815 ;
  assign n27817 = n26889 & ~n26890 ;
  assign n27818 = n26746 & ~n26890 ;
  assign n27819 = n27817 | n27818 ;
  assign n27820 = n4471 & n24770 ;
  assign n27821 = n4466 & n24167 ;
  assign n27822 = n4468 & ~n25054 ;
  assign n27823 = n27821 | n27822 ;
  assign n27824 = n27820 | n27823 ;
  assign n27825 = n4475 | n27824 ;
  assign n27826 = ( ~n25095 & n27824 ) | ( ~n25095 & n27825 ) | ( n27824 & n27825 ) ;
  assign n27827 = ~x17 & n27825 ;
  assign n27828 = ~x17 & n27824 ;
  assign n27829 = ( ~n25095 & n27827 ) | ( ~n25095 & n27828 ) | ( n27827 & n27828 ) ;
  assign n27830 = x17 | n27827 ;
  assign n27831 = x17 | n27828 ;
  assign n27832 = ( ~n25095 & n27830 ) | ( ~n25095 & n27831 ) | ( n27830 & n27831 ) ;
  assign n27833 = ( ~n27826 & n27829 ) | ( ~n27826 & n27832 ) | ( n27829 & n27832 ) ;
  assign n27834 = n27819 & n27833 ;
  assign n27835 = n27819 & ~n27834 ;
  assign n27836 = ~n27819 & n27833 ;
  assign n27837 = n27835 | n27836 ;
  assign n27838 = n26768 | n26862 ;
  assign n27839 = ~n26863 & n27838 ;
  assign n27840 = n4471 & n24167 ;
  assign n27841 = n4466 & n23316 ;
  assign n27842 = n4468 & n23614 ;
  assign n27843 = n27841 | n27842 ;
  assign n27844 = n27840 | n27843 ;
  assign n27845 = n4475 | n27844 ;
  assign n27846 = ( n24182 & n27844 ) | ( n24182 & n27845 ) | ( n27844 & n27845 ) ;
  assign n27847 = n27844 | n27845 ;
  assign n27848 = ( n24175 & n27846 ) | ( n24175 & n27847 ) | ( n27846 & n27847 ) ;
  assign n27849 = x17 & n27848 ;
  assign n27850 = x17 & ~n27848 ;
  assign n27851 = ( n27848 & ~n27849 ) | ( n27848 & n27850 ) | ( ~n27849 & n27850 ) ;
  assign n27852 = n27839 & n27851 ;
  assign n27853 = n26864 & n26887 ;
  assign n27854 = n26864 | n26887 ;
  assign n27855 = ~n27853 & n27854 ;
  assign n27856 = n4471 & ~n25054 ;
  assign n27857 = n4466 & n23614 ;
  assign n27858 = n4468 & n24167 ;
  assign n27859 = n27857 | n27858 ;
  assign n27860 = n27856 | n27859 ;
  assign n27861 = n4475 | n27856 ;
  assign n27862 = n27859 | n27861 ;
  assign n27863 = ( ~n25122 & n27860 ) | ( ~n25122 & n27862 ) | ( n27860 & n27862 ) ;
  assign n27864 = ~x17 & n27862 ;
  assign n27865 = ~x17 & n27860 ;
  assign n27866 = ( ~n25122 & n27864 ) | ( ~n25122 & n27865 ) | ( n27864 & n27865 ) ;
  assign n27867 = x17 | n27865 ;
  assign n27868 = x17 | n27864 ;
  assign n27869 = ( ~n25122 & n27867 ) | ( ~n25122 & n27868 ) | ( n27867 & n27868 ) ;
  assign n27870 = ( ~n27863 & n27866 ) | ( ~n27863 & n27869 ) | ( n27866 & n27869 ) ;
  assign n27871 = n27855 & n27870 ;
  assign n27872 = n27855 | n27870 ;
  assign n27873 = ~n27871 & n27872 ;
  assign n27874 = n27852 & n27873 ;
  assign n27875 = n27871 | n27873 ;
  assign n27876 = n26787 | n26860 ;
  assign n27877 = ~n26861 & n27876 ;
  assign n27878 = n4471 & n23614 ;
  assign n27879 = n4466 & n23620 ;
  assign n27880 = ( n4468 & n4503 ) | ( n4468 & n23620 ) | ( n4503 & n23620 ) ;
  assign n27881 = ( n23316 & n27879 ) | ( n23316 & n27880 ) | ( n27879 & n27880 ) ;
  assign n27883 = n4475 | n27881 ;
  assign n27884 = n27878 | n27883 ;
  assign n27882 = n27878 | n27881 ;
  assign n27885 = n27882 & n27884 ;
  assign n27886 = ( n23634 & n27884 ) | ( n23634 & n27885 ) | ( n27884 & n27885 ) ;
  assign n27887 = x17 & n27885 ;
  assign n27888 = x17 & n27884 ;
  assign n27889 = ( n23634 & n27887 ) | ( n23634 & n27888 ) | ( n27887 & n27888 ) ;
  assign n27890 = x17 & ~n27887 ;
  assign n27891 = x17 & ~n27888 ;
  assign n27892 = ( ~n23634 & n27890 ) | ( ~n23634 & n27891 ) | ( n27890 & n27891 ) ;
  assign n27893 = ( n27886 & ~n27889 ) | ( n27886 & n27892 ) | ( ~n27889 & n27892 ) ;
  assign n27894 = n27877 & n27893 ;
  assign n27895 = n27877 & ~n27894 ;
  assign n27896 = ~n27877 & n27893 ;
  assign n27897 = n27895 | n27896 ;
  assign n27898 = n26840 & n26854 ;
  assign n27899 = n26840 & ~n27898 ;
  assign n27900 = n4466 & ~n22385 ;
  assign n27901 = ( n4468 & n4503 ) | ( n4468 & ~n22385 ) | ( n4503 & ~n22385 ) ;
  assign n27902 = ( n22381 & n27900 ) | ( n22381 & n27901 ) | ( n27900 & n27901 ) ;
  assign n27903 = n4471 | n27902 ;
  assign n27904 = ( n23620 & n27902 ) | ( n23620 & n27903 ) | ( n27902 & n27903 ) ;
  assign n27905 = n4475 | n27904 ;
  assign n27906 = ( ~n23686 & n27904 ) | ( ~n23686 & n27905 ) | ( n27904 & n27905 ) ;
  assign n27907 = ~x17 & n27905 ;
  assign n27908 = ~x17 & n27904 ;
  assign n27909 = ( ~n23686 & n27907 ) | ( ~n23686 & n27908 ) | ( n27907 & n27908 ) ;
  assign n27910 = x17 | n27907 ;
  assign n27911 = x17 | n27908 ;
  assign n27912 = ( ~n23686 & n27910 ) | ( ~n23686 & n27911 ) | ( n27910 & n27911 ) ;
  assign n27913 = ( ~n27906 & n27909 ) | ( ~n27906 & n27912 ) | ( n27909 & n27912 ) ;
  assign n27914 = ~n26840 & n26854 ;
  assign n27915 = n27913 & n27914 ;
  assign n27916 = ( n27899 & n27913 ) | ( n27899 & n27915 ) | ( n27913 & n27915 ) ;
  assign n27917 = n27913 | n27914 ;
  assign n27918 = n27899 | n27917 ;
  assign n27919 = ~n27916 & n27918 ;
  assign n27920 = n26819 & n26837 ;
  assign n27921 = n26819 | n26837 ;
  assign n27922 = ~n27920 & n27921 ;
  assign n27923 = n4471 & n22381 ;
  assign n27924 = n4466 & ~n22398 ;
  assign n27925 = n4468 & ~n22385 ;
  assign n27926 = n27924 | n27925 ;
  assign n27927 = n27923 | n27926 ;
  assign n27928 = n4475 | n27927 ;
  assign n27929 = x17 & n27928 ;
  assign n27930 = x17 & n27927 ;
  assign n27931 = ( n22422 & n27929 ) | ( n22422 & n27930 ) | ( n27929 & n27930 ) ;
  assign n27932 = x17 | n27928 ;
  assign n27933 = x17 | n27927 ;
  assign n27934 = ( n22422 & n27932 ) | ( n22422 & n27933 ) | ( n27932 & n27933 ) ;
  assign n27935 = ~n27931 & n27934 ;
  assign n27936 = n27922 & n27935 ;
  assign n27937 = ~n27922 & n27935 ;
  assign n27938 = ( n27922 & ~n27936 ) | ( n27922 & n27937 ) | ( ~n27936 & n27937 ) ;
  assign n27939 = n26813 | n26815 ;
  assign n27940 = ~n26815 & n26817 ;
  assign n27941 = ( n26814 & n27939 ) | ( n26814 & ~n27940 ) | ( n27939 & ~n27940 ) ;
  assign n27942 = ~n26819 & n27941 ;
  assign n27943 = n4471 & ~n22385 ;
  assign n27944 = n4466 & n22393 ;
  assign n27945 = n4468 & ~n22398 ;
  assign n27946 = n27944 | n27945 ;
  assign n27947 = n27943 | n27946 ;
  assign n27948 = n4475 | n27943 ;
  assign n27949 = n27946 | n27948 ;
  assign n27950 = ( ~n22545 & n27947 ) | ( ~n22545 & n27949 ) | ( n27947 & n27949 ) ;
  assign n27951 = ~x17 & n27949 ;
  assign n27952 = ~x17 & n27947 ;
  assign n27953 = ( ~n22545 & n27951 ) | ( ~n22545 & n27952 ) | ( n27951 & n27952 ) ;
  assign n27954 = x17 | n27952 ;
  assign n27955 = x17 | n27951 ;
  assign n27956 = ( ~n22545 & n27954 ) | ( ~n22545 & n27955 ) | ( n27954 & n27955 ) ;
  assign n27957 = ( ~n27950 & n27953 ) | ( ~n27950 & n27956 ) | ( n27953 & n27956 ) ;
  assign n27958 = n27942 & n27957 ;
  assign n27959 = n4475 & n22474 ;
  assign n27960 = n4468 & ~n22409 ;
  assign n27961 = n4471 & ~n22406 ;
  assign n27962 = n27960 | n27961 ;
  assign n27963 = x17 | n27962 ;
  assign n27964 = n27959 | n27963 ;
  assign n27965 = ~x17 & n27964 ;
  assign n27966 = ( x17 & n16481 ) | ( x17 & n22409 ) | ( n16481 & n22409 ) ;
  assign n27967 = n27964 & n27966 ;
  assign n27968 = n27959 | n27962 ;
  assign n27969 = n27966 & ~n27968 ;
  assign n27970 = ( n27965 & n27967 ) | ( n27965 & n27969 ) | ( n27967 & n27969 ) ;
  assign n27971 = n4471 & n22393 ;
  assign n27972 = n4466 & ~n22409 ;
  assign n27973 = n4468 & ~n22406 ;
  assign n27974 = n27972 | n27973 ;
  assign n27975 = n27971 | n27974 ;
  assign n27976 = n22439 | n27975 ;
  assign n27977 = n4475 | n27971 ;
  assign n27978 = n27974 | n27977 ;
  assign n27979 = ~x17 & n27978 ;
  assign n27980 = n27976 & n27979 ;
  assign n27981 = x17 | n27980 ;
  assign n27982 = n3536 & ~n22409 ;
  assign n27983 = n27980 & n27982 ;
  assign n27984 = n27976 & n27978 ;
  assign n27985 = n27982 & ~n27984 ;
  assign n27986 = ( n27981 & n27983 ) | ( n27981 & n27985 ) | ( n27983 & n27985 ) ;
  assign n27987 = n27970 & n27986 ;
  assign n27988 = ( n27980 & n27981 ) | ( n27980 & ~n27984 ) | ( n27981 & ~n27984 ) ;
  assign n27989 = n27970 | n27982 ;
  assign n27990 = ( n27982 & n27988 ) | ( n27982 & n27989 ) | ( n27988 & n27989 ) ;
  assign n27991 = ~n27987 & n27990 ;
  assign n27992 = n4466 & ~n22406 ;
  assign n27993 = n4468 & n22393 ;
  assign n27994 = n27992 | n27993 ;
  assign n27995 = n4471 & ~n22398 ;
  assign n27996 = n4475 | n27995 ;
  assign n27997 = n27994 | n27996 ;
  assign n27998 = x17 & n27997 ;
  assign n27999 = n27994 | n27995 ;
  assign n28000 = x17 & n27999 ;
  assign n28001 = ( n22608 & n27998 ) | ( n22608 & n28000 ) | ( n27998 & n28000 ) ;
  assign n28002 = x17 | n27997 ;
  assign n28003 = x17 | n27999 ;
  assign n28004 = ( n22608 & n28002 ) | ( n22608 & n28003 ) | ( n28002 & n28003 ) ;
  assign n28005 = ~n28001 & n28004 ;
  assign n28006 = n27987 | n28005 ;
  assign n28007 = ( n27987 & n27991 ) | ( n27987 & n28006 ) | ( n27991 & n28006 ) ;
  assign n28008 = n27942 | n27957 ;
  assign n28009 = ~n27958 & n28008 ;
  assign n28010 = n27958 | n28009 ;
  assign n28011 = ( n27958 & n28007 ) | ( n27958 & n28010 ) | ( n28007 & n28010 ) ;
  assign n28012 = n27938 & n28011 ;
  assign n28013 = n27936 | n28012 ;
  assign n28014 = n27919 & n28013 ;
  assign n28015 = n27916 | n28014 ;
  assign n28016 = n4466 & n22381 ;
  assign n28017 = ( n4468 & n4503 ) | ( n4468 & n22381 ) | ( n4503 & n22381 ) ;
  assign n28018 = ( n23620 & n28016 ) | ( n23620 & n28017 ) | ( n28016 & n28017 ) ;
  assign n28019 = n4471 | n28017 ;
  assign n28020 = n4471 | n28016 ;
  assign n28021 = ( n23620 & n28019 ) | ( n23620 & n28020 ) | ( n28019 & n28020 ) ;
  assign n28022 = ( n23316 & n28018 ) | ( n23316 & n28021 ) | ( n28018 & n28021 ) ;
  assign n28023 = n4475 | n28022 ;
  assign n28024 = ~x17 & n28023 ;
  assign n28025 = ~x17 & n28022 ;
  assign n28026 = ( n23661 & n28024 ) | ( n23661 & n28025 ) | ( n28024 & n28025 ) ;
  assign n28027 = ( x17 & n16441 ) | ( x17 & n28022 ) | ( n16441 & n28022 ) ;
  assign n28028 = x17 & ~n28027 ;
  assign n28029 = x17 & n28022 ;
  assign n28030 = x17 & ~n28029 ;
  assign n28031 = ( ~n23661 & n28028 ) | ( ~n23661 & n28030 ) | ( n28028 & n28030 ) ;
  assign n28032 = n28026 | n28031 ;
  assign n28033 = n26856 & n26858 ;
  assign n28034 = n26856 | n26858 ;
  assign n28035 = ~n28033 & n28034 ;
  assign n28036 = n28032 & n28035 ;
  assign n28037 = n28032 | n28035 ;
  assign n28038 = ~n28036 & n28037 ;
  assign n28039 = n28036 | n28038 ;
  assign n28040 = ( n28015 & n28036 ) | ( n28015 & n28039 ) | ( n28036 & n28039 ) ;
  assign n28041 = n27897 & n28040 ;
  assign n28042 = n27894 | n28041 ;
  assign n28043 = ~n27839 & n27851 ;
  assign n28044 = ( n27839 & ~n27852 ) | ( n27839 & n28043 ) | ( ~n27852 & n28043 ) ;
  assign n28045 = n28042 & n28044 ;
  assign n28046 = n27871 | n28045 ;
  assign n28047 = ( n27874 & n27875 ) | ( n27874 & n28046 ) | ( n27875 & n28046 ) ;
  assign n28048 = n27834 | n28047 ;
  assign n28049 = ( n27834 & n27837 ) | ( n27834 & n28048 ) | ( n27837 & n28048 ) ;
  assign n28050 = n27816 & n28049 ;
  assign n28051 = n27812 | n28050 ;
  assign n28052 = ~n27777 & n27791 ;
  assign n28053 = ( n27777 & ~n27792 ) | ( n27777 & n28052 ) | ( ~n27792 & n28052 ) ;
  assign n28054 = n27792 | n28053 ;
  assign n28055 = ( n27792 & n28051 ) | ( n27792 & n28054 ) | ( n28051 & n28054 ) ;
  assign n28056 = n27770 | n28055 ;
  assign n28057 = ( n27770 & n27773 ) | ( n27770 & n28056 ) | ( n27773 & n28056 ) ;
  assign n28058 = n27735 | n27752 ;
  assign n28059 = ~n27753 & n28058 ;
  assign n28060 = n27753 | n28059 ;
  assign n28061 = ( n27753 & n28057 ) | ( n27753 & n28060 ) | ( n28057 & n28060 ) ;
  assign n28062 = n27732 & n28061 ;
  assign n28063 = ~n27716 & n27731 ;
  assign n28064 = n28061 | n28063 ;
  assign n28065 = n27716 | n28063 ;
  assign n28066 = ~n28063 & n28065 ;
  assign n28067 = ( n28062 & n28064 ) | ( n28062 & ~n28066 ) | ( n28064 & ~n28066 ) ;
  assign n28068 = n27709 | n28067 ;
  assign n28069 = ( n27709 & ~n27713 ) | ( n27709 & n28068 ) | ( ~n27713 & n28068 ) ;
  assign n28070 = n27674 | n28069 ;
  assign n28071 = ( n27674 & n27678 ) | ( n27674 & n28070 ) | ( n27678 & n28070 ) ;
  assign n28072 = n27644 & ~n28071 ;
  assign n28073 = ~n27644 & n28071 ;
  assign n28074 = n28072 | n28073 ;
  assign n28075 = n5231 | n5234 ;
  assign n28076 = ~n23234 & n28075 ;
  assign n28077 = n5237 | n28076 ;
  assign n28078 = ~n23235 & n28075 ;
  assign n28079 = n5237 | n28078 ;
  assign n28080 = ( ~n15882 & n28077 ) | ( ~n15882 & n28079 ) | ( n28077 & n28079 ) ;
  assign n28081 = n5227 | n28080 ;
  assign n28082 = ( ~n15882 & n28076 ) | ( ~n15882 & n28078 ) | ( n28076 & n28078 ) ;
  assign n28083 = n5227 | n28082 ;
  assign n28084 = ( ~n23240 & n28081 ) | ( ~n23240 & n28083 ) | ( n28081 & n28083 ) ;
  assign n28085 = ( ~n23240 & n28080 ) | ( ~n23240 & n28082 ) | ( n28080 & n28082 ) ;
  assign n28086 = n24135 & ~n28085 ;
  assign n28087 = n23240 & ~n28085 ;
  assign n28088 = ( n23575 & n28086 ) | ( n23575 & n28087 ) | ( n28086 & n28087 ) ;
  assign n28089 = ( n23577 & n28086 ) | ( n23577 & n28087 ) | ( n28086 & n28087 ) ;
  assign n28090 = ( ~n21554 & n28088 ) | ( ~n21554 & n28089 ) | ( n28088 & n28089 ) ;
  assign n28091 = n28084 & ~n28090 ;
  assign n28092 = x14 & ~n28091 ;
  assign n28093 = n28088 | n28089 ;
  assign n28094 = n28084 & ~n28093 ;
  assign n28095 = x14 & ~n28094 ;
  assign n28096 = ( n21584 & n28092 ) | ( n21584 & n28095 ) | ( n28092 & n28095 ) ;
  assign n28097 = ~x14 & n28091 ;
  assign n28098 = ~x14 & n28094 ;
  assign n28099 = ( ~n21584 & n28097 ) | ( ~n21584 & n28098 ) | ( n28097 & n28098 ) ;
  assign n28100 = n28096 | n28099 ;
  assign n28101 = n27502 | n27508 ;
  assign n28102 = n27477 | n27483 ;
  assign n28103 = n27427 | n27434 ;
  assign n28104 = n848 | n8052 ;
  assign n28105 = n7010 | n28104 ;
  assign n28106 = n289 | n333 ;
  assign n28107 = n735 | n28106 ;
  assign n28108 = n13834 | n28107 ;
  assign n28109 = n13005 | n28108 ;
  assign n28110 = n13843 | n28109 ;
  assign n28111 = n13831 | n28110 ;
  assign n28112 = n28105 | n28111 ;
  assign n28113 = n448 | n527 ;
  assign n28114 = n886 | n28113 ;
  assign n28115 = n3983 | n4374 ;
  assign n28116 = n4371 | n28115 ;
  assign n28117 = n124 | n387 ;
  assign n28118 = n1039 | n28117 ;
  assign n28119 = n5157 | n28118 ;
  assign n28120 = n28116 | n28119 ;
  assign n28121 = n28114 | n28120 ;
  assign n28122 = n28112 | n28121 ;
  assign n28123 = ( n27396 & ~n27398 ) | ( n27396 & n28122 ) | ( ~n27398 & n28122 ) ;
  assign n28124 = n27396 | n28122 ;
  assign n28125 = ( n27415 & n28123 ) | ( n27415 & n28124 ) | ( n28123 & n28124 ) ;
  assign n28126 = n27396 & ~n27398 ;
  assign n28127 = n28122 & n28126 ;
  assign n28128 = n27396 & n28122 ;
  assign n28129 = ( n27415 & n28127 ) | ( n27415 & n28128 ) | ( n28127 & n28128 ) ;
  assign n28130 = n28125 & ~n28129 ;
  assign n28131 = n1057 & n17111 ;
  assign n28132 = n1065 & ~n16069 ;
  assign n28133 = n1060 & n15886 ;
  assign n28134 = n28132 | n28133 ;
  assign n28135 = n28131 | n28134 ;
  assign n28136 = n28130 & n28135 ;
  assign n28137 = n1062 & ~n17194 ;
  assign n28138 = ~n17129 & n28137 ;
  assign n28139 = ( n28130 & n28136 ) | ( n28130 & n28138 ) | ( n28136 & n28138 ) ;
  assign n28140 = ( n1062 & n28130 ) | ( n1062 & n28136 ) | ( n28130 & n28136 ) ;
  assign n28141 = ( n17186 & n28139 ) | ( n17186 & n28140 ) | ( n28139 & n28140 ) ;
  assign n28142 = n28130 | n28135 ;
  assign n28143 = n28138 | n28142 ;
  assign n28144 = n1062 | n28142 ;
  assign n28145 = ( n17186 & n28143 ) | ( n17186 & n28144 ) | ( n28143 & n28144 ) ;
  assign n28146 = ~n28141 & n28145 ;
  assign n28147 = n28103 & n28146 ;
  assign n28148 = n28103 | n28146 ;
  assign n28149 = ~n28147 & n28148 ;
  assign n28151 = n1826 & n17100 ;
  assign n28152 = n1823 & ~n17092 ;
  assign n28153 = n28151 | n28152 ;
  assign n28150 = n1829 & n18037 ;
  assign n28155 = n1821 | n28150 ;
  assign n28156 = n28153 | n28155 ;
  assign n28154 = n28150 | n28153 ;
  assign n28157 = n28154 & n28156 ;
  assign n28158 = ( ~n18050 & n28156 ) | ( ~n18050 & n28157 ) | ( n28156 & n28157 ) ;
  assign n28159 = ~x29 & n28157 ;
  assign n28160 = ~x29 & n28156 ;
  assign n28161 = ( ~n18050 & n28159 ) | ( ~n18050 & n28160 ) | ( n28159 & n28160 ) ;
  assign n28162 = x29 | n28159 ;
  assign n28163 = x29 | n28160 ;
  assign n28164 = ( ~n18050 & n28162 ) | ( ~n18050 & n28163 ) | ( n28162 & n28163 ) ;
  assign n28165 = ( ~n28158 & n28161 ) | ( ~n28158 & n28164 ) | ( n28161 & n28164 ) ;
  assign n28166 = n28149 & n28165 ;
  assign n28167 = n28149 | n28165 ;
  assign n28168 = ~n28166 & n28167 ;
  assign n28169 = n27439 & n28168 ;
  assign n28170 = ( n27459 & n28168 ) | ( n27459 & n28169 ) | ( n28168 & n28169 ) ;
  assign n28171 = n27439 | n28168 ;
  assign n28172 = n27459 | n28171 ;
  assign n28173 = ~n28170 & n28172 ;
  assign n28174 = n2315 & n18576 ;
  assign n28175 = n2312 & ~n18585 ;
  assign n28176 = n2308 & n18410 ;
  assign n28177 = n28175 | n28176 ;
  assign n28178 = n28174 | n28177 ;
  assign n28179 = n2306 | n28174 ;
  assign n28180 = n28177 | n28179 ;
  assign n28181 = ( n18612 & n28178 ) | ( n18612 & n28180 ) | ( n28178 & n28180 ) ;
  assign n28182 = x26 & n28180 ;
  assign n28183 = x26 & n28178 ;
  assign n28184 = ( n18612 & n28182 ) | ( n18612 & n28183 ) | ( n28182 & n28183 ) ;
  assign n28185 = x26 & ~n28183 ;
  assign n28186 = x26 & ~n28182 ;
  assign n28187 = ( ~n18612 & n28185 ) | ( ~n18612 & n28186 ) | ( n28185 & n28186 ) ;
  assign n28188 = ( n28181 & ~n28184 ) | ( n28181 & n28187 ) | ( ~n28184 & n28187 ) ;
  assign n28189 = n28173 & ~n28188 ;
  assign n28190 = n28173 | n28188 ;
  assign n28191 = ( ~n28173 & n28189 ) | ( ~n28173 & n28190 ) | ( n28189 & n28190 ) ;
  assign n28192 = n28102 & n28191 ;
  assign n28193 = n28102 | n28191 ;
  assign n28194 = ~n28192 & n28193 ;
  assign n28195 = n2932 & n19631 ;
  assign n28196 = n2925 & n19352 ;
  assign n28197 = n2928 & n19494 ;
  assign n28198 = n28196 | n28197 ;
  assign n28199 = n28195 | n28198 ;
  assign n28200 = n2936 & n19652 ;
  assign n28201 = n2936 & n19655 ;
  assign n28202 = ( ~n18604 & n28200 ) | ( ~n18604 & n28201 ) | ( n28200 & n28201 ) ;
  assign n28203 = n28199 | n28202 ;
  assign n28204 = n2936 | n28199 ;
  assign n28205 = ( n19640 & n28203 ) | ( n19640 & n28204 ) | ( n28203 & n28204 ) ;
  assign n28206 = x23 | n28205 ;
  assign n28207 = ~x23 & n28205 ;
  assign n28208 = ( ~n28205 & n28206 ) | ( ~n28205 & n28207 ) | ( n28206 & n28207 ) ;
  assign n28209 = n28194 & ~n28208 ;
  assign n28210 = n28194 | n28208 ;
  assign n28211 = ( ~n28194 & n28209 ) | ( ~n28194 & n28210 ) | ( n28209 & n28210 ) ;
  assign n28212 = n28101 & n28211 ;
  assign n28213 = n28101 | n28211 ;
  assign n28214 = ~n28212 & n28213 ;
  assign n28215 = n3547 & n20609 ;
  assign n28216 = n3544 & ~n20630 ;
  assign n28217 = n3541 & ~n20618 ;
  assign n28218 = n28216 | n28217 ;
  assign n28219 = n28215 | n28218 ;
  assign n28220 = n3537 | n28215 ;
  assign n28221 = n28218 | n28220 ;
  assign n28222 = ( n20659 & n28219 ) | ( n20659 & n28221 ) | ( n28219 & n28221 ) ;
  assign n28223 = n28219 & n28221 ;
  assign n28224 = ( ~n20649 & n28222 ) | ( ~n20649 & n28223 ) | ( n28222 & n28223 ) ;
  assign n28225 = x20 & n28224 ;
  assign n28226 = x20 & ~n28224 ;
  assign n28227 = ( n28224 & ~n28225 ) | ( n28224 & n28226 ) | ( ~n28225 & n28226 ) ;
  assign n28228 = n28214 & n28227 ;
  assign n28229 = n28214 & ~n28228 ;
  assign n28231 = n27524 | n27528 ;
  assign n28232 = ~n27524 & n27525 ;
  assign n28233 = ( n27529 & n28231 ) | ( n27529 & ~n28232 ) | ( n28231 & ~n28232 ) ;
  assign n28230 = ~n28214 & n28227 ;
  assign n28234 = n28230 & n28233 ;
  assign n28235 = ( n28229 & n28233 ) | ( n28229 & n28234 ) | ( n28233 & n28234 ) ;
  assign n28236 = n28230 | n28233 ;
  assign n28237 = n28229 | n28236 ;
  assign n28238 = ~n28235 & n28237 ;
  assign n28239 = n4471 & ~n21551 ;
  assign n28240 = n4466 & ~n21563 ;
  assign n28241 = n4468 & ~n21517 ;
  assign n28242 = n28240 | n28241 ;
  assign n28243 = n28239 | n28242 ;
  assign n28244 = n4475 | n28239 ;
  assign n28245 = n28242 | n28244 ;
  assign n28246 = ( ~n21587 & n28243 ) | ( ~n21587 & n28245 ) | ( n28243 & n28245 ) ;
  assign n28247 = ~x17 & n28245 ;
  assign n28248 = ~x17 & n28243 ;
  assign n28249 = ( ~n21587 & n28247 ) | ( ~n21587 & n28248 ) | ( n28247 & n28248 ) ;
  assign n28250 = x17 | n28248 ;
  assign n28251 = x17 | n28247 ;
  assign n28252 = ( ~n21587 & n28250 ) | ( ~n21587 & n28251 ) | ( n28250 & n28251 ) ;
  assign n28253 = ( ~n28246 & n28249 ) | ( ~n28246 & n28252 ) | ( n28249 & n28252 ) ;
  assign n28254 = n28235 | n28253 ;
  assign n28255 = ( n28235 & n28238 ) | ( n28235 & n28254 ) | ( n28238 & n28254 ) ;
  assign n28256 = n28100 & n28255 ;
  assign n28257 = n28100 | n28255 ;
  assign n28258 = ~n28256 & n28257 ;
  assign n28259 = n1057 & n17100 ;
  assign n28260 = n1060 & ~n16069 ;
  assign n28261 = n1065 & n17111 ;
  assign n28262 = n28260 | n28261 ;
  assign n28263 = n28259 | n28262 ;
  assign n28264 = n1062 & n17169 ;
  assign n28265 = ~n17129 & n28264 ;
  assign n28266 = n28263 | n28265 ;
  assign n28267 = n1062 | n28263 ;
  assign n28268 = ( n17161 & n28266 ) | ( n17161 & n28267 ) | ( n28266 & n28267 ) ;
  assign n28269 = n4340 | n7016 ;
  assign n28270 = n11736 | n28269 ;
  assign n28271 = n407 | n22483 ;
  assign n28272 = n22482 | n28271 ;
  assign n28273 = n28270 | n28272 ;
  assign n28274 = n2147 | n4293 ;
  assign n28275 = n721 | n28274 ;
  assign n28276 = n442 | n5183 ;
  assign n28277 = n28275 | n28276 ;
  assign n28278 = n369 | n806 ;
  assign n28279 = n198 | n332 ;
  assign n28280 = n28278 | n28279 ;
  assign n28281 = n28277 | n28280 ;
  assign n28282 = n28273 | n28281 ;
  assign n28283 = n386 | n17701 ;
  assign n28284 = n18257 | n28283 ;
  assign n28285 = n17699 | n28284 ;
  assign n28286 = n1766 | n4246 ;
  assign n28287 = n28285 | n28286 ;
  assign n28288 = n28282 | n28287 ;
  assign n28289 = n702 | n4046 ;
  assign n28290 = n2265 | n28289 ;
  assign n28291 = n28288 | n28290 ;
  assign n28292 = n3330 | n15243 ;
  assign n28293 = n67 | n289 ;
  assign n28294 = n696 | n28293 ;
  assign n28295 = n28292 | n28294 ;
  assign n28296 = n270 | n310 ;
  assign n28297 = n280 | n28296 ;
  assign n28298 = n197 | n28297 ;
  assign n28299 = n28295 | n28298 ;
  assign n28300 = n333 | n28299 ;
  assign n28301 = n28291 | n28300 ;
  assign n28302 = n28122 & ~n28301 ;
  assign n28303 = ~n28122 & n28301 ;
  assign n28304 = n28302 | n28303 ;
  assign n28305 = n28259 & ~n28304 ;
  assign n28306 = ( n28262 & ~n28304 ) | ( n28262 & n28305 ) | ( ~n28304 & n28305 ) ;
  assign n28307 = ( n28265 & ~n28304 ) | ( n28265 & n28306 ) | ( ~n28304 & n28306 ) ;
  assign n28308 = ( n1062 & ~n28304 ) | ( n1062 & n28306 ) | ( ~n28304 & n28306 ) ;
  assign n28309 = ( n17161 & n28307 ) | ( n17161 & n28308 ) | ( n28307 & n28308 ) ;
  assign n28310 = n28268 & ~n28309 ;
  assign n28311 = n28125 & ~n28141 ;
  assign n28312 = n28304 | n28306 ;
  assign n28313 = n28265 | n28312 ;
  assign n28314 = n1062 | n28312 ;
  assign n28315 = ( n17161 & n28313 ) | ( n17161 & n28314 ) | ( n28313 & n28314 ) ;
  assign n28316 = n28311 | n28315 ;
  assign n28317 = ( ~n28310 & n28311 ) | ( ~n28310 & n28316 ) | ( n28311 & n28316 ) ;
  assign n28318 = n28311 & n28315 ;
  assign n28319 = ~n28310 & n28318 ;
  assign n28320 = n28317 & ~n28319 ;
  assign n28321 = n28147 | n28165 ;
  assign n28322 = ( n28147 & n28149 ) | ( n28147 & n28321 ) | ( n28149 & n28321 ) ;
  assign n28323 = n28320 & n28322 ;
  assign n28324 = n28320 | n28322 ;
  assign n28325 = ~n28323 & n28324 ;
  assign n28326 = n1829 & ~n18585 ;
  assign n28327 = n1826 & ~n17092 ;
  assign n28328 = n1823 & n18037 ;
  assign n28329 = n28327 | n28328 ;
  assign n28330 = n28326 | n28329 ;
  assign n28331 = n1821 & ~n18675 ;
  assign n28332 = ( n1821 & n18672 ) | ( n1821 & n28331 ) | ( n18672 & n28331 ) ;
  assign n28333 = n28330 | n28332 ;
  assign n28334 = x29 | n28330 ;
  assign n28335 = n28332 | n28334 ;
  assign n28336 = ~x29 & n28334 ;
  assign n28337 = ( ~x29 & n28332 ) | ( ~x29 & n28336 ) | ( n28332 & n28336 ) ;
  assign n28338 = ( ~n28333 & n28335 ) | ( ~n28333 & n28337 ) | ( n28335 & n28337 ) ;
  assign n28339 = n28325 & n28338 ;
  assign n28340 = n28325 & ~n28339 ;
  assign n28341 = n2315 & n19352 ;
  assign n28342 = n2312 & n18410 ;
  assign n28343 = n2308 & n18576 ;
  assign n28344 = n28342 | n28343 ;
  assign n28345 = n28341 | n28344 ;
  assign n28346 = n2306 | n28341 ;
  assign n28347 = n28344 | n28346 ;
  assign n28348 = ( n19674 & n28345 ) | ( n19674 & n28347 ) | ( n28345 & n28347 ) ;
  assign n28349 = x26 & n28347 ;
  assign n28350 = x26 & n28345 ;
  assign n28351 = ( n19674 & n28349 ) | ( n19674 & n28350 ) | ( n28349 & n28350 ) ;
  assign n28352 = x26 & ~n28350 ;
  assign n28353 = x26 & ~n28349 ;
  assign n28354 = ( ~n19674 & n28352 ) | ( ~n19674 & n28353 ) | ( n28352 & n28353 ) ;
  assign n28355 = ( n28348 & ~n28351 ) | ( n28348 & n28354 ) | ( ~n28351 & n28354 ) ;
  assign n28356 = ~n28325 & n28338 ;
  assign n28357 = n28355 & n28356 ;
  assign n28358 = ( n28340 & n28355 ) | ( n28340 & n28357 ) | ( n28355 & n28357 ) ;
  assign n28359 = n28355 | n28356 ;
  assign n28360 = n28340 | n28359 ;
  assign n28361 = ~n28358 & n28360 ;
  assign n28362 = n28170 | n28188 ;
  assign n28363 = ( n28170 & n28173 ) | ( n28170 & n28362 ) | ( n28173 & n28362 ) ;
  assign n28364 = n28361 & n28363 ;
  assign n28365 = n28361 | n28363 ;
  assign n28366 = ~n28364 & n28365 ;
  assign n28367 = n2932 & ~n20630 ;
  assign n28368 = n2925 & n19494 ;
  assign n28369 = n2928 & n19631 ;
  assign n28370 = n28368 | n28369 ;
  assign n28371 = n28367 | n28370 ;
  assign n28372 = n2936 | n28367 ;
  assign n28373 = n28370 | n28372 ;
  assign n28374 = ( ~n20709 & n28371 ) | ( ~n20709 & n28373 ) | ( n28371 & n28373 ) ;
  assign n28375 = ~x23 & n28373 ;
  assign n28376 = ~x23 & n28371 ;
  assign n28377 = ( ~n20709 & n28375 ) | ( ~n20709 & n28376 ) | ( n28375 & n28376 ) ;
  assign n28378 = x23 | n28376 ;
  assign n28379 = x23 | n28375 ;
  assign n28380 = ( ~n20709 & n28378 ) | ( ~n20709 & n28379 ) | ( n28378 & n28379 ) ;
  assign n28381 = ( ~n28374 & n28377 ) | ( ~n28374 & n28380 ) | ( n28377 & n28380 ) ;
  assign n28382 = n28366 & ~n28381 ;
  assign n28383 = n28366 | n28381 ;
  assign n28384 = ( ~n28366 & n28382 ) | ( ~n28366 & n28383 ) | ( n28382 & n28383 ) ;
  assign n28385 = n28192 | n28208 ;
  assign n28386 = ( n28192 & n28194 ) | ( n28192 & n28385 ) | ( n28194 & n28385 ) ;
  assign n28387 = n28384 & n28386 ;
  assign n28388 = n28384 | n28386 ;
  assign n28389 = ~n28387 & n28388 ;
  assign n28390 = n3547 & ~n21563 ;
  assign n28391 = n3544 & ~n20618 ;
  assign n28392 = n3541 & n20609 ;
  assign n28393 = n28391 | n28392 ;
  assign n28394 = n28390 | n28393 ;
  assign n28395 = n3537 & ~n21570 ;
  assign n28396 = n22270 & n28395 ;
  assign n28397 = ( n3537 & n22304 ) | ( n3537 & n28396 ) | ( n22304 & n28396 ) ;
  assign n28398 = n28394 | n28397 ;
  assign n28399 = x20 | n28394 ;
  assign n28400 = n28397 | n28399 ;
  assign n28401 = ~x20 & n28399 ;
  assign n28402 = ( ~x20 & n28397 ) | ( ~x20 & n28401 ) | ( n28397 & n28401 ) ;
  assign n28403 = ( ~n28398 & n28400 ) | ( ~n28398 & n28402 ) | ( n28400 & n28402 ) ;
  assign n28404 = n28389 & ~n28403 ;
  assign n28405 = n28389 | n28403 ;
  assign n28406 = ( ~n28389 & n28404 ) | ( ~n28389 & n28405 ) | ( n28404 & n28405 ) ;
  assign n28407 = n28212 | n28227 ;
  assign n28408 = ( n28212 & n28214 ) | ( n28212 & n28407 ) | ( n28214 & n28407 ) ;
  assign n28409 = n28406 & n28408 ;
  assign n28410 = n28406 | n28408 ;
  assign n28411 = ~n28409 & n28410 ;
  assign n28412 = n4466 & ~n21517 ;
  assign n28413 = n4468 & ~n21551 ;
  assign n28414 = n28412 | n28413 ;
  assign n28415 = n4471 & n23227 ;
  assign n28416 = ( n4471 & n23217 ) | ( n4471 & n28415 ) | ( n23217 & n28415 ) ;
  assign n28417 = n28414 | n28416 ;
  assign n28418 = n4475 & n23299 ;
  assign n28419 = n4475 & n23298 ;
  assign n28420 = ( n21584 & n28418 ) | ( n21584 & n28419 ) | ( n28418 & n28419 ) ;
  assign n28421 = n28417 | n28420 ;
  assign n28422 = n4475 | n28417 ;
  assign n28423 = ( n23289 & n28421 ) | ( n23289 & n28422 ) | ( n28421 & n28422 ) ;
  assign n28424 = x17 | n28423 ;
  assign n28425 = ~x17 & n28423 ;
  assign n28426 = ( ~n28423 & n28424 ) | ( ~n28423 & n28425 ) | ( n28424 & n28425 ) ;
  assign n28427 = n28411 & ~n28426 ;
  assign n28428 = n28411 | n28426 ;
  assign n28429 = ( ~n28411 & n28427 ) | ( ~n28411 & n28428 ) | ( n28427 & n28428 ) ;
  assign n28430 = n28258 & n28429 ;
  assign n28431 = ~n28258 & n28429 ;
  assign n28432 = ( n28258 & ~n28430 ) | ( n28258 & n28431 ) | ( ~n28430 & n28431 ) ;
  assign n28433 = n28238 & n28253 ;
  assign n28434 = n28238 & ~n28433 ;
  assign n28436 = n27547 | n27552 ;
  assign n28437 = ( n27547 & ~n27550 ) | ( n27547 & n28436 ) | ( ~n27550 & n28436 ) ;
  assign n28435 = ~n28238 & n28253 ;
  assign n28438 = n28435 & n28437 ;
  assign n28439 = ( n28434 & n28437 ) | ( n28434 & n28438 ) | ( n28437 & n28438 ) ;
  assign n28440 = n28435 | n28437 ;
  assign n28441 = n28434 | n28440 ;
  assign n28442 = ~n28439 & n28441 ;
  assign n28443 = n5231 & ~n23240 ;
  assign n28444 = n5237 & n23227 ;
  assign n28445 = ( n5237 & n23217 ) | ( n5237 & n28444 ) | ( n23217 & n28444 ) ;
  assign n28446 = n28443 | n28445 ;
  assign n28447 = n5234 & ~n23234 ;
  assign n28448 = n5234 & ~n23235 ;
  assign n28449 = ( ~n15882 & n28447 ) | ( ~n15882 & n28448 ) | ( n28447 & n28448 ) ;
  assign n28450 = n28446 | n28449 ;
  assign n28451 = n5227 | n28449 ;
  assign n28452 = n28446 | n28451 ;
  assign n28453 = ( ~n23587 & n28450 ) | ( ~n23587 & n28452 ) | ( n28450 & n28452 ) ;
  assign n28454 = ~x14 & n28452 ;
  assign n28455 = ~x14 & n28450 ;
  assign n28456 = ( ~n23587 & n28454 ) | ( ~n23587 & n28455 ) | ( n28454 & n28455 ) ;
  assign n28457 = x14 | n28455 ;
  assign n28458 = x14 | n28454 ;
  assign n28459 = ( ~n23587 & n28457 ) | ( ~n23587 & n28458 ) | ( n28457 & n28458 ) ;
  assign n28460 = ( ~n28453 & n28456 ) | ( ~n28453 & n28459 ) | ( n28456 & n28459 ) ;
  assign n28461 = n28439 | n28460 ;
  assign n28462 = ( n28439 & n28442 ) | ( n28439 & n28461 ) | ( n28442 & n28461 ) ;
  assign n28463 = n28432 & n28462 ;
  assign n28464 = n28432 | n28462 ;
  assign n28465 = ~n28463 & n28464 ;
  assign n28466 = n28442 & ~n28460 ;
  assign n28467 = n28442 | n28460 ;
  assign n28468 = ( ~n28442 & n28466 ) | ( ~n28442 & n28467 ) | ( n28466 & n28467 ) ;
  assign n28469 = n27574 | n27577 ;
  assign n28470 = n27555 & ~n27574 ;
  assign n28471 = ( n27575 & n28469 ) | ( n27575 & ~n28470 ) | ( n28469 & ~n28470 ) ;
  assign n28472 = n28468 & n28471 ;
  assign n28473 = n28471 & ~n28472 ;
  assign n28474 = n28468 & ~n28471 ;
  assign n28475 = n28473 | n28474 ;
  assign n28476 = n27585 & n28475 ;
  assign n28477 = n28472 | n28476 ;
  assign n28478 = n28472 | n28475 ;
  assign n28479 = ( n27600 & n28477 ) | ( n27600 & n28478 ) | ( n28477 & n28478 ) ;
  assign n28480 = n27585 | n27601 ;
  assign n28481 = n28475 & n28480 ;
  assign n28482 = n28472 | n28481 ;
  assign n28483 = ~n27585 & n27602 ;
  assign n28484 = n28475 & ~n28483 ;
  assign n28485 = n28472 | n28484 ;
  assign n28486 = ( n27130 & n28482 ) | ( n27130 & n28485 ) | ( n28482 & n28485 ) ;
  assign n28487 = ( n26009 & n28479 ) | ( n26009 & n28486 ) | ( n28479 & n28486 ) ;
  assign n28488 = ( n26011 & n28479 ) | ( n26011 & n28486 ) | ( n28479 & n28486 ) ;
  assign n28489 = ( n24765 & n28487 ) | ( n24765 & n28488 ) | ( n28487 & n28488 ) ;
  assign n28490 = n28465 & n28489 ;
  assign n28491 = n28465 | n28489 ;
  assign n28492 = ~n28490 & n28491 ;
  assign n28493 = n27585 | n27600 ;
  assign n28494 = ( n27130 & n28480 ) | ( n27130 & ~n28483 ) | ( n28480 & ~n28483 ) ;
  assign n28495 = ( n26009 & n28493 ) | ( n26009 & n28494 ) | ( n28493 & n28494 ) ;
  assign n28496 = ( n26011 & n28493 ) | ( n26011 & n28494 ) | ( n28493 & n28494 ) ;
  assign n28497 = ( n24765 & n28495 ) | ( n24765 & n28496 ) | ( n28495 & n28496 ) ;
  assign n28498 = n28475 | n28497 ;
  assign n28499 = ( n27600 & n28475 ) | ( n27600 & n28476 ) | ( n28475 & n28476 ) ;
  assign n28500 = ( n27130 & n28481 ) | ( n27130 & n28484 ) | ( n28481 & n28484 ) ;
  assign n28501 = ( n26009 & n28499 ) | ( n26009 & n28500 ) | ( n28499 & n28500 ) ;
  assign n28502 = ( n26011 & n28499 ) | ( n26011 & n28500 ) | ( n28499 & n28500 ) ;
  assign n28503 = ( n24765 & n28501 ) | ( n24765 & n28502 ) | ( n28501 & n28502 ) ;
  assign n28504 = n28498 & ~n28503 ;
  assign n28505 = n28492 & n28504 ;
  assign n28506 = n28492 | n28504 ;
  assign n28507 = ~n28505 & n28506 ;
  assign n28508 = ~n27626 & n28504 ;
  assign n28509 = n27626 & ~n28504 ;
  assign n28510 = n27627 | n28509 ;
  assign n28511 = ( ~n27629 & n28509 ) | ( ~n27629 & n28510 ) | ( n28509 & n28510 ) ;
  assign n28512 = ~n28508 & n28511 ;
  assign n28513 = ~n28508 & n28510 ;
  assign n28514 = n28512 & n28513 ;
  assign n28515 = n28507 & ~n28514 ;
  assign n28516 = ( n27612 & n28512 ) | ( n27612 & n28513 ) | ( n28512 & n28513 ) ;
  assign n28517 = n28507 & ~n28516 ;
  assign n28518 = ( n27625 & n28515 ) | ( n27625 & n28517 ) | ( n28515 & n28517 ) ;
  assign n28519 = n28505 | n28518 ;
  assign n28520 = n1607 | n3431 ;
  assign n28521 = n88 | n469 ;
  assign n28522 = n600 | n28521 ;
  assign n28523 = n28520 | n28522 ;
  assign n28524 = n390 | n28523 ;
  assign n28525 = n4144 | n24262 ;
  assign n28526 = n14388 | n28525 ;
  assign n28527 = n5962 | n18089 ;
  assign n28528 = n28526 | n28527 ;
  assign n28529 = n28524 | n28528 ;
  assign n28530 = n2731 & ~n28529 ;
  assign n28531 = ~n9170 & n28530 ;
  assign n28532 = n223 | n696 ;
  assign n28533 = n179 | n721 ;
  assign n28534 = n92 | n28533 ;
  assign n28535 = n594 | n28534 ;
  assign n28536 = n2742 | n28535 ;
  assign n28537 = ( ~n3355 & n28532 ) | ( ~n3355 & n28536 ) | ( n28532 & n28536 ) ;
  assign n28538 = n3355 | n28537 ;
  assign n28539 = n3355 & ~n28532 ;
  assign n28540 = ~n3355 & n28539 ;
  assign n28541 = ( n28531 & ~n28538 ) | ( n28531 & n28540 ) | ( ~n28538 & n28540 ) ;
  assign n28542 = n28122 & ~n28541 ;
  assign n28543 = ~n28122 & n28541 ;
  assign n28544 = n28542 | n28543 ;
  assign n28545 = n5237 | n28075 ;
  assign n28546 = n5227 | n28545 ;
  assign n28547 = ~n23229 & n28546 ;
  assign n28548 = ( n23154 & n28546 ) | ( n23154 & n28547 ) | ( n28546 & n28547 ) ;
  assign n28549 = ~n23232 & n28546 ;
  assign n28550 = ~n23231 & n28546 ;
  assign n28551 = ( n9072 & n28549 ) | ( n9072 & n28550 ) | ( n28549 & n28550 ) ;
  assign n28552 = ( ~n21543 & n28548 ) | ( ~n21543 & n28551 ) | ( n28548 & n28551 ) ;
  assign n28553 = ( ~n21545 & n28548 ) | ( ~n21545 & n28551 ) | ( n28548 & n28551 ) ;
  assign n28554 = ( ~n15882 & n28552 ) | ( ~n15882 & n28553 ) | ( n28552 & n28553 ) ;
  assign n28555 = ~x14 & n28552 ;
  assign n28556 = ~x14 & n28553 ;
  assign n28557 = ( ~n15882 & n28555 ) | ( ~n15882 & n28556 ) | ( n28555 & n28556 ) ;
  assign n28558 = x14 | n28555 ;
  assign n28559 = x14 | n28556 ;
  assign n28560 = ( ~n15882 & n28558 ) | ( ~n15882 & n28559 ) | ( n28558 & n28559 ) ;
  assign n28561 = ( ~n28554 & n28557 ) | ( ~n28554 & n28560 ) | ( n28557 & n28560 ) ;
  assign n28562 = n28544 | n28561 ;
  assign n28563 = n28544 & n28561 ;
  assign n28564 = n28562 & ~n28563 ;
  assign n28565 = n28303 | n28306 ;
  assign n28566 = ~n28303 & n28304 ;
  assign n28567 = ( n28265 & n28565 ) | ( n28265 & ~n28566 ) | ( n28565 & ~n28566 ) ;
  assign n28568 = ( n1062 & n28565 ) | ( n1062 & ~n28566 ) | ( n28565 & ~n28566 ) ;
  assign n28569 = ( n17161 & n28567 ) | ( n17161 & n28568 ) | ( n28567 & n28568 ) ;
  assign n28570 = n28564 & n28569 ;
  assign n28571 = n28564 | n28569 ;
  assign n28572 = ~n28570 & n28571 ;
  assign n28573 = n1057 & ~n17092 ;
  assign n28574 = n1060 & n17111 ;
  assign n28575 = n1065 & n17100 ;
  assign n28576 = n28574 | n28575 ;
  assign n28577 = n28573 | n28576 ;
  assign n28578 = n1062 | n28573 ;
  assign n28579 = n28576 | n28578 ;
  assign n28580 = ( ~n17134 & n28577 ) | ( ~n17134 & n28579 ) | ( n28577 & n28579 ) ;
  assign n28581 = ~n28572 & n28580 ;
  assign n28582 = n28572 & ~n28580 ;
  assign n28583 = n28581 | n28582 ;
  assign n28584 = n1829 & n18410 ;
  assign n28585 = n1826 & n18037 ;
  assign n28586 = n1823 & ~n18585 ;
  assign n28587 = n28585 | n28586 ;
  assign n28588 = n28584 | n28587 ;
  assign n28589 = n1821 & ~n18586 ;
  assign n28590 = ~n18609 & n28589 ;
  assign n28591 = ( n1821 & n18650 ) | ( n1821 & n28590 ) | ( n18650 & n28590 ) ;
  assign n28592 = n28588 | n28591 ;
  assign n28593 = x29 | n28588 ;
  assign n28594 = n28591 | n28593 ;
  assign n28595 = ~x29 & n28593 ;
  assign n28596 = ( ~x29 & n28591 ) | ( ~x29 & n28595 ) | ( n28591 & n28595 ) ;
  assign n28597 = ( ~n28592 & n28594 ) | ( ~n28592 & n28596 ) | ( n28594 & n28596 ) ;
  assign n28598 = n28583 & n28597 ;
  assign n28599 = n28583 & ~n28598 ;
  assign n28601 = n28317 & ~n28320 ;
  assign n28602 = ( n28317 & ~n28322 ) | ( n28317 & n28601 ) | ( ~n28322 & n28601 ) ;
  assign n28600 = ~n28583 & n28597 ;
  assign n28603 = n28600 & ~n28602 ;
  assign n28604 = ( n28599 & ~n28602 ) | ( n28599 & n28603 ) | ( ~n28602 & n28603 ) ;
  assign n28605 = ~n28600 & n28602 ;
  assign n28606 = ~n28599 & n28605 ;
  assign n28607 = n28604 | n28606 ;
  assign n28608 = n2315 & n19494 ;
  assign n28609 = n2312 & n18576 ;
  assign n28610 = n2308 & n19352 ;
  assign n28611 = n28609 | n28610 ;
  assign n28612 = n28608 | n28611 ;
  assign n28613 = n2306 | n28608 ;
  assign n28614 = n28611 | n28613 ;
  assign n28615 = ( n20320 & n28612 ) | ( n20320 & n28614 ) | ( n28612 & n28614 ) ;
  assign n28616 = x26 & n28614 ;
  assign n28617 = x26 & n28612 ;
  assign n28618 = ( n20320 & n28616 ) | ( n20320 & n28617 ) | ( n28616 & n28617 ) ;
  assign n28619 = x26 & ~n28617 ;
  assign n28620 = x26 & ~n28616 ;
  assign n28621 = ( ~n20320 & n28619 ) | ( ~n20320 & n28620 ) | ( n28619 & n28620 ) ;
  assign n28622 = ( n28615 & ~n28618 ) | ( n28615 & n28621 ) | ( ~n28618 & n28621 ) ;
  assign n28623 = ~n28607 & n28622 ;
  assign n28624 = n28607 | n28623 ;
  assign n28625 = n28607 & n28622 ;
  assign n28626 = n28624 & ~n28625 ;
  assign n28627 = n28339 | n28358 ;
  assign n28628 = ~n28626 & n28627 ;
  assign n28629 = n28626 & ~n28627 ;
  assign n28630 = n28628 | n28629 ;
  assign n28631 = n2936 & n20680 ;
  assign n28632 = n2932 & ~n20618 ;
  assign n28633 = n2925 & n19631 ;
  assign n28634 = n2928 & ~n20630 ;
  assign n28635 = n28633 | n28634 ;
  assign n28636 = n28632 | n28635 ;
  assign n28637 = n20689 | n28636 ;
  assign n28638 = n2936 | n28636 ;
  assign n28639 = ( n28631 & n28637 ) | ( n28631 & n28638 ) | ( n28637 & n28638 ) ;
  assign n28640 = x23 | n28639 ;
  assign n28641 = ~x23 & n28639 ;
  assign n28642 = ( ~n28639 & n28640 ) | ( ~n28639 & n28641 ) | ( n28640 & n28641 ) ;
  assign n28643 = ~n28630 & n28642 ;
  assign n28644 = n28630 | n28643 ;
  assign n28646 = n28364 | n28381 ;
  assign n28647 = ( n28364 & n28366 ) | ( n28364 & n28646 ) | ( n28366 & n28646 ) ;
  assign n28645 = n28630 & n28642 ;
  assign n28648 = n28645 & n28647 ;
  assign n28649 = ( ~n28644 & n28647 ) | ( ~n28644 & n28648 ) | ( n28647 & n28648 ) ;
  assign n28650 = n28645 | n28647 ;
  assign n28651 = n28644 & ~n28650 ;
  assign n28652 = n28649 | n28651 ;
  assign n28653 = n3547 & ~n21517 ;
  assign n28654 = n3544 & n20609 ;
  assign n28655 = n3541 & ~n21563 ;
  assign n28656 = n28654 | n28655 ;
  assign n28657 = n28653 | n28656 ;
  assign n28658 = n3537 | n28653 ;
  assign n28659 = n28656 | n28658 ;
  assign n28660 = ( ~n22283 & n28657 ) | ( ~n22283 & n28659 ) | ( n28657 & n28659 ) ;
  assign n28661 = n28657 & n28659 ;
  assign n28662 = ( ~n22271 & n28660 ) | ( ~n22271 & n28661 ) | ( n28660 & n28661 ) ;
  assign n28663 = ~x20 & n28662 ;
  assign n28664 = x20 | n28662 ;
  assign n28665 = ( ~n28662 & n28663 ) | ( ~n28662 & n28664 ) | ( n28663 & n28664 ) ;
  assign n28666 = ~n28652 & n28665 ;
  assign n28667 = n28652 | n28666 ;
  assign n28668 = n28387 | n28403 ;
  assign n28669 = ( n28387 & n28389 ) | ( n28387 & n28668 ) | ( n28389 & n28668 ) ;
  assign n28670 = n28652 & n28665 ;
  assign n28671 = n28669 & n28670 ;
  assign n28672 = ( ~n28667 & n28669 ) | ( ~n28667 & n28671 ) | ( n28669 & n28671 ) ;
  assign n28673 = n28669 | n28670 ;
  assign n28674 = n28667 & ~n28673 ;
  assign n28675 = n28672 | n28674 ;
  assign n28692 = n28409 | n28426 ;
  assign n28693 = ( n28409 & n28411 ) | ( n28409 & n28692 ) | ( n28411 & n28692 ) ;
  assign n28676 = n4471 & ~n23240 ;
  assign n28677 = n4466 & ~n21551 ;
  assign n28678 = n4468 & n23227 ;
  assign n28679 = ( n4468 & n23217 ) | ( n4468 & n28678 ) | ( n23217 & n28678 ) ;
  assign n28680 = n28677 | n28679 ;
  assign n28681 = n28676 | n28680 ;
  assign n28682 = n4475 | n28676 ;
  assign n28683 = n28680 | n28682 ;
  assign n28684 = ( n23260 & n28681 ) | ( n23260 & n28683 ) | ( n28681 & n28683 ) ;
  assign n28685 = x17 & n28683 ;
  assign n28686 = x17 & n28681 ;
  assign n28687 = ( n23260 & n28685 ) | ( n23260 & n28686 ) | ( n28685 & n28686 ) ;
  assign n28688 = x17 & ~n28686 ;
  assign n28689 = x17 & ~n28685 ;
  assign n28690 = ( ~n23260 & n28688 ) | ( ~n23260 & n28689 ) | ( n28688 & n28689 ) ;
  assign n28691 = ( n28684 & ~n28687 ) | ( n28684 & n28690 ) | ( ~n28687 & n28690 ) ;
  assign n28694 = n28691 & n28693 ;
  assign n28695 = n28693 & ~n28694 ;
  assign n28696 = n28691 & ~n28693 ;
  assign n28697 = ~n28675 & n28696 ;
  assign n28698 = ( ~n28675 & n28695 ) | ( ~n28675 & n28697 ) | ( n28695 & n28697 ) ;
  assign n28699 = n28675 & ~n28696 ;
  assign n28700 = ~n28695 & n28699 ;
  assign n28701 = n28698 | n28700 ;
  assign n28702 = n28256 | n28429 ;
  assign n28703 = ( n28256 & n28258 ) | ( n28256 & n28702 ) | ( n28258 & n28702 ) ;
  assign n28704 = ~n28701 & n28703 ;
  assign n28705 = n28701 & ~n28703 ;
  assign n28706 = n28704 | n28705 ;
  assign n28707 = n28463 & ~n28706 ;
  assign n28708 = ( n28465 & ~n28706 ) | ( n28465 & n28707 ) | ( ~n28706 & n28707 ) ;
  assign n28709 = ~n28706 & n28707 ;
  assign n28710 = ( n28489 & n28708 ) | ( n28489 & n28709 ) | ( n28708 & n28709 ) ;
  assign n28711 = ~n28463 & n28706 ;
  assign n28712 = ~n28465 & n28711 ;
  assign n28713 = ( ~n28489 & n28711 ) | ( ~n28489 & n28712 ) | ( n28711 & n28712 ) ;
  assign n28714 = n28710 | n28713 ;
  assign n28715 = n28492 & ~n28714 ;
  assign n28716 = ~n28492 & n28714 ;
  assign n28717 = n28715 | n28716 ;
  assign n28718 = n28505 & ~n28717 ;
  assign n28719 = ( n28518 & ~n28717 ) | ( n28518 & n28718 ) | ( ~n28717 & n28718 ) ;
  assign n28720 = n28519 & ~n28719 ;
  assign n28721 = n5231 & n28492 ;
  assign n28722 = n5237 & ~n28503 ;
  assign n28723 = n28498 & n28722 ;
  assign n28724 = n28721 | n28723 ;
  assign n28725 = n5234 & ~n28714 ;
  assign n28726 = n5227 | n28725 ;
  assign n28727 = n28724 | n28726 ;
  assign n28728 = n28724 | n28725 ;
  assign n28729 = n28505 | n28715 ;
  assign n28730 = ( n28715 & ~n28717 ) | ( n28715 & n28729 ) | ( ~n28717 & n28729 ) ;
  assign n28731 = n28716 | n28730 ;
  assign n28732 = ~n28728 & n28731 ;
  assign n28733 = ( n28518 & ~n28728 ) | ( n28518 & n28732 ) | ( ~n28728 & n28732 ) ;
  assign n28734 = n28727 & ~n28733 ;
  assign n28735 = ( n28720 & n28727 ) | ( n28720 & n28734 ) | ( n28727 & n28734 ) ;
  assign n28736 = x14 & n28735 ;
  assign n28737 = x14 & ~n28735 ;
  assign n28738 = ( n28735 & ~n28736 ) | ( n28735 & n28737 ) | ( ~n28736 & n28737 ) ;
  assign n28739 = ~n28074 & n28738 ;
  assign n28740 = n28074 | n28739 ;
  assign n28741 = n28074 & n28738 ;
  assign n28742 = n28740 & ~n28741 ;
  assign n28743 = n27678 & n28069 ;
  assign n28744 = n27678 | n28069 ;
  assign n28745 = ~n28743 & n28744 ;
  assign n28746 = ~n28507 & n28514 ;
  assign n28747 = ~n28507 & n28516 ;
  assign n28748 = ( ~n27625 & n28746 ) | ( ~n27625 & n28747 ) | ( n28746 & n28747 ) ;
  assign n28749 = n28518 | n28748 ;
  assign n28750 = n5234 & n28492 ;
  assign n28751 = n5237 & ~n27606 ;
  assign n28752 = ~n27597 & n28751 ;
  assign n28753 = n5231 & ~n28503 ;
  assign n28754 = n28498 & n28753 ;
  assign n28755 = n28752 | n28754 ;
  assign n28756 = n28750 | n28755 ;
  assign n28757 = n5227 | n28756 ;
  assign n28758 = n28756 & n28757 ;
  assign n28759 = ( ~n28749 & n28757 ) | ( ~n28749 & n28758 ) | ( n28757 & n28758 ) ;
  assign n28760 = ~x14 & n28758 ;
  assign n28761 = ~x14 & n28757 ;
  assign n28762 = ( ~n28749 & n28760 ) | ( ~n28749 & n28761 ) | ( n28760 & n28761 ) ;
  assign n28763 = x14 | n28760 ;
  assign n28764 = x14 | n28761 ;
  assign n28765 = ( ~n28749 & n28763 ) | ( ~n28749 & n28764 ) | ( n28763 & n28764 ) ;
  assign n28766 = ( ~n28759 & n28762 ) | ( ~n28759 & n28765 ) | ( n28762 & n28765 ) ;
  assign n28767 = n28745 & n28766 ;
  assign n28768 = n28745 & ~n28767 ;
  assign n28769 = ~n28745 & n28766 ;
  assign n28770 = n28768 | n28769 ;
  assign n28771 = ~n27713 & n28067 ;
  assign n28772 = n27713 & ~n28067 ;
  assign n28773 = n28771 | n28772 ;
  assign n28774 = n27627 & ~n27629 ;
  assign n28775 = ( n27612 & n27627 ) | ( n27612 & n28774 ) | ( n27627 & n28774 ) ;
  assign n28776 = n27627 & n28774 ;
  assign n28777 = ( ~n27625 & n28775 ) | ( ~n27625 & n28776 ) | ( n28775 & n28776 ) ;
  assign n28778 = n28508 | n28511 ;
  assign n28779 = n28508 | n28510 ;
  assign n28780 = ( n27612 & n28778 ) | ( n27612 & n28779 ) | ( n28778 & n28779 ) ;
  assign n28781 = n28778 & n28779 ;
  assign n28782 = ( ~n27625 & n28780 ) | ( ~n27625 & n28781 ) | ( n28780 & n28781 ) ;
  assign n28783 = ~n28777 & n28782 ;
  assign n28784 = n5237 & ~n27371 ;
  assign n28785 = ~n27363 & n28784 ;
  assign n28786 = n5231 & ~n27606 ;
  assign n28787 = ~n27597 & n28786 ;
  assign n28788 = n28785 | n28787 ;
  assign n28789 = n5234 & ~n28503 ;
  assign n28790 = n28498 & n28789 ;
  assign n28791 = n28788 | n28790 ;
  assign n28792 = ~n28509 & n28514 ;
  assign n28793 = ~n28509 & n28516 ;
  assign n28794 = ( ~n27625 & n28792 ) | ( ~n27625 & n28793 ) | ( n28792 & n28793 ) ;
  assign n28795 = n28791 | n28794 ;
  assign n28796 = n28783 | n28795 ;
  assign n28797 = n5227 | n28790 ;
  assign n28798 = n28788 | n28797 ;
  assign n28799 = n28796 & n28798 ;
  assign n28800 = ~x14 & n28798 ;
  assign n28801 = n28796 & n28800 ;
  assign n28802 = x14 | n28800 ;
  assign n28803 = ( x14 & n28796 ) | ( x14 & n28802 ) | ( n28796 & n28802 ) ;
  assign n28804 = ( ~n28799 & n28801 ) | ( ~n28799 & n28803 ) | ( n28801 & n28803 ) ;
  assign n28805 = ~n28773 & n28804 ;
  assign n28806 = n28773 | n28805 ;
  assign n28807 = n28773 & n28804 ;
  assign n28808 = n28806 & ~n28807 ;
  assign n28809 = ( n28061 & n28062 ) | ( n28061 & ~n28065 ) | ( n28062 & ~n28065 ) ;
  assign n28810 = n27732 | n28061 ;
  assign n28811 = n28065 & ~n28810 ;
  assign n28812 = n28809 | n28811 ;
  assign n28813 = n5237 & ~n27133 ;
  assign n28814 = ~n27125 & n28813 ;
  assign n28815 = n5231 & ~n27371 ;
  assign n28816 = ~n27363 & n28815 ;
  assign n28817 = n28814 | n28816 ;
  assign n28818 = n5234 & ~n27606 ;
  assign n28819 = ~n27597 & n28818 ;
  assign n28820 = n28817 | n28819 ;
  assign n28821 = n27630 | n28820 ;
  assign n28822 = ( ~n27625 & n28820 ) | ( ~n27625 & n28821 ) | ( n28820 & n28821 ) ;
  assign n28823 = n27634 & ~n28822 ;
  assign n28824 = n5227 | n28819 ;
  assign n28825 = n28817 | n28824 ;
  assign n28826 = ~n28823 & n28825 ;
  assign n28827 = x14 & n28825 ;
  assign n28828 = ~n28823 & n28827 ;
  assign n28829 = x14 & ~n28827 ;
  assign n28830 = ( x14 & n28823 ) | ( x14 & n28829 ) | ( n28823 & n28829 ) ;
  assign n28831 = ( n28826 & ~n28828 ) | ( n28826 & n28830 ) | ( ~n28828 & n28830 ) ;
  assign n28832 = ~n28812 & n28831 ;
  assign n28833 = n28812 | n28832 ;
  assign n28834 = n28812 & n28831 ;
  assign n28835 = n28833 & ~n28834 ;
  assign n28836 = n28057 & n28059 ;
  assign n28837 = n28057 | n28059 ;
  assign n28838 = ~n28836 & n28837 ;
  assign n28839 = n5237 & ~n26526 ;
  assign n28840 = ~n26520 & n28839 ;
  assign n28841 = n5231 & ~n27133 ;
  assign n28842 = ~n27125 & n28841 ;
  assign n28843 = n28840 | n28842 ;
  assign n28844 = n5234 & ~n27371 ;
  assign n28845 = ~n27363 & n28844 ;
  assign n28846 = n28843 | n28845 ;
  assign n28847 = n5227 | n28845 ;
  assign n28848 = n28843 | n28847 ;
  assign n28849 = ( ~n27654 & n28846 ) | ( ~n27654 & n28848 ) | ( n28846 & n28848 ) ;
  assign n28850 = ~x14 & n28848 ;
  assign n28851 = ~x14 & n28846 ;
  assign n28852 = ( ~n27654 & n28850 ) | ( ~n27654 & n28851 ) | ( n28850 & n28851 ) ;
  assign n28853 = x14 | n28851 ;
  assign n28854 = x14 | n28850 ;
  assign n28855 = ( ~n27654 & n28853 ) | ( ~n27654 & n28854 ) | ( n28853 & n28854 ) ;
  assign n28856 = ( ~n28849 & n28852 ) | ( ~n28849 & n28855 ) | ( n28852 & n28855 ) ;
  assign n28857 = n28838 & n28856 ;
  assign n28858 = ~n27773 & n28055 ;
  assign n28859 = n27773 & ~n28055 ;
  assign n28860 = n28858 | n28859 ;
  assign n28861 = n5237 & ~n26270 ;
  assign n28862 = ~n26263 & n28861 ;
  assign n28863 = n5231 & ~n26526 ;
  assign n28864 = ~n26520 & n28863 ;
  assign n28865 = n28862 | n28864 ;
  assign n28866 = n5234 & ~n27133 ;
  assign n28867 = ~n27125 & n28866 ;
  assign n28868 = n28865 | n28867 ;
  assign n28869 = n5227 & n27699 ;
  assign n28870 = ( n5227 & ~n27696 ) | ( n5227 & n28869 ) | ( ~n27696 & n28869 ) ;
  assign n28871 = n28868 | n28870 ;
  assign n28872 = x14 | n28868 ;
  assign n28873 = n28870 | n28872 ;
  assign n28874 = ~x14 & n28872 ;
  assign n28875 = ( ~x14 & n28870 ) | ( ~x14 & n28874 ) | ( n28870 & n28874 ) ;
  assign n28876 = ( ~n28871 & n28873 ) | ( ~n28871 & n28875 ) | ( n28873 & n28875 ) ;
  assign n28877 = n28860 & n28876 ;
  assign n28878 = n28860 | n28876 ;
  assign n28879 = ~n28877 & n28878 ;
  assign n28880 = n28051 & n28053 ;
  assign n28881 = n28051 | n28053 ;
  assign n28882 = ~n28880 & n28881 ;
  assign n28883 = n5237 & n26017 ;
  assign n28884 = n5231 & ~n26270 ;
  assign n28885 = ~n26263 & n28884 ;
  assign n28886 = n28883 | n28885 ;
  assign n28887 = n5234 & ~n26526 ;
  assign n28888 = ~n26520 & n28887 ;
  assign n28890 = n5227 | n28888 ;
  assign n28891 = n28886 | n28890 ;
  assign n28889 = n28886 | n28888 ;
  assign n28892 = n28889 & n28891 ;
  assign n28893 = ( ~n26555 & n28891 ) | ( ~n26555 & n28892 ) | ( n28891 & n28892 ) ;
  assign n28894 = ( n26528 & n28891 ) | ( n26528 & n28892 ) | ( n28891 & n28892 ) ;
  assign n28895 = ( ~n26543 & n28893 ) | ( ~n26543 & n28894 ) | ( n28893 & n28894 ) ;
  assign n28896 = ~x14 & n28895 ;
  assign n28897 = x14 | n28895 ;
  assign n28898 = ( ~n28895 & n28896 ) | ( ~n28895 & n28897 ) | ( n28896 & n28897 ) ;
  assign n28899 = n28882 & n28898 ;
  assign n28900 = n27816 | n28049 ;
  assign n28901 = ~n28050 & n28900 ;
  assign n28902 = n5237 & ~n25728 ;
  assign n28903 = n5231 & n26017 ;
  assign n28904 = n28902 | n28903 ;
  assign n28905 = n5234 & ~n26270 ;
  assign n28906 = ~n26263 & n28905 ;
  assign n28908 = n5227 | n28906 ;
  assign n28909 = n28904 | n28908 ;
  assign n28907 = n28904 | n28906 ;
  assign n28910 = n28907 & n28909 ;
  assign n28911 = ( n26571 & n28909 ) | ( n26571 & n28910 ) | ( n28909 & n28910 ) ;
  assign n28912 = x14 & n28910 ;
  assign n28913 = x14 & n28909 ;
  assign n28914 = ( n26571 & n28912 ) | ( n26571 & n28913 ) | ( n28912 & n28913 ) ;
  assign n28915 = x14 & ~n28912 ;
  assign n28916 = x14 & ~n28913 ;
  assign n28917 = ( ~n26571 & n28915 ) | ( ~n26571 & n28916 ) | ( n28915 & n28916 ) ;
  assign n28918 = ( n28911 & ~n28914 ) | ( n28911 & n28917 ) | ( ~n28914 & n28917 ) ;
  assign n28919 = n28901 & n28918 ;
  assign n28920 = n28901 & ~n28919 ;
  assign n28921 = ~n28901 & n28918 ;
  assign n28922 = n28920 | n28921 ;
  assign n28923 = n27837 & n28047 ;
  assign n28924 = n27837 | n28047 ;
  assign n28925 = ~n28923 & n28924 ;
  assign n28926 = n5234 & n26017 ;
  assign n28927 = n5237 & ~n25046 ;
  assign n28928 = n5231 & ~n25728 ;
  assign n28929 = n28927 | n28928 ;
  assign n28930 = n28926 | n28929 ;
  assign n28931 = n5227 | n28926 ;
  assign n28932 = n28929 | n28931 ;
  assign n28933 = ( n26613 & n28930 ) | ( n26613 & n28932 ) | ( n28930 & n28932 ) ;
  assign n28934 = n28930 | n28932 ;
  assign n28935 = ( n26605 & n28933 ) | ( n26605 & n28934 ) | ( n28933 & n28934 ) ;
  assign n28936 = x14 & n28935 ;
  assign n28937 = x14 & ~n28935 ;
  assign n28938 = ( n28935 & ~n28936 ) | ( n28935 & n28937 ) | ( ~n28936 & n28937 ) ;
  assign n28939 = n28925 & n28938 ;
  assign n28940 = n28925 & ~n28939 ;
  assign n28941 = ~n28925 & n28938 ;
  assign n28942 = n28940 | n28941 ;
  assign n28943 = ( n27873 & n27874 ) | ( n27873 & n28045 ) | ( n27874 & n28045 ) ;
  assign n28944 = n27852 | n27873 ;
  assign n28945 = n28045 | n28944 ;
  assign n28946 = ~n28943 & n28945 ;
  assign n28947 = n5234 & ~n25728 ;
  assign n28948 = n5237 & n24770 ;
  assign n28949 = n5231 & ~n25046 ;
  assign n28950 = n28948 | n28949 ;
  assign n28951 = n28947 | n28950 ;
  assign n28952 = n5227 & n25740 ;
  assign n28953 = n5227 & n25731 ;
  assign n28954 = ( ~n25441 & n28952 ) | ( ~n25441 & n28953 ) | ( n28952 & n28953 ) ;
  assign n28955 = n28951 | n28954 ;
  assign n28956 = n5227 | n28951 ;
  assign n28957 = ( n25733 & n28955 ) | ( n25733 & n28956 ) | ( n28955 & n28956 ) ;
  assign n28958 = x14 | n28957 ;
  assign n28959 = ~x14 & n28957 ;
  assign n28960 = ( ~n28957 & n28958 ) | ( ~n28957 & n28959 ) | ( n28958 & n28959 ) ;
  assign n28961 = n28946 & n28960 ;
  assign n28962 = n28042 & ~n28045 ;
  assign n28965 = n5234 & ~n25046 ;
  assign n28966 = n5237 & ~n25054 ;
  assign n28967 = n5231 & n24770 ;
  assign n28968 = n28966 | n28967 ;
  assign n28969 = n28965 | n28968 ;
  assign n28970 = n5227 | n28965 ;
  assign n28971 = n28968 | n28970 ;
  assign n28972 = ( ~n25069 & n28969 ) | ( ~n25069 & n28971 ) | ( n28969 & n28971 ) ;
  assign n28973 = ~x14 & n28971 ;
  assign n28974 = ~x14 & n28969 ;
  assign n28975 = ( ~n25069 & n28973 ) | ( ~n25069 & n28974 ) | ( n28973 & n28974 ) ;
  assign n28976 = x14 | n28974 ;
  assign n28977 = x14 | n28973 ;
  assign n28978 = ( ~n25069 & n28976 ) | ( ~n25069 & n28977 ) | ( n28976 & n28977 ) ;
  assign n28979 = ( ~n28972 & n28975 ) | ( ~n28972 & n28978 ) | ( n28975 & n28978 ) ;
  assign n28963 = ~n28042 & n28044 ;
  assign n28980 = n28963 & n28979 ;
  assign n28981 = ( n28962 & n28979 ) | ( n28962 & n28980 ) | ( n28979 & n28980 ) ;
  assign n28964 = n28962 | n28963 ;
  assign n28982 = n28964 & ~n28981 ;
  assign n28983 = ~n28963 & n28979 ;
  assign n28984 = ~n28962 & n28983 ;
  assign n28985 = n28982 | n28984 ;
  assign n28986 = n28040 & ~n28041 ;
  assign n28987 = n27897 & ~n28041 ;
  assign n28988 = n28986 | n28987 ;
  assign n28989 = n5234 & n24770 ;
  assign n28990 = n5237 & n24167 ;
  assign n28991 = n5231 & ~n25054 ;
  assign n28992 = n28990 | n28991 ;
  assign n28993 = n28989 | n28992 ;
  assign n28994 = n5227 | n28993 ;
  assign n28995 = ( ~n25095 & n28993 ) | ( ~n25095 & n28994 ) | ( n28993 & n28994 ) ;
  assign n28996 = ~x14 & n28994 ;
  assign n28997 = ~x14 & n28993 ;
  assign n28998 = ( ~n25095 & n28996 ) | ( ~n25095 & n28997 ) | ( n28996 & n28997 ) ;
  assign n28999 = x14 | n28996 ;
  assign n29000 = x14 | n28997 ;
  assign n29001 = ( ~n25095 & n28999 ) | ( ~n25095 & n29000 ) | ( n28999 & n29000 ) ;
  assign n29002 = ( ~n28995 & n28998 ) | ( ~n28995 & n29001 ) | ( n28998 & n29001 ) ;
  assign n29003 = n28988 & n29002 ;
  assign n29004 = n28988 & ~n29003 ;
  assign n29005 = ~n28988 & n29002 ;
  assign n29006 = n29004 | n29005 ;
  assign n29007 = n27919 | n28013 ;
  assign n29008 = ~n28014 & n29007 ;
  assign n29009 = n5234 & n24167 ;
  assign n29010 = n5237 & n23316 ;
  assign n29011 = n5231 & n23614 ;
  assign n29012 = n29010 | n29011 ;
  assign n29013 = n29009 | n29012 ;
  assign n29014 = n5227 | n29013 ;
  assign n29015 = ( n24182 & n29013 ) | ( n24182 & n29014 ) | ( n29013 & n29014 ) ;
  assign n29016 = n29013 | n29014 ;
  assign n29017 = ( n24175 & n29015 ) | ( n24175 & n29016 ) | ( n29015 & n29016 ) ;
  assign n29018 = x14 & n29017 ;
  assign n29019 = x14 & ~n29017 ;
  assign n29020 = ( n29017 & ~n29018 ) | ( n29017 & n29019 ) | ( ~n29018 & n29019 ) ;
  assign n29021 = n29008 & n29020 ;
  assign n29022 = n28015 & n28038 ;
  assign n29023 = n28015 | n28038 ;
  assign n29024 = ~n29022 & n29023 ;
  assign n29025 = n5234 & ~n25054 ;
  assign n29026 = n5237 & n23614 ;
  assign n29027 = n5231 & n24167 ;
  assign n29028 = n29026 | n29027 ;
  assign n29029 = n29025 | n29028 ;
  assign n29030 = n5227 | n29025 ;
  assign n29031 = n29028 | n29030 ;
  assign n29032 = ( ~n25122 & n29029 ) | ( ~n25122 & n29031 ) | ( n29029 & n29031 ) ;
  assign n29033 = ~x14 & n29031 ;
  assign n29034 = ~x14 & n29029 ;
  assign n29035 = ( ~n25122 & n29033 ) | ( ~n25122 & n29034 ) | ( n29033 & n29034 ) ;
  assign n29036 = x14 | n29034 ;
  assign n29037 = x14 | n29033 ;
  assign n29038 = ( ~n25122 & n29036 ) | ( ~n25122 & n29037 ) | ( n29036 & n29037 ) ;
  assign n29039 = ( ~n29032 & n29035 ) | ( ~n29032 & n29038 ) | ( n29035 & n29038 ) ;
  assign n29040 = n29024 & n29039 ;
  assign n29041 = n29024 | n29039 ;
  assign n29042 = ~n29040 & n29041 ;
  assign n29043 = n29021 & n29042 ;
  assign n29044 = n29040 | n29042 ;
  assign n29045 = n27938 | n28011 ;
  assign n29046 = ~n28012 & n29045 ;
  assign n29047 = n5234 & n23614 ;
  assign n29048 = n5237 & n23620 ;
  assign n29049 = ( n5231 & n5357 ) | ( n5231 & n23620 ) | ( n5357 & n23620 ) ;
  assign n29050 = ( n23316 & n29048 ) | ( n23316 & n29049 ) | ( n29048 & n29049 ) ;
  assign n29052 = n5227 | n29050 ;
  assign n29053 = n29047 | n29052 ;
  assign n29051 = n29047 | n29050 ;
  assign n29054 = n29051 & n29053 ;
  assign n29055 = ( n23634 & n29053 ) | ( n23634 & n29054 ) | ( n29053 & n29054 ) ;
  assign n29056 = x14 & n29054 ;
  assign n29057 = x14 & n29053 ;
  assign n29058 = ( n23634 & n29056 ) | ( n23634 & n29057 ) | ( n29056 & n29057 ) ;
  assign n29059 = x14 & ~n29056 ;
  assign n29060 = x14 & ~n29057 ;
  assign n29061 = ( ~n23634 & n29059 ) | ( ~n23634 & n29060 ) | ( n29059 & n29060 ) ;
  assign n29062 = ( n29055 & ~n29058 ) | ( n29055 & n29061 ) | ( ~n29058 & n29061 ) ;
  assign n29063 = n29046 & n29062 ;
  assign n29064 = n29046 & ~n29063 ;
  assign n29065 = ~n29046 & n29062 ;
  assign n29066 = n29064 | n29065 ;
  assign n29067 = n27991 & n28005 ;
  assign n29068 = n27991 & ~n29067 ;
  assign n29069 = n5237 & ~n22385 ;
  assign n29070 = ( n5231 & n5357 ) | ( n5231 & ~n22385 ) | ( n5357 & ~n22385 ) ;
  assign n29071 = ( n22381 & n29069 ) | ( n22381 & n29070 ) | ( n29069 & n29070 ) ;
  assign n29072 = n5234 | n29071 ;
  assign n29073 = ( n23620 & n29071 ) | ( n23620 & n29072 ) | ( n29071 & n29072 ) ;
  assign n29074 = n5227 | n29073 ;
  assign n29075 = ( ~n23686 & n29073 ) | ( ~n23686 & n29074 ) | ( n29073 & n29074 ) ;
  assign n29076 = ~x14 & n29074 ;
  assign n29077 = ~x14 & n29073 ;
  assign n29078 = ( ~n23686 & n29076 ) | ( ~n23686 & n29077 ) | ( n29076 & n29077 ) ;
  assign n29079 = x14 | n29076 ;
  assign n29080 = x14 | n29077 ;
  assign n29081 = ( ~n23686 & n29079 ) | ( ~n23686 & n29080 ) | ( n29079 & n29080 ) ;
  assign n29082 = ( ~n29075 & n29078 ) | ( ~n29075 & n29081 ) | ( n29078 & n29081 ) ;
  assign n29083 = ~n27991 & n28005 ;
  assign n29084 = n29082 & n29083 ;
  assign n29085 = ( n29068 & n29082 ) | ( n29068 & n29084 ) | ( n29082 & n29084 ) ;
  assign n29086 = n29082 | n29083 ;
  assign n29087 = n29068 | n29086 ;
  assign n29088 = ~n29085 & n29087 ;
  assign n29089 = n27970 & n27988 ;
  assign n29090 = n27970 | n27988 ;
  assign n29091 = ~n29089 & n29090 ;
  assign n29092 = n5234 & n22381 ;
  assign n29093 = n5237 & ~n22398 ;
  assign n29094 = n5231 & ~n22385 ;
  assign n29095 = n29093 | n29094 ;
  assign n29096 = n29092 | n29095 ;
  assign n29097 = n5227 | n29096 ;
  assign n29098 = x14 & n29097 ;
  assign n29099 = x14 & n29096 ;
  assign n29100 = ( n22422 & n29098 ) | ( n22422 & n29099 ) | ( n29098 & n29099 ) ;
  assign n29101 = x14 | n29097 ;
  assign n29102 = x14 | n29096 ;
  assign n29103 = ( n22422 & n29101 ) | ( n22422 & n29102 ) | ( n29101 & n29102 ) ;
  assign n29104 = ~n29100 & n29103 ;
  assign n29105 = n29091 & n29104 ;
  assign n29106 = ~n29091 & n29104 ;
  assign n29107 = ( n29091 & ~n29105 ) | ( n29091 & n29106 ) | ( ~n29105 & n29106 ) ;
  assign n29108 = n27964 | n27966 ;
  assign n29109 = ~n27966 & n27968 ;
  assign n29110 = ( n27965 & n29108 ) | ( n27965 & ~n29109 ) | ( n29108 & ~n29109 ) ;
  assign n29111 = ~n27970 & n29110 ;
  assign n29112 = n5234 & ~n22385 ;
  assign n29113 = n5237 & n22393 ;
  assign n29114 = n5231 & ~n22398 ;
  assign n29115 = n29113 | n29114 ;
  assign n29116 = n29112 | n29115 ;
  assign n29117 = n5227 | n29112 ;
  assign n29118 = n29115 | n29117 ;
  assign n29119 = ( ~n22545 & n29116 ) | ( ~n22545 & n29118 ) | ( n29116 & n29118 ) ;
  assign n29120 = ~x14 & n29118 ;
  assign n29121 = ~x14 & n29116 ;
  assign n29122 = ( ~n22545 & n29120 ) | ( ~n22545 & n29121 ) | ( n29120 & n29121 ) ;
  assign n29123 = x14 | n29121 ;
  assign n29124 = x14 | n29120 ;
  assign n29125 = ( ~n22545 & n29123 ) | ( ~n22545 & n29124 ) | ( n29123 & n29124 ) ;
  assign n29126 = ( ~n29119 & n29122 ) | ( ~n29119 & n29125 ) | ( n29122 & n29125 ) ;
  assign n29127 = n29111 & n29126 ;
  assign n29128 = n5227 & n22474 ;
  assign n29129 = n5231 & ~n22409 ;
  assign n29130 = n5234 & ~n22406 ;
  assign n29131 = n29129 | n29130 ;
  assign n29132 = x14 | n29131 ;
  assign n29133 = n29128 | n29132 ;
  assign n29134 = ~x14 & n29133 ;
  assign n29135 = ( x14 & n17563 ) | ( x14 & n22409 ) | ( n17563 & n22409 ) ;
  assign n29136 = n29133 & n29135 ;
  assign n29137 = n29128 | n29131 ;
  assign n29138 = n29135 & ~n29137 ;
  assign n29139 = ( n29134 & n29136 ) | ( n29134 & n29138 ) | ( n29136 & n29138 ) ;
  assign n29140 = n5234 & n22393 ;
  assign n29141 = n5237 & ~n22409 ;
  assign n29142 = n5231 & ~n22406 ;
  assign n29143 = n29141 | n29142 ;
  assign n29144 = n29140 | n29143 ;
  assign n29145 = n22439 | n29144 ;
  assign n29146 = n5227 | n29140 ;
  assign n29147 = n29143 | n29146 ;
  assign n29148 = ~x14 & n29147 ;
  assign n29149 = n29145 & n29148 ;
  assign n29150 = x14 | n29149 ;
  assign n29151 = n4461 & ~n22409 ;
  assign n29152 = n29149 & n29151 ;
  assign n29153 = n29145 & n29147 ;
  assign n29154 = n29151 & ~n29153 ;
  assign n29155 = ( n29150 & n29152 ) | ( n29150 & n29154 ) | ( n29152 & n29154 ) ;
  assign n29156 = n29139 & n29155 ;
  assign n29157 = ( n29149 & n29150 ) | ( n29149 & ~n29153 ) | ( n29150 & ~n29153 ) ;
  assign n29158 = n29139 | n29151 ;
  assign n29159 = ( n29151 & n29157 ) | ( n29151 & n29158 ) | ( n29157 & n29158 ) ;
  assign n29160 = ~n29156 & n29159 ;
  assign n29161 = n5237 & ~n22406 ;
  assign n29162 = n5231 & n22393 ;
  assign n29163 = n29161 | n29162 ;
  assign n29164 = n5234 & ~n22398 ;
  assign n29165 = n5227 | n29164 ;
  assign n29166 = n29163 | n29165 ;
  assign n29167 = x14 & n29166 ;
  assign n29168 = n29163 | n29164 ;
  assign n29169 = x14 & n29168 ;
  assign n29170 = ( n22608 & n29167 ) | ( n22608 & n29169 ) | ( n29167 & n29169 ) ;
  assign n29171 = x14 | n29166 ;
  assign n29172 = x14 | n29168 ;
  assign n29173 = ( n22608 & n29171 ) | ( n22608 & n29172 ) | ( n29171 & n29172 ) ;
  assign n29174 = ~n29170 & n29173 ;
  assign n29175 = n29156 | n29174 ;
  assign n29176 = ( n29156 & n29160 ) | ( n29156 & n29175 ) | ( n29160 & n29175 ) ;
  assign n29177 = n29111 | n29126 ;
  assign n29178 = ~n29127 & n29177 ;
  assign n29179 = n29127 | n29178 ;
  assign n29180 = ( n29127 & n29176 ) | ( n29127 & n29179 ) | ( n29176 & n29179 ) ;
  assign n29181 = n29107 & n29180 ;
  assign n29182 = n29105 | n29181 ;
  assign n29183 = n29088 & n29182 ;
  assign n29184 = n29085 | n29183 ;
  assign n29185 = n5237 & n22381 ;
  assign n29186 = ( n5231 & n5357 ) | ( n5231 & n22381 ) | ( n5357 & n22381 ) ;
  assign n29187 = ( n23620 & n29185 ) | ( n23620 & n29186 ) | ( n29185 & n29186 ) ;
  assign n29188 = n5234 | n29186 ;
  assign n29189 = n5234 | n29185 ;
  assign n29190 = ( n23620 & n29188 ) | ( n23620 & n29189 ) | ( n29188 & n29189 ) ;
  assign n29191 = ( n23316 & n29187 ) | ( n23316 & n29190 ) | ( n29187 & n29190 ) ;
  assign n29192 = n5227 | n29191 ;
  assign n29193 = ~x14 & n29192 ;
  assign n29194 = ~x14 & n29191 ;
  assign n29195 = ( n23661 & n29193 ) | ( n23661 & n29194 ) | ( n29193 & n29194 ) ;
  assign n29196 = ( x14 & n17523 ) | ( x14 & n29191 ) | ( n17523 & n29191 ) ;
  assign n29197 = x14 & ~n29196 ;
  assign n29198 = x14 & n29191 ;
  assign n29199 = x14 & ~n29198 ;
  assign n29200 = ( ~n23661 & n29197 ) | ( ~n23661 & n29199 ) | ( n29197 & n29199 ) ;
  assign n29201 = n29195 | n29200 ;
  assign n29202 = n28007 & n28009 ;
  assign n29203 = n28007 | n28009 ;
  assign n29204 = ~n29202 & n29203 ;
  assign n29205 = n29201 & n29204 ;
  assign n29206 = n29201 | n29204 ;
  assign n29207 = ~n29205 & n29206 ;
  assign n29208 = n29205 | n29207 ;
  assign n29209 = ( n29184 & n29205 ) | ( n29184 & n29208 ) | ( n29205 & n29208 ) ;
  assign n29210 = n29066 & n29209 ;
  assign n29211 = n29063 | n29210 ;
  assign n29212 = ~n29008 & n29020 ;
  assign n29213 = ( n29008 & ~n29021 ) | ( n29008 & n29212 ) | ( ~n29021 & n29212 ) ;
  assign n29214 = n29211 & n29213 ;
  assign n29215 = n29040 | n29214 ;
  assign n29216 = ( n29043 & n29044 ) | ( n29043 & n29215 ) | ( n29044 & n29215 ) ;
  assign n29217 = n29003 | n29216 ;
  assign n29218 = ( n29003 & n29006 ) | ( n29003 & n29217 ) | ( n29006 & n29217 ) ;
  assign n29219 = n28985 & n29218 ;
  assign n29220 = n28981 | n29219 ;
  assign n29221 = ~n28946 & n28960 ;
  assign n29222 = ( n28946 & ~n28961 ) | ( n28946 & n29221 ) | ( ~n28961 & n29221 ) ;
  assign n29223 = n28961 | n29222 ;
  assign n29224 = ( n28961 & n29220 ) | ( n28961 & n29223 ) | ( n29220 & n29223 ) ;
  assign n29225 = n28939 | n29224 ;
  assign n29226 = ( n28939 & n28942 ) | ( n28939 & n29225 ) | ( n28942 & n29225 ) ;
  assign n29227 = n28922 & n29226 ;
  assign n29228 = n28919 | n29227 ;
  assign n29229 = n28882 | n28898 ;
  assign n29230 = ~n28899 & n29229 ;
  assign n29231 = n28899 | n29230 ;
  assign n29232 = ( n28899 & n29228 ) | ( n28899 & n29231 ) | ( n29228 & n29231 ) ;
  assign n29233 = n28879 & n29232 ;
  assign n29234 = n28877 | n29233 ;
  assign n29235 = ~n28838 & n28856 ;
  assign n29236 = ( n28838 & ~n28857 ) | ( n28838 & n29235 ) | ( ~n28857 & n29235 ) ;
  assign n29237 = n28857 | n29236 ;
  assign n29238 = ( n28857 & n29234 ) | ( n28857 & n29237 ) | ( n29234 & n29237 ) ;
  assign n29239 = n28832 | n29238 ;
  assign n29240 = ( n28832 & ~n28835 ) | ( n28832 & n29239 ) | ( ~n28835 & n29239 ) ;
  assign n29241 = n28805 | n29240 ;
  assign n29242 = ( n28805 & ~n28808 ) | ( n28805 & n29241 ) | ( ~n28808 & n29241 ) ;
  assign n29243 = n28767 | n29242 ;
  assign n29244 = ( n28767 & n28770 ) | ( n28767 & n29243 ) | ( n28770 & n29243 ) ;
  assign n29245 = ~n28742 & n29244 ;
  assign n29246 = n28739 | n29245 ;
  assign n29247 = ~n26565 & n26908 ;
  assign n29248 = n26562 | n29247 ;
  assign n29357 = ~n25431 & n25434 ;
  assign n29358 = ( n25329 & n25431 ) | ( n25329 & ~n29357 ) | ( n25431 & ~n29357 ) ;
  assign n29249 = n1829 & n23614 ;
  assign n29250 = n1826 & n23620 ;
  assign n29251 = ( n1823 & n13998 ) | ( n1823 & n23620 ) | ( n13998 & n23620 ) ;
  assign n29252 = ( n23316 & n29250 ) | ( n23316 & n29251 ) | ( n29250 & n29251 ) ;
  assign n29253 = n1821 | n29252 ;
  assign n29254 = n29249 | n29253 ;
  assign n29255 = ~x29 & n29254 ;
  assign n29256 = n29249 | n29252 ;
  assign n29257 = ~x29 & n29256 ;
  assign n29258 = ( n23634 & n29255 ) | ( n23634 & n29257 ) | ( n29255 & n29257 ) ;
  assign n29259 = x29 & n29254 ;
  assign n29260 = x29 & ~n29259 ;
  assign n29261 = x29 & n29252 ;
  assign n29262 = ( x29 & n29249 ) | ( x29 & n29261 ) | ( n29249 & n29261 ) ;
  assign n29263 = x29 & ~n29262 ;
  assign n29264 = ( ~n23634 & n29260 ) | ( ~n23634 & n29263 ) | ( n29260 & n29263 ) ;
  assign n29265 = n29258 | n29264 ;
  assign n29266 = ~n25402 & n25404 ;
  assign n29267 = n25397 | n29266 ;
  assign n29268 = n1057 & n22381 ;
  assign n29269 = n1065 & ~n22385 ;
  assign n29270 = n1060 & ~n22398 ;
  assign n29271 = n29269 | n29270 ;
  assign n29272 = n29268 | n29271 ;
  assign n29273 = n1062 | n29271 ;
  assign n29274 = n29268 | n29273 ;
  assign n29275 = ( n22422 & n29272 ) | ( n22422 & n29274 ) | ( n29272 & n29274 ) ;
  assign n29276 = n213 | n284 ;
  assign n29277 = n64 | n416 ;
  assign n29278 = n29276 | n29277 ;
  assign n29279 = n413 | n468 ;
  assign n29280 = n878 | n29279 ;
  assign n29281 = n29278 | n29280 ;
  assign n29282 = n581 | n29281 ;
  assign n29283 = n12274 | n22450 ;
  assign n29284 = n317 | n806 ;
  assign n29285 = n387 | n457 ;
  assign n29286 = n29284 | n29285 ;
  assign n29287 = n356 | n518 ;
  assign n29288 = n29286 | n29287 ;
  assign n29289 = ( ~n14381 & n29283 ) | ( ~n14381 & n29288 ) | ( n29283 & n29288 ) ;
  assign n29290 = n648 | n3431 ;
  assign n29291 = n179 | n29290 ;
  assign n29292 = n11407 | n29291 ;
  assign n29293 = n14381 | n29292 ;
  assign n29294 = n29289 | n29293 ;
  assign n29295 = n29282 | n29294 ;
  assign n29296 = n261 | n412 ;
  assign n29297 = n926 & ~n29296 ;
  assign n29298 = n85 | n341 ;
  assign n29299 = n123 | n29298 ;
  assign n29300 = n29297 & ~n29299 ;
  assign n29301 = ~n99 & n29300 ;
  assign n29302 = n110 | n18434 ;
  assign n29303 = n15234 | n29302 ;
  assign n29304 = n371 | n1577 ;
  assign n29305 = n29303 | n29304 ;
  assign n29306 = n29301 & ~n29305 ;
  assign n29307 = ~n14401 & n29306 ;
  assign n29308 = n663 | n1657 ;
  assign n29309 = n967 | n29308 ;
  assign n29310 = n1251 | n29309 ;
  assign n29311 = n17914 | n29310 ;
  assign n29312 = n29307 & ~n29311 ;
  assign n29313 = ~n29295 & n29312 ;
  assign n29314 = n395 | n638 ;
  assign n29315 = n277 | n375 ;
  assign n29316 = n29314 | n29315 ;
  assign n29317 = n29313 & ~n29316 ;
  assign n29318 = n29272 & ~n29317 ;
  assign n29319 = n29268 & ~n29317 ;
  assign n29320 = ( n29273 & ~n29317 ) | ( n29273 & n29319 ) | ( ~n29317 & n29319 ) ;
  assign n29321 = ( n22422 & n29318 ) | ( n22422 & n29320 ) | ( n29318 & n29320 ) ;
  assign n29322 = n29275 & ~n29321 ;
  assign n29323 = n29274 | n29317 ;
  assign n29324 = n29272 | n29317 ;
  assign n29325 = ( n22422 & n29323 ) | ( n22422 & n29324 ) | ( n29323 & n29324 ) ;
  assign n29326 = ~n29322 & n29325 ;
  assign n29327 = n29267 & ~n29326 ;
  assign n29328 = n29267 & ~n29327 ;
  assign n29329 = n29267 | n29326 ;
  assign n29330 = ~n29328 & n29329 ;
  assign n29331 = n29265 & ~n29330 ;
  assign n29332 = ~n29265 & n29330 ;
  assign n29333 = n29331 | n29332 ;
  assign n29334 = ~n25408 & n25410 ;
  assign n29335 = ( n25408 & n25412 ) | ( n25408 & ~n29334 ) | ( n25412 & ~n29334 ) ;
  assign n29336 = n29333 & ~n29335 ;
  assign n29337 = ~n29333 & n29335 ;
  assign n29338 = n29336 | n29337 ;
  assign n29339 = n2315 & n24770 ;
  assign n29340 = n2312 & n24167 ;
  assign n29341 = n2308 & ~n25054 ;
  assign n29342 = n29340 | n29341 ;
  assign n29343 = n29339 | n29342 ;
  assign n29344 = n2306 | n29343 ;
  assign n29345 = ( ~n25095 & n29343 ) | ( ~n25095 & n29344 ) | ( n29343 & n29344 ) ;
  assign n29346 = ~x26 & n29344 ;
  assign n29347 = ~x26 & n29343 ;
  assign n29348 = ( ~n25095 & n29346 ) | ( ~n25095 & n29347 ) | ( n29346 & n29347 ) ;
  assign n29349 = x26 | n29346 ;
  assign n29350 = x26 | n29347 ;
  assign n29351 = ( ~n25095 & n29349 ) | ( ~n25095 & n29350 ) | ( n29349 & n29350 ) ;
  assign n29352 = ( ~n29345 & n29348 ) | ( ~n29345 & n29351 ) | ( n29348 & n29351 ) ;
  assign n29353 = ~n29338 & n29352 ;
  assign n29354 = n29338 | n29353 ;
  assign n29355 = n29338 & n29352 ;
  assign n29356 = n29354 & ~n29355 ;
  assign n29359 = ~n29356 & n29358 ;
  assign n29360 = n29358 & ~n29359 ;
  assign n29361 = n29356 | n29358 ;
  assign n29362 = ~n29360 & n29361 ;
  assign n29363 = n2932 & n26017 ;
  assign n29364 = n2925 & ~n25046 ;
  assign n29365 = n2928 & ~n25728 ;
  assign n29366 = n29364 | n29365 ;
  assign n29367 = n29363 | n29366 ;
  assign n29368 = n2936 | n29363 ;
  assign n29369 = n29366 | n29368 ;
  assign n29370 = ( n26613 & n29367 ) | ( n26613 & n29369 ) | ( n29367 & n29369 ) ;
  assign n29371 = n29367 | n29369 ;
  assign n29372 = ( n26605 & n29370 ) | ( n26605 & n29371 ) | ( n29370 & n29371 ) ;
  assign n29373 = x23 & n29372 ;
  assign n29374 = x23 & ~n29372 ;
  assign n29375 = ( n29372 & ~n29373 ) | ( n29372 & n29374 ) | ( ~n29373 & n29374 ) ;
  assign n29376 = ~n29361 & n29375 ;
  assign n29377 = ( n29360 & n29375 ) | ( n29360 & n29376 ) | ( n29375 & n29376 ) ;
  assign n29378 = n29362 | n29377 ;
  assign n29379 = n29361 & n29375 ;
  assign n29380 = ~n29360 & n29379 ;
  assign n29381 = n29378 & ~n29380 ;
  assign n29382 = n25750 | n25756 ;
  assign n29383 = n29381 & ~n29382 ;
  assign n29384 = ~n29381 & n29382 ;
  assign n29385 = n29383 | n29384 ;
  assign n29386 = n3544 & ~n26270 ;
  assign n29387 = ~n26263 & n29386 ;
  assign n29388 = n3541 & ~n26526 ;
  assign n29389 = ~n26520 & n29388 ;
  assign n29390 = n29387 | n29389 ;
  assign n29391 = n3547 & ~n27133 ;
  assign n29392 = ~n27125 & n29391 ;
  assign n29393 = n29390 | n29392 ;
  assign n29394 = n27699 | n29393 ;
  assign n29395 = n27696 & ~n29394 ;
  assign n29396 = n3537 | n29392 ;
  assign n29397 = n29390 | n29396 ;
  assign n29398 = ~n29395 & n29397 ;
  assign n29399 = x20 & n29397 ;
  assign n29400 = ~n29395 & n29399 ;
  assign n29401 = x20 & ~n29399 ;
  assign n29402 = ( x20 & n29395 ) | ( x20 & n29401 ) | ( n29395 & n29401 ) ;
  assign n29403 = ( n29398 & ~n29400 ) | ( n29398 & n29402 ) | ( ~n29400 & n29402 ) ;
  assign n29404 = ~n29385 & n29403 ;
  assign n29405 = n29385 | n29404 ;
  assign n29406 = n29385 & n29403 ;
  assign n29407 = n29405 & ~n29406 ;
  assign n29408 = n29248 & ~n29407 ;
  assign n29409 = n29248 & ~n29408 ;
  assign n29410 = n29407 | n29408 ;
  assign n29411 = ~n29409 & n29410 ;
  assign n29412 = n4466 & ~n27371 ;
  assign n29413 = ~n27363 & n29412 ;
  assign n29414 = n4468 & ~n27606 ;
  assign n29415 = ~n27597 & n29414 ;
  assign n29416 = n29413 | n29415 ;
  assign n29417 = n4471 & ~n28503 ;
  assign n29418 = n28498 & n29417 ;
  assign n29419 = n29416 | n29418 ;
  assign n29420 = n4475 & n28794 ;
  assign n29421 = ( n4475 & n28783 ) | ( n4475 & n29420 ) | ( n28783 & n29420 ) ;
  assign n29422 = n29419 | n29421 ;
  assign n29423 = x17 | n29419 ;
  assign n29424 = n29421 | n29423 ;
  assign n29425 = ~x17 & n29423 ;
  assign n29426 = ( ~x17 & n29421 ) | ( ~x17 & n29425 ) | ( n29421 & n29425 ) ;
  assign n29427 = ( ~n29422 & n29424 ) | ( ~n29422 & n29426 ) | ( n29424 & n29426 ) ;
  assign n29428 = ~n29411 & n29427 ;
  assign n29429 = n29411 | n29428 ;
  assign n29430 = n29411 & n29427 ;
  assign n29431 = ~n27642 & n27644 ;
  assign n29432 = ( n27642 & n28071 ) | ( n27642 & ~n29431 ) | ( n28071 & ~n29431 ) ;
  assign n29433 = n29430 | n29432 ;
  assign n29434 = n29429 & ~n29433 ;
  assign n29435 = n29430 & n29432 ;
  assign n29436 = ( ~n29429 & n29432 ) | ( ~n29429 & n29435 ) | ( n29432 & n29435 ) ;
  assign n29437 = n29434 | n29436 ;
  assign n29438 = ~n28715 & n28717 ;
  assign n29439 = ( n28518 & n28730 ) | ( n28518 & ~n29438 ) | ( n28730 & ~n29438 ) ;
  assign n29440 = n28694 | n28698 ;
  assign n29441 = n28643 | n28649 ;
  assign n29442 = n858 | n2639 ;
  assign n29443 = n1239 | n29442 ;
  assign n29444 = n11750 | n29443 ;
  assign n29445 = n984 | n29444 ;
  assign n29446 = n1001 | n1013 ;
  assign n29447 = n539 | n703 ;
  assign n29448 = n29446 | n29447 ;
  assign n29449 = n190 | n197 ;
  assign n29450 = n263 | n29449 ;
  assign n29451 = n162 | n588 ;
  assign n29452 = n176 | n330 ;
  assign n29453 = n29451 | n29452 ;
  assign n29454 = n29450 | n29453 ;
  assign n29455 = n29448 | n29454 ;
  assign n29456 = n271 | n3495 ;
  assign n29457 = n679 | n29456 ;
  assign n29458 = n1307 | n29457 ;
  assign n29459 = n29455 | n29458 ;
  assign n29460 = n29445 | n29459 ;
  assign n29461 = n29295 | n29460 ;
  assign n29462 = n167 | n602 ;
  assign n29463 = n134 | n451 ;
  assign n29464 = n29462 | n29463 ;
  assign n29465 = n363 | n381 ;
  assign n29466 = n694 | n29465 ;
  assign n29467 = n29464 | n29466 ;
  assign n29468 = n29461 | n29467 ;
  assign n29469 = ( ~n28542 & n28544 ) | ( ~n28542 & n29468 ) | ( n28544 & n29468 ) ;
  assign n29470 = n28542 & ~n29468 ;
  assign n29471 = ( n28561 & n29469 ) | ( n28561 & ~n29470 ) | ( n29469 & ~n29470 ) ;
  assign n29472 = ~n28542 & n28544 ;
  assign n29473 = n29468 & n29472 ;
  assign n29474 = ~n28542 & n29468 ;
  assign n29475 = ( n28561 & n29473 ) | ( n28561 & n29474 ) | ( n29473 & n29474 ) ;
  assign n29476 = n29471 & ~n29475 ;
  assign n29477 = n1065 & ~n17092 ;
  assign n29478 = n1060 & n17100 ;
  assign n29479 = n29477 | n29478 ;
  assign n29480 = n1057 & n18037 ;
  assign n29481 = n1062 | n29480 ;
  assign n29482 = n29479 | n29481 ;
  assign n29483 = n29476 & n29482 ;
  assign n29484 = n29479 | n29480 ;
  assign n29485 = n29476 & n29484 ;
  assign n29486 = ( ~n18050 & n29483 ) | ( ~n18050 & n29485 ) | ( n29483 & n29485 ) ;
  assign n29487 = n29476 | n29482 ;
  assign n29488 = n29476 | n29484 ;
  assign n29489 = ( ~n18050 & n29487 ) | ( ~n18050 & n29488 ) | ( n29487 & n29488 ) ;
  assign n29490 = ~n29486 & n29489 ;
  assign n29491 = n28570 | n28580 ;
  assign n29492 = ( n28570 & n28572 ) | ( n28570 & n29491 ) | ( n28572 & n29491 ) ;
  assign n29493 = n29490 & n29492 ;
  assign n29494 = n29490 | n29492 ;
  assign n29495 = ~n29493 & n29494 ;
  assign n29497 = n1826 & ~n18585 ;
  assign n29498 = n1823 & n18410 ;
  assign n29499 = n29497 | n29498 ;
  assign n29496 = n1829 & n18576 ;
  assign n29501 = n1821 | n29496 ;
  assign n29502 = n29499 | n29501 ;
  assign n29500 = n29496 | n29499 ;
  assign n29503 = n29500 & n29502 ;
  assign n29504 = ( n18612 & n29502 ) | ( n18612 & n29503 ) | ( n29502 & n29503 ) ;
  assign n29505 = x29 & n29503 ;
  assign n29506 = x29 & n29502 ;
  assign n29507 = ( n18612 & n29505 ) | ( n18612 & n29506 ) | ( n29505 & n29506 ) ;
  assign n29508 = x29 & ~n29505 ;
  assign n29509 = x29 & ~n29506 ;
  assign n29510 = ( ~n18612 & n29508 ) | ( ~n18612 & n29509 ) | ( n29508 & n29509 ) ;
  assign n29511 = ( n29504 & ~n29507 ) | ( n29504 & n29510 ) | ( ~n29507 & n29510 ) ;
  assign n29512 = n29495 & n29511 ;
  assign n29513 = n29495 | n29511 ;
  assign n29514 = ~n29512 & n29513 ;
  assign n29515 = n28598 & n29514 ;
  assign n29516 = ( n28604 & n29514 ) | ( n28604 & n29515 ) | ( n29514 & n29515 ) ;
  assign n29517 = n28598 | n29514 ;
  assign n29518 = n28604 | n29517 ;
  assign n29519 = ~n29516 & n29518 ;
  assign n29520 = n2315 & n19631 ;
  assign n29521 = n2312 & n19352 ;
  assign n29522 = n2308 & n19494 ;
  assign n29523 = n29521 | n29522 ;
  assign n29524 = n29520 | n29523 ;
  assign n29525 = n2306 & n19652 ;
  assign n29526 = n2306 & n19655 ;
  assign n29527 = ( ~n18604 & n29525 ) | ( ~n18604 & n29526 ) | ( n29525 & n29526 ) ;
  assign n29528 = n29524 | n29527 ;
  assign n29529 = n2306 | n29524 ;
  assign n29530 = ( n19640 & n29528 ) | ( n19640 & n29529 ) | ( n29528 & n29529 ) ;
  assign n29531 = x26 | n29530 ;
  assign n29532 = ~x26 & n29530 ;
  assign n29533 = ( ~n29530 & n29531 ) | ( ~n29530 & n29532 ) | ( n29531 & n29532 ) ;
  assign n29534 = n29519 & ~n29533 ;
  assign n29535 = n29519 | n29533 ;
  assign n29536 = ( ~n29519 & n29534 ) | ( ~n29519 & n29535 ) | ( n29534 & n29535 ) ;
  assign n29537 = n28623 | n28627 ;
  assign n29538 = ( n28623 & ~n28626 ) | ( n28623 & n29537 ) | ( ~n28626 & n29537 ) ;
  assign n29539 = n29536 & n29538 ;
  assign n29540 = n29536 | n29538 ;
  assign n29541 = ~n29539 & n29540 ;
  assign n29542 = n2932 & n20609 ;
  assign n29543 = n2925 & ~n20630 ;
  assign n29544 = n2928 & ~n20618 ;
  assign n29545 = n29543 | n29544 ;
  assign n29546 = n29542 | n29545 ;
  assign n29547 = n2936 | n29542 ;
  assign n29548 = n29545 | n29547 ;
  assign n29549 = ( n20659 & n29546 ) | ( n20659 & n29548 ) | ( n29546 & n29548 ) ;
  assign n29550 = n29546 & n29548 ;
  assign n29551 = ( ~n20649 & n29549 ) | ( ~n20649 & n29550 ) | ( n29549 & n29550 ) ;
  assign n29552 = x23 & n29551 ;
  assign n29553 = x23 & ~n29551 ;
  assign n29554 = ( n29551 & ~n29552 ) | ( n29551 & n29553 ) | ( ~n29552 & n29553 ) ;
  assign n29555 = n29541 & ~n29554 ;
  assign n29556 = n29541 | n29554 ;
  assign n29557 = ( ~n29541 & n29555 ) | ( ~n29541 & n29556 ) | ( n29555 & n29556 ) ;
  assign n29558 = n29441 & n29557 ;
  assign n29559 = n29441 | n29557 ;
  assign n29560 = ~n29558 & n29559 ;
  assign n29561 = n3547 & ~n21551 ;
  assign n29562 = n3544 & ~n21563 ;
  assign n29563 = n3541 & ~n21517 ;
  assign n29564 = n29562 | n29563 ;
  assign n29565 = n29561 | n29564 ;
  assign n29566 = n3537 | n29561 ;
  assign n29567 = n29564 | n29566 ;
  assign n29568 = ( ~n21587 & n29565 ) | ( ~n21587 & n29567 ) | ( n29565 & n29567 ) ;
  assign n29569 = ~x20 & n29567 ;
  assign n29570 = ~x20 & n29565 ;
  assign n29571 = ( ~n21587 & n29569 ) | ( ~n21587 & n29570 ) | ( n29569 & n29570 ) ;
  assign n29572 = x20 | n29570 ;
  assign n29573 = x20 | n29569 ;
  assign n29574 = ( ~n21587 & n29572 ) | ( ~n21587 & n29573 ) | ( n29572 & n29573 ) ;
  assign n29575 = ( ~n29568 & n29571 ) | ( ~n29568 & n29574 ) | ( n29571 & n29574 ) ;
  assign n29576 = n29560 & ~n29575 ;
  assign n29577 = n29560 | n29575 ;
  assign n29578 = ( ~n29560 & n29576 ) | ( ~n29560 & n29577 ) | ( n29576 & n29577 ) ;
  assign n29579 = n28666 | n28672 ;
  assign n29580 = n29578 & n29579 ;
  assign n29581 = n29578 | n29579 ;
  assign n29582 = ~n29580 & n29581 ;
  assign n29583 = n4468 & ~n23240 ;
  assign n29584 = n4466 & n23227 ;
  assign n29585 = ( n4466 & n23217 ) | ( n4466 & n29584 ) | ( n23217 & n29584 ) ;
  assign n29586 = n29583 | n29585 ;
  assign n29587 = n4471 & ~n23234 ;
  assign n29588 = n4471 & ~n23235 ;
  assign n29589 = ( ~n15882 & n29587 ) | ( ~n15882 & n29588 ) | ( n29587 & n29588 ) ;
  assign n29590 = n29586 | n29589 ;
  assign n29591 = n4475 | n29589 ;
  assign n29592 = n29586 | n29591 ;
  assign n29593 = ( ~n23587 & n29590 ) | ( ~n23587 & n29592 ) | ( n29590 & n29592 ) ;
  assign n29594 = ~x17 & n29592 ;
  assign n29595 = ~x17 & n29590 ;
  assign n29596 = ( ~n23587 & n29594 ) | ( ~n23587 & n29595 ) | ( n29594 & n29595 ) ;
  assign n29597 = x17 | n29595 ;
  assign n29598 = x17 | n29594 ;
  assign n29599 = ( ~n23587 & n29597 ) | ( ~n23587 & n29598 ) | ( n29597 & n29598 ) ;
  assign n29600 = ( ~n29593 & n29596 ) | ( ~n29593 & n29599 ) | ( n29596 & n29599 ) ;
  assign n29601 = n29582 & ~n29600 ;
  assign n29602 = n29582 | n29600 ;
  assign n29603 = ( ~n29582 & n29601 ) | ( ~n29582 & n29602 ) | ( n29601 & n29602 ) ;
  assign n29604 = n29440 & n29603 ;
  assign n29605 = n29440 & ~n29604 ;
  assign n29606 = ~n29440 & n29603 ;
  assign n29607 = n29605 | n29606 ;
  assign n29608 = ~n28704 & n28706 ;
  assign n29609 = ( n28463 & n28704 ) | ( n28463 & ~n29608 ) | ( n28704 & ~n29608 ) ;
  assign n29610 = n29607 & n29609 ;
  assign n29611 = n29607 & ~n29608 ;
  assign n29612 = ( n28465 & n29610 ) | ( n28465 & n29611 ) | ( n29610 & n29611 ) ;
  assign n29613 = n29610 & n29611 ;
  assign n29614 = ( n28489 & n29612 ) | ( n28489 & n29613 ) | ( n29612 & n29613 ) ;
  assign n29615 = ~n29608 & n29609 ;
  assign n29616 = n29607 | n29615 ;
  assign n29617 = ( n28465 & ~n29608 ) | ( n28465 & n29609 ) | ( ~n29608 & n29609 ) ;
  assign n29618 = n29607 | n29617 ;
  assign n29619 = ( n28489 & n29616 ) | ( n28489 & n29618 ) | ( n29616 & n29618 ) ;
  assign n29620 = ~n29614 & n29619 ;
  assign n29621 = ~n28714 & n29620 ;
  assign n29622 = n28714 & ~n29620 ;
  assign n29623 = n28715 & ~n29622 ;
  assign n29624 = ( n28717 & n29622 ) | ( n28717 & ~n29623 ) | ( n29622 & ~n29623 ) ;
  assign n29625 = n29621 | n29624 ;
  assign n29626 = n29621 | n29622 ;
  assign n29627 = n28730 & ~n29626 ;
  assign n29628 = ( n28518 & ~n29625 ) | ( n28518 & n29627 ) | ( ~n29625 & n29627 ) ;
  assign n29629 = n29439 & ~n29628 ;
  assign n29631 = n5237 & n28492 ;
  assign n29632 = n5231 & ~n28714 ;
  assign n29633 = n29631 | n29632 ;
  assign n29630 = n5234 & n29620 ;
  assign n29635 = n5227 | n29630 ;
  assign n29636 = n29633 | n29635 ;
  assign n29634 = n29630 | n29633 ;
  assign n29637 = n29634 & n29636 ;
  assign n29638 = ~n29621 & n29625 ;
  assign n29639 = ~n29622 & n29638 ;
  assign n29640 = n29621 | n29627 ;
  assign n29641 = n29622 | n29640 ;
  assign n29642 = ( n28518 & ~n29639 ) | ( n28518 & n29641 ) | ( ~n29639 & n29641 ) ;
  assign n29643 = ( n29636 & n29637 ) | ( n29636 & ~n29642 ) | ( n29637 & ~n29642 ) ;
  assign n29644 = n29636 | n29637 ;
  assign n29645 = ( n29629 & n29643 ) | ( n29629 & n29644 ) | ( n29643 & n29644 ) ;
  assign n29646 = ~x14 & n29645 ;
  assign n29647 = x14 | n29645 ;
  assign n29648 = ( ~n29645 & n29646 ) | ( ~n29645 & n29647 ) | ( n29646 & n29647 ) ;
  assign n29649 = ~n29437 & n29648 ;
  assign n29650 = n29437 | n29649 ;
  assign n29651 = n29437 & n29648 ;
  assign n29652 = n29650 & ~n29651 ;
  assign n29653 = n29246 & ~n29652 ;
  assign n29654 = n29246 & ~n29653 ;
  assign n29655 = n29652 | n29653 ;
  assign n29656 = ~n29654 & n29655 ;
  assign n29657 = n29604 | n29607 ;
  assign n29658 = ( n29604 & n29609 ) | ( n29604 & n29657 ) | ( n29609 & n29657 ) ;
  assign n29659 = n29471 & ~n29476 ;
  assign n29660 = ( n29471 & ~n29482 ) | ( n29471 & n29659 ) | ( ~n29482 & n29659 ) ;
  assign n29661 = ( n29471 & ~n29484 ) | ( n29471 & n29659 ) | ( ~n29484 & n29659 ) ;
  assign n29662 = ( n18050 & n29660 ) | ( n18050 & n29661 ) | ( n29660 & n29661 ) ;
  assign n29663 = n331 | n477 ;
  assign n29664 = n12268 | n29663 ;
  assign n29665 = n206 | n280 ;
  assign n29666 = n103 | n29665 ;
  assign n29667 = n29664 | n29666 ;
  assign n29668 = n263 | n29667 ;
  assign n29669 = n1222 | n1335 ;
  assign n29670 = n242 | n29669 ;
  assign n29671 = ( n1756 & n29301 ) | ( n1756 & ~n29670 ) | ( n29301 & ~n29670 ) ;
  assign n29672 = n636 | n1756 ;
  assign n29673 = n29671 & ~n29672 ;
  assign n29674 = n1146 | n10379 ;
  assign n29675 = n575 | n29674 ;
  assign n29676 = n319 | n29675 ;
  assign n29677 = n13017 | n29676 ;
  assign n29678 = n16808 | n29677 ;
  assign n29679 = n29673 & ~n29678 ;
  assign n29680 = ~n29668 & n29679 ;
  assign n29681 = n29468 & n29680 ;
  assign n29682 = n29468 | n29680 ;
  assign n29683 = ~n29681 & n29682 ;
  assign n29684 = ~n29660 & n29683 ;
  assign n29685 = ~n29661 & n29683 ;
  assign n29686 = ( ~n18050 & n29684 ) | ( ~n18050 & n29685 ) | ( n29684 & n29685 ) ;
  assign n29687 = n29662 | n29686 ;
  assign n29688 = n29681 | n29683 ;
  assign n29689 = ( ~n29661 & n29681 ) | ( ~n29661 & n29688 ) | ( n29681 & n29688 ) ;
  assign n29690 = n29682 & ~n29689 ;
  assign n29691 = ( ~n29660 & n29681 ) | ( ~n29660 & n29688 ) | ( n29681 & n29688 ) ;
  assign n29692 = n29682 & ~n29691 ;
  assign n29693 = ( n18050 & n29690 ) | ( n18050 & n29692 ) | ( n29690 & n29692 ) ;
  assign n29694 = n29687 & ~n29693 ;
  assign n29695 = n1057 & ~n18585 ;
  assign n29696 = n1060 & ~n17092 ;
  assign n29697 = n1065 & n18037 ;
  assign n29698 = n29696 | n29697 ;
  assign n29699 = n29695 | n29698 ;
  assign n29700 = n1062 & ~n18675 ;
  assign n29701 = ( n1062 & n18672 ) | ( n1062 & n29700 ) | ( n18672 & n29700 ) ;
  assign n29702 = n29699 | n29701 ;
  assign n29703 = ~n29694 & n29702 ;
  assign n29704 = n29694 | n29703 ;
  assign n29706 = n1826 & n18410 ;
  assign n29707 = n1823 & n18576 ;
  assign n29708 = n29706 | n29707 ;
  assign n29705 = n1829 & n19352 ;
  assign n29710 = n1821 | n29705 ;
  assign n29711 = n29708 | n29710 ;
  assign n29709 = n29705 | n29708 ;
  assign n29712 = n29709 & n29711 ;
  assign n29713 = ( n19674 & n29711 ) | ( n19674 & n29712 ) | ( n29711 & n29712 ) ;
  assign n29714 = x29 & n29712 ;
  assign n29715 = x29 & n29711 ;
  assign n29716 = ( n19674 & n29714 ) | ( n19674 & n29715 ) | ( n29714 & n29715 ) ;
  assign n29717 = x29 & ~n29714 ;
  assign n29718 = x29 & ~n29715 ;
  assign n29719 = ( ~n19674 & n29717 ) | ( ~n19674 & n29718 ) | ( n29717 & n29718 ) ;
  assign n29720 = ( n29713 & ~n29716 ) | ( n29713 & n29719 ) | ( ~n29716 & n29719 ) ;
  assign n29721 = n29694 & n29702 ;
  assign n29722 = n29720 & n29721 ;
  assign n29723 = ( ~n29704 & n29720 ) | ( ~n29704 & n29722 ) | ( n29720 & n29722 ) ;
  assign n29724 = n29703 | n29723 ;
  assign n29725 = ( ~n18050 & n29689 ) | ( ~n18050 & n29691 ) | ( n29689 & n29691 ) ;
  assign n29726 = n1057 & n18410 ;
  assign n29727 = n1060 & n18037 ;
  assign n29728 = n1065 & ~n18585 ;
  assign n29729 = n29727 | n29728 ;
  assign n29730 = n29726 | n29729 ;
  assign n29731 = n1062 & ~n18586 ;
  assign n29732 = ~n18609 & n29731 ;
  assign n29733 = ( n1062 & n18650 ) | ( n1062 & n29732 ) | ( n18650 & n29732 ) ;
  assign n29734 = n29730 | n29733 ;
  assign n29735 = n988 | n25779 ;
  assign n29736 = n1265 | n20374 ;
  assign n29737 = n29735 | n29736 ;
  assign n29738 = n20370 | n29737 ;
  assign n29739 = n1364 | n13301 ;
  assign n29740 = n3995 | n18246 ;
  assign n29741 = n46 | n29740 ;
  assign n29742 = n29739 | n29741 ;
  assign n29743 = n720 | n895 ;
  assign n29744 = n154 | n374 ;
  assign n29745 = n29743 | n29744 ;
  assign n29746 = n676 | n29745 ;
  assign n29747 = n247 | n477 ;
  assign n29748 = n131 | n254 ;
  assign n29749 = n29747 | n29748 ;
  assign n29750 = n29746 | n29749 ;
  assign n29751 = n29742 | n29750 ;
  assign n29752 = n572 | n29751 ;
  assign n29753 = n29738 | n29752 ;
  assign n29754 = n15215 | n29753 ;
  assign n29755 = n498 | n3495 ;
  assign n29756 = n282 | n438 ;
  assign n29757 = n29755 | n29756 ;
  assign n29758 = n171 | n289 ;
  assign n29759 = n295 | n29758 ;
  assign n29760 = n758 | n29759 ;
  assign n29761 = n29757 | n29760 ;
  assign n29762 = n29754 | n29761 ;
  assign n29763 = ~n29680 & n29762 ;
  assign n29764 = n29680 & ~n29762 ;
  assign n29765 = n29763 | n29764 ;
  assign n29766 = n4468 | n4471 ;
  assign n29767 = n4466 | n29766 ;
  assign n29768 = n4475 | n29767 ;
  assign n29769 = ~n23229 & n29768 ;
  assign n29770 = ( n23154 & n29768 ) | ( n23154 & n29769 ) | ( n29768 & n29769 ) ;
  assign n29771 = ~n23232 & n29768 ;
  assign n29772 = ~n23231 & n29768 ;
  assign n29773 = ( n9072 & n29771 ) | ( n9072 & n29772 ) | ( n29771 & n29772 ) ;
  assign n29774 = ( ~n21543 & n29770 ) | ( ~n21543 & n29773 ) | ( n29770 & n29773 ) ;
  assign n29775 = ( ~n21545 & n29770 ) | ( ~n21545 & n29773 ) | ( n29770 & n29773 ) ;
  assign n29776 = ( ~n15882 & n29774 ) | ( ~n15882 & n29775 ) | ( n29774 & n29775 ) ;
  assign n29777 = ~x17 & n29774 ;
  assign n29778 = ~x17 & n29775 ;
  assign n29779 = ( ~n15882 & n29777 ) | ( ~n15882 & n29778 ) | ( n29777 & n29778 ) ;
  assign n29780 = x17 | n29777 ;
  assign n29781 = x17 | n29778 ;
  assign n29782 = ( ~n15882 & n29780 ) | ( ~n15882 & n29781 ) | ( n29780 & n29781 ) ;
  assign n29783 = ( ~n29776 & n29779 ) | ( ~n29776 & n29782 ) | ( n29779 & n29782 ) ;
  assign n29784 = n29765 | n29783 ;
  assign n29785 = n29765 & n29783 ;
  assign n29786 = n29784 & ~n29785 ;
  assign n29787 = n29730 & n29786 ;
  assign n29788 = ( n29733 & n29786 ) | ( n29733 & n29787 ) | ( n29786 & n29787 ) ;
  assign n29789 = n29734 & ~n29788 ;
  assign n29790 = ~n29730 & n29786 ;
  assign n29791 = ~n29733 & n29790 ;
  assign n29792 = n29725 & n29791 ;
  assign n29793 = ( n29725 & n29789 ) | ( n29725 & n29792 ) | ( n29789 & n29792 ) ;
  assign n29794 = n29725 | n29791 ;
  assign n29795 = n29789 | n29794 ;
  assign n29796 = ~n29793 & n29795 ;
  assign n29797 = n29703 & n29796 ;
  assign n29798 = ( n29723 & n29796 ) | ( n29723 & n29797 ) | ( n29796 & n29797 ) ;
  assign n29799 = n29724 & ~n29798 ;
  assign n29800 = n29796 & ~n29798 ;
  assign n29801 = n29799 | n29800 ;
  assign n29802 = n1829 & n19494 ;
  assign n29803 = n1826 & n18576 ;
  assign n29804 = n1823 & n19352 ;
  assign n29805 = n29803 | n29804 ;
  assign n29806 = n29802 | n29805 ;
  assign n29807 = n1821 | n29802 ;
  assign n29808 = n29805 | n29807 ;
  assign n29809 = ( n20320 & n29806 ) | ( n20320 & n29808 ) | ( n29806 & n29808 ) ;
  assign n29810 = x29 & n29808 ;
  assign n29811 = x29 & n29806 ;
  assign n29812 = ( n20320 & n29810 ) | ( n20320 & n29811 ) | ( n29810 & n29811 ) ;
  assign n29813 = x29 & ~n29811 ;
  assign n29814 = x29 & ~n29810 ;
  assign n29815 = ( ~n20320 & n29813 ) | ( ~n20320 & n29814 ) | ( n29813 & n29814 ) ;
  assign n29816 = ( n29809 & ~n29812 ) | ( n29809 & n29815 ) | ( ~n29812 & n29815 ) ;
  assign n29817 = ~n29801 & n29816 ;
  assign n29818 = n29801 & ~n29816 ;
  assign n29819 = n29817 | n29818 ;
  assign n29820 = n2306 & n20680 ;
  assign n29821 = n2315 & ~n20618 ;
  assign n29822 = n2312 & n19631 ;
  assign n29823 = n2308 & ~n20630 ;
  assign n29824 = n29822 | n29823 ;
  assign n29825 = n29821 | n29824 ;
  assign n29826 = n20689 | n29825 ;
  assign n29827 = n2306 | n29825 ;
  assign n29828 = ( n29820 & n29826 ) | ( n29820 & n29827 ) | ( n29826 & n29827 ) ;
  assign n29829 = x26 | n29828 ;
  assign n29830 = ~x26 & n29828 ;
  assign n29831 = ( ~n29828 & n29829 ) | ( ~n29828 & n29830 ) | ( n29829 & n29830 ) ;
  assign n29832 = n29819 & n29831 ;
  assign n29833 = n29819 | n29831 ;
  assign n29834 = ~n29832 & n29833 ;
  assign n29835 = n29720 | n29721 ;
  assign n29836 = n29704 & ~n29835 ;
  assign n29837 = n29723 | n29836 ;
  assign n29838 = n29493 | n29511 ;
  assign n29839 = ( n29493 & n29495 ) | ( n29493 & n29838 ) | ( n29495 & n29838 ) ;
  assign n29840 = ~n29837 & n29839 ;
  assign n29841 = n29837 & ~n29839 ;
  assign n29842 = n29840 | n29841 ;
  assign n29843 = n2315 & ~n20630 ;
  assign n29844 = n2312 & n19494 ;
  assign n29845 = n2308 & n19631 ;
  assign n29846 = n29844 | n29845 ;
  assign n29847 = n29843 | n29846 ;
  assign n29848 = n2306 | n29843 ;
  assign n29849 = n29846 | n29848 ;
  assign n29850 = ( ~n20709 & n29847 ) | ( ~n20709 & n29849 ) | ( n29847 & n29849 ) ;
  assign n29851 = ~x26 & n29849 ;
  assign n29852 = ~x26 & n29847 ;
  assign n29853 = ( ~n20709 & n29851 ) | ( ~n20709 & n29852 ) | ( n29851 & n29852 ) ;
  assign n29854 = x26 | n29852 ;
  assign n29855 = x26 | n29851 ;
  assign n29856 = ( ~n20709 & n29854 ) | ( ~n20709 & n29855 ) | ( n29854 & n29855 ) ;
  assign n29857 = ( ~n29850 & n29853 ) | ( ~n29850 & n29856 ) | ( n29853 & n29856 ) ;
  assign n29858 = n29840 | n29857 ;
  assign n29859 = ( n29840 & ~n29842 ) | ( n29840 & n29858 ) | ( ~n29842 & n29858 ) ;
  assign n29860 = n29834 & n29859 ;
  assign n29861 = n29834 | n29859 ;
  assign n29862 = ~n29860 & n29861 ;
  assign n29863 = n2932 & ~n21517 ;
  assign n29864 = n2925 & n20609 ;
  assign n29865 = n2928 & ~n21563 ;
  assign n29866 = n29864 | n29865 ;
  assign n29867 = n29863 | n29866 ;
  assign n29868 = n2936 | n29863 ;
  assign n29869 = n29866 | n29868 ;
  assign n29870 = ( ~n22283 & n29867 ) | ( ~n22283 & n29869 ) | ( n29867 & n29869 ) ;
  assign n29871 = n29867 & n29869 ;
  assign n29872 = ( ~n22271 & n29870 ) | ( ~n22271 & n29871 ) | ( n29870 & n29871 ) ;
  assign n29873 = ~x23 & n29872 ;
  assign n29874 = x23 | n29872 ;
  assign n29875 = ( ~n29872 & n29873 ) | ( ~n29872 & n29874 ) | ( n29873 & n29874 ) ;
  assign n29876 = n29862 & n29875 ;
  assign n29877 = n29862 & ~n29876 ;
  assign n29879 = n29842 | n29857 ;
  assign n29880 = n29842 & ~n29857 ;
  assign n29881 = ( ~n29842 & n29879 ) | ( ~n29842 & n29880 ) | ( n29879 & n29880 ) ;
  assign n29882 = n29516 | n29533 ;
  assign n29883 = ( n29516 & n29519 ) | ( n29516 & n29882 ) | ( n29519 & n29882 ) ;
  assign n29884 = ~n29881 & n29883 ;
  assign n29885 = n29881 & ~n29883 ;
  assign n29886 = n29884 | n29885 ;
  assign n29887 = n2932 & ~n21563 ;
  assign n29888 = n2925 & ~n20618 ;
  assign n29889 = n2928 & n20609 ;
  assign n29890 = n29888 | n29889 ;
  assign n29891 = n29887 | n29890 ;
  assign n29892 = n2936 & ~n21570 ;
  assign n29893 = n22270 & n29892 ;
  assign n29894 = ( n2936 & n22304 ) | ( n2936 & n29893 ) | ( n22304 & n29893 ) ;
  assign n29895 = n29891 | n29894 ;
  assign n29896 = x23 | n29891 ;
  assign n29897 = n29894 | n29896 ;
  assign n29898 = ~x23 & n29896 ;
  assign n29899 = ( ~x23 & n29894 ) | ( ~x23 & n29898 ) | ( n29894 & n29898 ) ;
  assign n29900 = ( ~n29895 & n29897 ) | ( ~n29895 & n29899 ) | ( n29897 & n29899 ) ;
  assign n29901 = n29884 | n29900 ;
  assign n29902 = ( n29884 & ~n29886 ) | ( n29884 & n29901 ) | ( ~n29886 & n29901 ) ;
  assign n29878 = ~n29862 & n29875 ;
  assign n29903 = n29878 & n29902 ;
  assign n29904 = ( n29877 & n29902 ) | ( n29877 & n29903 ) | ( n29902 & n29903 ) ;
  assign n29905 = n29876 | n29904 ;
  assign n29906 = n261 | n5038 ;
  assign n29907 = n13289 | n29906 ;
  assign n29908 = n133 | n330 ;
  assign n29909 = n1445 | n29908 ;
  assign n29910 = n381 | n401 ;
  assign n29911 = n347 | n29910 ;
  assign n29912 = n29909 | n29911 ;
  assign n29913 = n289 | n12280 ;
  assign n29914 = n29912 | n29913 ;
  assign n29915 = ( ~n25383 & n29907 ) | ( ~n25383 & n29914 ) | ( n29907 & n29914 ) ;
  assign n29916 = n25383 | n29915 ;
  assign n29917 = n441 | n839 ;
  assign n29918 = n458 | n29917 ;
  assign n29919 = ~n967 & n5878 ;
  assign n29920 = ~n29918 & n29919 ;
  assign n29921 = ~n448 & n29920 ;
  assign n29922 = n776 | n852 ;
  assign n29923 = n307 | n1483 ;
  assign n29924 = n29922 | n29923 ;
  assign n29925 = n1690 | n29924 ;
  assign n29926 = n29921 & ~n29925 ;
  assign n29927 = ( n528 & ~n29916 ) | ( n528 & n29926 ) | ( ~n29916 & n29926 ) ;
  assign n29928 = n29916 & ~n29926 ;
  assign n29929 = ( n586 & n29927 ) | ( n586 & ~n29928 ) | ( n29927 & ~n29928 ) ;
  assign n29930 = ~n587 & n29929 ;
  assign n29931 = n214 | n591 ;
  assign n29932 = n416 | n29931 ;
  assign n29933 = n29742 | n29746 ;
  assign n29934 = n1380 | n25375 ;
  assign n29935 = n29933 | n29934 ;
  assign n29936 = n168 | n14392 ;
  assign n29937 = n29935 | n29936 ;
  assign n29938 = n29932 | n29937 ;
  assign n29939 = n29930 & ~n29938 ;
  assign n29940 = ( n29763 & ~n29765 ) | ( n29763 & n29939 ) | ( ~n29765 & n29939 ) ;
  assign n29941 = n29763 & n29939 ;
  assign n29942 = ( ~n29783 & n29940 ) | ( ~n29783 & n29941 ) | ( n29940 & n29941 ) ;
  assign n29943 = ~n29763 & n29765 ;
  assign n29944 = ~n29939 & n29943 ;
  assign n29945 = n29763 | n29939 ;
  assign n29946 = ( n29783 & n29944 ) | ( n29783 & ~n29945 ) | ( n29944 & ~n29945 ) ;
  assign n29947 = n29942 | n29946 ;
  assign n29948 = n1065 & n18410 ;
  assign n29949 = n1060 & ~n18585 ;
  assign n29950 = n29948 | n29949 ;
  assign n29951 = n1057 & n18576 ;
  assign n29952 = n1062 | n29951 ;
  assign n29953 = n29950 | n29952 ;
  assign n29954 = ~n29947 & n29953 ;
  assign n29955 = n29950 | n29951 ;
  assign n29956 = ~n29947 & n29955 ;
  assign n29957 = ( n18612 & n29954 ) | ( n18612 & n29956 ) | ( n29954 & n29956 ) ;
  assign n29958 = n29947 & ~n29953 ;
  assign n29959 = n29947 & ~n29955 ;
  assign n29960 = ( ~n18612 & n29958 ) | ( ~n18612 & n29959 ) | ( n29958 & n29959 ) ;
  assign n29961 = n29957 | n29960 ;
  assign n29962 = n29788 & ~n29961 ;
  assign n29963 = ( n29793 & ~n29961 ) | ( n29793 & n29962 ) | ( ~n29961 & n29962 ) ;
  assign n29964 = ~n29788 & n29961 ;
  assign n29965 = ~n29793 & n29964 ;
  assign n29966 = n29963 | n29965 ;
  assign n29967 = n1826 & n19352 ;
  assign n29968 = n1823 & n19494 ;
  assign n29969 = n29967 | n29968 ;
  assign n29970 = n1829 & n19631 ;
  assign n29971 = n1821 | n29970 ;
  assign n29972 = n29969 | n29971 ;
  assign n29973 = n29969 | n29970 ;
  assign n29974 = n19652 | n29973 ;
  assign n29975 = n19655 | n29973 ;
  assign n29976 = ( ~n18604 & n29974 ) | ( ~n18604 & n29975 ) | ( n29974 & n29975 ) ;
  assign n29977 = n29972 & n29976 ;
  assign n29978 = ( n19640 & n29972 ) | ( n19640 & n29977 ) | ( n29972 & n29977 ) ;
  assign n29979 = ~x29 & n29978 ;
  assign n29980 = x29 | n29978 ;
  assign n29981 = ( ~n29978 & n29979 ) | ( ~n29978 & n29980 ) | ( n29979 & n29980 ) ;
  assign n29982 = ~n29966 & n29981 ;
  assign n29983 = n29966 & ~n29981 ;
  assign n29984 = n29982 | n29983 ;
  assign n29985 = n29798 | n29816 ;
  assign n29986 = ~n29984 & n29985 ;
  assign n29987 = n29798 & ~n29984 ;
  assign n29988 = ( n29801 & n29986 ) | ( n29801 & n29987 ) | ( n29986 & n29987 ) ;
  assign n29989 = n29984 & ~n29985 ;
  assign n29990 = ~n29798 & n29984 ;
  assign n29991 = ( ~n29801 & n29989 ) | ( ~n29801 & n29990 ) | ( n29989 & n29990 ) ;
  assign n29992 = n29988 | n29991 ;
  assign n29993 = n2315 & n20609 ;
  assign n29994 = n2312 & ~n20630 ;
  assign n29995 = n2308 & ~n20618 ;
  assign n29996 = n29994 | n29995 ;
  assign n29997 = n29993 | n29996 ;
  assign n29998 = n2306 | n29993 ;
  assign n29999 = n29996 | n29998 ;
  assign n30000 = ( n20659 & n29997 ) | ( n20659 & n29999 ) | ( n29997 & n29999 ) ;
  assign n30001 = n29997 & n29999 ;
  assign n30002 = ( ~n20649 & n30000 ) | ( ~n20649 & n30001 ) | ( n30000 & n30001 ) ;
  assign n30003 = x26 & n30002 ;
  assign n30004 = x26 & ~n30002 ;
  assign n30005 = ( n30002 & ~n30003 ) | ( n30002 & n30004 ) | ( ~n30003 & n30004 ) ;
  assign n30006 = n29992 | n30005 ;
  assign n30007 = n29992 & ~n30005 ;
  assign n30008 = ( ~n29992 & n30006 ) | ( ~n29992 & n30007 ) | ( n30006 & n30007 ) ;
  assign n30009 = n29832 | n29859 ;
  assign n30010 = ( n29832 & n29834 ) | ( n29832 & n30009 ) | ( n29834 & n30009 ) ;
  assign n30011 = ~n30008 & n30010 ;
  assign n30012 = n30008 & ~n30010 ;
  assign n30013 = n30011 | n30012 ;
  assign n30014 = n2932 & ~n21551 ;
  assign n30015 = n2925 & ~n21563 ;
  assign n30016 = n2928 & ~n21517 ;
  assign n30017 = n30015 | n30016 ;
  assign n30018 = n30014 | n30017 ;
  assign n30019 = n2936 | n30014 ;
  assign n30020 = n30017 | n30019 ;
  assign n30021 = ( ~n21587 & n30018 ) | ( ~n21587 & n30020 ) | ( n30018 & n30020 ) ;
  assign n30022 = ~x23 & n30020 ;
  assign n30023 = ~x23 & n30018 ;
  assign n30024 = ( ~n21587 & n30022 ) | ( ~n21587 & n30023 ) | ( n30022 & n30023 ) ;
  assign n30025 = x23 | n30023 ;
  assign n30026 = x23 | n30022 ;
  assign n30027 = ( ~n21587 & n30025 ) | ( ~n21587 & n30026 ) | ( n30025 & n30026 ) ;
  assign n30028 = ( ~n30021 & n30024 ) | ( ~n30021 & n30027 ) | ( n30024 & n30027 ) ;
  assign n30029 = n30013 | n30028 ;
  assign n30030 = n30013 & ~n30028 ;
  assign n30031 = ( ~n30013 & n30029 ) | ( ~n30013 & n30030 ) | ( n30029 & n30030 ) ;
  assign n30032 = n29905 & ~n30031 ;
  assign n30033 = ~n29905 & n30031 ;
  assign n30034 = n30032 | n30033 ;
  assign n30035 = n3541 & ~n23240 ;
  assign n30036 = n3544 & n23227 ;
  assign n30037 = ( n3544 & n23217 ) | ( n3544 & n30036 ) | ( n23217 & n30036 ) ;
  assign n30038 = n30035 | n30037 ;
  assign n30039 = n3547 & ~n23234 ;
  assign n30040 = n3547 & ~n23235 ;
  assign n30041 = ( ~n15882 & n30039 ) | ( ~n15882 & n30040 ) | ( n30039 & n30040 ) ;
  assign n30042 = n30038 | n30041 ;
  assign n30043 = n3537 | n30041 ;
  assign n30044 = n30038 | n30043 ;
  assign n30045 = ( ~n23587 & n30042 ) | ( ~n23587 & n30044 ) | ( n30042 & n30044 ) ;
  assign n30046 = ~x20 & n30044 ;
  assign n30047 = ~x20 & n30042 ;
  assign n30048 = ( ~n23587 & n30046 ) | ( ~n23587 & n30047 ) | ( n30046 & n30047 ) ;
  assign n30049 = x20 | n30047 ;
  assign n30050 = x20 | n30046 ;
  assign n30051 = ( ~n23587 & n30049 ) | ( ~n23587 & n30050 ) | ( n30049 & n30050 ) ;
  assign n30052 = ( ~n30045 & n30048 ) | ( ~n30045 & n30051 ) | ( n30048 & n30051 ) ;
  assign n30053 = n30034 | n30052 ;
  assign n30054 = n30034 & ~n30052 ;
  assign n30055 = ( ~n30034 & n30053 ) | ( ~n30034 & n30054 ) | ( n30053 & n30054 ) ;
  assign n30072 = n29886 | n29900 ;
  assign n30073 = n29886 & ~n29900 ;
  assign n30074 = ( ~n29886 & n30072 ) | ( ~n29886 & n30073 ) | ( n30072 & n30073 ) ;
  assign n30075 = n29539 | n29554 ;
  assign n30076 = ( n29539 & n29541 ) | ( n29539 & n30075 ) | ( n29541 & n30075 ) ;
  assign n30077 = ~n30074 & n30076 ;
  assign n30078 = n30074 & ~n30076 ;
  assign n30079 = n30077 | n30078 ;
  assign n30080 = n3544 & ~n21517 ;
  assign n30081 = n3541 & ~n21551 ;
  assign n30082 = n30080 | n30081 ;
  assign n30083 = n3547 & n23227 ;
  assign n30084 = ( n3547 & n23217 ) | ( n3547 & n30083 ) | ( n23217 & n30083 ) ;
  assign n30085 = n30082 | n30084 ;
  assign n30086 = n3537 & n23299 ;
  assign n30087 = n3537 & n23298 ;
  assign n30088 = ( n21584 & n30086 ) | ( n21584 & n30087 ) | ( n30086 & n30087 ) ;
  assign n30089 = n30085 | n30088 ;
  assign n30090 = n3537 | n30085 ;
  assign n30091 = ( n23289 & n30089 ) | ( n23289 & n30090 ) | ( n30089 & n30090 ) ;
  assign n30092 = x20 | n30091 ;
  assign n30093 = ~x20 & n30091 ;
  assign n30094 = ( ~n30091 & n30092 ) | ( ~n30091 & n30093 ) | ( n30092 & n30093 ) ;
  assign n30095 = n30077 | n30094 ;
  assign n30096 = ( n30077 & ~n30079 ) | ( n30077 & n30095 ) | ( ~n30079 & n30095 ) ;
  assign n30056 = n3547 & ~n23240 ;
  assign n30057 = n3544 & ~n21551 ;
  assign n30058 = n3541 & n23227 ;
  assign n30059 = ( n3541 & n23217 ) | ( n3541 & n30058 ) | ( n23217 & n30058 ) ;
  assign n30060 = n30057 | n30059 ;
  assign n30061 = n30056 | n30060 ;
  assign n30062 = n3537 | n30056 ;
  assign n30063 = n30060 | n30062 ;
  assign n30064 = ( n23260 & n30061 ) | ( n23260 & n30063 ) | ( n30061 & n30063 ) ;
  assign n30065 = x20 & n30063 ;
  assign n30066 = x20 & n30061 ;
  assign n30067 = ( n23260 & n30065 ) | ( n23260 & n30066 ) | ( n30065 & n30066 ) ;
  assign n30068 = x20 & ~n30066 ;
  assign n30069 = x20 & ~n30065 ;
  assign n30070 = ( ~n23260 & n30068 ) | ( ~n23260 & n30069 ) | ( n30068 & n30069 ) ;
  assign n30071 = ( n30064 & ~n30067 ) | ( n30064 & n30070 ) | ( ~n30067 & n30070 ) ;
  assign n30097 = n30071 & n30096 ;
  assign n30098 = n30096 & ~n30097 ;
  assign n30099 = n29878 | n29902 ;
  assign n30100 = n29877 | n30099 ;
  assign n30101 = ~n29904 & n30100 ;
  assign n30102 = n30071 & n30101 ;
  assign n30103 = ~n30096 & n30102 ;
  assign n30104 = n30097 | n30103 ;
  assign n30105 = n30097 | n30101 ;
  assign n30106 = ( n30098 & n30104 ) | ( n30098 & n30105 ) | ( n30104 & n30105 ) ;
  assign n30107 = ~n30055 & n30106 ;
  assign n30108 = n30055 | n30107 ;
  assign n30109 = n30055 & n30106 ;
  assign n30110 = n30108 & ~n30109 ;
  assign n30111 = ( n30098 & n30101 ) | ( n30098 & n30103 ) | ( n30101 & n30103 ) ;
  assign n30112 = n30071 | n30101 ;
  assign n30113 = ( ~n30096 & n30101 ) | ( ~n30096 & n30112 ) | ( n30101 & n30112 ) ;
  assign n30114 = n30098 | n30113 ;
  assign n30115 = ~n30111 & n30114 ;
  assign n30116 = ~n23234 & n29766 ;
  assign n30117 = n4466 | n30116 ;
  assign n30118 = ~n23235 & n29766 ;
  assign n30119 = n4466 | n30118 ;
  assign n30120 = ( ~n15882 & n30117 ) | ( ~n15882 & n30119 ) | ( n30117 & n30119 ) ;
  assign n30121 = n4475 | n30120 ;
  assign n30122 = ( ~n15882 & n30116 ) | ( ~n15882 & n30118 ) | ( n30116 & n30118 ) ;
  assign n30123 = n4475 | n30122 ;
  assign n30124 = ( ~n23240 & n30121 ) | ( ~n23240 & n30123 ) | ( n30121 & n30123 ) ;
  assign n30125 = ( ~n23240 & n30120 ) | ( ~n23240 & n30122 ) | ( n30120 & n30122 ) ;
  assign n30126 = n24135 & ~n30125 ;
  assign n30127 = n23240 & ~n30125 ;
  assign n30128 = ( n23575 & n30126 ) | ( n23575 & n30127 ) | ( n30126 & n30127 ) ;
  assign n30129 = ( n23577 & n30126 ) | ( n23577 & n30127 ) | ( n30126 & n30127 ) ;
  assign n30130 = ( ~n21554 & n30128 ) | ( ~n21554 & n30129 ) | ( n30128 & n30129 ) ;
  assign n30131 = n30124 & ~n30130 ;
  assign n30132 = x17 & ~n30131 ;
  assign n30133 = n30128 | n30129 ;
  assign n30134 = n30124 & ~n30133 ;
  assign n30135 = x17 & ~n30134 ;
  assign n30136 = ( n21584 & n30132 ) | ( n21584 & n30135 ) | ( n30132 & n30135 ) ;
  assign n30137 = ~x17 & n30131 ;
  assign n30138 = ~x17 & n30134 ;
  assign n30139 = ( ~n21584 & n30137 ) | ( ~n21584 & n30138 ) | ( n30137 & n30138 ) ;
  assign n30140 = n30136 | n30139 ;
  assign n30141 = n29558 | n29575 ;
  assign n30142 = ( n29558 & n29560 ) | ( n29558 & n30141 ) | ( n29560 & n30141 ) ;
  assign n30143 = n30140 & n30142 ;
  assign n30144 = n30140 | n30142 ;
  assign n30145 = ~n30143 & n30144 ;
  assign n30146 = n30079 | n30094 ;
  assign n30147 = n30079 & ~n30094 ;
  assign n30148 = ( ~n30079 & n30146 ) | ( ~n30079 & n30147 ) | ( n30146 & n30147 ) ;
  assign n30149 = ~n30143 & n30148 ;
  assign n30150 = ( n30143 & n30145 ) | ( n30143 & ~n30149 ) | ( n30145 & ~n30149 ) ;
  assign n30151 = n30115 & n30150 ;
  assign n30152 = n30115 | n30150 ;
  assign n30153 = ~n30151 & n30152 ;
  assign n30154 = n30145 & ~n30148 ;
  assign n30155 = n30145 | n30148 ;
  assign n30156 = ( ~n30145 & n30154 ) | ( ~n30145 & n30155 ) | ( n30154 & n30155 ) ;
  assign n30157 = n29580 | n29600 ;
  assign n30158 = ( n29580 & n29582 ) | ( n29580 & n30157 ) | ( n29582 & n30157 ) ;
  assign n30159 = ~n30156 & n30158 ;
  assign n30160 = n30156 & ~n30158 ;
  assign n30161 = n30159 | n30160 ;
  assign n30162 = ~n30159 & n30161 ;
  assign n30163 = n30153 & ~n30162 ;
  assign n30164 = n30151 | n30163 ;
  assign n30165 = ~n30110 & n30164 ;
  assign n30166 = n30153 & n30159 ;
  assign n30167 = n30151 | n30166 ;
  assign n30168 = ~n30110 & n30167 ;
  assign n30169 = ( n29658 & n30165 ) | ( n29658 & n30168 ) | ( n30165 & n30168 ) ;
  assign n30170 = n29604 & ~n30161 ;
  assign n30171 = n30159 | n30170 ;
  assign n30172 = n30153 & n30171 ;
  assign n30173 = ( n29611 & n30163 ) | ( n29611 & n30172 ) | ( n30163 & n30172 ) ;
  assign n30174 = ~n30110 & n30151 ;
  assign n30175 = ( ~n30110 & n30173 ) | ( ~n30110 & n30174 ) | ( n30173 & n30174 ) ;
  assign n30176 = ( n28465 & n30169 ) | ( n28465 & n30175 ) | ( n30169 & n30175 ) ;
  assign n30177 = n30169 & n30175 ;
  assign n30178 = ( n28489 & n30176 ) | ( n28489 & n30177 ) | ( n30176 & n30177 ) ;
  assign n30179 = n30151 | n30173 ;
  assign n30180 = ( n29658 & n30164 ) | ( n29658 & n30167 ) | ( n30164 & n30167 ) ;
  assign n30181 = n30179 & n30180 ;
  assign n30182 = n30110 & ~n30181 ;
  assign n30183 = ( n28465 & n30179 ) | ( n28465 & n30180 ) | ( n30179 & n30180 ) ;
  assign n30184 = n30110 & ~n30183 ;
  assign n30185 = ( ~n28489 & n30182 ) | ( ~n28489 & n30184 ) | ( n30182 & n30184 ) ;
  assign n30186 = n30178 | n30185 ;
  assign n30187 = n6122 & ~n30186 ;
  assign n30188 = n29658 & ~n30161 ;
  assign n30189 = ( n29611 & ~n30161 ) | ( n29611 & n30170 ) | ( ~n30161 & n30170 ) ;
  assign n30190 = ( n28465 & n30188 ) | ( n28465 & n30189 ) | ( n30188 & n30189 ) ;
  assign n30191 = n30188 & n30189 ;
  assign n30192 = ( n28489 & n30190 ) | ( n28489 & n30191 ) | ( n30190 & n30191 ) ;
  assign n30193 = n29604 | n29611 ;
  assign n30194 = n29658 & n30193 ;
  assign n30195 = n30161 & ~n30194 ;
  assign n30196 = ( n28465 & n29658 ) | ( n28465 & n30193 ) | ( n29658 & n30193 ) ;
  assign n30197 = n30161 & ~n30196 ;
  assign n30198 = ( ~n28489 & n30195 ) | ( ~n28489 & n30197 ) | ( n30195 & n30197 ) ;
  assign n30199 = n30192 | n30198 ;
  assign n30200 = n6125 & ~n30199 ;
  assign n30201 = ( n29658 & n30163 ) | ( n29658 & n30166 ) | ( n30163 & n30166 ) ;
  assign n30202 = ( n28465 & n30173 ) | ( n28465 & n30201 ) | ( n30173 & n30201 ) ;
  assign n30203 = n30173 & n30201 ;
  assign n30204 = ( n28489 & n30202 ) | ( n28489 & n30203 ) | ( n30202 & n30203 ) ;
  assign n30205 = ( n29658 & n30159 ) | ( n29658 & ~n30162 ) | ( n30159 & ~n30162 ) ;
  assign n30206 = ( n29611 & ~n30162 ) | ( n29611 & n30171 ) | ( ~n30162 & n30171 ) ;
  assign n30207 = n30205 & n30206 ;
  assign n30208 = n30153 | n30207 ;
  assign n30209 = ( n28465 & n30205 ) | ( n28465 & n30206 ) | ( n30205 & n30206 ) ;
  assign n30210 = n30153 | n30209 ;
  assign n30211 = ( n28489 & n30208 ) | ( n28489 & n30210 ) | ( n30208 & n30210 ) ;
  assign n30212 = ~n30204 & n30211 ;
  assign n30213 = n6119 & n30212 ;
  assign n30214 = n30200 | n30213 ;
  assign n30215 = n30187 | n30214 ;
  assign n30216 = ~n30186 & n30212 ;
  assign n30217 = n30186 & ~n30212 ;
  assign n30218 = n30199 & ~n30212 ;
  assign n30219 = n29620 & ~n30199 ;
  assign n30220 = ~n29620 & n30199 ;
  assign n30221 = n30219 | n30220 ;
  assign n30222 = ~n30218 & n30219 ;
  assign n30223 = ( n30218 & n30221 ) | ( n30218 & ~n30222 ) | ( n30221 & ~n30222 ) ;
  assign n30224 = ~n30199 & n30212 ;
  assign n30225 = ~n30217 & n30224 ;
  assign n30226 = ( n30217 & n30223 ) | ( n30217 & ~n30225 ) | ( n30223 & ~n30225 ) ;
  assign n30227 = ( ~n30217 & n30222 ) | ( ~n30217 & n30225 ) | ( n30222 & n30225 ) ;
  assign n30228 = ( n29640 & ~n30226 ) | ( n29640 & n30227 ) | ( ~n30226 & n30227 ) ;
  assign n30229 = ~n30216 & n30228 ;
  assign n30230 = ( n29638 & n30226 ) | ( n29638 & ~n30227 ) | ( n30226 & ~n30227 ) ;
  assign n30231 = n30216 | n30230 ;
  assign n30232 = ( n28518 & n30229 ) | ( n28518 & ~n30231 ) | ( n30229 & ~n30231 ) ;
  assign n30233 = n30216 | n30217 ;
  assign n30234 = n30223 & ~n30224 ;
  assign n30235 = n30222 | n30224 ;
  assign n30236 = ( n29640 & ~n30234 ) | ( n29640 & n30235 ) | ( ~n30234 & n30235 ) ;
  assign n30237 = n30233 & ~n30236 ;
  assign n30238 = ( n29638 & n30234 ) | ( n29638 & ~n30235 ) | ( n30234 & ~n30235 ) ;
  assign n30239 = n30233 & n30238 ;
  assign n30240 = ( ~n28518 & n30237 ) | ( ~n28518 & n30239 ) | ( n30237 & n30239 ) ;
  assign n30241 = n30232 | n30240 ;
  assign n30242 = n6115 | n30187 ;
  assign n30243 = n30214 | n30242 ;
  assign n30244 = ( n30215 & ~n30241 ) | ( n30215 & n30243 ) | ( ~n30241 & n30243 ) ;
  assign n30245 = ~x11 & n30243 ;
  assign n30246 = ~x11 & n30215 ;
  assign n30247 = ( ~n30241 & n30245 ) | ( ~n30241 & n30246 ) | ( n30245 & n30246 ) ;
  assign n30248 = x11 | n30246 ;
  assign n30249 = x11 | n30245 ;
  assign n30250 = ( ~n30241 & n30248 ) | ( ~n30241 & n30249 ) | ( n30248 & n30249 ) ;
  assign n30251 = ( ~n30244 & n30247 ) | ( ~n30244 & n30250 ) | ( n30247 & n30250 ) ;
  assign n30252 = ~n29656 & n30251 ;
  assign n30253 = n29656 | n30252 ;
  assign n30254 = n29656 & n30251 ;
  assign n30255 = n30253 & ~n30254 ;
  assign n30256 = n29244 & ~n29245 ;
  assign n30257 = n28742 | n29245 ;
  assign n30258 = ~n30256 & n30257 ;
  assign n30259 = n6122 & n30212 ;
  assign n30260 = n6125 & n29620 ;
  assign n30261 = n6119 & ~n30199 ;
  assign n30262 = n30260 | n30261 ;
  assign n30263 = n30259 | n30262 ;
  assign n30264 = n30218 | n30236 ;
  assign n30265 = ~n30218 & n30238 ;
  assign n30266 = ( n28518 & n30264 ) | ( n28518 & ~n30265 ) | ( n30264 & ~n30265 ) ;
  assign n30267 = n6115 & ~n30266 ;
  assign n30268 = n30223 | n30224 ;
  assign n30269 = n30222 & ~n30224 ;
  assign n30270 = ( n29638 & n30268 ) | ( n29638 & ~n30269 ) | ( n30268 & ~n30269 ) ;
  assign n30271 = ( n29640 & ~n30268 ) | ( n29640 & n30269 ) | ( ~n30268 & n30269 ) ;
  assign n30272 = ( n28518 & ~n30270 ) | ( n28518 & n30271 ) | ( ~n30270 & n30271 ) ;
  assign n30273 = n29638 | n30221 ;
  assign n30274 = n29640 & ~n30221 ;
  assign n30275 = ( n28518 & ~n30273 ) | ( n28518 & n30274 ) | ( ~n30273 & n30274 ) ;
  assign n30276 = ( n30219 & ~n30272 ) | ( n30219 & n30275 ) | ( ~n30272 & n30275 ) ;
  assign n30277 = ( n6115 & n30267 ) | ( n6115 & n30276 ) | ( n30267 & n30276 ) ;
  assign n30278 = n30263 | n30277 ;
  assign n30279 = x11 | n30263 ;
  assign n30280 = n30277 | n30279 ;
  assign n30281 = ~x11 & n30279 ;
  assign n30282 = ( ~x11 & n30277 ) | ( ~x11 & n30281 ) | ( n30277 & n30281 ) ;
  assign n30283 = ( ~n30278 & n30280 ) | ( ~n30278 & n30282 ) | ( n30280 & n30282 ) ;
  assign n30284 = ~n30258 & n30283 ;
  assign n30285 = n30258 | n30284 ;
  assign n30286 = n30258 & n30283 ;
  assign n30287 = n30285 & ~n30286 ;
  assign n30288 = ~n28770 & n29242 ;
  assign n30289 = n28770 & ~n29242 ;
  assign n30290 = n30288 | n30289 ;
  assign n30291 = n6122 & ~n30199 ;
  assign n30292 = n6125 & ~n28714 ;
  assign n30293 = n6119 & n29620 ;
  assign n30294 = n30292 | n30293 ;
  assign n30295 = n30291 | n30294 ;
  assign n30296 = n29638 & n30221 ;
  assign n30297 = ~n29640 & n30221 ;
  assign n30298 = ( ~n28518 & n30296 ) | ( ~n28518 & n30297 ) | ( n30296 & n30297 ) ;
  assign n30299 = n30275 | n30298 ;
  assign n30300 = n6115 | n30291 ;
  assign n30301 = n30294 | n30300 ;
  assign n30302 = ( n30295 & ~n30299 ) | ( n30295 & n30301 ) | ( ~n30299 & n30301 ) ;
  assign n30303 = ~x11 & n30301 ;
  assign n30304 = ~x11 & n30295 ;
  assign n30305 = ( ~n30299 & n30303 ) | ( ~n30299 & n30304 ) | ( n30303 & n30304 ) ;
  assign n30306 = x11 | n30304 ;
  assign n30307 = x11 | n30303 ;
  assign n30308 = ( ~n30299 & n30306 ) | ( ~n30299 & n30307 ) | ( n30306 & n30307 ) ;
  assign n30309 = ( ~n30302 & n30305 ) | ( ~n30302 & n30308 ) | ( n30305 & n30308 ) ;
  assign n30310 = n30290 & n30309 ;
  assign n30311 = n30290 | n30309 ;
  assign n30312 = ~n30310 & n30311 ;
  assign n30313 = n28808 & n29240 ;
  assign n30314 = n28808 | n29240 ;
  assign n30315 = ~n30313 & n30314 ;
  assign n30316 = n6122 & n29620 ;
  assign n30317 = n6125 & n28492 ;
  assign n30318 = n6119 & ~n28714 ;
  assign n30319 = n30317 | n30318 ;
  assign n30320 = n30316 | n30319 ;
  assign n30321 = n6115 | n30316 ;
  assign n30322 = n30319 | n30321 ;
  assign n30323 = ( ~n29642 & n30320 ) | ( ~n29642 & n30322 ) | ( n30320 & n30322 ) ;
  assign n30324 = n30320 | n30322 ;
  assign n30325 = ( n29629 & n30323 ) | ( n29629 & n30324 ) | ( n30323 & n30324 ) ;
  assign n30326 = ~x11 & n30325 ;
  assign n30327 = x11 | n30325 ;
  assign n30328 = ( ~n30325 & n30326 ) | ( ~n30325 & n30327 ) | ( n30326 & n30327 ) ;
  assign n30329 = ~n30315 & n30328 ;
  assign n30330 = n30315 & ~n30328 ;
  assign n30331 = n30329 | n30330 ;
  assign n30332 = ~n28835 & n29238 ;
  assign n30333 = n28835 | n30332 ;
  assign n30336 = n6122 & ~n28714 ;
  assign n30337 = n6119 & n28492 ;
  assign n30338 = n6125 & ~n28503 ;
  assign n30339 = n28498 & n30338 ;
  assign n30340 = n30337 | n30339 ;
  assign n30341 = n30336 | n30340 ;
  assign n30342 = n6115 & ~n28731 ;
  assign n30343 = ~n28518 & n30342 ;
  assign n30344 = n30341 | n30343 ;
  assign n30345 = n6115 | n30341 ;
  assign n30346 = ( n28720 & n30344 ) | ( n28720 & n30345 ) | ( n30344 & n30345 ) ;
  assign n30347 = x11 | n30346 ;
  assign n30348 = ~x11 & n30346 ;
  assign n30349 = ( ~n30346 & n30347 ) | ( ~n30346 & n30348 ) | ( n30347 & n30348 ) ;
  assign n30334 = n28835 & n29238 ;
  assign n30350 = n30334 & n30349 ;
  assign n30351 = ( ~n30333 & n30349 ) | ( ~n30333 & n30350 ) | ( n30349 & n30350 ) ;
  assign n30335 = n30333 & ~n30334 ;
  assign n30352 = n30335 | n30351 ;
  assign n30353 = ~n30334 & n30349 ;
  assign n30354 = n30333 & n30353 ;
  assign n30355 = n30352 & ~n30354 ;
  assign n30356 = n28879 | n29232 ;
  assign n30357 = ~n29233 & n30356 ;
  assign n30358 = n6125 & ~n27371 ;
  assign n30359 = ~n27363 & n30358 ;
  assign n30360 = n6119 & ~n27606 ;
  assign n30361 = ~n27597 & n30360 ;
  assign n30362 = n30359 | n30361 ;
  assign n30363 = n6122 & ~n28503 ;
  assign n30364 = n28498 & n30363 ;
  assign n30365 = n30362 | n30364 ;
  assign n30366 = n28794 | n30365 ;
  assign n30367 = n28783 | n30366 ;
  assign n30368 = n6115 | n30364 ;
  assign n30369 = n30362 | n30368 ;
  assign n30370 = n30367 & n30369 ;
  assign n30371 = ~x11 & n30369 ;
  assign n30372 = n30367 & n30371 ;
  assign n30373 = x11 | n30371 ;
  assign n30374 = ( x11 & n30367 ) | ( x11 & n30373 ) | ( n30367 & n30373 ) ;
  assign n30375 = ( ~n30370 & n30372 ) | ( ~n30370 & n30374 ) | ( n30372 & n30374 ) ;
  assign n30376 = n30357 & n30375 ;
  assign n30377 = n29234 & n29236 ;
  assign n30378 = n29234 | n29236 ;
  assign n30379 = ~n30377 & n30378 ;
  assign n30380 = n6122 & n28492 ;
  assign n30381 = n6125 & ~n27606 ;
  assign n30382 = ~n27597 & n30381 ;
  assign n30383 = n6119 & ~n28503 ;
  assign n30384 = n28498 & n30383 ;
  assign n30385 = n30382 | n30384 ;
  assign n30386 = n30380 | n30385 ;
  assign n30387 = n6115 | n30386 ;
  assign n30388 = n30386 & n30387 ;
  assign n30389 = ( ~n28749 & n30387 ) | ( ~n28749 & n30388 ) | ( n30387 & n30388 ) ;
  assign n30390 = ~x11 & n30388 ;
  assign n30391 = ~x11 & n30387 ;
  assign n30392 = ( ~n28749 & n30390 ) | ( ~n28749 & n30391 ) | ( n30390 & n30391 ) ;
  assign n30393 = x11 | n30390 ;
  assign n30394 = x11 | n30391 ;
  assign n30395 = ( ~n28749 & n30393 ) | ( ~n28749 & n30394 ) | ( n30393 & n30394 ) ;
  assign n30396 = ( ~n30389 & n30392 ) | ( ~n30389 & n30395 ) | ( n30392 & n30395 ) ;
  assign n30397 = n30379 & n30396 ;
  assign n30398 = n30379 | n30396 ;
  assign n30399 = ~n30397 & n30398 ;
  assign n30400 = n30376 & n30399 ;
  assign n30401 = n30397 | n30399 ;
  assign n30402 = n29228 & n29230 ;
  assign n30403 = n29228 | n29230 ;
  assign n30404 = ~n30402 & n30403 ;
  assign n30405 = n6125 & ~n27133 ;
  assign n30406 = ~n27125 & n30405 ;
  assign n30407 = n6119 & ~n27371 ;
  assign n30408 = ~n27363 & n30407 ;
  assign n30409 = n30406 | n30408 ;
  assign n30410 = n6122 & ~n27606 ;
  assign n30411 = ~n27597 & n30410 ;
  assign n30412 = n30409 | n30411 ;
  assign n30413 = n6115 & n27630 ;
  assign n30414 = ~n27625 & n30413 ;
  assign n30415 = ( n6115 & ~n27634 ) | ( n6115 & n30414 ) | ( ~n27634 & n30414 ) ;
  assign n30416 = n30412 | n30415 ;
  assign n30417 = x11 | n30412 ;
  assign n30418 = n30415 | n30417 ;
  assign n30419 = ~x11 & n30417 ;
  assign n30420 = ( ~x11 & n30415 ) | ( ~x11 & n30419 ) | ( n30415 & n30419 ) ;
  assign n30421 = ( ~n30416 & n30418 ) | ( ~n30416 & n30420 ) | ( n30418 & n30420 ) ;
  assign n30422 = n30404 & n30421 ;
  assign n30423 = ~n30404 & n30421 ;
  assign n30424 = ( n30404 & ~n30422 ) | ( n30404 & n30423 ) | ( ~n30422 & n30423 ) ;
  assign n30425 = ~n28922 & n29226 ;
  assign n30426 = n28922 & ~n29226 ;
  assign n30427 = n30425 | n30426 ;
  assign n30428 = n6125 & ~n26526 ;
  assign n30429 = ~n26520 & n30428 ;
  assign n30430 = n6119 & ~n27133 ;
  assign n30431 = ~n27125 & n30430 ;
  assign n30432 = n30429 | n30431 ;
  assign n30433 = n6122 & ~n27371 ;
  assign n30434 = ~n27363 & n30433 ;
  assign n30435 = n30432 | n30434 ;
  assign n30436 = n6115 | n30434 ;
  assign n30437 = n30432 | n30436 ;
  assign n30438 = ( ~n27654 & n30435 ) | ( ~n27654 & n30437 ) | ( n30435 & n30437 ) ;
  assign n30439 = ~x11 & n30437 ;
  assign n30440 = ~x11 & n30435 ;
  assign n30441 = ( ~n27654 & n30439 ) | ( ~n27654 & n30440 ) | ( n30439 & n30440 ) ;
  assign n30442 = x11 | n30440 ;
  assign n30443 = x11 | n30439 ;
  assign n30444 = ( ~n27654 & n30442 ) | ( ~n27654 & n30443 ) | ( n30442 & n30443 ) ;
  assign n30445 = ( ~n30438 & n30441 ) | ( ~n30438 & n30444 ) | ( n30441 & n30444 ) ;
  assign n30446 = n30427 & n30445 ;
  assign n30447 = ~n28942 & n29224 ;
  assign n30448 = n28942 & ~n29224 ;
  assign n30449 = n30447 | n30448 ;
  assign n30450 = n6125 & ~n26270 ;
  assign n30451 = ~n26263 & n30450 ;
  assign n30452 = n6119 & ~n26526 ;
  assign n30453 = ~n26520 & n30452 ;
  assign n30454 = n30451 | n30453 ;
  assign n30455 = n6122 & ~n27133 ;
  assign n30456 = ~n27125 & n30455 ;
  assign n30457 = n30454 | n30456 ;
  assign n30458 = n6115 & n27699 ;
  assign n30459 = ( n6115 & ~n27696 ) | ( n6115 & n30458 ) | ( ~n27696 & n30458 ) ;
  assign n30460 = n30457 | n30459 ;
  assign n30461 = x11 | n30457 ;
  assign n30462 = n30459 | n30461 ;
  assign n30463 = ~x11 & n30461 ;
  assign n30464 = ( ~x11 & n30459 ) | ( ~x11 & n30463 ) | ( n30459 & n30463 ) ;
  assign n30465 = ( ~n30460 & n30462 ) | ( ~n30460 & n30464 ) | ( n30462 & n30464 ) ;
  assign n30466 = n30449 & n30465 ;
  assign n30467 = n30449 | n30465 ;
  assign n30468 = ~n30466 & n30467 ;
  assign n30469 = n29220 & n29222 ;
  assign n30470 = n29220 | n29222 ;
  assign n30471 = ~n30469 & n30470 ;
  assign n30472 = n6125 & n26017 ;
  assign n30473 = n6119 & ~n26270 ;
  assign n30474 = ~n26263 & n30473 ;
  assign n30475 = n30472 | n30474 ;
  assign n30476 = n6122 & ~n26526 ;
  assign n30477 = ~n26520 & n30476 ;
  assign n30479 = n6115 | n30477 ;
  assign n30480 = n30475 | n30479 ;
  assign n30478 = n30475 | n30477 ;
  assign n30481 = n30478 & n30480 ;
  assign n30482 = ( ~n26555 & n30480 ) | ( ~n26555 & n30481 ) | ( n30480 & n30481 ) ;
  assign n30483 = ( n26528 & n30480 ) | ( n26528 & n30481 ) | ( n30480 & n30481 ) ;
  assign n30484 = ( ~n26543 & n30482 ) | ( ~n26543 & n30483 ) | ( n30482 & n30483 ) ;
  assign n30485 = ~x11 & n30484 ;
  assign n30486 = x11 | n30484 ;
  assign n30487 = ( ~n30484 & n30485 ) | ( ~n30484 & n30486 ) | ( n30485 & n30486 ) ;
  assign n30488 = n30471 & n30487 ;
  assign n30489 = n28985 | n29218 ;
  assign n30490 = ~n29219 & n30489 ;
  assign n30491 = n6125 & ~n25728 ;
  assign n30492 = n6119 & n26017 ;
  assign n30493 = n30491 | n30492 ;
  assign n30494 = n6122 & ~n26270 ;
  assign n30495 = ~n26263 & n30494 ;
  assign n30497 = n6115 | n30495 ;
  assign n30498 = n30493 | n30497 ;
  assign n30496 = n30493 | n30495 ;
  assign n30499 = n30496 & n30498 ;
  assign n30500 = ( n26571 & n30498 ) | ( n26571 & n30499 ) | ( n30498 & n30499 ) ;
  assign n30501 = x11 & n30499 ;
  assign n30502 = x11 & n30498 ;
  assign n30503 = ( n26571 & n30501 ) | ( n26571 & n30502 ) | ( n30501 & n30502 ) ;
  assign n30504 = x11 & ~n30501 ;
  assign n30505 = x11 & ~n30502 ;
  assign n30506 = ( ~n26571 & n30504 ) | ( ~n26571 & n30505 ) | ( n30504 & n30505 ) ;
  assign n30507 = ( n30500 & ~n30503 ) | ( n30500 & n30506 ) | ( ~n30503 & n30506 ) ;
  assign n30508 = n30490 & n30507 ;
  assign n30509 = n30490 & ~n30508 ;
  assign n30510 = ~n30490 & n30507 ;
  assign n30511 = n30509 | n30510 ;
  assign n30512 = n29006 & n29216 ;
  assign n30513 = n29006 | n29216 ;
  assign n30514 = ~n30512 & n30513 ;
  assign n30515 = n6122 & n26017 ;
  assign n30516 = n6125 & ~n25046 ;
  assign n30517 = n6119 & ~n25728 ;
  assign n30518 = n30516 | n30517 ;
  assign n30519 = n30515 | n30518 ;
  assign n30520 = n6115 | n30515 ;
  assign n30521 = n30518 | n30520 ;
  assign n30522 = ( n26613 & n30519 ) | ( n26613 & n30521 ) | ( n30519 & n30521 ) ;
  assign n30523 = n30519 | n30521 ;
  assign n30524 = ( n26605 & n30522 ) | ( n26605 & n30523 ) | ( n30522 & n30523 ) ;
  assign n30525 = x11 & n30524 ;
  assign n30526 = x11 & ~n30524 ;
  assign n30527 = ( n30524 & ~n30525 ) | ( n30524 & n30526 ) | ( ~n30525 & n30526 ) ;
  assign n30528 = n30514 & n30527 ;
  assign n30529 = n30514 & ~n30528 ;
  assign n30530 = ~n30514 & n30527 ;
  assign n30531 = n30529 | n30530 ;
  assign n30532 = ( n29042 & n29043 ) | ( n29042 & n29214 ) | ( n29043 & n29214 ) ;
  assign n30533 = n29021 | n29042 ;
  assign n30534 = n29214 | n30533 ;
  assign n30535 = ~n30532 & n30534 ;
  assign n30536 = n6122 & ~n25728 ;
  assign n30537 = n6125 & n24770 ;
  assign n30538 = n6119 & ~n25046 ;
  assign n30539 = n30537 | n30538 ;
  assign n30540 = n30536 | n30539 ;
  assign n30541 = n6115 & n25740 ;
  assign n30542 = n6115 & n25731 ;
  assign n30543 = ( ~n25441 & n30541 ) | ( ~n25441 & n30542 ) | ( n30541 & n30542 ) ;
  assign n30544 = n30540 | n30543 ;
  assign n30545 = n6115 | n30540 ;
  assign n30546 = ( n25733 & n30544 ) | ( n25733 & n30545 ) | ( n30544 & n30545 ) ;
  assign n30547 = x11 | n30546 ;
  assign n30548 = ~x11 & n30546 ;
  assign n30549 = ( ~n30546 & n30547 ) | ( ~n30546 & n30548 ) | ( n30547 & n30548 ) ;
  assign n30550 = n30535 & n30549 ;
  assign n30551 = n29211 & ~n29214 ;
  assign n30554 = n6122 & ~n25046 ;
  assign n30555 = n6125 & ~n25054 ;
  assign n30556 = n6119 & n24770 ;
  assign n30557 = n30555 | n30556 ;
  assign n30558 = n30554 | n30557 ;
  assign n30559 = n6115 | n30554 ;
  assign n30560 = n30557 | n30559 ;
  assign n30561 = ( ~n25069 & n30558 ) | ( ~n25069 & n30560 ) | ( n30558 & n30560 ) ;
  assign n30562 = ~x11 & n30560 ;
  assign n30563 = ~x11 & n30558 ;
  assign n30564 = ( ~n25069 & n30562 ) | ( ~n25069 & n30563 ) | ( n30562 & n30563 ) ;
  assign n30565 = x11 | n30563 ;
  assign n30566 = x11 | n30562 ;
  assign n30567 = ( ~n25069 & n30565 ) | ( ~n25069 & n30566 ) | ( n30565 & n30566 ) ;
  assign n30568 = ( ~n30561 & n30564 ) | ( ~n30561 & n30567 ) | ( n30564 & n30567 ) ;
  assign n30552 = ~n29211 & n29213 ;
  assign n30569 = n30552 & n30568 ;
  assign n30570 = ( n30551 & n30568 ) | ( n30551 & n30569 ) | ( n30568 & n30569 ) ;
  assign n30553 = n30551 | n30552 ;
  assign n30571 = n30553 & ~n30570 ;
  assign n30572 = ~n30552 & n30568 ;
  assign n30573 = ~n30551 & n30572 ;
  assign n30574 = n30571 | n30573 ;
  assign n30575 = n29209 & ~n29210 ;
  assign n30576 = n29066 & ~n29210 ;
  assign n30577 = n30575 | n30576 ;
  assign n30578 = n6122 & n24770 ;
  assign n30579 = n6125 & n24167 ;
  assign n30580 = n6119 & ~n25054 ;
  assign n30581 = n30579 | n30580 ;
  assign n30582 = n30578 | n30581 ;
  assign n30583 = n6115 | n30582 ;
  assign n30584 = ( ~n25095 & n30582 ) | ( ~n25095 & n30583 ) | ( n30582 & n30583 ) ;
  assign n30585 = ~x11 & n30583 ;
  assign n30586 = ~x11 & n30582 ;
  assign n30587 = ( ~n25095 & n30585 ) | ( ~n25095 & n30586 ) | ( n30585 & n30586 ) ;
  assign n30588 = x11 | n30585 ;
  assign n30589 = x11 | n30586 ;
  assign n30590 = ( ~n25095 & n30588 ) | ( ~n25095 & n30589 ) | ( n30588 & n30589 ) ;
  assign n30591 = ( ~n30584 & n30587 ) | ( ~n30584 & n30590 ) | ( n30587 & n30590 ) ;
  assign n30592 = n30577 & n30591 ;
  assign n30593 = n30577 & ~n30592 ;
  assign n30594 = ~n30577 & n30591 ;
  assign n30595 = n30593 | n30594 ;
  assign n30596 = n29088 | n29182 ;
  assign n30597 = ~n29183 & n30596 ;
  assign n30598 = n6122 & n24167 ;
  assign n30599 = n6125 & n23316 ;
  assign n30600 = n6119 & n23614 ;
  assign n30601 = n30599 | n30600 ;
  assign n30602 = n30598 | n30601 ;
  assign n30603 = n6115 | n30602 ;
  assign n30604 = ( n24182 & n30602 ) | ( n24182 & n30603 ) | ( n30602 & n30603 ) ;
  assign n30605 = n30602 | n30603 ;
  assign n30606 = ( n24175 & n30604 ) | ( n24175 & n30605 ) | ( n30604 & n30605 ) ;
  assign n30607 = x11 & n30606 ;
  assign n30608 = x11 & ~n30606 ;
  assign n30609 = ( n30606 & ~n30607 ) | ( n30606 & n30608 ) | ( ~n30607 & n30608 ) ;
  assign n30610 = n30597 & n30609 ;
  assign n30611 = n29184 & n29207 ;
  assign n30612 = n29184 | n29207 ;
  assign n30613 = ~n30611 & n30612 ;
  assign n30614 = n6122 & ~n25054 ;
  assign n30615 = n6125 & n23614 ;
  assign n30616 = n6119 & n24167 ;
  assign n30617 = n30615 | n30616 ;
  assign n30618 = n30614 | n30617 ;
  assign n30619 = n6115 | n30614 ;
  assign n30620 = n30617 | n30619 ;
  assign n30621 = ( ~n25122 & n30618 ) | ( ~n25122 & n30620 ) | ( n30618 & n30620 ) ;
  assign n30622 = ~x11 & n30620 ;
  assign n30623 = ~x11 & n30618 ;
  assign n30624 = ( ~n25122 & n30622 ) | ( ~n25122 & n30623 ) | ( n30622 & n30623 ) ;
  assign n30625 = x11 | n30623 ;
  assign n30626 = x11 | n30622 ;
  assign n30627 = ( ~n25122 & n30625 ) | ( ~n25122 & n30626 ) | ( n30625 & n30626 ) ;
  assign n30628 = ( ~n30621 & n30624 ) | ( ~n30621 & n30627 ) | ( n30624 & n30627 ) ;
  assign n30629 = n30613 & n30628 ;
  assign n30630 = n30613 | n30628 ;
  assign n30631 = ~n30629 & n30630 ;
  assign n30632 = n30610 & n30631 ;
  assign n30633 = n30629 | n30631 ;
  assign n30634 = n29107 | n29180 ;
  assign n30635 = ~n29181 & n30634 ;
  assign n30636 = n6122 & n23614 ;
  assign n30637 = n6125 & n23620 ;
  assign n30638 = ( n6119 & n6294 ) | ( n6119 & n23620 ) | ( n6294 & n23620 ) ;
  assign n30639 = ( n23316 & n30637 ) | ( n23316 & n30638 ) | ( n30637 & n30638 ) ;
  assign n30641 = n6115 | n30639 ;
  assign n30642 = n30636 | n30641 ;
  assign n30640 = n30636 | n30639 ;
  assign n30643 = n30640 & n30642 ;
  assign n30644 = ( n23634 & n30642 ) | ( n23634 & n30643 ) | ( n30642 & n30643 ) ;
  assign n30645 = x11 & n30643 ;
  assign n30646 = x11 & n30642 ;
  assign n30647 = ( n23634 & n30645 ) | ( n23634 & n30646 ) | ( n30645 & n30646 ) ;
  assign n30648 = x11 & ~n30645 ;
  assign n30649 = x11 & ~n30646 ;
  assign n30650 = ( ~n23634 & n30648 ) | ( ~n23634 & n30649 ) | ( n30648 & n30649 ) ;
  assign n30651 = ( n30644 & ~n30647 ) | ( n30644 & n30650 ) | ( ~n30647 & n30650 ) ;
  assign n30652 = n30635 & n30651 ;
  assign n30653 = n30635 & ~n30652 ;
  assign n30654 = ~n30635 & n30651 ;
  assign n30655 = n30653 | n30654 ;
  assign n30656 = n29160 & n29174 ;
  assign n30657 = n29160 & ~n30656 ;
  assign n30658 = n6125 & ~n22385 ;
  assign n30659 = ( n6119 & n6294 ) | ( n6119 & ~n22385 ) | ( n6294 & ~n22385 ) ;
  assign n30660 = ( n22381 & n30658 ) | ( n22381 & n30659 ) | ( n30658 & n30659 ) ;
  assign n30661 = n6122 | n30660 ;
  assign n30662 = ( n23620 & n30660 ) | ( n23620 & n30661 ) | ( n30660 & n30661 ) ;
  assign n30663 = n6115 | n30662 ;
  assign n30664 = ( ~n23686 & n30662 ) | ( ~n23686 & n30663 ) | ( n30662 & n30663 ) ;
  assign n30665 = ~x11 & n30663 ;
  assign n30666 = ~x11 & n30662 ;
  assign n30667 = ( ~n23686 & n30665 ) | ( ~n23686 & n30666 ) | ( n30665 & n30666 ) ;
  assign n30668 = x11 | n30665 ;
  assign n30669 = x11 | n30666 ;
  assign n30670 = ( ~n23686 & n30668 ) | ( ~n23686 & n30669 ) | ( n30668 & n30669 ) ;
  assign n30671 = ( ~n30664 & n30667 ) | ( ~n30664 & n30670 ) | ( n30667 & n30670 ) ;
  assign n30672 = ~n29160 & n29174 ;
  assign n30673 = n30671 & n30672 ;
  assign n30674 = ( n30657 & n30671 ) | ( n30657 & n30673 ) | ( n30671 & n30673 ) ;
  assign n30675 = n30671 | n30672 ;
  assign n30676 = n30657 | n30675 ;
  assign n30677 = ~n30674 & n30676 ;
  assign n30678 = n29139 & n29157 ;
  assign n30679 = n29139 | n29157 ;
  assign n30680 = ~n30678 & n30679 ;
  assign n30681 = n6122 & n22381 ;
  assign n30682 = n6125 & ~n22398 ;
  assign n30683 = n6119 & ~n22385 ;
  assign n30684 = n30682 | n30683 ;
  assign n30685 = n30681 | n30684 ;
  assign n30686 = n6115 | n30685 ;
  assign n30687 = x11 & n30686 ;
  assign n30688 = x11 & n30685 ;
  assign n30689 = ( n22422 & n30687 ) | ( n22422 & n30688 ) | ( n30687 & n30688 ) ;
  assign n30690 = x11 | n30686 ;
  assign n30691 = x11 | n30685 ;
  assign n30692 = ( n22422 & n30690 ) | ( n22422 & n30691 ) | ( n30690 & n30691 ) ;
  assign n30693 = ~n30689 & n30692 ;
  assign n30694 = n30680 & n30693 ;
  assign n30695 = ~n30680 & n30693 ;
  assign n30696 = ( n30680 & ~n30694 ) | ( n30680 & n30695 ) | ( ~n30694 & n30695 ) ;
  assign n30697 = n29133 | n29135 ;
  assign n30698 = ~n29135 & n29137 ;
  assign n30699 = ( n29134 & n30697 ) | ( n29134 & ~n30698 ) | ( n30697 & ~n30698 ) ;
  assign n30700 = ~n29139 & n30699 ;
  assign n30701 = n6122 & ~n22385 ;
  assign n30702 = n6125 & n22393 ;
  assign n30703 = n6119 & ~n22398 ;
  assign n30704 = n30702 | n30703 ;
  assign n30705 = n30701 | n30704 ;
  assign n30706 = n6115 | n30701 ;
  assign n30707 = n30704 | n30706 ;
  assign n30708 = ( ~n22545 & n30705 ) | ( ~n22545 & n30707 ) | ( n30705 & n30707 ) ;
  assign n30709 = ~x11 & n30707 ;
  assign n30710 = ~x11 & n30705 ;
  assign n30711 = ( ~n22545 & n30709 ) | ( ~n22545 & n30710 ) | ( n30709 & n30710 ) ;
  assign n30712 = x11 | n30710 ;
  assign n30713 = x11 | n30709 ;
  assign n30714 = ( ~n22545 & n30712 ) | ( ~n22545 & n30713 ) | ( n30712 & n30713 ) ;
  assign n30715 = ( ~n30708 & n30711 ) | ( ~n30708 & n30714 ) | ( n30711 & n30714 ) ;
  assign n30716 = n30700 & n30715 ;
  assign n30717 = n6115 & n22474 ;
  assign n30718 = n6119 & ~n22409 ;
  assign n30719 = n6122 & ~n22406 ;
  assign n30720 = n30718 | n30719 ;
  assign n30721 = x11 | n30720 ;
  assign n30722 = n30717 | n30721 ;
  assign n30723 = ~x11 & n30722 ;
  assign n30724 = ( x11 & n19122 ) | ( x11 & n22409 ) | ( n19122 & n22409 ) ;
  assign n30725 = n30722 & n30724 ;
  assign n30726 = n30717 | n30720 ;
  assign n30727 = n30724 & ~n30726 ;
  assign n30728 = ( n30723 & n30725 ) | ( n30723 & n30727 ) | ( n30725 & n30727 ) ;
  assign n30729 = n6122 & n22393 ;
  assign n30730 = n6125 & ~n22409 ;
  assign n30731 = n6119 & ~n22406 ;
  assign n30732 = n30730 | n30731 ;
  assign n30733 = n30729 | n30732 ;
  assign n30734 = n22439 | n30733 ;
  assign n30735 = n6115 | n30729 ;
  assign n30736 = n30732 | n30735 ;
  assign n30737 = ~x11 & n30736 ;
  assign n30738 = n30734 & n30737 ;
  assign n30739 = x11 | n30738 ;
  assign n30740 = n5223 & ~n22409 ;
  assign n30741 = n30738 & n30740 ;
  assign n30742 = n30734 & n30736 ;
  assign n30743 = n30740 & ~n30742 ;
  assign n30744 = ( n30739 & n30741 ) | ( n30739 & n30743 ) | ( n30741 & n30743 ) ;
  assign n30745 = n30728 & n30744 ;
  assign n30746 = ( n30738 & n30739 ) | ( n30738 & ~n30742 ) | ( n30739 & ~n30742 ) ;
  assign n30747 = n30728 | n30740 ;
  assign n30748 = ( n30740 & n30746 ) | ( n30740 & n30747 ) | ( n30746 & n30747 ) ;
  assign n30749 = ~n30745 & n30748 ;
  assign n30750 = n6125 & ~n22406 ;
  assign n30751 = n6119 & n22393 ;
  assign n30752 = n30750 | n30751 ;
  assign n30753 = n6122 & ~n22398 ;
  assign n30754 = n6115 | n30753 ;
  assign n30755 = n30752 | n30754 ;
  assign n30756 = x11 & n30755 ;
  assign n30757 = n30752 | n30753 ;
  assign n30758 = x11 & n30757 ;
  assign n30759 = ( n22608 & n30756 ) | ( n22608 & n30758 ) | ( n30756 & n30758 ) ;
  assign n30760 = x11 | n30755 ;
  assign n30761 = x11 | n30757 ;
  assign n30762 = ( n22608 & n30760 ) | ( n22608 & n30761 ) | ( n30760 & n30761 ) ;
  assign n30763 = ~n30759 & n30762 ;
  assign n30764 = n30745 | n30763 ;
  assign n30765 = ( n30745 & n30749 ) | ( n30745 & n30764 ) | ( n30749 & n30764 ) ;
  assign n30766 = n30700 | n30715 ;
  assign n30767 = ~n30716 & n30766 ;
  assign n30768 = n30716 | n30767 ;
  assign n30769 = ( n30716 & n30765 ) | ( n30716 & n30768 ) | ( n30765 & n30768 ) ;
  assign n30770 = n30696 & n30769 ;
  assign n30771 = n30694 | n30770 ;
  assign n30772 = n30677 & n30771 ;
  assign n30773 = n30674 | n30772 ;
  assign n30774 = n6125 & n22381 ;
  assign n30775 = ( n6119 & n6294 ) | ( n6119 & n22381 ) | ( n6294 & n22381 ) ;
  assign n30776 = ( n23620 & n30774 ) | ( n23620 & n30775 ) | ( n30774 & n30775 ) ;
  assign n30777 = n6122 | n30775 ;
  assign n30778 = n6122 | n30774 ;
  assign n30779 = ( n23620 & n30777 ) | ( n23620 & n30778 ) | ( n30777 & n30778 ) ;
  assign n30780 = ( n23316 & n30776 ) | ( n23316 & n30779 ) | ( n30776 & n30779 ) ;
  assign n30781 = n6115 | n30780 ;
  assign n30782 = ~x11 & n30781 ;
  assign n30783 = ~x11 & n30780 ;
  assign n30784 = ( n23661 & n30782 ) | ( n23661 & n30783 ) | ( n30782 & n30783 ) ;
  assign n30785 = ( x11 & n19082 ) | ( x11 & n30780 ) | ( n19082 & n30780 ) ;
  assign n30786 = x11 & ~n30785 ;
  assign n30787 = x11 & n30780 ;
  assign n30788 = x11 & ~n30787 ;
  assign n30789 = ( ~n23661 & n30786 ) | ( ~n23661 & n30788 ) | ( n30786 & n30788 ) ;
  assign n30790 = n30784 | n30789 ;
  assign n30791 = n29176 & n29178 ;
  assign n30792 = n29176 | n29178 ;
  assign n30793 = ~n30791 & n30792 ;
  assign n30794 = n30790 & n30793 ;
  assign n30795 = n30790 | n30793 ;
  assign n30796 = ~n30794 & n30795 ;
  assign n30797 = n30794 | n30796 ;
  assign n30798 = ( n30773 & n30794 ) | ( n30773 & n30797 ) | ( n30794 & n30797 ) ;
  assign n30799 = n30655 & n30798 ;
  assign n30800 = n30652 | n30799 ;
  assign n30801 = ~n30597 & n30609 ;
  assign n30802 = ( n30597 & ~n30610 ) | ( n30597 & n30801 ) | ( ~n30610 & n30801 ) ;
  assign n30803 = n30800 & n30802 ;
  assign n30804 = n30629 | n30803 ;
  assign n30805 = ( n30632 & n30633 ) | ( n30632 & n30804 ) | ( n30633 & n30804 ) ;
  assign n30806 = n30592 | n30805 ;
  assign n30807 = ( n30592 & n30595 ) | ( n30592 & n30806 ) | ( n30595 & n30806 ) ;
  assign n30808 = n30574 & n30807 ;
  assign n30809 = n30570 | n30808 ;
  assign n30810 = ~n30535 & n30549 ;
  assign n30811 = ( n30535 & ~n30550 ) | ( n30535 & n30810 ) | ( ~n30550 & n30810 ) ;
  assign n30812 = n30550 | n30811 ;
  assign n30813 = ( n30550 & n30809 ) | ( n30550 & n30812 ) | ( n30809 & n30812 ) ;
  assign n30814 = n30528 | n30813 ;
  assign n30815 = ( n30528 & n30531 ) | ( n30528 & n30814 ) | ( n30531 & n30814 ) ;
  assign n30816 = n30511 & n30815 ;
  assign n30817 = n30508 | n30816 ;
  assign n30818 = n30471 | n30487 ;
  assign n30819 = ~n30488 & n30818 ;
  assign n30820 = n30488 | n30819 ;
  assign n30821 = ( n30488 & n30817 ) | ( n30488 & n30820 ) | ( n30817 & n30820 ) ;
  assign n30822 = n30468 & n30821 ;
  assign n30823 = n30466 | n30822 ;
  assign n30824 = n30427 | n30445 ;
  assign n30825 = ~n30446 & n30824 ;
  assign n30826 = n30446 | n30825 ;
  assign n30827 = ( n30446 & n30823 ) | ( n30446 & n30826 ) | ( n30823 & n30826 ) ;
  assign n30828 = n30424 & n30827 ;
  assign n30829 = n30422 | n30828 ;
  assign n30830 = n30357 & ~n30376 ;
  assign n30831 = ~n30357 & n30375 ;
  assign n30832 = n30830 | n30831 ;
  assign n30833 = n30829 & n30832 ;
  assign n30834 = n30397 | n30833 ;
  assign n30835 = ( n30400 & n30401 ) | ( n30400 & n30834 ) | ( n30401 & n30834 ) ;
  assign n30836 = n30351 | n30835 ;
  assign n30837 = ( n30351 & ~n30355 ) | ( n30351 & n30836 ) | ( ~n30355 & n30836 ) ;
  assign n30838 = ~n30331 & n30837 ;
  assign n30839 = n30329 | n30838 ;
  assign n30840 = n30312 & n30839 ;
  assign n30841 = n30310 | n30840 ;
  assign n30842 = n30284 | n30841 ;
  assign n30843 = ( n30284 & ~n30287 ) | ( n30284 & n30842 ) | ( ~n30287 & n30842 ) ;
  assign n30844 = n30255 & ~n30843 ;
  assign n30845 = ~n30255 & n30843 ;
  assign n30846 = n30844 | n30845 ;
  assign n30847 = n3541 | n3547 ;
  assign n31218 = ~n23234 & n30847 ;
  assign n31219 = n3544 | n31218 ;
  assign n31220 = ~n23235 & n30847 ;
  assign n31221 = n3544 | n31220 ;
  assign n31222 = ( ~n15882 & n31219 ) | ( ~n15882 & n31221 ) | ( n31219 & n31221 ) ;
  assign n31223 = n3537 | n31222 ;
  assign n31224 = ( ~n15882 & n31218 ) | ( ~n15882 & n31220 ) | ( n31218 & n31220 ) ;
  assign n31225 = n3537 | n31224 ;
  assign n31226 = ( ~n23240 & n31223 ) | ( ~n23240 & n31225 ) | ( n31223 & n31225 ) ;
  assign n31227 = ( ~n23240 & n31222 ) | ( ~n23240 & n31224 ) | ( n31222 & n31224 ) ;
  assign n31228 = n24135 & ~n31227 ;
  assign n31229 = n23240 & ~n31227 ;
  assign n31230 = ( n23575 & n31228 ) | ( n23575 & n31229 ) | ( n31228 & n31229 ) ;
  assign n31231 = ( n23577 & n31228 ) | ( n23577 & n31229 ) | ( n31228 & n31229 ) ;
  assign n31232 = ( ~n21554 & n31230 ) | ( ~n21554 & n31231 ) | ( n31230 & n31231 ) ;
  assign n31233 = n31226 & ~n31232 ;
  assign n31234 = x20 & ~n31233 ;
  assign n31235 = n31230 | n31231 ;
  assign n31236 = n31226 & ~n31235 ;
  assign n31237 = x20 & ~n31236 ;
  assign n31238 = ( n21584 & n31234 ) | ( n21584 & n31237 ) | ( n31234 & n31237 ) ;
  assign n31239 = ~x20 & n31233 ;
  assign n31240 = ~x20 & n31236 ;
  assign n31241 = ( ~n21584 & n31239 ) | ( ~n21584 & n31240 ) | ( n31239 & n31240 ) ;
  assign n31242 = n31238 | n31241 ;
  assign n31243 = n30011 | n30028 ;
  assign n31244 = ( n30011 & ~n30013 ) | ( n30011 & n31243 ) | ( ~n30013 & n31243 ) ;
  assign n31245 = n31242 & n31244 ;
  assign n31246 = n31242 | n31244 ;
  assign n31247 = ~n31245 & n31246 ;
  assign n31009 = n29963 | n29981 ;
  assign n31010 = ( n29963 & ~n29966 ) | ( n29963 & n31009 ) | ( ~n29966 & n31009 ) ;
  assign n30958 = n1060 & n18410 ;
  assign n30959 = n1065 & n18576 ;
  assign n30960 = n30958 | n30959 ;
  assign n30961 = n1057 & n19352 ;
  assign n30968 = n1062 | n30961 ;
  assign n30969 = n30960 | n30968 ;
  assign n31011 = n30960 | n30961 ;
  assign n31012 = ( n19674 & n30969 ) | ( n19674 & n31011 ) | ( n30969 & n31011 ) ;
  assign n30931 = n448 | n623 ;
  assign n30932 = n2134 | n2138 ;
  assign n30933 = n175 | n959 ;
  assign n30934 = n331 | n510 ;
  assign n30935 = n30933 | n30934 ;
  assign n30936 = n182 | n30935 ;
  assign n30937 = n7927 | n14362 ;
  assign n30938 = n30936 | n30937 ;
  assign n30939 = n1133 | n4406 ;
  assign n30940 = n30938 | n30939 ;
  assign n30941 = n30932 | n30940 ;
  assign n30942 = n1113 & ~n30941 ;
  assign n30943 = n24222 | n24231 ;
  assign n30944 = n24227 | n30943 ;
  assign n30945 = n1287 | n30944 ;
  assign n30946 = n661 | n1675 ;
  assign n30947 = n112 | n1785 ;
  assign n30948 = n30946 | n30947 ;
  assign n30949 = n284 | n441 ;
  assign n30950 = n762 | n30949 ;
  assign n30951 = n1417 | n30950 ;
  assign n30952 = n30948 | n30951 ;
  assign n30953 = n600 | n30952 ;
  assign n30954 = n30945 | n30953 ;
  assign n30955 = n30942 & ~n30954 ;
  assign n30956 = ~n30931 & n30955 ;
  assign n30957 = n29939 & ~n30956 ;
  assign n30962 = ~n30957 & n30961 ;
  assign n30963 = ( ~n30957 & n30960 ) | ( ~n30957 & n30962 ) | ( n30960 & n30962 ) ;
  assign n30964 = ~n29939 & n30956 ;
  assign n31013 = n30963 & ~n30964 ;
  assign n30970 = n30957 | n30964 ;
  assign n31014 = n30969 & ~n30970 ;
  assign n31015 = ( n19674 & n31013 ) | ( n19674 & n31014 ) | ( n31013 & n31014 ) ;
  assign n31016 = n31012 & ~n31015 ;
  assign n31017 = n29942 | n29956 ;
  assign n31018 = n29942 | n29954 ;
  assign n31019 = ( n18612 & n31017 ) | ( n18612 & n31018 ) | ( n31017 & n31018 ) ;
  assign n30965 = ~n30957 & n30964 ;
  assign n30966 = ( n30957 & n30963 ) | ( n30957 & ~n30965 ) | ( n30963 & ~n30965 ) ;
  assign n31020 = n30964 | n30966 ;
  assign n30971 = ~n30957 & n30970 ;
  assign n30972 = ( n30957 & n30969 ) | ( n30957 & ~n30971 ) | ( n30969 & ~n30971 ) ;
  assign n31021 = n30964 | n30972 ;
  assign n31022 = ( n19674 & n31020 ) | ( n19674 & n31021 ) | ( n31020 & n31021 ) ;
  assign n31023 = n31019 & ~n31022 ;
  assign n31024 = ( n31016 & n31019 ) | ( n31016 & n31023 ) | ( n31019 & n31023 ) ;
  assign n31025 = ~n31019 & n31022 ;
  assign n31026 = ~n31016 & n31025 ;
  assign n31027 = n31024 | n31026 ;
  assign n31074 = n31010 & ~n31027 ;
  assign n31075 = ~n31010 & n31027 ;
  assign n31076 = n31074 | n31075 ;
  assign n31077 = n1829 & ~n20630 ;
  assign n31078 = n1826 & n19494 ;
  assign n31079 = n1823 & n19631 ;
  assign n31080 = n31078 | n31079 ;
  assign n31081 = n31077 | n31080 ;
  assign n31082 = n1821 | n31077 ;
  assign n31083 = n31080 | n31082 ;
  assign n31084 = ( ~n20709 & n31081 ) | ( ~n20709 & n31083 ) | ( n31081 & n31083 ) ;
  assign n31085 = ~x29 & n31083 ;
  assign n31086 = ~x29 & n31081 ;
  assign n31087 = ( ~n20709 & n31085 ) | ( ~n20709 & n31086 ) | ( n31085 & n31086 ) ;
  assign n31088 = x29 | n31086 ;
  assign n31089 = x29 | n31085 ;
  assign n31090 = ( ~n20709 & n31088 ) | ( ~n20709 & n31089 ) | ( n31088 & n31089 ) ;
  assign n31091 = ( ~n31084 & n31087 ) | ( ~n31084 & n31090 ) | ( n31087 & n31090 ) ;
  assign n31092 = ~n31076 & n31091 ;
  assign n31093 = n31076 | n31092 ;
  assign n31094 = n2315 & ~n21563 ;
  assign n31095 = n2312 & ~n20618 ;
  assign n31096 = n2308 & n20609 ;
  assign n31097 = n31095 | n31096 ;
  assign n31098 = n31094 | n31097 ;
  assign n31099 = n2306 & ~n21570 ;
  assign n31100 = n22270 & n31099 ;
  assign n31101 = ( n2306 & n22304 ) | ( n2306 & n31100 ) | ( n22304 & n31100 ) ;
  assign n31102 = n31098 | n31101 ;
  assign n31103 = x26 | n31098 ;
  assign n31104 = n31101 | n31103 ;
  assign n31105 = ~x26 & n31103 ;
  assign n31106 = ( ~x26 & n31101 ) | ( ~x26 & n31105 ) | ( n31101 & n31105 ) ;
  assign n31107 = ( ~n31102 & n31104 ) | ( ~n31102 & n31106 ) | ( n31104 & n31106 ) ;
  assign n31108 = n31076 & n31091 ;
  assign n31109 = n31107 & n31108 ;
  assign n31110 = ( ~n31093 & n31107 ) | ( ~n31093 & n31109 ) | ( n31107 & n31109 ) ;
  assign n31175 = n31107 | n31108 ;
  assign n31176 = n31093 & ~n31175 ;
  assign n31177 = n31110 | n31176 ;
  assign n31178 = n29988 | n30005 ;
  assign n31179 = ( n29988 & ~n29992 ) | ( n29988 & n31178 ) | ( ~n29992 & n31178 ) ;
  assign n31180 = ~n31177 & n31179 ;
  assign n31181 = n31177 & ~n31179 ;
  assign n31182 = n31180 | n31181 ;
  assign n31183 = n2925 & ~n21517 ;
  assign n31184 = n2928 & ~n21551 ;
  assign n31185 = n31183 | n31184 ;
  assign n31186 = n2932 & n23227 ;
  assign n31187 = ( n2932 & n23217 ) | ( n2932 & n31186 ) | ( n23217 & n31186 ) ;
  assign n31188 = n31185 | n31187 ;
  assign n31189 = n2936 & n23299 ;
  assign n31190 = n2936 & n23298 ;
  assign n31191 = ( n21584 & n31189 ) | ( n21584 & n31190 ) | ( n31189 & n31190 ) ;
  assign n31192 = n31188 | n31191 ;
  assign n31193 = n2936 | n31188 ;
  assign n31194 = ( n23289 & n31192 ) | ( n23289 & n31193 ) | ( n31192 & n31193 ) ;
  assign n31195 = x23 | n31194 ;
  assign n31196 = ~x23 & n31194 ;
  assign n31197 = ( ~n31194 & n31195 ) | ( ~n31194 & n31196 ) | ( n31195 & n31196 ) ;
  assign n31248 = n31182 | n31197 ;
  assign n31249 = n31182 & ~n31197 ;
  assign n31250 = ( ~n31182 & n31248 ) | ( ~n31182 & n31249 ) | ( n31248 & n31249 ) ;
  assign n31256 = n31247 & ~n31250 ;
  assign n31257 = n31247 | n31250 ;
  assign n31258 = ( ~n31247 & n31256 ) | ( ~n31247 & n31257 ) | ( n31256 & n31257 ) ;
  assign n31259 = n30032 | n30052 ;
  assign n31260 = ( n30032 & ~n30034 ) | ( n30032 & n31259 ) | ( ~n30034 & n31259 ) ;
  assign n31261 = ~n31258 & n31260 ;
  assign n31262 = n31258 & ~n31260 ;
  assign n31263 = n31261 | n31262 ;
  assign n31276 = n30107 & ~n31263 ;
  assign n31297 = ( n30169 & ~n31263 ) | ( n30169 & n31276 ) | ( ~n31263 & n31276 ) ;
  assign n31264 = n30107 | n30174 ;
  assign n31265 = ~n31263 & n31264 ;
  assign n31269 = ~n30107 & n30110 ;
  assign n31270 = n31263 | n31269 ;
  assign n31298 = ( n30173 & n31265 ) | ( n30173 & ~n31270 ) | ( n31265 & ~n31270 ) ;
  assign n31299 = ( n28465 & n31297 ) | ( n28465 & n31298 ) | ( n31297 & n31298 ) ;
  assign n31300 = n31297 & n31298 ;
  assign n31301 = ( n28489 & n31299 ) | ( n28489 & n31300 ) | ( n31299 & n31300 ) ;
  assign n31302 = n30107 | n30169 ;
  assign n31303 = ( n30173 & n31264 ) | ( n30173 & ~n31269 ) | ( n31264 & ~n31269 ) ;
  assign n31304 = n31302 & n31303 ;
  assign n31305 = n31263 & ~n31304 ;
  assign n31306 = ( n28465 & n31302 ) | ( n28465 & n31303 ) | ( n31302 & n31303 ) ;
  assign n31307 = n31263 & ~n31306 ;
  assign n31308 = ( ~n28489 & n31305 ) | ( ~n28489 & n31307 ) | ( n31305 & n31307 ) ;
  assign n31309 = n31301 | n31308 ;
  assign n31310 = n7074 & ~n31309 ;
  assign n31198 = n31180 | n31197 ;
  assign n31199 = ( n31180 & ~n31182 ) | ( n31180 & n31198 ) | ( ~n31182 & n31198 ) ;
  assign n31159 = n2932 & ~n23240 ;
  assign n31160 = n2925 & ~n21551 ;
  assign n31161 = n2928 & n23227 ;
  assign n31162 = ( n2928 & n23217 ) | ( n2928 & n31161 ) | ( n23217 & n31161 ) ;
  assign n31163 = n31160 | n31162 ;
  assign n31164 = n31159 | n31163 ;
  assign n31165 = n2936 | n31159 ;
  assign n31166 = n31163 | n31165 ;
  assign n31167 = ( n23260 & n31164 ) | ( n23260 & n31166 ) | ( n31164 & n31166 ) ;
  assign n31168 = x23 & n31166 ;
  assign n31169 = x23 & n31164 ;
  assign n31170 = ( n23260 & n31168 ) | ( n23260 & n31169 ) | ( n31168 & n31169 ) ;
  assign n31171 = x23 & ~n31169 ;
  assign n31172 = x23 & ~n31168 ;
  assign n31173 = ( ~n23260 & n31171 ) | ( ~n23260 & n31172 ) | ( n31171 & n31172 ) ;
  assign n31174 = ( n31167 & ~n31170 ) | ( n31167 & n31173 ) | ( ~n31170 & n31173 ) ;
  assign n31200 = n31174 & n31199 ;
  assign n31201 = n31199 & ~n31200 ;
  assign n31111 = n31092 | n31110 ;
  assign n30848 = n3544 | n30847 ;
  assign n30849 = n3537 | n30848 ;
  assign n30850 = ~n23229 & n30849 ;
  assign n30851 = ( n23154 & n30849 ) | ( n23154 & n30850 ) | ( n30849 & n30850 ) ;
  assign n30852 = ~n23232 & n30849 ;
  assign n30853 = ~n23231 & n30849 ;
  assign n30854 = ( n9072 & n30852 ) | ( n9072 & n30853 ) | ( n30852 & n30853 ) ;
  assign n30855 = ( ~n21543 & n30851 ) | ( ~n21543 & n30854 ) | ( n30851 & n30854 ) ;
  assign n30856 = ( ~n21545 & n30851 ) | ( ~n21545 & n30854 ) | ( n30851 & n30854 ) ;
  assign n30857 = ( ~n15882 & n30855 ) | ( ~n15882 & n30856 ) | ( n30855 & n30856 ) ;
  assign n30858 = ~x20 & n30855 ;
  assign n30859 = ~x20 & n30856 ;
  assign n30860 = ( ~n15882 & n30858 ) | ( ~n15882 & n30859 ) | ( n30858 & n30859 ) ;
  assign n30861 = x20 | n30858 ;
  assign n30862 = x20 | n30859 ;
  assign n30863 = ( ~n15882 & n30861 ) | ( ~n15882 & n30862 ) | ( n30861 & n30862 ) ;
  assign n30864 = ( ~n30857 & n30860 ) | ( ~n30857 & n30863 ) | ( n30860 & n30863 ) ;
  assign n30865 = ( ~n948 & n2874 ) | ( ~n948 & n10851 ) | ( n2874 & n10851 ) ;
  assign n30866 = n784 | n4263 ;
  assign n30867 = n4260 | n30866 ;
  assign n30868 = n948 | n30867 ;
  assign n30869 = n30865 | n30868 ;
  assign n30870 = n624 | n30869 ;
  assign n30871 = n164 | n13310 ;
  assign n30872 = n553 | n30871 ;
  assign n30873 = n240 | n2614 ;
  assign n30874 = n6823 | n30873 ;
  assign n30875 = n30872 | n30874 ;
  assign n30876 = n1785 | n3467 ;
  assign n30877 = n179 | n602 ;
  assign n30878 = n117 | n30877 ;
  assign n30879 = n30876 | n30878 ;
  assign n30880 = n363 | n30879 ;
  assign n30881 = n1725 | n4157 ;
  assign n30882 = n4155 | n30881 ;
  assign n30883 = n30880 | n30882 ;
  assign n30884 = n30875 | n30883 ;
  assign n30885 = n30870 | n30884 ;
  assign n30886 = n259 | n4046 ;
  assign n30887 = n85 | n1523 ;
  assign n30888 = n30886 | n30887 ;
  assign n30889 = n283 | n318 ;
  assign n30890 = n374 | n30889 ;
  assign n30891 = n225 | n30890 ;
  assign n30892 = n30888 | n30891 ;
  assign n30893 = n245 | n30892 ;
  assign n30894 = ~n2818 & n2822 ;
  assign n30895 = ~n2802 & n30894 ;
  assign n30896 = ~n30893 & n30895 ;
  assign n30897 = ~n30885 & n30896 ;
  assign n30898 = ~n577 & n30897 ;
  assign n30899 = n29939 | n30898 ;
  assign n30900 = n29939 & n30898 ;
  assign n30901 = n30899 & ~n30900 ;
  assign n30928 = ~n30864 & n30901 ;
  assign n30929 = n30864 & ~n30901 ;
  assign n30930 = n30928 | n30929 ;
  assign n30967 = ~n30930 & n30966 ;
  assign n30973 = ~n30930 & n30972 ;
  assign n30974 = ( n19674 & n30967 ) | ( n19674 & n30973 ) | ( n30967 & n30973 ) ;
  assign n30975 = n30930 & ~n30966 ;
  assign n30976 = n30930 & ~n30972 ;
  assign n30977 = ( ~n19674 & n30975 ) | ( ~n19674 & n30976 ) | ( n30975 & n30976 ) ;
  assign n30978 = n30974 | n30977 ;
  assign n30979 = n1057 & n19494 ;
  assign n30980 = n1060 & n18576 ;
  assign n30981 = n1065 & n19352 ;
  assign n30982 = n30980 | n30981 ;
  assign n30983 = n30979 | n30982 ;
  assign n30984 = n1062 | n30979 ;
  assign n30985 = n30982 | n30984 ;
  assign n30986 = ( n20320 & n30983 ) | ( n20320 & n30985 ) | ( n30983 & n30985 ) ;
  assign n31028 = n30978 & n30986 ;
  assign n31029 = n30978 | n30986 ;
  assign n31030 = ~n31028 & n31029 ;
  assign n31031 = ( ~n31024 & n31027 ) | ( ~n31024 & n31030 ) | ( n31027 & n31030 ) ;
  assign n31032 = n31024 & ~n31030 ;
  assign n31033 = ( n31010 & ~n31031 ) | ( n31010 & n31032 ) | ( ~n31031 & n31032 ) ;
  assign n31034 = ~n31024 & n31027 ;
  assign n31035 = n31030 & n31034 ;
  assign n31036 = ~n31024 & n31030 ;
  assign n31037 = ( ~n31010 & n31035 ) | ( ~n31010 & n31036 ) | ( n31035 & n31036 ) ;
  assign n31038 = n31033 | n31037 ;
  assign n31039 = n1821 & n20680 ;
  assign n31040 = n1829 & ~n20618 ;
  assign n31041 = n1826 & n19631 ;
  assign n31042 = n1823 & ~n20630 ;
  assign n31043 = n31041 | n31042 ;
  assign n31044 = n31040 | n31043 ;
  assign n31045 = n20689 | n31044 ;
  assign n31046 = n1821 | n31044 ;
  assign n31047 = ( n31039 & n31045 ) | ( n31039 & n31046 ) | ( n31045 & n31046 ) ;
  assign n31048 = x29 | n31047 ;
  assign n31049 = ~x29 & n31047 ;
  assign n31050 = ( ~n31047 & n31048 ) | ( ~n31047 & n31049 ) | ( n31048 & n31049 ) ;
  assign n31112 = ~n31038 & n31050 ;
  assign n31113 = n31038 | n31112 ;
  assign n31114 = n2315 & ~n21517 ;
  assign n31115 = n2312 & n20609 ;
  assign n31116 = n2308 & ~n21563 ;
  assign n31117 = n31115 | n31116 ;
  assign n31118 = n31114 | n31117 ;
  assign n31119 = n2306 | n31114 ;
  assign n31120 = n31117 | n31119 ;
  assign n31121 = ( ~n22283 & n31118 ) | ( ~n22283 & n31120 ) | ( n31118 & n31120 ) ;
  assign n31122 = n31118 & n31120 ;
  assign n31123 = ( ~n22271 & n31121 ) | ( ~n22271 & n31122 ) | ( n31121 & n31122 ) ;
  assign n31124 = ~x26 & n31123 ;
  assign n31125 = x26 | n31123 ;
  assign n31126 = ( ~n31123 & n31124 ) | ( ~n31123 & n31125 ) | ( n31124 & n31125 ) ;
  assign n31127 = n31038 & n31050 ;
  assign n31128 = n31126 & n31127 ;
  assign n31129 = ( ~n31113 & n31126 ) | ( ~n31113 & n31128 ) | ( n31126 & n31128 ) ;
  assign n31130 = n31126 | n31127 ;
  assign n31131 = n31113 & ~n31130 ;
  assign n31132 = n31129 | n31131 ;
  assign n31133 = n31111 & ~n31132 ;
  assign n31202 = ~n31111 & n31132 ;
  assign n31203 = n31133 | n31202 ;
  assign n31204 = n31174 & ~n31203 ;
  assign n31205 = ~n31199 & n31204 ;
  assign n31213 = ( n31201 & ~n31203 ) | ( n31201 & n31205 ) | ( ~n31203 & n31205 ) ;
  assign n31214 = ~n31174 & n31203 ;
  assign n31215 = ( n31199 & n31203 ) | ( n31199 & n31214 ) | ( n31203 & n31214 ) ;
  assign n31216 = ~n31201 & n31215 ;
  assign n31217 = n31213 | n31216 ;
  assign n31251 = ~n31245 & n31250 ;
  assign n31252 = ( n31245 & n31247 ) | ( n31245 & ~n31251 ) | ( n31247 & ~n31251 ) ;
  assign n31253 = ~n31217 & n31252 ;
  assign n31254 = n31217 & ~n31252 ;
  assign n31255 = n31253 | n31254 ;
  assign n31277 = n31261 | n31276 ;
  assign n31278 = ~n31255 & n31277 ;
  assign n31281 = ~n31261 & n31263 ;
  assign n31282 = n31255 | n31281 ;
  assign n31311 = ( n30169 & n31278 ) | ( n30169 & ~n31282 ) | ( n31278 & ~n31282 ) ;
  assign n31266 = n31261 | n31265 ;
  assign n31267 = ~n31255 & n31266 ;
  assign n31271 = ~n31261 & n31270 ;
  assign n31272 = n31255 | n31271 ;
  assign n31312 = ( n30173 & n31267 ) | ( n30173 & ~n31272 ) | ( n31267 & ~n31272 ) ;
  assign n31313 = ( n28465 & n31311 ) | ( n28465 & n31312 ) | ( n31311 & n31312 ) ;
  assign n31314 = n31311 & n31312 ;
  assign n31315 = ( n28489 & n31313 ) | ( n28489 & n31314 ) | ( n31313 & n31314 ) ;
  assign n31316 = ( n30169 & n31277 ) | ( n30169 & ~n31281 ) | ( n31277 & ~n31281 ) ;
  assign n31317 = ( n30173 & n31266 ) | ( n30173 & ~n31271 ) | ( n31266 & ~n31271 ) ;
  assign n31318 = n31316 & n31317 ;
  assign n31319 = n31255 & ~n31318 ;
  assign n31320 = ( n28465 & n31316 ) | ( n28465 & n31317 ) | ( n31316 & n31317 ) ;
  assign n31321 = n31255 & ~n31320 ;
  assign n31322 = ( ~n28489 & n31319 ) | ( ~n28489 & n31321 ) | ( n31319 & n31321 ) ;
  assign n31323 = n31315 | n31322 ;
  assign n31324 = n7068 & ~n31323 ;
  assign n31325 = n31310 | n31324 ;
  assign n31206 = n31200 | n31205 ;
  assign n31207 = ~n31200 & n31203 ;
  assign n31208 = ( n31201 & n31206 ) | ( n31201 & ~n31207 ) | ( n31206 & ~n31207 ) ;
  assign n30902 = n23167 | n23191 ;
  assign n30903 = ( n30899 & ~n30901 ) | ( n30899 & n30902 ) | ( ~n30901 & n30902 ) ;
  assign n30904 = n30899 | n30902 ;
  assign n30905 = ( n30864 & n30903 ) | ( n30864 & n30904 ) | ( n30903 & n30904 ) ;
  assign n30906 = n30899 & ~n30901 ;
  assign n30907 = n30902 & n30906 ;
  assign n30908 = n30899 & n30902 ;
  assign n30909 = ( n30864 & n30907 ) | ( n30864 & n30908 ) | ( n30907 & n30908 ) ;
  assign n30910 = n30905 & ~n30909 ;
  assign n30911 = n1057 & n19631 ;
  assign n30912 = n1065 & n19494 ;
  assign n30913 = n1060 & n19352 ;
  assign n30914 = n30912 | n30913 ;
  assign n30915 = n30911 | n30914 ;
  assign n30916 = n30910 & n30915 ;
  assign n30917 = n1062 & n19652 ;
  assign n30918 = n1062 & n19655 ;
  assign n30919 = ( ~n18604 & n30917 ) | ( ~n18604 & n30918 ) | ( n30917 & n30918 ) ;
  assign n30920 = ( n30910 & n30916 ) | ( n30910 & n30919 ) | ( n30916 & n30919 ) ;
  assign n30921 = ( n1062 & n30910 ) | ( n1062 & n30916 ) | ( n30910 & n30916 ) ;
  assign n30922 = ( n19640 & n30920 ) | ( n19640 & n30921 ) | ( n30920 & n30921 ) ;
  assign n30923 = n30910 | n30915 ;
  assign n30924 = n30919 | n30923 ;
  assign n30925 = n1062 | n30923 ;
  assign n30926 = ( n19640 & n30924 ) | ( n19640 & n30925 ) | ( n30924 & n30925 ) ;
  assign n30927 = ~n30922 & n30926 ;
  assign n30987 = n30974 | n30986 ;
  assign n30988 = ( n30974 & ~n30978 ) | ( n30974 & n30987 ) | ( ~n30978 & n30987 ) ;
  assign n30989 = n30927 & n30988 ;
  assign n30990 = n30927 | n30988 ;
  assign n30991 = ~n30989 & n30990 ;
  assign n30993 = n1826 & ~n20630 ;
  assign n30994 = n1823 & ~n20618 ;
  assign n30995 = n30993 | n30994 ;
  assign n30992 = n1829 & n20609 ;
  assign n30997 = n1821 | n30992 ;
  assign n30998 = n30995 | n30997 ;
  assign n30996 = n30992 | n30995 ;
  assign n30999 = n30996 & n30998 ;
  assign n31000 = ( n20659 & n30998 ) | ( n20659 & n30999 ) | ( n30998 & n30999 ) ;
  assign n31001 = n30998 & n30999 ;
  assign n31002 = ( ~n20649 & n31000 ) | ( ~n20649 & n31001 ) | ( n31000 & n31001 ) ;
  assign n31003 = x29 & n31002 ;
  assign n31004 = x29 & ~n31002 ;
  assign n31005 = ( n31002 & ~n31003 ) | ( n31002 & n31004 ) | ( ~n31003 & n31004 ) ;
  assign n31006 = n30991 & n31005 ;
  assign n31007 = n30991 | n31005 ;
  assign n31008 = ~n31006 & n31007 ;
  assign n31051 = n31033 | n31050 ;
  assign n31052 = ( n31033 & ~n31038 ) | ( n31033 & n31051 ) | ( ~n31038 & n31051 ) ;
  assign n31053 = n31008 & n31052 ;
  assign n31054 = n31008 | n31052 ;
  assign n31055 = ~n31053 & n31054 ;
  assign n31056 = n2315 & ~n21551 ;
  assign n31057 = n2312 & ~n21563 ;
  assign n31058 = n2308 & ~n21517 ;
  assign n31059 = n31057 | n31058 ;
  assign n31060 = n31056 | n31059 ;
  assign n31061 = n2306 | n31056 ;
  assign n31062 = n31059 | n31061 ;
  assign n31063 = ( ~n21587 & n31060 ) | ( ~n21587 & n31062 ) | ( n31060 & n31062 ) ;
  assign n31064 = ~x26 & n31062 ;
  assign n31065 = ~x26 & n31060 ;
  assign n31066 = ( ~n21587 & n31064 ) | ( ~n21587 & n31065 ) | ( n31064 & n31065 ) ;
  assign n31067 = x26 | n31065 ;
  assign n31068 = x26 | n31064 ;
  assign n31069 = ( ~n21587 & n31067 ) | ( ~n21587 & n31068 ) | ( n31067 & n31068 ) ;
  assign n31070 = ( ~n31063 & n31066 ) | ( ~n31063 & n31069 ) | ( n31066 & n31069 ) ;
  assign n31071 = n31055 & ~n31070 ;
  assign n31072 = n31055 | n31070 ;
  assign n31073 = ( ~n31055 & n31071 ) | ( ~n31055 & n31072 ) | ( n31071 & n31072 ) ;
  assign n31134 = n31129 | n31133 ;
  assign n31135 = n31073 & n31134 ;
  assign n31136 = n31073 | n31134 ;
  assign n31137 = ~n31135 & n31136 ;
  assign n31138 = n2928 & ~n23240 ;
  assign n31139 = n2925 & n23227 ;
  assign n31140 = ( n2925 & n23217 ) | ( n2925 & n31139 ) | ( n23217 & n31139 ) ;
  assign n31141 = n31138 | n31140 ;
  assign n31142 = n2932 & ~n23234 ;
  assign n31143 = n2932 & ~n23235 ;
  assign n31144 = ( ~n15882 & n31142 ) | ( ~n15882 & n31143 ) | ( n31142 & n31143 ) ;
  assign n31145 = n31141 | n31144 ;
  assign n31146 = n2936 | n31144 ;
  assign n31147 = n31141 | n31146 ;
  assign n31148 = ( ~n23587 & n31145 ) | ( ~n23587 & n31147 ) | ( n31145 & n31147 ) ;
  assign n31149 = ~x23 & n31147 ;
  assign n31150 = ~x23 & n31145 ;
  assign n31151 = ( ~n23587 & n31149 ) | ( ~n23587 & n31150 ) | ( n31149 & n31150 ) ;
  assign n31152 = x23 | n31150 ;
  assign n31153 = x23 | n31149 ;
  assign n31154 = ( ~n23587 & n31152 ) | ( ~n23587 & n31153 ) | ( n31152 & n31153 ) ;
  assign n31155 = ( ~n31148 & n31151 ) | ( ~n31148 & n31154 ) | ( n31151 & n31154 ) ;
  assign n31156 = n31137 & ~n31155 ;
  assign n31157 = n31137 | n31155 ;
  assign n31158 = ( ~n31137 & n31156 ) | ( ~n31137 & n31157 ) | ( n31156 & n31157 ) ;
  assign n31209 = n31158 & n31208 ;
  assign n31210 = n31208 & ~n31209 ;
  assign n31211 = n31158 & ~n31208 ;
  assign n31212 = n31210 | n31211 ;
  assign n31268 = n31253 | n31267 ;
  assign n31273 = ~n31253 & n31272 ;
  assign n31274 = ( n30173 & n31268 ) | ( n30173 & ~n31273 ) | ( n31268 & ~n31273 ) ;
  assign n31275 = n31212 & n31274 ;
  assign n31279 = n31253 | n31278 ;
  assign n31280 = n31212 & n31279 ;
  assign n31283 = ~n31253 & n31282 ;
  assign n31284 = n31212 & ~n31283 ;
  assign n31285 = ( n30169 & n31280 ) | ( n30169 & n31284 ) | ( n31280 & n31284 ) ;
  assign n31286 = ( n28465 & n31275 ) | ( n28465 & n31285 ) | ( n31275 & n31285 ) ;
  assign n31287 = n31275 & n31285 ;
  assign n31288 = ( n28489 & n31286 ) | ( n28489 & n31287 ) | ( n31286 & n31287 ) ;
  assign n31289 = ( n30169 & n31279 ) | ( n30169 & ~n31283 ) | ( n31279 & ~n31283 ) ;
  assign n31290 = n31274 & n31289 ;
  assign n31291 = n31212 | n31290 ;
  assign n31292 = ( n28465 & n31274 ) | ( n28465 & n31289 ) | ( n31274 & n31289 ) ;
  assign n31293 = n31212 | n31292 ;
  assign n31294 = ( n28489 & n31291 ) | ( n28489 & n31293 ) | ( n31291 & n31293 ) ;
  assign n31295 = ~n31288 & n31294 ;
  assign n31296 = n7079 & n31295 ;
  assign n31327 = n7078 | n31296 ;
  assign n31328 = n31325 | n31327 ;
  assign n31326 = n31296 | n31325 ;
  assign n31329 = n31326 & n31328 ;
  assign n31330 = n31295 & ~n31323 ;
  assign n31331 = ~n31295 & n31323 ;
  assign n31332 = n31309 | n31323 ;
  assign n31333 = n30186 | n31309 ;
  assign n31334 = n30186 & n31309 ;
  assign n31335 = n31333 & ~n31334 ;
  assign n31336 = ~n30216 & n31333 ;
  assign n31337 = ( n31333 & ~n31335 ) | ( n31333 & n31336 ) | ( ~n31335 & n31336 ) ;
  assign n31338 = n31309 & n31323 ;
  assign n31339 = n31332 & ~n31338 ;
  assign n31340 = n31332 & ~n31339 ;
  assign n31341 = ( n31332 & n31337 ) | ( n31332 & n31340 ) | ( n31337 & n31340 ) ;
  assign n31342 = n31331 | n31341 ;
  assign n31343 = n31330 | n31342 ;
  assign n31344 = n31333 | n31338 ;
  assign n31345 = ( ~n31335 & n31338 ) | ( ~n31335 & n31344 ) | ( n31338 & n31344 ) ;
  assign n31346 = n31331 | n31332 ;
  assign n31347 = ( n31331 & n31345 ) | ( n31331 & n31346 ) | ( n31345 & n31346 ) ;
  assign n31348 = n31330 | n31347 ;
  assign n31349 = ( ~n30232 & n31343 ) | ( ~n30232 & n31348 ) | ( n31343 & n31348 ) ;
  assign n31350 = n31330 | n31331 ;
  assign n31351 = n31332 & n31345 ;
  assign n31352 = n31350 & n31351 ;
  assign n31353 = n31341 & n31350 ;
  assign n31354 = ( ~n30232 & n31352 ) | ( ~n30232 & n31353 ) | ( n31352 & n31353 ) ;
  assign n31355 = n31349 & ~n31354 ;
  assign n31356 = ( n31328 & n31329 ) | ( n31328 & n31355 ) | ( n31329 & n31355 ) ;
  assign n31357 = x8 & n31329 ;
  assign n31358 = x8 & n31328 ;
  assign n31359 = ( n31355 & n31357 ) | ( n31355 & n31358 ) | ( n31357 & n31358 ) ;
  assign n31360 = x8 & ~n31357 ;
  assign n31361 = x8 & ~n31358 ;
  assign n31362 = ( ~n31355 & n31360 ) | ( ~n31355 & n31361 ) | ( n31360 & n31361 ) ;
  assign n31363 = ( n31356 & ~n31359 ) | ( n31356 & n31362 ) | ( ~n31359 & n31362 ) ;
  assign n31364 = ~n30846 & n31363 ;
  assign n31365 = n30846 | n31364 ;
  assign n31366 = n30846 & n31363 ;
  assign n31367 = n31365 & ~n31366 ;
  assign n31368 = ~n30287 & n30841 ;
  assign n31369 = n30287 & ~n30841 ;
  assign n31370 = n31368 | n31369 ;
  assign n31371 = n31333 & ~n31335 ;
  assign n31372 = ( ~n30232 & n31337 ) | ( ~n30232 & n31371 ) | ( n31337 & n31371 ) ;
  assign n31373 = n31332 & ~n31345 ;
  assign n31374 = ~n31337 & n31339 ;
  assign n31375 = ( n30232 & n31373 ) | ( n30232 & n31374 ) | ( n31373 & n31374 ) ;
  assign n31376 = n31372 | n31375 ;
  assign n31377 = n7074 & ~n30186 ;
  assign n31378 = n7068 & ~n31309 ;
  assign n31379 = n31377 | n31378 ;
  assign n31380 = n7079 & ~n31323 ;
  assign n31381 = n7078 | n31380 ;
  assign n31382 = n31379 | n31381 ;
  assign n31383 = n31379 | n31380 ;
  assign n31384 = ~n31338 & n31341 ;
  assign n31385 = n31383 | n31384 ;
  assign n31386 = ~n31338 & n31351 ;
  assign n31387 = n31383 | n31386 ;
  assign n31388 = ( ~n30232 & n31385 ) | ( ~n30232 & n31387 ) | ( n31385 & n31387 ) ;
  assign n31389 = n31382 & n31388 ;
  assign n31390 = ( ~n31376 & n31382 ) | ( ~n31376 & n31389 ) | ( n31382 & n31389 ) ;
  assign n31391 = x8 & n31390 ;
  assign n31392 = x8 & ~n31390 ;
  assign n31393 = ( n31390 & ~n31391 ) | ( n31390 & n31392 ) | ( ~n31391 & n31392 ) ;
  assign n31394 = ~n31370 & n31393 ;
  assign n31395 = n31370 | n31394 ;
  assign n31396 = n31370 & n31393 ;
  assign n31397 = n31395 & ~n31396 ;
  assign n31398 = n30312 | n30839 ;
  assign n31399 = ~n30840 & n31398 ;
  assign n31400 = n30216 & n31335 ;
  assign n31401 = ( n30232 & n31335 ) | ( n30232 & n31400 ) | ( n31335 & n31400 ) ;
  assign n31402 = n30216 | n31335 ;
  assign n31403 = n30232 | n31402 ;
  assign n31404 = ~n31401 & n31403 ;
  assign n31406 = n7074 & n30212 ;
  assign n31407 = n7068 & ~n30186 ;
  assign n31408 = n31406 | n31407 ;
  assign n31405 = n7079 & ~n31309 ;
  assign n31410 = n7078 | n31405 ;
  assign n31411 = n31408 | n31410 ;
  assign n31409 = n31405 | n31408 ;
  assign n31412 = n31409 & n31411 ;
  assign n31413 = ( n31404 & n31411 ) | ( n31404 & n31412 ) | ( n31411 & n31412 ) ;
  assign n31414 = x8 & n31412 ;
  assign n31415 = x8 & n31411 ;
  assign n31416 = ( n31404 & n31414 ) | ( n31404 & n31415 ) | ( n31414 & n31415 ) ;
  assign n31417 = x8 & ~n31414 ;
  assign n31418 = x8 & ~n31415 ;
  assign n31419 = ( ~n31404 & n31417 ) | ( ~n31404 & n31418 ) | ( n31417 & n31418 ) ;
  assign n31420 = ( n31413 & ~n31416 ) | ( n31413 & n31419 ) | ( ~n31416 & n31419 ) ;
  assign n31421 = n31399 & n31420 ;
  assign n31422 = n31399 & ~n31421 ;
  assign n31423 = ~n31399 & n31420 ;
  assign n31424 = n31422 | n31423 ;
  assign n31425 = n30331 & ~n30837 ;
  assign n31426 = n30838 | n31425 ;
  assign n31428 = n7074 & ~n30199 ;
  assign n31429 = n7068 & n30212 ;
  assign n31430 = n31428 | n31429 ;
  assign n31427 = n7079 & ~n30186 ;
  assign n31432 = n7078 | n31427 ;
  assign n31433 = n31430 | n31432 ;
  assign n31431 = n31427 | n31430 ;
  assign n31434 = n31431 & n31433 ;
  assign n31435 = ( ~n30241 & n31433 ) | ( ~n30241 & n31434 ) | ( n31433 & n31434 ) ;
  assign n31436 = ~x8 & n31434 ;
  assign n31437 = ~x8 & n31433 ;
  assign n31438 = ( ~n30241 & n31436 ) | ( ~n30241 & n31437 ) | ( n31436 & n31437 ) ;
  assign n31439 = x8 | n31436 ;
  assign n31440 = x8 | n31437 ;
  assign n31441 = ( ~n30241 & n31439 ) | ( ~n30241 & n31440 ) | ( n31439 & n31440 ) ;
  assign n31442 = ( ~n31435 & n31438 ) | ( ~n31435 & n31441 ) | ( n31438 & n31441 ) ;
  assign n31443 = ~n31426 & n31442 ;
  assign n31444 = n31426 | n31443 ;
  assign n31445 = n31426 & n31442 ;
  assign n31446 = n31444 & ~n31445 ;
  assign n31447 = ~n30355 & n30835 ;
  assign n31448 = n30355 & ~n30835 ;
  assign n31449 = n31447 | n31448 ;
  assign n31450 = n7079 & n30212 ;
  assign n31451 = n7074 & n29620 ;
  assign n31452 = n7068 & ~n30199 ;
  assign n31453 = n31451 | n31452 ;
  assign n31454 = n31450 | n31453 ;
  assign n31455 = n30266 & ~n31454 ;
  assign n31456 = ~n30276 & n31455 ;
  assign n31457 = n7078 | n31450 ;
  assign n31458 = n31453 | n31457 ;
  assign n31459 = ~n31456 & n31458 ;
  assign n31460 = x8 & n31458 ;
  assign n31461 = ~n31456 & n31460 ;
  assign n31462 = x8 & ~n31460 ;
  assign n31463 = ( x8 & n31456 ) | ( x8 & n31462 ) | ( n31456 & n31462 ) ;
  assign n31464 = ( n31459 & ~n31461 ) | ( n31459 & n31463 ) | ( ~n31461 & n31463 ) ;
  assign n31465 = ~n31449 & n31464 ;
  assign n31466 = n31449 | n31465 ;
  assign n31467 = n31449 & n31464 ;
  assign n31468 = n31466 & ~n31467 ;
  assign n31469 = ( n30399 & n30400 ) | ( n30399 & n30833 ) | ( n30400 & n30833 ) ;
  assign n31470 = n30376 | n30399 ;
  assign n31471 = n30833 | n31470 ;
  assign n31472 = ~n31469 & n31471 ;
  assign n31473 = n7079 & ~n30199 ;
  assign n31474 = n7074 & ~n28714 ;
  assign n31475 = n7068 & n29620 ;
  assign n31476 = n31474 | n31475 ;
  assign n31477 = n31473 | n31476 ;
  assign n31478 = n7078 | n31473 ;
  assign n31479 = n31476 | n31478 ;
  assign n31480 = ( ~n30299 & n31477 ) | ( ~n30299 & n31479 ) | ( n31477 & n31479 ) ;
  assign n31481 = ~x8 & n31479 ;
  assign n31482 = ~x8 & n31477 ;
  assign n31483 = ( ~n30299 & n31481 ) | ( ~n30299 & n31482 ) | ( n31481 & n31482 ) ;
  assign n31484 = x8 | n31482 ;
  assign n31485 = x8 | n31481 ;
  assign n31486 = ( ~n30299 & n31484 ) | ( ~n30299 & n31485 ) | ( n31484 & n31485 ) ;
  assign n31487 = ( ~n31480 & n31483 ) | ( ~n31480 & n31486 ) | ( n31483 & n31486 ) ;
  assign n31488 = n31472 & n31487 ;
  assign n31489 = n30829 & ~n30833 ;
  assign n31490 = n30832 & ~n30833 ;
  assign n31491 = n31489 | n31490 ;
  assign n31492 = n7079 & n29620 ;
  assign n31493 = n7074 & n28492 ;
  assign n31494 = n7068 & ~n28714 ;
  assign n31495 = n31493 | n31494 ;
  assign n31496 = n31492 | n31495 ;
  assign n31497 = n7078 | n31492 ;
  assign n31498 = n31495 | n31497 ;
  assign n31499 = ( ~n29642 & n31496 ) | ( ~n29642 & n31498 ) | ( n31496 & n31498 ) ;
  assign n31500 = n31496 | n31498 ;
  assign n31501 = ( n29629 & n31499 ) | ( n29629 & n31500 ) | ( n31499 & n31500 ) ;
  assign n31502 = ~x8 & n31501 ;
  assign n31503 = x8 | n31501 ;
  assign n31504 = ( ~n31501 & n31502 ) | ( ~n31501 & n31503 ) | ( n31502 & n31503 ) ;
  assign n31505 = n31491 & n31504 ;
  assign n31506 = n31491 & ~n31505 ;
  assign n31507 = ~n31491 & n31504 ;
  assign n31508 = n31506 | n31507 ;
  assign n31509 = n30424 | n30827 ;
  assign n31510 = ~n30828 & n31509 ;
  assign n31511 = n7068 & n28492 ;
  assign n31512 = n7074 & ~n28503 ;
  assign n31513 = n28498 & n31512 ;
  assign n31514 = n31511 | n31513 ;
  assign n31515 = n7079 & ~n28714 ;
  assign n31516 = n7078 | n31515 ;
  assign n31517 = n31514 | n31516 ;
  assign n31518 = n31514 | n31515 ;
  assign n31519 = n28731 & ~n31518 ;
  assign n31520 = ( n28518 & ~n31518 ) | ( n28518 & n31519 ) | ( ~n31518 & n31519 ) ;
  assign n31521 = n31517 & ~n31520 ;
  assign n31522 = ( n28720 & n31517 ) | ( n28720 & n31521 ) | ( n31517 & n31521 ) ;
  assign n31523 = x8 & n31522 ;
  assign n31524 = x8 & ~n31522 ;
  assign n31525 = ( n31522 & ~n31523 ) | ( n31522 & n31524 ) | ( ~n31523 & n31524 ) ;
  assign n31526 = n31510 & n31525 ;
  assign n31527 = n30468 | n30821 ;
  assign n31528 = ~n30822 & n31527 ;
  assign n31529 = n7074 & ~n27371 ;
  assign n31530 = ~n27363 & n31529 ;
  assign n31531 = n7068 & ~n27606 ;
  assign n31532 = ~n27597 & n31531 ;
  assign n31533 = n31530 | n31532 ;
  assign n31534 = n7079 & ~n28503 ;
  assign n31535 = n28498 & n31534 ;
  assign n31536 = n31533 | n31535 ;
  assign n31537 = n28794 | n31536 ;
  assign n31538 = n28783 | n31537 ;
  assign n31539 = n7078 | n31535 ;
  assign n31540 = n31533 | n31539 ;
  assign n31541 = n31538 & n31540 ;
  assign n31542 = ~x8 & n31540 ;
  assign n31543 = n31538 & n31542 ;
  assign n31544 = x8 | n31542 ;
  assign n31545 = ( x8 & n31538 ) | ( x8 & n31544 ) | ( n31538 & n31544 ) ;
  assign n31546 = ( ~n31541 & n31543 ) | ( ~n31541 & n31545 ) | ( n31543 & n31545 ) ;
  assign n31547 = n31528 & n31546 ;
  assign n31548 = n30817 & n30819 ;
  assign n31549 = n30817 | n30819 ;
  assign n31550 = ~n31548 & n31549 ;
  assign n31551 = n7074 & ~n27133 ;
  assign n31552 = ~n27125 & n31551 ;
  assign n31553 = n7068 & ~n27371 ;
  assign n31554 = ~n27363 & n31553 ;
  assign n31555 = n31552 | n31554 ;
  assign n31556 = n7079 & ~n27606 ;
  assign n31557 = ~n27597 & n31556 ;
  assign n31558 = n31555 | n31557 ;
  assign n31559 = n7078 & n27630 ;
  assign n31560 = ~n27625 & n31559 ;
  assign n31561 = ( n7078 & ~n27634 ) | ( n7078 & n31560 ) | ( ~n27634 & n31560 ) ;
  assign n31562 = n31558 | n31561 ;
  assign n31563 = x8 | n31558 ;
  assign n31564 = n31561 | n31563 ;
  assign n31565 = ~x8 & n31563 ;
  assign n31566 = ( ~x8 & n31561 ) | ( ~x8 & n31565 ) | ( n31561 & n31565 ) ;
  assign n31567 = ( ~n31562 & n31564 ) | ( ~n31562 & n31566 ) | ( n31564 & n31566 ) ;
  assign n31568 = n31550 & n31567 ;
  assign n31569 = ~n31550 & n31567 ;
  assign n31570 = ( n31550 & ~n31568 ) | ( n31550 & n31569 ) | ( ~n31568 & n31569 ) ;
  assign n31571 = ~n30511 & n30815 ;
  assign n31572 = n30511 & ~n30815 ;
  assign n31573 = n31571 | n31572 ;
  assign n31574 = n7074 & ~n26526 ;
  assign n31575 = ~n26520 & n31574 ;
  assign n31576 = n7068 & ~n27133 ;
  assign n31577 = ~n27125 & n31576 ;
  assign n31578 = n31575 | n31577 ;
  assign n31579 = n7079 & ~n27371 ;
  assign n31580 = ~n27363 & n31579 ;
  assign n31581 = n31578 | n31580 ;
  assign n31582 = n7078 | n31580 ;
  assign n31583 = n31578 | n31582 ;
  assign n31584 = ( ~n27654 & n31581 ) | ( ~n27654 & n31583 ) | ( n31581 & n31583 ) ;
  assign n31585 = ~x8 & n31583 ;
  assign n31586 = ~x8 & n31581 ;
  assign n31587 = ( ~n27654 & n31585 ) | ( ~n27654 & n31586 ) | ( n31585 & n31586 ) ;
  assign n31588 = x8 | n31586 ;
  assign n31589 = x8 | n31585 ;
  assign n31590 = ( ~n27654 & n31588 ) | ( ~n27654 & n31589 ) | ( n31588 & n31589 ) ;
  assign n31591 = ( ~n31584 & n31587 ) | ( ~n31584 & n31590 ) | ( n31587 & n31590 ) ;
  assign n31592 = n31573 & n31591 ;
  assign n31593 = ~n30531 & n30813 ;
  assign n31594 = n30531 & ~n30813 ;
  assign n31595 = n31593 | n31594 ;
  assign n31596 = n7074 & ~n26270 ;
  assign n31597 = ~n26263 & n31596 ;
  assign n31598 = n7068 & ~n26526 ;
  assign n31599 = ~n26520 & n31598 ;
  assign n31600 = n31597 | n31599 ;
  assign n31601 = n7079 & ~n27133 ;
  assign n31602 = ~n27125 & n31601 ;
  assign n31603 = n31600 | n31602 ;
  assign n31604 = n7078 & n27699 ;
  assign n31605 = ( n7078 & ~n27696 ) | ( n7078 & n31604 ) | ( ~n27696 & n31604 ) ;
  assign n31606 = n31603 | n31605 ;
  assign n31607 = x8 | n31603 ;
  assign n31608 = n31605 | n31607 ;
  assign n31609 = ~x8 & n31607 ;
  assign n31610 = ( ~x8 & n31605 ) | ( ~x8 & n31609 ) | ( n31605 & n31609 ) ;
  assign n31611 = ( ~n31606 & n31608 ) | ( ~n31606 & n31610 ) | ( n31608 & n31610 ) ;
  assign n31612 = n31595 & n31611 ;
  assign n31613 = n31595 | n31611 ;
  assign n31614 = ~n31612 & n31613 ;
  assign n31615 = n30809 & n30811 ;
  assign n31616 = n30809 | n30811 ;
  assign n31617 = ~n31615 & n31616 ;
  assign n31618 = n7074 & n26017 ;
  assign n31619 = n7068 & ~n26270 ;
  assign n31620 = ~n26263 & n31619 ;
  assign n31621 = n31618 | n31620 ;
  assign n31622 = n7079 & ~n26526 ;
  assign n31623 = ~n26520 & n31622 ;
  assign n31625 = n7078 | n31623 ;
  assign n31626 = n31621 | n31625 ;
  assign n31624 = n31621 | n31623 ;
  assign n31627 = n31624 & n31626 ;
  assign n31628 = ( ~n26555 & n31626 ) | ( ~n26555 & n31627 ) | ( n31626 & n31627 ) ;
  assign n31629 = ( n26528 & n31626 ) | ( n26528 & n31627 ) | ( n31626 & n31627 ) ;
  assign n31630 = ( ~n26543 & n31628 ) | ( ~n26543 & n31629 ) | ( n31628 & n31629 ) ;
  assign n31631 = ~x8 & n31630 ;
  assign n31632 = x8 | n31630 ;
  assign n31633 = ( ~n31630 & n31631 ) | ( ~n31630 & n31632 ) | ( n31631 & n31632 ) ;
  assign n31634 = n31617 & n31633 ;
  assign n31635 = n30574 | n30807 ;
  assign n31636 = ~n30808 & n31635 ;
  assign n31637 = n7074 & ~n25728 ;
  assign n31638 = n7068 & n26017 ;
  assign n31639 = n31637 | n31638 ;
  assign n31640 = n7079 & ~n26270 ;
  assign n31641 = ~n26263 & n31640 ;
  assign n31643 = n7078 | n31641 ;
  assign n31644 = n31639 | n31643 ;
  assign n31642 = n31639 | n31641 ;
  assign n31645 = n31642 & n31644 ;
  assign n31646 = ( n26571 & n31644 ) | ( n26571 & n31645 ) | ( n31644 & n31645 ) ;
  assign n31647 = x8 & n31645 ;
  assign n31648 = x8 & n31644 ;
  assign n31649 = ( n26571 & n31647 ) | ( n26571 & n31648 ) | ( n31647 & n31648 ) ;
  assign n31650 = x8 & ~n31647 ;
  assign n31651 = x8 & ~n31648 ;
  assign n31652 = ( ~n26571 & n31650 ) | ( ~n26571 & n31651 ) | ( n31650 & n31651 ) ;
  assign n31653 = ( n31646 & ~n31649 ) | ( n31646 & n31652 ) | ( ~n31649 & n31652 ) ;
  assign n31654 = n31636 & n31653 ;
  assign n31655 = n31636 & ~n31654 ;
  assign n31656 = ~n31636 & n31653 ;
  assign n31657 = n31655 | n31656 ;
  assign n31658 = n30595 & n30805 ;
  assign n31659 = n30595 | n30805 ;
  assign n31660 = ~n31658 & n31659 ;
  assign n31661 = n7079 & n26017 ;
  assign n31662 = n7074 & ~n25046 ;
  assign n31663 = n7068 & ~n25728 ;
  assign n31664 = n31662 | n31663 ;
  assign n31665 = n31661 | n31664 ;
  assign n31666 = n7078 | n31661 ;
  assign n31667 = n31664 | n31666 ;
  assign n31668 = ( n26613 & n31665 ) | ( n26613 & n31667 ) | ( n31665 & n31667 ) ;
  assign n31669 = n31665 | n31667 ;
  assign n31670 = ( n26605 & n31668 ) | ( n26605 & n31669 ) | ( n31668 & n31669 ) ;
  assign n31671 = x8 & n31670 ;
  assign n31672 = x8 & ~n31670 ;
  assign n31673 = ( n31670 & ~n31671 ) | ( n31670 & n31672 ) | ( ~n31671 & n31672 ) ;
  assign n31674 = n31660 & n31673 ;
  assign n31675 = n31660 & ~n31674 ;
  assign n31676 = ~n31660 & n31673 ;
  assign n31677 = n31675 | n31676 ;
  assign n31678 = ( n30631 & n30632 ) | ( n30631 & n30803 ) | ( n30632 & n30803 ) ;
  assign n31679 = n30610 | n30631 ;
  assign n31680 = n30803 | n31679 ;
  assign n31681 = ~n31678 & n31680 ;
  assign n31682 = n7079 & ~n25728 ;
  assign n31683 = n7074 & n24770 ;
  assign n31684 = n7068 & ~n25046 ;
  assign n31685 = n31683 | n31684 ;
  assign n31686 = n31682 | n31685 ;
  assign n31687 = n7078 & n25740 ;
  assign n31688 = n7078 & n25731 ;
  assign n31689 = ( ~n25441 & n31687 ) | ( ~n25441 & n31688 ) | ( n31687 & n31688 ) ;
  assign n31690 = n31686 | n31689 ;
  assign n31691 = n7078 | n31686 ;
  assign n31692 = ( n25733 & n31690 ) | ( n25733 & n31691 ) | ( n31690 & n31691 ) ;
  assign n31693 = x8 | n31692 ;
  assign n31694 = ~x8 & n31692 ;
  assign n31695 = ( ~n31692 & n31693 ) | ( ~n31692 & n31694 ) | ( n31693 & n31694 ) ;
  assign n31696 = n31681 & n31695 ;
  assign n31697 = n30800 & ~n30803 ;
  assign n31700 = n7079 & ~n25046 ;
  assign n31701 = n7074 & ~n25054 ;
  assign n31702 = n7068 & n24770 ;
  assign n31703 = n31701 | n31702 ;
  assign n31704 = n31700 | n31703 ;
  assign n31705 = n7078 | n31700 ;
  assign n31706 = n31703 | n31705 ;
  assign n31707 = ( ~n25069 & n31704 ) | ( ~n25069 & n31706 ) | ( n31704 & n31706 ) ;
  assign n31708 = ~x8 & n31706 ;
  assign n31709 = ~x8 & n31704 ;
  assign n31710 = ( ~n25069 & n31708 ) | ( ~n25069 & n31709 ) | ( n31708 & n31709 ) ;
  assign n31711 = x8 | n31709 ;
  assign n31712 = x8 | n31708 ;
  assign n31713 = ( ~n25069 & n31711 ) | ( ~n25069 & n31712 ) | ( n31711 & n31712 ) ;
  assign n31714 = ( ~n31707 & n31710 ) | ( ~n31707 & n31713 ) | ( n31710 & n31713 ) ;
  assign n31698 = ~n30800 & n30802 ;
  assign n31715 = n31698 & n31714 ;
  assign n31716 = ( n31697 & n31714 ) | ( n31697 & n31715 ) | ( n31714 & n31715 ) ;
  assign n31699 = n31697 | n31698 ;
  assign n31717 = n31699 & ~n31716 ;
  assign n31718 = ~n31698 & n31714 ;
  assign n31719 = ~n31697 & n31718 ;
  assign n31720 = n31717 | n31719 ;
  assign n31721 = n30798 & ~n30799 ;
  assign n31722 = n30655 & ~n30799 ;
  assign n31723 = n31721 | n31722 ;
  assign n31724 = n7079 & n24770 ;
  assign n31725 = n7074 & n24167 ;
  assign n31726 = n7068 & ~n25054 ;
  assign n31727 = n31725 | n31726 ;
  assign n31728 = n31724 | n31727 ;
  assign n31729 = n7078 | n31728 ;
  assign n31730 = ( ~n25095 & n31728 ) | ( ~n25095 & n31729 ) | ( n31728 & n31729 ) ;
  assign n31731 = ~x8 & n31729 ;
  assign n31732 = ~x8 & n31728 ;
  assign n31733 = ( ~n25095 & n31731 ) | ( ~n25095 & n31732 ) | ( n31731 & n31732 ) ;
  assign n31734 = x8 | n31731 ;
  assign n31735 = x8 | n31732 ;
  assign n31736 = ( ~n25095 & n31734 ) | ( ~n25095 & n31735 ) | ( n31734 & n31735 ) ;
  assign n31737 = ( ~n31730 & n31733 ) | ( ~n31730 & n31736 ) | ( n31733 & n31736 ) ;
  assign n31738 = n31723 & n31737 ;
  assign n31739 = n31723 & ~n31738 ;
  assign n31740 = ~n31723 & n31737 ;
  assign n31741 = n31739 | n31740 ;
  assign n31742 = n30677 | n30771 ;
  assign n31743 = ~n30772 & n31742 ;
  assign n31744 = n7079 & n24167 ;
  assign n31745 = n7074 & n23316 ;
  assign n31746 = n7068 & n23614 ;
  assign n31747 = n31745 | n31746 ;
  assign n31748 = n31744 | n31747 ;
  assign n31749 = n7078 | n31748 ;
  assign n31750 = ( n24182 & n31748 ) | ( n24182 & n31749 ) | ( n31748 & n31749 ) ;
  assign n31751 = n31748 | n31749 ;
  assign n31752 = ( n24175 & n31750 ) | ( n24175 & n31751 ) | ( n31750 & n31751 ) ;
  assign n31753 = x8 & n31752 ;
  assign n31754 = x8 & ~n31752 ;
  assign n31755 = ( n31752 & ~n31753 ) | ( n31752 & n31754 ) | ( ~n31753 & n31754 ) ;
  assign n31756 = n31743 & n31755 ;
  assign n31757 = n30773 & n30796 ;
  assign n31758 = n30773 | n30796 ;
  assign n31759 = ~n31757 & n31758 ;
  assign n31760 = n7079 & ~n25054 ;
  assign n31761 = n7074 & n23614 ;
  assign n31762 = n7068 & n24167 ;
  assign n31763 = n31761 | n31762 ;
  assign n31764 = n31760 | n31763 ;
  assign n31765 = n7078 | n31760 ;
  assign n31766 = n31763 | n31765 ;
  assign n31767 = ( ~n25122 & n31764 ) | ( ~n25122 & n31766 ) | ( n31764 & n31766 ) ;
  assign n31768 = ~x8 & n31766 ;
  assign n31769 = ~x8 & n31764 ;
  assign n31770 = ( ~n25122 & n31768 ) | ( ~n25122 & n31769 ) | ( n31768 & n31769 ) ;
  assign n31771 = x8 | n31769 ;
  assign n31772 = x8 | n31768 ;
  assign n31773 = ( ~n25122 & n31771 ) | ( ~n25122 & n31772 ) | ( n31771 & n31772 ) ;
  assign n31774 = ( ~n31767 & n31770 ) | ( ~n31767 & n31773 ) | ( n31770 & n31773 ) ;
  assign n31775 = n31759 & n31774 ;
  assign n31776 = n31759 | n31774 ;
  assign n31777 = ~n31775 & n31776 ;
  assign n31778 = n31756 & n31777 ;
  assign n31779 = n31775 | n31777 ;
  assign n31780 = n30696 | n30769 ;
  assign n31781 = ~n30770 & n31780 ;
  assign n31782 = n7079 & n23614 ;
  assign n31783 = n7074 & n23620 ;
  assign n31784 = ( n7068 & n7314 ) | ( n7068 & n23620 ) | ( n7314 & n23620 ) ;
  assign n31785 = ( n23316 & n31783 ) | ( n23316 & n31784 ) | ( n31783 & n31784 ) ;
  assign n31787 = n7078 | n31785 ;
  assign n31788 = n31782 | n31787 ;
  assign n31786 = n31782 | n31785 ;
  assign n31789 = n31786 & n31788 ;
  assign n31790 = ( n23634 & n31788 ) | ( n23634 & n31789 ) | ( n31788 & n31789 ) ;
  assign n31791 = x8 & n31789 ;
  assign n31792 = x8 & n31788 ;
  assign n31793 = ( n23634 & n31791 ) | ( n23634 & n31792 ) | ( n31791 & n31792 ) ;
  assign n31794 = x8 & ~n31791 ;
  assign n31795 = x8 & ~n31792 ;
  assign n31796 = ( ~n23634 & n31794 ) | ( ~n23634 & n31795 ) | ( n31794 & n31795 ) ;
  assign n31797 = ( n31790 & ~n31793 ) | ( n31790 & n31796 ) | ( ~n31793 & n31796 ) ;
  assign n31798 = n31781 & n31797 ;
  assign n31799 = n31781 & ~n31798 ;
  assign n31800 = ~n31781 & n31797 ;
  assign n31801 = n31799 | n31800 ;
  assign n31802 = n30749 & n30763 ;
  assign n31803 = n30749 & ~n31802 ;
  assign n31804 = n7074 & ~n22385 ;
  assign n31805 = ( n7068 & n7314 ) | ( n7068 & ~n22385 ) | ( n7314 & ~n22385 ) ;
  assign n31806 = ( n22381 & n31804 ) | ( n22381 & n31805 ) | ( n31804 & n31805 ) ;
  assign n31807 = n7079 | n31806 ;
  assign n31808 = ( n23620 & n31806 ) | ( n23620 & n31807 ) | ( n31806 & n31807 ) ;
  assign n31809 = n7078 | n31808 ;
  assign n31810 = ( ~n23686 & n31808 ) | ( ~n23686 & n31809 ) | ( n31808 & n31809 ) ;
  assign n31811 = ~x8 & n31809 ;
  assign n31812 = ~x8 & n31808 ;
  assign n31813 = ( ~n23686 & n31811 ) | ( ~n23686 & n31812 ) | ( n31811 & n31812 ) ;
  assign n31814 = x8 | n31811 ;
  assign n31815 = x8 | n31812 ;
  assign n31816 = ( ~n23686 & n31814 ) | ( ~n23686 & n31815 ) | ( n31814 & n31815 ) ;
  assign n31817 = ( ~n31810 & n31813 ) | ( ~n31810 & n31816 ) | ( n31813 & n31816 ) ;
  assign n31818 = ~n30749 & n30763 ;
  assign n31819 = n31817 & n31818 ;
  assign n31820 = ( n31803 & n31817 ) | ( n31803 & n31819 ) | ( n31817 & n31819 ) ;
  assign n31821 = n31817 | n31818 ;
  assign n31822 = n31803 | n31821 ;
  assign n31823 = ~n31820 & n31822 ;
  assign n31824 = n30728 & n30746 ;
  assign n31825 = n30728 | n30746 ;
  assign n31826 = ~n31824 & n31825 ;
  assign n31827 = n7079 & n22381 ;
  assign n31828 = n7074 & ~n22398 ;
  assign n31829 = n7068 & ~n22385 ;
  assign n31830 = n31828 | n31829 ;
  assign n31831 = n31827 | n31830 ;
  assign n31832 = n7078 | n31831 ;
  assign n31833 = x8 & n31832 ;
  assign n31834 = x8 & n31831 ;
  assign n31835 = ( n22422 & n31833 ) | ( n22422 & n31834 ) | ( n31833 & n31834 ) ;
  assign n31836 = x8 | n31832 ;
  assign n31837 = x8 | n31831 ;
  assign n31838 = ( n22422 & n31836 ) | ( n22422 & n31837 ) | ( n31836 & n31837 ) ;
  assign n31839 = ~n31835 & n31838 ;
  assign n31840 = n31826 & n31839 ;
  assign n31841 = ~n31826 & n31839 ;
  assign n31842 = ( n31826 & ~n31840 ) | ( n31826 & n31841 ) | ( ~n31840 & n31841 ) ;
  assign n31843 = n30722 | n30724 ;
  assign n31844 = ~n30724 & n30726 ;
  assign n31845 = ( n30723 & n31843 ) | ( n30723 & ~n31844 ) | ( n31843 & ~n31844 ) ;
  assign n31846 = ~n30728 & n31845 ;
  assign n31847 = n7079 & ~n22385 ;
  assign n31848 = n7074 & n22393 ;
  assign n31849 = n7068 & ~n22398 ;
  assign n31850 = n31848 | n31849 ;
  assign n31851 = n31847 | n31850 ;
  assign n31852 = n7078 | n31847 ;
  assign n31853 = n31850 | n31852 ;
  assign n31854 = ( ~n22545 & n31851 ) | ( ~n22545 & n31853 ) | ( n31851 & n31853 ) ;
  assign n31855 = ~x8 & n31853 ;
  assign n31856 = ~x8 & n31851 ;
  assign n31857 = ( ~n22545 & n31855 ) | ( ~n22545 & n31856 ) | ( n31855 & n31856 ) ;
  assign n31858 = x8 | n31856 ;
  assign n31859 = x8 | n31855 ;
  assign n31860 = ( ~n22545 & n31858 ) | ( ~n22545 & n31859 ) | ( n31858 & n31859 ) ;
  assign n31861 = ( ~n31854 & n31857 ) | ( ~n31854 & n31860 ) | ( n31857 & n31860 ) ;
  assign n31862 = n31846 & n31861 ;
  assign n31863 = n7078 & n22474 ;
  assign n31864 = n7068 & ~n22409 ;
  assign n31865 = n7079 & ~n22406 ;
  assign n31866 = n31864 | n31865 ;
  assign n31867 = x8 | n31866 ;
  assign n31868 = n31863 | n31867 ;
  assign n31869 = ~x8 & n31868 ;
  assign n31870 = ( x8 & n20190 ) | ( x8 & n22409 ) | ( n20190 & n22409 ) ;
  assign n31871 = n31868 & n31870 ;
  assign n31872 = n31863 | n31866 ;
  assign n31873 = n31870 & ~n31872 ;
  assign n31874 = ( n31869 & n31871 ) | ( n31869 & n31873 ) | ( n31871 & n31873 ) ;
  assign n31875 = n7079 & n22393 ;
  assign n31876 = n7074 & ~n22409 ;
  assign n31877 = n7068 & ~n22406 ;
  assign n31878 = n31876 | n31877 ;
  assign n31879 = n31875 | n31878 ;
  assign n31880 = n22439 | n31879 ;
  assign n31881 = n7078 | n31875 ;
  assign n31882 = n31878 | n31881 ;
  assign n31883 = ~x8 & n31882 ;
  assign n31884 = n31880 & n31883 ;
  assign n31885 = x8 | n31884 ;
  assign n31886 = n6114 & ~n22409 ;
  assign n31887 = n31884 & n31886 ;
  assign n31888 = n31880 & n31882 ;
  assign n31889 = n31886 & ~n31888 ;
  assign n31890 = ( n31885 & n31887 ) | ( n31885 & n31889 ) | ( n31887 & n31889 ) ;
  assign n31891 = n31874 & n31890 ;
  assign n31892 = ( n31884 & n31885 ) | ( n31884 & ~n31888 ) | ( n31885 & ~n31888 ) ;
  assign n31893 = n31874 | n31886 ;
  assign n31894 = ( n31886 & n31892 ) | ( n31886 & n31893 ) | ( n31892 & n31893 ) ;
  assign n31895 = ~n31891 & n31894 ;
  assign n31896 = n7074 & ~n22406 ;
  assign n31897 = n7068 & n22393 ;
  assign n31898 = n31896 | n31897 ;
  assign n31899 = n7079 & ~n22398 ;
  assign n31900 = n7078 | n31899 ;
  assign n31901 = n31898 | n31900 ;
  assign n31902 = x8 & n31901 ;
  assign n31903 = n31898 | n31899 ;
  assign n31904 = x8 & n31903 ;
  assign n31905 = ( n22608 & n31902 ) | ( n22608 & n31904 ) | ( n31902 & n31904 ) ;
  assign n31906 = x8 | n31901 ;
  assign n31907 = x8 | n31903 ;
  assign n31908 = ( n22608 & n31906 ) | ( n22608 & n31907 ) | ( n31906 & n31907 ) ;
  assign n31909 = ~n31905 & n31908 ;
  assign n31910 = n31891 | n31909 ;
  assign n31911 = ( n31891 & n31895 ) | ( n31891 & n31910 ) | ( n31895 & n31910 ) ;
  assign n31912 = n31846 | n31861 ;
  assign n31913 = ~n31862 & n31912 ;
  assign n31914 = n31862 | n31913 ;
  assign n31915 = ( n31862 & n31911 ) | ( n31862 & n31914 ) | ( n31911 & n31914 ) ;
  assign n31916 = n31842 & n31915 ;
  assign n31917 = n31840 | n31916 ;
  assign n31918 = n31823 & n31917 ;
  assign n31919 = n31820 | n31918 ;
  assign n31920 = n7074 & n22381 ;
  assign n31921 = ( n7068 & n7314 ) | ( n7068 & n22381 ) | ( n7314 & n22381 ) ;
  assign n31922 = ( n23620 & n31920 ) | ( n23620 & n31921 ) | ( n31920 & n31921 ) ;
  assign n31923 = n7079 | n31921 ;
  assign n31924 = n7079 | n31920 ;
  assign n31925 = ( n23620 & n31923 ) | ( n23620 & n31924 ) | ( n31923 & n31924 ) ;
  assign n31926 = ( n23316 & n31922 ) | ( n23316 & n31925 ) | ( n31922 & n31925 ) ;
  assign n31927 = n7078 | n31926 ;
  assign n31928 = ~x8 & n31927 ;
  assign n31929 = ~x8 & n31926 ;
  assign n31930 = ( n23661 & n31928 ) | ( n23661 & n31929 ) | ( n31928 & n31929 ) ;
  assign n31931 = ( x8 & n20150 ) | ( x8 & n31926 ) | ( n20150 & n31926 ) ;
  assign n31932 = x8 & ~n31931 ;
  assign n31933 = x8 & n31926 ;
  assign n31934 = x8 & ~n31933 ;
  assign n31935 = ( ~n23661 & n31932 ) | ( ~n23661 & n31934 ) | ( n31932 & n31934 ) ;
  assign n31936 = n31930 | n31935 ;
  assign n31937 = n30765 & n30767 ;
  assign n31938 = n30765 | n30767 ;
  assign n31939 = ~n31937 & n31938 ;
  assign n31940 = n31936 & n31939 ;
  assign n31941 = n31936 | n31939 ;
  assign n31942 = ~n31940 & n31941 ;
  assign n31943 = n31940 | n31942 ;
  assign n31944 = ( n31919 & n31940 ) | ( n31919 & n31943 ) | ( n31940 & n31943 ) ;
  assign n31945 = n31801 & n31944 ;
  assign n31946 = n31798 | n31945 ;
  assign n31947 = ~n31743 & n31755 ;
  assign n31948 = ( n31743 & ~n31756 ) | ( n31743 & n31947 ) | ( ~n31756 & n31947 ) ;
  assign n31949 = n31946 & n31948 ;
  assign n31950 = n31775 | n31949 ;
  assign n31951 = ( n31778 & n31779 ) | ( n31778 & n31950 ) | ( n31779 & n31950 ) ;
  assign n31952 = n31738 | n31951 ;
  assign n31953 = ( n31738 & n31741 ) | ( n31738 & n31952 ) | ( n31741 & n31952 ) ;
  assign n31954 = n31720 & n31953 ;
  assign n31955 = n31716 | n31954 ;
  assign n31956 = ~n31681 & n31695 ;
  assign n31957 = ( n31681 & ~n31696 ) | ( n31681 & n31956 ) | ( ~n31696 & n31956 ) ;
  assign n31958 = n31696 | n31957 ;
  assign n31959 = ( n31696 & n31955 ) | ( n31696 & n31958 ) | ( n31955 & n31958 ) ;
  assign n31960 = n31674 | n31959 ;
  assign n31961 = ( n31674 & n31677 ) | ( n31674 & n31960 ) | ( n31677 & n31960 ) ;
  assign n31962 = n31657 & n31961 ;
  assign n31963 = n31654 | n31962 ;
  assign n31964 = n31617 | n31633 ;
  assign n31965 = ~n31634 & n31964 ;
  assign n31966 = n31634 | n31965 ;
  assign n31967 = ( n31634 & n31963 ) | ( n31634 & n31966 ) | ( n31963 & n31966 ) ;
  assign n31968 = n31614 & n31967 ;
  assign n31969 = n31612 | n31968 ;
  assign n31970 = n31573 | n31591 ;
  assign n31971 = ~n31592 & n31970 ;
  assign n31972 = n31592 | n31971 ;
  assign n31973 = ( n31592 & n31969 ) | ( n31592 & n31972 ) | ( n31969 & n31972 ) ;
  assign n31974 = n31570 & n31973 ;
  assign n31975 = n31568 | n31974 ;
  assign n31976 = n31528 & ~n31547 ;
  assign n31977 = ~n31528 & n31546 ;
  assign n31978 = n31976 | n31977 ;
  assign n31979 = n31975 & n31978 ;
  assign n31980 = n31547 | n31979 ;
  assign n31981 = n30823 & n30825 ;
  assign n31982 = n30823 | n30825 ;
  assign n31983 = ~n31981 & n31982 ;
  assign n31984 = n7079 & n28492 ;
  assign n31985 = n7074 & ~n27606 ;
  assign n31986 = ~n27597 & n31985 ;
  assign n31987 = n7068 & ~n28503 ;
  assign n31988 = n28498 & n31987 ;
  assign n31989 = n31986 | n31988 ;
  assign n31990 = n31984 | n31989 ;
  assign n31991 = n7078 | n31990 ;
  assign n31992 = n31990 & n31991 ;
  assign n31993 = ( ~n28749 & n31991 ) | ( ~n28749 & n31992 ) | ( n31991 & n31992 ) ;
  assign n31994 = ~x8 & n31992 ;
  assign n31995 = ~x8 & n31991 ;
  assign n31996 = ( ~n28749 & n31994 ) | ( ~n28749 & n31995 ) | ( n31994 & n31995 ) ;
  assign n31997 = x8 | n31994 ;
  assign n31998 = x8 | n31995 ;
  assign n31999 = ( ~n28749 & n31997 ) | ( ~n28749 & n31998 ) | ( n31997 & n31998 ) ;
  assign n32000 = ( ~n31993 & n31996 ) | ( ~n31993 & n31999 ) | ( n31996 & n31999 ) ;
  assign n32001 = n31983 & n32000 ;
  assign n32002 = n31983 & ~n32001 ;
  assign n32003 = ~n31983 & n32000 ;
  assign n32004 = n32002 | n32003 ;
  assign n32005 = n31980 & n32004 ;
  assign n32006 = n31510 | n31525 ;
  assign n32007 = ~n31526 & n32006 ;
  assign n32008 = n32001 & n32007 ;
  assign n32009 = ( n32005 & n32007 ) | ( n32005 & n32008 ) | ( n32007 & n32008 ) ;
  assign n32010 = n31526 | n32009 ;
  assign n32011 = n31505 | n32010 ;
  assign n32012 = ( n31505 & n31508 ) | ( n31505 & n32011 ) | ( n31508 & n32011 ) ;
  assign n32013 = ~n31472 & n31487 ;
  assign n32014 = ( n31472 & ~n31488 ) | ( n31472 & n32013 ) | ( ~n31488 & n32013 ) ;
  assign n32015 = n31488 | n32014 ;
  assign n32016 = ( n31488 & n32012 ) | ( n31488 & n32015 ) | ( n32012 & n32015 ) ;
  assign n32017 = n31465 | n32016 ;
  assign n32018 = ( n31465 & ~n31468 ) | ( n31465 & n32017 ) | ( ~n31468 & n32017 ) ;
  assign n32019 = ~n31446 & n32018 ;
  assign n32020 = n31443 | n32019 ;
  assign n32021 = n31424 & n32020 ;
  assign n32022 = n31421 | n32021 ;
  assign n32023 = n31394 | n32022 ;
  assign n32024 = ( n31394 & ~n31397 ) | ( n31394 & n32023 ) | ( ~n31397 & n32023 ) ;
  assign n32025 = n31367 & n32024 ;
  assign n32026 = n31367 | n32024 ;
  assign n32027 = ~n32025 & n32026 ;
  assign n32028 = n99 | n18477 ;
  assign n32029 = n262 | n1283 ;
  assign n32030 = n12687 | n32029 ;
  assign n32031 = n32028 | n32030 ;
  assign n32032 = n1690 | n6844 ;
  assign n32033 = n32031 | n32032 ;
  assign n32034 = n25367 | n32033 ;
  assign n32035 = n29916 | n32034 ;
  assign n32036 = n14423 | n32035 ;
  assign n32037 = n256 | n411 ;
  assign n32038 = n543 | n1398 ;
  assign n32039 = n32037 | n32038 ;
  assign n32040 = n344 | n356 ;
  assign n32041 = n59 | n32040 ;
  assign n32042 = n32039 | n32041 ;
  assign n32043 = n32036 | n32042 ;
  assign n32044 = n333 | n758 ;
  assign n32045 = n29278 | n29279 ;
  assign n32046 = n29294 | n32045 ;
  assign n32047 = n1482 | n18102 ;
  assign n32048 = n4004 | n32047 ;
  assign n32049 = n15222 | n32048 ;
  assign n32050 = n15221 | n32049 ;
  assign n32051 = n10748 | n25788 ;
  assign n32052 = n32050 | n32051 ;
  assign n32053 = n721 | n5946 ;
  assign n32054 = n3430 | n32053 ;
  assign n32055 = n7851 | n32054 ;
  assign n32056 = n291 | n412 ;
  assign n32057 = n340 | n32056 ;
  assign n32058 = n801 | n32057 ;
  assign n32059 = n32055 | n32058 ;
  assign n32060 = n32052 | n32059 ;
  assign n32061 = n32046 | n32060 ;
  assign n32062 = n32044 | n32061 ;
  assign n32063 = n32043 | n32062 ;
  assign n32064 = n32043 & n32062 ;
  assign n32065 = n32063 & ~n32064 ;
  assign n32066 = n2928 | n2932 ;
  assign n32067 = n2925 | n32066 ;
  assign n32068 = n2936 | n32067 ;
  assign n32069 = ~n23229 & n32068 ;
  assign n32070 = ( n23154 & n32068 ) | ( n23154 & n32069 ) | ( n32068 & n32069 ) ;
  assign n32071 = ~n23232 & n32068 ;
  assign n32072 = ~n23231 & n32068 ;
  assign n32073 = ( n9072 & n32071 ) | ( n9072 & n32072 ) | ( n32071 & n32072 ) ;
  assign n32074 = ( ~n21543 & n32070 ) | ( ~n21543 & n32073 ) | ( n32070 & n32073 ) ;
  assign n32075 = ( ~n21545 & n32070 ) | ( ~n21545 & n32073 ) | ( n32070 & n32073 ) ;
  assign n32076 = ( ~n15882 & n32074 ) | ( ~n15882 & n32075 ) | ( n32074 & n32075 ) ;
  assign n32077 = ~x23 & n32074 ;
  assign n32078 = ~x23 & n32075 ;
  assign n32079 = ( ~n15882 & n32077 ) | ( ~n15882 & n32078 ) | ( n32077 & n32078 ) ;
  assign n32080 = x23 | n32077 ;
  assign n32081 = x23 | n32078 ;
  assign n32082 = ( ~n15882 & n32080 ) | ( ~n15882 & n32081 ) | ( n32080 & n32081 ) ;
  assign n32083 = ( ~n32076 & n32079 ) | ( ~n32076 & n32082 ) | ( n32079 & n32082 ) ;
  assign n32084 = n32065 & ~n32083 ;
  assign n32085 = ~n32065 & n32083 ;
  assign n32086 = n32084 | n32085 ;
  assign n32087 = n30902 & ~n32043 ;
  assign n32088 = n30905 & ~n30910 ;
  assign n32089 = ( n30905 & ~n30915 ) | ( n30905 & n32088 ) | ( ~n30915 & n32088 ) ;
  assign n32090 = ~n30902 & n32043 ;
  assign n32091 = n32087 | n32090 ;
  assign n32092 = ~n32087 & n32091 ;
  assign n32093 = ( ~n32087 & n32089 ) | ( ~n32087 & n32092 ) | ( n32089 & n32092 ) ;
  assign n32094 = n30905 | n32090 ;
  assign n32095 = ( ~n30910 & n32090 ) | ( ~n30910 & n32094 ) | ( n32090 & n32094 ) ;
  assign n32096 = ~n32087 & n32095 ;
  assign n32097 = ( ~n30919 & n32093 ) | ( ~n30919 & n32096 ) | ( n32093 & n32096 ) ;
  assign n32098 = ( ~n1062 & n32093 ) | ( ~n1062 & n32096 ) | ( n32093 & n32096 ) ;
  assign n32099 = ( ~n19640 & n32097 ) | ( ~n19640 & n32098 ) | ( n32097 & n32098 ) ;
  assign n32100 = n32086 | n32099 ;
  assign n32101 = n32086 & n32099 ;
  assign n32102 = n32100 & ~n32101 ;
  assign n32103 = n1062 & n20680 ;
  assign n32104 = n1057 & ~n20618 ;
  assign n32105 = n1060 & n19631 ;
  assign n32106 = n1065 & ~n20630 ;
  assign n32107 = n32105 | n32106 ;
  assign n32108 = n32104 | n32107 ;
  assign n32109 = n20689 | n32108 ;
  assign n32110 = n1062 | n32108 ;
  assign n32111 = ( n32103 & n32109 ) | ( n32103 & n32110 ) | ( n32109 & n32110 ) ;
  assign n32112 = n32102 & n32111 ;
  assign n32113 = n32102 & ~n32112 ;
  assign n32114 = ~n32102 & n32111 ;
  assign n32115 = n32113 | n32114 ;
  assign n32116 = ( ~n30919 & n32088 ) | ( ~n30919 & n32089 ) | ( n32088 & n32089 ) ;
  assign n32117 = ( ~n1062 & n32088 ) | ( ~n1062 & n32089 ) | ( n32088 & n32089 ) ;
  assign n32118 = ( ~n19640 & n32116 ) | ( ~n19640 & n32117 ) | ( n32116 & n32117 ) ;
  assign n32119 = n32087 | n32095 ;
  assign n32120 = n32089 | n32091 ;
  assign n32121 = ( ~n30919 & n32119 ) | ( ~n30919 & n32120 ) | ( n32119 & n32120 ) ;
  assign n32122 = ( ~n1062 & n32119 ) | ( ~n1062 & n32120 ) | ( n32119 & n32120 ) ;
  assign n32123 = ( ~n19640 & n32121 ) | ( ~n19640 & n32122 ) | ( n32121 & n32122 ) ;
  assign n32124 = ~n32118 & n32123 ;
  assign n32125 = ~n32090 & n32099 ;
  assign n32126 = n32124 | n32125 ;
  assign n32127 = n1057 & ~n20630 ;
  assign n32128 = n1060 & n19494 ;
  assign n32129 = n1065 & n19631 ;
  assign n32130 = n32128 | n32129 ;
  assign n32131 = n32127 | n32130 ;
  assign n32132 = n1062 | n32127 ;
  assign n32133 = n32130 | n32132 ;
  assign n32134 = ( ~n20709 & n32131 ) | ( ~n20709 & n32133 ) | ( n32131 & n32133 ) ;
  assign n32135 = n32126 & n32134 ;
  assign n32136 = n32126 | n32134 ;
  assign n32137 = ~n32135 & n32136 ;
  assign n32138 = n1829 & ~n21563 ;
  assign n32139 = n1826 & ~n20618 ;
  assign n32140 = n1823 & n20609 ;
  assign n32141 = n32139 | n32140 ;
  assign n32142 = n32138 | n32141 ;
  assign n32143 = n21570 & ~n32142 ;
  assign n32144 = ( n22270 & n32142 ) | ( n22270 & ~n32143 ) | ( n32142 & ~n32143 ) ;
  assign n32145 = n22304 | n32144 ;
  assign n32146 = n1821 | n32138 ;
  assign n32147 = n32141 | n32146 ;
  assign n32148 = n32145 & n32147 ;
  assign n32149 = ~x29 & n32147 ;
  assign n32150 = n32145 & n32149 ;
  assign n32151 = x29 | n32149 ;
  assign n32152 = ( x29 & n32145 ) | ( x29 & n32151 ) | ( n32145 & n32151 ) ;
  assign n32153 = ( ~n32148 & n32150 ) | ( ~n32148 & n32152 ) | ( n32150 & n32152 ) ;
  assign n32154 = n32135 | n32153 ;
  assign n32155 = ( n32135 & n32137 ) | ( n32135 & n32154 ) | ( n32137 & n32154 ) ;
  assign n32156 = n32115 | n32155 ;
  assign n32157 = n32115 & n32155 ;
  assign n32158 = n32156 & ~n32157 ;
  assign n32159 = n1829 & ~n21517 ;
  assign n32160 = n1826 & n20609 ;
  assign n32161 = n1823 & ~n21563 ;
  assign n32162 = n32160 | n32161 ;
  assign n32163 = n32159 | n32162 ;
  assign n32164 = n1821 | n32159 ;
  assign n32165 = n32162 | n32164 ;
  assign n32166 = ( ~n22283 & n32163 ) | ( ~n22283 & n32165 ) | ( n32163 & n32165 ) ;
  assign n32167 = n32163 & n32165 ;
  assign n32168 = ( ~n22271 & n32166 ) | ( ~n22271 & n32167 ) | ( n32166 & n32167 ) ;
  assign n32169 = ~x29 & n32168 ;
  assign n32170 = x29 | n32168 ;
  assign n32171 = ( ~n32168 & n32169 ) | ( ~n32168 & n32170 ) | ( n32169 & n32170 ) ;
  assign n32172 = ~n32158 & n32171 ;
  assign n32173 = n32157 | n32171 ;
  assign n32174 = n32156 & ~n32173 ;
  assign n32175 = n32172 | n32174 ;
  assign n32176 = n2315 & ~n23240 ;
  assign n32177 = n2312 & ~n21551 ;
  assign n32178 = n2308 & n23227 ;
  assign n32179 = ( n2308 & n23217 ) | ( n2308 & n32178 ) | ( n23217 & n32178 ) ;
  assign n32180 = n32177 | n32179 ;
  assign n32181 = n32176 | n32180 ;
  assign n32182 = n2306 | n32176 ;
  assign n32183 = n32180 | n32182 ;
  assign n32184 = ( n23260 & n32181 ) | ( n23260 & n32183 ) | ( n32181 & n32183 ) ;
  assign n32185 = x26 & n32183 ;
  assign n32186 = x26 & n32181 ;
  assign n32187 = ( n23260 & n32185 ) | ( n23260 & n32186 ) | ( n32185 & n32186 ) ;
  assign n32188 = x26 & ~n32186 ;
  assign n32189 = x26 & ~n32185 ;
  assign n32190 = ( ~n23260 & n32188 ) | ( ~n23260 & n32189 ) | ( n32188 & n32189 ) ;
  assign n32191 = ( n32184 & ~n32187 ) | ( n32184 & n32190 ) | ( ~n32187 & n32190 ) ;
  assign n32192 = n32137 & n32153 ;
  assign n32193 = n32137 | n32153 ;
  assign n32194 = ~n32192 & n32193 ;
  assign n32195 = n30989 | n31005 ;
  assign n32196 = ( n30989 & n30991 ) | ( n30989 & n32195 ) | ( n30991 & n32195 ) ;
  assign n32197 = n32194 & n32196 ;
  assign n32198 = n32194 | n32196 ;
  assign n32199 = ~n32197 & n32198 ;
  assign n32200 = n2312 & ~n21517 ;
  assign n32201 = n2308 & ~n21551 ;
  assign n32202 = n32200 | n32201 ;
  assign n32203 = n2315 & n23227 ;
  assign n32204 = ( n2315 & n23217 ) | ( n2315 & n32203 ) | ( n23217 & n32203 ) ;
  assign n32205 = n32202 | n32204 ;
  assign n32206 = n2306 & n23299 ;
  assign n32207 = n2306 & n23298 ;
  assign n32208 = ( n21584 & n32206 ) | ( n21584 & n32207 ) | ( n32206 & n32207 ) ;
  assign n32209 = n32205 | n32208 ;
  assign n32210 = n2306 | n32205 ;
  assign n32211 = ( n23289 & n32209 ) | ( n23289 & n32210 ) | ( n32209 & n32210 ) ;
  assign n32212 = x26 | n32211 ;
  assign n32213 = ~x26 & n32211 ;
  assign n32214 = ( ~n32211 & n32212 ) | ( ~n32211 & n32213 ) | ( n32212 & n32213 ) ;
  assign n32215 = n32197 | n32214 ;
  assign n32216 = ( n32197 & n32199 ) | ( n32197 & n32215 ) | ( n32199 & n32215 ) ;
  assign n32217 = ( n32175 & n32191 ) | ( n32175 & ~n32216 ) | ( n32191 & ~n32216 ) ;
  assign n32218 = ( ~n32191 & n32216 ) | ( ~n32191 & n32217 ) | ( n32216 & n32217 ) ;
  assign n32219 = ( ~n32175 & n32217 ) | ( ~n32175 & n32218 ) | ( n32217 & n32218 ) ;
  assign n32220 = ~n23234 & n32066 ;
  assign n32221 = n2925 | n32220 ;
  assign n32222 = ~n23235 & n32066 ;
  assign n32223 = n2925 | n32222 ;
  assign n32224 = ( ~n15882 & n32221 ) | ( ~n15882 & n32223 ) | ( n32221 & n32223 ) ;
  assign n32225 = n2936 | n32224 ;
  assign n32226 = ( ~n15882 & n32220 ) | ( ~n15882 & n32222 ) | ( n32220 & n32222 ) ;
  assign n32227 = n2936 | n32226 ;
  assign n32228 = ( ~n23240 & n32225 ) | ( ~n23240 & n32227 ) | ( n32225 & n32227 ) ;
  assign n32229 = ( ~n23240 & n32224 ) | ( ~n23240 & n32226 ) | ( n32224 & n32226 ) ;
  assign n32230 = n24135 & ~n32229 ;
  assign n32231 = n23240 & ~n32229 ;
  assign n32232 = ( n23575 & n32230 ) | ( n23575 & n32231 ) | ( n32230 & n32231 ) ;
  assign n32233 = ( n23577 & n32230 ) | ( n23577 & n32231 ) | ( n32230 & n32231 ) ;
  assign n32234 = ( ~n21554 & n32232 ) | ( ~n21554 & n32233 ) | ( n32232 & n32233 ) ;
  assign n32235 = n32228 & ~n32234 ;
  assign n32236 = x23 & ~n32235 ;
  assign n32237 = n32232 | n32233 ;
  assign n32238 = n32228 & ~n32237 ;
  assign n32239 = x23 & ~n32238 ;
  assign n32240 = ( n21584 & n32236 ) | ( n21584 & n32239 ) | ( n32236 & n32239 ) ;
  assign n32241 = ~x23 & n32235 ;
  assign n32242 = ~x23 & n32238 ;
  assign n32243 = ( ~n21584 & n32241 ) | ( ~n21584 & n32242 ) | ( n32241 & n32242 ) ;
  assign n32244 = n32240 | n32243 ;
  assign n32245 = n31053 | n31070 ;
  assign n32246 = ( n31053 & n31055 ) | ( n31053 & n32245 ) | ( n31055 & n32245 ) ;
  assign n32247 = n32244 & n32246 ;
  assign n32248 = n32244 | n32246 ;
  assign n32249 = ~n32247 & n32248 ;
  assign n32250 = n32199 & ~n32214 ;
  assign n32251 = n32199 | n32214 ;
  assign n32252 = ( ~n32199 & n32250 ) | ( ~n32199 & n32251 ) | ( n32250 & n32251 ) ;
  assign n32253 = n32247 | n32252 ;
  assign n32254 = ( n32247 & n32249 ) | ( n32247 & n32253 ) | ( n32249 & n32253 ) ;
  assign n32255 = n32219 & n32254 ;
  assign n32256 = n32219 | n32254 ;
  assign n32257 = ~n32255 & n32256 ;
  assign n32258 = n32249 & ~n32252 ;
  assign n32259 = n32249 | n32252 ;
  assign n32260 = ( ~n32249 & n32258 ) | ( ~n32249 & n32259 ) | ( n32258 & n32259 ) ;
  assign n32261 = n31135 | n31155 ;
  assign n32262 = ( n31135 & n31137 ) | ( n31135 & n32261 ) | ( n31137 & n32261 ) ;
  assign n32263 = n32260 & n32262 ;
  assign n32264 = n32260 | n32262 ;
  assign n32265 = ~n32263 & n32264 ;
  assign n32266 = n31209 | n31280 ;
  assign n32267 = n32265 & n32266 ;
  assign n32268 = n32263 | n32267 ;
  assign n32269 = n32257 & n32268 ;
  assign n32270 = n31209 | n31284 ;
  assign n32271 = n32265 & n32270 ;
  assign n32272 = n32263 | n32271 ;
  assign n32273 = n32257 & n32272 ;
  assign n32274 = ( n30169 & n32269 ) | ( n30169 & n32273 ) | ( n32269 & n32273 ) ;
  assign n32275 = n31209 | n31212 ;
  assign n32276 = n32265 & n32275 ;
  assign n32277 = n32263 | n32276 ;
  assign n32278 = n32257 & n32277 ;
  assign n32279 = n31209 & n32265 ;
  assign n32280 = n32263 | n32279 ;
  assign n32281 = n32257 & n32280 ;
  assign n32282 = ( n31274 & n32278 ) | ( n31274 & n32281 ) | ( n32278 & n32281 ) ;
  assign n32283 = ( n28465 & n32274 ) | ( n28465 & n32282 ) | ( n32274 & n32282 ) ;
  assign n32284 = n32274 & n32282 ;
  assign n32285 = ( n28489 & n32283 ) | ( n28489 & n32284 ) | ( n32283 & n32284 ) ;
  assign n32286 = ( n30169 & n32268 ) | ( n30169 & n32272 ) | ( n32268 & n32272 ) ;
  assign n32287 = ( n31274 & n32277 ) | ( n31274 & n32280 ) | ( n32277 & n32280 ) ;
  assign n32288 = n32286 & n32287 ;
  assign n32289 = n32257 | n32288 ;
  assign n32290 = ( n28465 & n32286 ) | ( n28465 & n32287 ) | ( n32286 & n32287 ) ;
  assign n32291 = n32257 | n32290 ;
  assign n32292 = ( n28489 & n32289 ) | ( n28489 & n32291 ) | ( n32289 & n32291 ) ;
  assign n32293 = ~n32285 & n32292 ;
  assign n32294 = ( n30169 & n32267 ) | ( n30169 & n32271 ) | ( n32267 & n32271 ) ;
  assign n32295 = ( n31274 & n32276 ) | ( n31274 & n32279 ) | ( n32276 & n32279 ) ;
  assign n32296 = ( n28465 & n32294 ) | ( n28465 & n32295 ) | ( n32294 & n32295 ) ;
  assign n32297 = n32294 & n32295 ;
  assign n32298 = ( n28489 & n32296 ) | ( n28489 & n32297 ) | ( n32296 & n32297 ) ;
  assign n32299 = ( n30169 & n32266 ) | ( n30169 & n32270 ) | ( n32266 & n32270 ) ;
  assign n32300 = ( n31209 & n31274 ) | ( n31209 & n32275 ) | ( n31274 & n32275 ) ;
  assign n32301 = n32299 & n32300 ;
  assign n32302 = n32265 | n32301 ;
  assign n32303 = ( n28465 & n32299 ) | ( n28465 & n32300 ) | ( n32299 & n32300 ) ;
  assign n32304 = n32265 | n32303 ;
  assign n32305 = ( n28489 & n32302 ) | ( n28489 & n32304 ) | ( n32302 & n32304 ) ;
  assign n32306 = ~n32298 & n32305 ;
  assign n32307 = n32293 & n32306 ;
  assign n32308 = n31295 & n32306 ;
  assign n32309 = n31295 | n32306 ;
  assign n32310 = ~n32308 & n32309 ;
  assign n32311 = n31330 | n32308 ;
  assign n32312 = ( n32308 & n32310 ) | ( n32308 & n32311 ) | ( n32310 & n32311 ) ;
  assign n32313 = n32293 | n32306 ;
  assign n32314 = ~n32307 & n32313 ;
  assign n32315 = n32307 | n32314 ;
  assign n32316 = ( n32307 & n32312 ) | ( n32307 & n32315 ) | ( n32312 & n32315 ) ;
  assign n32317 = n32308 & n32313 ;
  assign n32318 = ( n32310 & n32313 ) | ( n32310 & n32317 ) | ( n32313 & n32317 ) ;
  assign n32319 = n32307 | n32318 ;
  assign n32320 = ( ~n31343 & n32316 ) | ( ~n31343 & n32319 ) | ( n32316 & n32319 ) ;
  assign n32321 = ( ~n31348 & n32316 ) | ( ~n31348 & n32319 ) | ( n32316 & n32319 ) ;
  assign n32322 = ( n30232 & n32320 ) | ( n30232 & n32321 ) | ( n32320 & n32321 ) ;
  assign n32323 = n32191 & n32216 ;
  assign n32324 = n32216 & ~n32323 ;
  assign n32325 = n32191 & ~n32216 ;
  assign n32326 = n32175 & ~n32325 ;
  assign n32327 = ~n32324 & n32326 ;
  assign n32328 = ( n32175 & n32323 ) | ( n32175 & ~n32327 ) | ( n32323 & ~n32327 ) ;
  assign n32329 = n4410 | n20360 ;
  assign n32330 = n8004 | n32329 ;
  assign n32331 = n6839 | n32330 ;
  assign n32332 = n6821 | n32331 ;
  assign n32333 = n7895 | n7896 ;
  assign n32334 = n6868 & ~n32333 ;
  assign n32335 = n721 | n1146 ;
  assign n32336 = n1387 | n32335 ;
  assign n32337 = n96 | n623 ;
  assign n32338 = n257 | n434 ;
  assign n32339 = n1398 | n32338 ;
  assign n32340 = n32337 | n32339 ;
  assign n32341 = n32336 | n32340 ;
  assign n32342 = n1034 | n2651 ;
  assign n32343 = n3425 | n32342 ;
  assign n32344 = n228 | n32343 ;
  assign n32345 = n32341 | n32344 ;
  assign n32346 = n32334 & ~n32345 ;
  assign n32347 = ~n32332 & n32346 ;
  assign n32348 = ~n4174 & n32347 ;
  assign n32349 = ( n32064 & n32065 ) | ( n32064 & n32348 ) | ( n32065 & n32348 ) ;
  assign n32350 = n32064 & n32348 ;
  assign n32351 = ( ~n32083 & n32349 ) | ( ~n32083 & n32350 ) | ( n32349 & n32350 ) ;
  assign n32352 = n32064 | n32065 ;
  assign n32353 = n32348 | n32352 ;
  assign n32354 = n32064 | n32348 ;
  assign n32355 = ( ~n32083 & n32353 ) | ( ~n32083 & n32354 ) | ( n32353 & n32354 ) ;
  assign n32356 = ~n32351 & n32355 ;
  assign n32357 = n1057 & n20609 ;
  assign n32358 = n1065 & ~n20618 ;
  assign n32359 = n1060 & ~n20630 ;
  assign n32360 = n32358 | n32359 ;
  assign n32361 = n32357 | n32360 ;
  assign n32362 = n1062 | n32357 ;
  assign n32363 = n32360 | n32362 ;
  assign n32364 = ( n20659 & n32361 ) | ( n20659 & n32363 ) | ( n32361 & n32363 ) ;
  assign n32365 = n32361 & n32363 ;
  assign n32366 = ( ~n20649 & n32364 ) | ( ~n20649 & n32365 ) | ( n32364 & n32365 ) ;
  assign n32367 = n32356 | n32366 ;
  assign n32368 = n32356 & n32363 ;
  assign n32369 = n32356 & n32361 ;
  assign n32370 = ( n20659 & n32368 ) | ( n20659 & n32369 ) | ( n32368 & n32369 ) ;
  assign n32371 = n32368 & n32369 ;
  assign n32372 = ( ~n20649 & n32370 ) | ( ~n20649 & n32371 ) | ( n32370 & n32371 ) ;
  assign n32373 = n32367 & ~n32372 ;
  assign n32374 = n32100 & ~n32373 ;
  assign n32375 = ~n32112 & n32374 ;
  assign n32376 = ( ~n32100 & n32112 ) | ( ~n32100 & n32373 ) | ( n32112 & n32373 ) ;
  assign n32377 = n32375 | n32376 ;
  assign n32378 = n1829 & ~n21551 ;
  assign n32379 = n1826 & ~n21563 ;
  assign n32380 = n1823 & ~n21517 ;
  assign n32381 = n32379 | n32380 ;
  assign n32382 = n32378 | n32381 ;
  assign n32383 = n1821 | n32378 ;
  assign n32384 = n32381 | n32383 ;
  assign n32385 = ( ~n21587 & n32382 ) | ( ~n21587 & n32384 ) | ( n32382 & n32384 ) ;
  assign n32386 = ~x29 & n32384 ;
  assign n32387 = ~x29 & n32382 ;
  assign n32388 = ( ~n21587 & n32386 ) | ( ~n21587 & n32387 ) | ( n32386 & n32387 ) ;
  assign n32389 = x29 | n32387 ;
  assign n32390 = x29 | n32386 ;
  assign n32391 = ( ~n21587 & n32389 ) | ( ~n21587 & n32390 ) | ( n32389 & n32390 ) ;
  assign n32392 = ( ~n32385 & n32388 ) | ( ~n32385 & n32391 ) | ( n32388 & n32391 ) ;
  assign n32393 = ~n32377 & n32392 ;
  assign n32394 = n32377 & ~n32392 ;
  assign n32395 = n32393 | n32394 ;
  assign n32396 = ( n32157 & n32158 ) | ( n32157 & n32173 ) | ( n32158 & n32173 ) ;
  assign n32397 = ~n32395 & n32396 ;
  assign n32398 = n32395 & ~n32396 ;
  assign n32399 = n32397 | n32398 ;
  assign n32400 = n2308 & ~n23240 ;
  assign n32401 = n2312 & n23227 ;
  assign n32402 = ( n2312 & n23217 ) | ( n2312 & n32401 ) | ( n23217 & n32401 ) ;
  assign n32403 = n32400 | n32402 ;
  assign n32404 = n2315 & ~n23234 ;
  assign n32405 = n2315 & ~n23235 ;
  assign n32406 = ( ~n15882 & n32404 ) | ( ~n15882 & n32405 ) | ( n32404 & n32405 ) ;
  assign n32407 = n32403 | n32406 ;
  assign n32408 = n2306 | n32406 ;
  assign n32409 = n32403 | n32408 ;
  assign n32410 = ( ~n23587 & n32407 ) | ( ~n23587 & n32409 ) | ( n32407 & n32409 ) ;
  assign n32411 = ~x26 & n32409 ;
  assign n32412 = ~x26 & n32407 ;
  assign n32413 = ( ~n23587 & n32411 ) | ( ~n23587 & n32412 ) | ( n32411 & n32412 ) ;
  assign n32414 = x26 | n32412 ;
  assign n32415 = x26 | n32411 ;
  assign n32416 = ( ~n23587 & n32414 ) | ( ~n23587 & n32415 ) | ( n32414 & n32415 ) ;
  assign n32417 = ( ~n32410 & n32413 ) | ( ~n32410 & n32416 ) | ( n32413 & n32416 ) ;
  assign n32418 = n32399 | n32417 ;
  assign n32419 = n32399 & ~n32417 ;
  assign n32420 = ( ~n32399 & n32418 ) | ( ~n32399 & n32419 ) | ( n32418 & n32419 ) ;
  assign n32421 = n32328 & ~n32420 ;
  assign n32422 = n32328 & ~n32421 ;
  assign n32423 = n32328 | n32420 ;
  assign n32424 = ~n32422 & n32423 ;
  assign n32425 = n32255 & ~n32424 ;
  assign n32426 = ( n32274 & ~n32424 ) | ( n32274 & n32425 ) | ( ~n32424 & n32425 ) ;
  assign n32427 = n32255 | n32278 ;
  assign n32428 = ~n32424 & n32427 ;
  assign n32429 = n32255 | n32281 ;
  assign n32430 = ~n32424 & n32429 ;
  assign n32431 = ( n31274 & n32428 ) | ( n31274 & n32430 ) | ( n32428 & n32430 ) ;
  assign n32432 = ( n28465 & n32426 ) | ( n28465 & n32431 ) | ( n32426 & n32431 ) ;
  assign n32433 = n32426 & n32431 ;
  assign n32434 = ( n28489 & n32432 ) | ( n28489 & n32433 ) | ( n32432 & n32433 ) ;
  assign n32435 = n32255 | n32274 ;
  assign n32436 = ( n31274 & n32427 ) | ( n31274 & n32429 ) | ( n32427 & n32429 ) ;
  assign n32437 = n32435 & n32436 ;
  assign n32438 = n32424 & ~n32437 ;
  assign n32439 = ( n28465 & n32435 ) | ( n28465 & n32436 ) | ( n32435 & n32436 ) ;
  assign n32440 = n32424 & ~n32439 ;
  assign n32441 = ( ~n28489 & n32438 ) | ( ~n28489 & n32440 ) | ( n32438 & n32440 ) ;
  assign n32442 = n32434 | n32441 ;
  assign n32443 = n32293 & ~n32442 ;
  assign n32444 = ~n32293 & n32442 ;
  assign n32445 = n32443 | n32444 ;
  assign n32446 = n32316 & ~n32445 ;
  assign n32447 = n32307 & ~n32444 ;
  assign n32448 = ~n32443 & n32447 ;
  assign n32449 = ( n32318 & ~n32445 ) | ( n32318 & n32448 ) | ( ~n32445 & n32448 ) ;
  assign n32450 = ( ~n31343 & n32446 ) | ( ~n31343 & n32449 ) | ( n32446 & n32449 ) ;
  assign n32451 = ( ~n31348 & n32446 ) | ( ~n31348 & n32449 ) | ( n32446 & n32449 ) ;
  assign n32452 = ( n30232 & n32450 ) | ( n30232 & n32451 ) | ( n32450 & n32451 ) ;
  assign n32453 = n32322 & ~n32452 ;
  assign n32454 = n32443 | n32450 ;
  assign n32455 = n32443 | n32451 ;
  assign n32456 = ( n30232 & n32454 ) | ( n30232 & n32455 ) | ( n32454 & n32455 ) ;
  assign n32457 = n32444 | n32456 ;
  assign n32458 = ~n32453 & n32457 ;
  assign n32459 = n8122 & ~n32442 ;
  assign n32460 = n8115 & n32306 ;
  assign n32461 = n8118 & n32293 ;
  assign n32462 = n32460 | n32461 ;
  assign n32463 = n32459 | n32462 ;
  assign n32464 = n8125 | n32459 ;
  assign n32465 = n32462 | n32464 ;
  assign n32466 = ( ~n32458 & n32463 ) | ( ~n32458 & n32465 ) | ( n32463 & n32465 ) ;
  assign n32467 = ~x5 & n32465 ;
  assign n32468 = ~x5 & n32463 ;
  assign n32469 = ( ~n32458 & n32467 ) | ( ~n32458 & n32468 ) | ( n32467 & n32468 ) ;
  assign n32470 = x5 | n32468 ;
  assign n32471 = x5 | n32467 ;
  assign n32472 = ( ~n32458 & n32470 ) | ( ~n32458 & n32471 ) | ( n32470 & n32471 ) ;
  assign n32473 = ( ~n32466 & n32469 ) | ( ~n32466 & n32472 ) | ( n32469 & n32472 ) ;
  assign n32474 = ~n32027 & n32473 ;
  assign n32475 = n32027 & ~n32473 ;
  assign n32476 = n32474 | n32475 ;
  assign n32477 = n31397 & n32022 ;
  assign n32478 = n31397 | n32022 ;
  assign n32479 = ~n32477 & n32478 ;
  assign n32480 = n8122 & n32293 ;
  assign n32481 = n8115 & n31295 ;
  assign n32482 = n8118 & n32306 ;
  assign n32483 = n32481 | n32482 ;
  assign n32484 = n32480 | n32483 ;
  assign n32485 = n32308 | n32310 ;
  assign n32486 = ( ~n31343 & n32312 ) | ( ~n31343 & n32485 ) | ( n32312 & n32485 ) ;
  assign n32487 = ( ~n31348 & n32312 ) | ( ~n31348 & n32485 ) | ( n32312 & n32485 ) ;
  assign n32488 = ( n30232 & n32486 ) | ( n30232 & n32487 ) | ( n32486 & n32487 ) ;
  assign n32489 = ~n32307 & n32318 ;
  assign n32490 = n32312 & n32314 ;
  assign n32491 = ( ~n31343 & n32489 ) | ( ~n31343 & n32490 ) | ( n32489 & n32490 ) ;
  assign n32492 = ( ~n31348 & n32489 ) | ( ~n31348 & n32490 ) | ( n32489 & n32490 ) ;
  assign n32493 = ( n30232 & n32491 ) | ( n30232 & n32492 ) | ( n32491 & n32492 ) ;
  assign n32494 = n32488 & ~n32493 ;
  assign n32495 = n32313 & ~n32320 ;
  assign n32496 = n32313 & ~n32321 ;
  assign n32497 = ( ~n30232 & n32495 ) | ( ~n30232 & n32496 ) | ( n32495 & n32496 ) ;
  assign n32498 = n8125 & n32497 ;
  assign n32499 = ( n8125 & n32494 ) | ( n8125 & n32498 ) | ( n32494 & n32498 ) ;
  assign n32500 = n32484 | n32499 ;
  assign n32501 = x5 | n32484 ;
  assign n32502 = n32499 | n32501 ;
  assign n32503 = ~x5 & n32501 ;
  assign n32504 = ( ~x5 & n32499 ) | ( ~x5 & n32503 ) | ( n32499 & n32503 ) ;
  assign n32505 = ( ~n32500 & n32502 ) | ( ~n32500 & n32504 ) | ( n32502 & n32504 ) ;
  assign n32506 = ~n32479 & n32505 ;
  assign n32507 = n32479 & ~n32505 ;
  assign n32508 = n32506 | n32507 ;
  assign n32509 = ~n31424 & n32020 ;
  assign n32510 = n31424 & ~n32020 ;
  assign n32511 = n32509 | n32510 ;
  assign n32512 = n8122 & n32306 ;
  assign n32513 = n8115 & ~n31323 ;
  assign n32514 = n8118 & n31295 ;
  assign n32515 = n32513 | n32514 ;
  assign n32516 = n32512 | n32515 ;
  assign n32517 = n31330 & n32310 ;
  assign n32518 = ( ~n31343 & n32310 ) | ( ~n31343 & n32517 ) | ( n32310 & n32517 ) ;
  assign n32519 = ( ~n31348 & n32310 ) | ( ~n31348 & n32517 ) | ( n32310 & n32517 ) ;
  assign n32520 = ( n30232 & n32518 ) | ( n30232 & n32519 ) | ( n32518 & n32519 ) ;
  assign n32521 = n31330 | n32310 ;
  assign n32522 = n31343 & ~n32521 ;
  assign n32523 = n31348 & ~n32521 ;
  assign n32524 = ( ~n30232 & n32522 ) | ( ~n30232 & n32523 ) | ( n32522 & n32523 ) ;
  assign n32525 = n32520 | n32524 ;
  assign n32526 = n8125 | n32512 ;
  assign n32527 = n32515 | n32526 ;
  assign n32528 = ( n32516 & ~n32525 ) | ( n32516 & n32527 ) | ( ~n32525 & n32527 ) ;
  assign n32529 = ~x5 & n32527 ;
  assign n32530 = ~x5 & n32516 ;
  assign n32531 = ( ~n32525 & n32529 ) | ( ~n32525 & n32530 ) | ( n32529 & n32530 ) ;
  assign n32532 = x5 | n32530 ;
  assign n32533 = x5 | n32529 ;
  assign n32534 = ( ~n32525 & n32532 ) | ( ~n32525 & n32533 ) | ( n32532 & n32533 ) ;
  assign n32535 = ( ~n32528 & n32531 ) | ( ~n32528 & n32534 ) | ( n32531 & n32534 ) ;
  assign n32536 = n32511 & n32535 ;
  assign n32537 = n32511 | n32535 ;
  assign n32538 = ~n32536 & n32537 ;
  assign n32539 = n31446 & n32018 ;
  assign n32540 = n31446 | n32018 ;
  assign n32541 = ~n32539 & n32540 ;
  assign n32542 = n8122 & n31295 ;
  assign n32543 = n8115 & ~n31309 ;
  assign n32544 = n8118 & ~n31323 ;
  assign n32545 = n32543 | n32544 ;
  assign n32546 = n32542 | n32545 ;
  assign n32547 = n8125 | n32542 ;
  assign n32548 = n32545 | n32547 ;
  assign n32549 = ( n31355 & n32546 ) | ( n31355 & n32548 ) | ( n32546 & n32548 ) ;
  assign n32550 = x5 & n32548 ;
  assign n32551 = x5 & n32546 ;
  assign n32552 = ( n31355 & n32550 ) | ( n31355 & n32551 ) | ( n32550 & n32551 ) ;
  assign n32553 = x5 & ~n32551 ;
  assign n32554 = x5 & ~n32550 ;
  assign n32555 = ( ~n31355 & n32553 ) | ( ~n31355 & n32554 ) | ( n32553 & n32554 ) ;
  assign n32556 = ( n32549 & ~n32552 ) | ( n32549 & n32555 ) | ( ~n32552 & n32555 ) ;
  assign n32557 = ~n32541 & n32556 ;
  assign n32558 = n31468 & n32016 ;
  assign n32559 = n31468 | n32016 ;
  assign n32560 = ~n32558 & n32559 ;
  assign n32561 = n8122 & ~n31323 ;
  assign n32562 = n8115 & ~n30186 ;
  assign n32563 = n8118 & ~n31309 ;
  assign n32564 = n32562 | n32563 ;
  assign n32565 = n32561 | n32564 ;
  assign n32566 = n8125 & n31384 ;
  assign n32567 = n8125 & n31386 ;
  assign n32568 = ( ~n30232 & n32566 ) | ( ~n30232 & n32567 ) | ( n32566 & n32567 ) ;
  assign n32569 = n32565 | n32568 ;
  assign n32570 = n8125 | n32565 ;
  assign n32571 = ( ~n31376 & n32569 ) | ( ~n31376 & n32570 ) | ( n32569 & n32570 ) ;
  assign n32572 = x5 | n32571 ;
  assign n32573 = ~x5 & n32571 ;
  assign n32574 = ( ~n32571 & n32572 ) | ( ~n32571 & n32573 ) | ( n32572 & n32573 ) ;
  assign n32575 = ~n32560 & n32574 ;
  assign n32576 = n32560 & ~n32574 ;
  assign n32577 = n32575 | n32576 ;
  assign n32578 = n32012 & n32014 ;
  assign n32579 = n32012 | n32014 ;
  assign n32580 = ~n32578 & n32579 ;
  assign n32582 = n8115 & n30212 ;
  assign n32583 = n8118 & ~n30186 ;
  assign n32584 = n32582 | n32583 ;
  assign n32581 = n8122 & ~n31309 ;
  assign n32586 = n8125 | n32581 ;
  assign n32587 = n32584 | n32586 ;
  assign n32585 = n32581 | n32584 ;
  assign n32588 = n32585 & n32587 ;
  assign n32589 = ( n31404 & n32587 ) | ( n31404 & n32588 ) | ( n32587 & n32588 ) ;
  assign n32590 = x5 & n32588 ;
  assign n32591 = x5 & n32587 ;
  assign n32592 = ( n31404 & n32590 ) | ( n31404 & n32591 ) | ( n32590 & n32591 ) ;
  assign n32593 = x5 & ~n32590 ;
  assign n32594 = x5 & ~n32591 ;
  assign n32595 = ( ~n31404 & n32593 ) | ( ~n31404 & n32594 ) | ( n32593 & n32594 ) ;
  assign n32596 = ( n32589 & ~n32592 ) | ( n32589 & n32595 ) | ( ~n32592 & n32595 ) ;
  assign n32597 = n32580 & n32596 ;
  assign n32598 = n31508 & n32010 ;
  assign n32599 = n31508 | n32010 ;
  assign n32600 = ~n32598 & n32599 ;
  assign n32602 = n8115 & ~n30199 ;
  assign n32603 = n8118 & n30212 ;
  assign n32604 = n32602 | n32603 ;
  assign n32601 = n8122 & ~n30186 ;
  assign n32606 = n8125 | n32601 ;
  assign n32607 = n32604 | n32606 ;
  assign n32605 = n32601 | n32604 ;
  assign n32608 = n32605 & n32607 ;
  assign n32609 = ( ~n30241 & n32607 ) | ( ~n30241 & n32608 ) | ( n32607 & n32608 ) ;
  assign n32610 = ~x5 & n32608 ;
  assign n32611 = ~x5 & n32607 ;
  assign n32612 = ( ~n30241 & n32610 ) | ( ~n30241 & n32611 ) | ( n32610 & n32611 ) ;
  assign n32613 = x5 | n32610 ;
  assign n32614 = x5 | n32611 ;
  assign n32615 = ( ~n30241 & n32613 ) | ( ~n30241 & n32614 ) | ( n32613 & n32614 ) ;
  assign n32616 = ( ~n32609 & n32612 ) | ( ~n32609 & n32615 ) | ( n32612 & n32615 ) ;
  assign n32617 = n32600 & n32616 ;
  assign n32618 = n32600 & ~n32617 ;
  assign n32619 = ~n32600 & n32616 ;
  assign n32620 = n32618 | n32619 ;
  assign n32621 = n32001 | n32007 ;
  assign n32622 = n32005 | n32621 ;
  assign n32623 = ~n32009 & n32622 ;
  assign n32624 = n8122 & n30212 ;
  assign n32625 = n8115 & n29620 ;
  assign n32626 = n8118 & ~n30199 ;
  assign n32627 = n32625 | n32626 ;
  assign n32628 = n32624 | n32627 ;
  assign n32629 = n8125 & ~n30266 ;
  assign n32630 = ( n8125 & n30276 ) | ( n8125 & n32629 ) | ( n30276 & n32629 ) ;
  assign n32631 = n32628 | n32630 ;
  assign n32632 = x5 | n32628 ;
  assign n32633 = n32630 | n32632 ;
  assign n32634 = ~x5 & n32632 ;
  assign n32635 = ( ~x5 & n32630 ) | ( ~x5 & n32634 ) | ( n32630 & n32634 ) ;
  assign n32636 = ( ~n32631 & n32633 ) | ( ~n32631 & n32635 ) | ( n32633 & n32635 ) ;
  assign n32637 = n32623 & n32636 ;
  assign n32638 = n31980 & ~n32005 ;
  assign n32639 = n32004 & ~n32005 ;
  assign n32640 = n32638 | n32639 ;
  assign n32641 = n8122 & ~n30199 ;
  assign n32642 = n8115 & ~n28714 ;
  assign n32643 = n8118 & n29620 ;
  assign n32644 = n32642 | n32643 ;
  assign n32645 = n32641 | n32644 ;
  assign n32646 = n8125 | n32641 ;
  assign n32647 = n32644 | n32646 ;
  assign n32648 = ( ~n30299 & n32645 ) | ( ~n30299 & n32647 ) | ( n32645 & n32647 ) ;
  assign n32649 = ~x5 & n32647 ;
  assign n32650 = ~x5 & n32645 ;
  assign n32651 = ( ~n30299 & n32649 ) | ( ~n30299 & n32650 ) | ( n32649 & n32650 ) ;
  assign n32652 = x5 | n32650 ;
  assign n32653 = x5 | n32649 ;
  assign n32654 = ( ~n30299 & n32652 ) | ( ~n30299 & n32653 ) | ( n32652 & n32653 ) ;
  assign n32655 = ( ~n32648 & n32651 ) | ( ~n32648 & n32654 ) | ( n32651 & n32654 ) ;
  assign n32656 = n32640 & n32655 ;
  assign n32657 = n32640 & ~n32656 ;
  assign n32658 = ~n32640 & n32655 ;
  assign n32659 = n32657 | n32658 ;
  assign n32660 = n31975 & ~n31979 ;
  assign n32661 = n31978 & ~n31979 ;
  assign n32662 = n32660 | n32661 ;
  assign n32663 = n8122 & n29620 ;
  assign n32664 = n8115 & n28492 ;
  assign n32665 = n8118 & ~n28714 ;
  assign n32666 = n32664 | n32665 ;
  assign n32667 = n32663 | n32666 ;
  assign n32668 = n8125 | n32663 ;
  assign n32669 = n32666 | n32668 ;
  assign n32670 = ( ~n29642 & n32667 ) | ( ~n29642 & n32669 ) | ( n32667 & n32669 ) ;
  assign n32671 = n32667 | n32669 ;
  assign n32672 = ( n29629 & n32670 ) | ( n29629 & n32671 ) | ( n32670 & n32671 ) ;
  assign n32673 = ~x5 & n32672 ;
  assign n32674 = x5 | n32672 ;
  assign n32675 = ( ~n32672 & n32673 ) | ( ~n32672 & n32674 ) | ( n32673 & n32674 ) ;
  assign n32676 = n32662 & n32675 ;
  assign n32677 = n32662 & ~n32676 ;
  assign n32678 = ~n32662 & n32675 ;
  assign n32679 = n32677 | n32678 ;
  assign n32680 = n31570 | n31973 ;
  assign n32681 = ~n31974 & n32680 ;
  assign n32682 = n8118 & n28492 ;
  assign n32683 = n8115 & ~n28503 ;
  assign n32684 = n28498 & n32683 ;
  assign n32685 = n32682 | n32684 ;
  assign n32686 = n8122 & ~n28714 ;
  assign n32687 = n8125 | n32686 ;
  assign n32688 = n32685 | n32687 ;
  assign n32689 = n32685 | n32686 ;
  assign n32690 = n28731 & ~n32689 ;
  assign n32691 = ( n28518 & ~n32689 ) | ( n28518 & n32690 ) | ( ~n32689 & n32690 ) ;
  assign n32692 = n32688 & ~n32691 ;
  assign n32693 = ( n28720 & n32688 ) | ( n28720 & n32692 ) | ( n32688 & n32692 ) ;
  assign n32694 = x5 & n32693 ;
  assign n32695 = x5 & ~n32693 ;
  assign n32696 = ( n32693 & ~n32694 ) | ( n32693 & n32695 ) | ( ~n32694 & n32695 ) ;
  assign n32697 = n32681 & n32696 ;
  assign n32698 = n31614 | n31967 ;
  assign n32699 = ~n31968 & n32698 ;
  assign n32700 = n8115 & ~n27371 ;
  assign n32701 = ~n27363 & n32700 ;
  assign n32702 = n8118 & ~n27606 ;
  assign n32703 = ~n27597 & n32702 ;
  assign n32704 = n32701 | n32703 ;
  assign n32705 = n8122 & ~n28503 ;
  assign n32706 = n28498 & n32705 ;
  assign n32707 = n32704 | n32706 ;
  assign n32708 = n28794 | n32707 ;
  assign n32709 = n28783 | n32708 ;
  assign n32710 = n8125 | n32706 ;
  assign n32711 = n32704 | n32710 ;
  assign n32712 = n32709 & n32711 ;
  assign n32713 = ~x5 & n32711 ;
  assign n32714 = n32709 & n32713 ;
  assign n32715 = x5 | n32713 ;
  assign n32716 = ( x5 & n32709 ) | ( x5 & n32715 ) | ( n32709 & n32715 ) ;
  assign n32717 = ( ~n32712 & n32714 ) | ( ~n32712 & n32716 ) | ( n32714 & n32716 ) ;
  assign n32718 = n32699 & n32717 ;
  assign n32719 = n31963 & n31965 ;
  assign n32720 = n31963 | n31965 ;
  assign n32721 = ~n32719 & n32720 ;
  assign n32722 = n8115 & ~n27133 ;
  assign n32723 = ~n27125 & n32722 ;
  assign n32724 = n8118 & ~n27371 ;
  assign n32725 = ~n27363 & n32724 ;
  assign n32726 = n32723 | n32725 ;
  assign n32727 = n8122 & ~n27606 ;
  assign n32728 = ~n27597 & n32727 ;
  assign n32729 = n32726 | n32728 ;
  assign n32730 = n8125 & n27630 ;
  assign n32731 = ~n27625 & n32730 ;
  assign n32732 = ( n8125 & ~n27634 ) | ( n8125 & n32731 ) | ( ~n27634 & n32731 ) ;
  assign n32733 = n32729 | n32732 ;
  assign n32734 = x5 | n32729 ;
  assign n32735 = n32732 | n32734 ;
  assign n32736 = ~x5 & n32734 ;
  assign n32737 = ( ~x5 & n32732 ) | ( ~x5 & n32736 ) | ( n32732 & n32736 ) ;
  assign n32738 = ( ~n32733 & n32735 ) | ( ~n32733 & n32737 ) | ( n32735 & n32737 ) ;
  assign n32739 = n32721 & n32738 ;
  assign n32740 = ~n32721 & n32738 ;
  assign n32741 = ( n32721 & ~n32739 ) | ( n32721 & n32740 ) | ( ~n32739 & n32740 ) ;
  assign n32742 = ~n31657 & n31961 ;
  assign n32743 = n31657 & ~n31961 ;
  assign n32744 = n32742 | n32743 ;
  assign n32745 = n8115 & ~n26526 ;
  assign n32746 = ~n26520 & n32745 ;
  assign n32747 = n8118 & ~n27133 ;
  assign n32748 = ~n27125 & n32747 ;
  assign n32749 = n32746 | n32748 ;
  assign n32750 = n8122 & ~n27371 ;
  assign n32751 = ~n27363 & n32750 ;
  assign n32752 = n32749 | n32751 ;
  assign n32753 = n8125 | n32751 ;
  assign n32754 = n32749 | n32753 ;
  assign n32755 = ( ~n27654 & n32752 ) | ( ~n27654 & n32754 ) | ( n32752 & n32754 ) ;
  assign n32756 = ~x5 & n32754 ;
  assign n32757 = ~x5 & n32752 ;
  assign n32758 = ( ~n27654 & n32756 ) | ( ~n27654 & n32757 ) | ( n32756 & n32757 ) ;
  assign n32759 = x5 | n32757 ;
  assign n32760 = x5 | n32756 ;
  assign n32761 = ( ~n27654 & n32759 ) | ( ~n27654 & n32760 ) | ( n32759 & n32760 ) ;
  assign n32762 = ( ~n32755 & n32758 ) | ( ~n32755 & n32761 ) | ( n32758 & n32761 ) ;
  assign n32763 = n32744 & n32762 ;
  assign n32764 = ~n31677 & n31959 ;
  assign n32765 = n31677 & ~n31959 ;
  assign n32766 = n32764 | n32765 ;
  assign n32767 = n8115 & ~n26270 ;
  assign n32768 = ~n26263 & n32767 ;
  assign n32769 = n8118 & ~n26526 ;
  assign n32770 = ~n26520 & n32769 ;
  assign n32771 = n32768 | n32770 ;
  assign n32772 = n8122 & ~n27133 ;
  assign n32773 = ~n27125 & n32772 ;
  assign n32774 = n32771 | n32773 ;
  assign n32775 = n8125 & n27699 ;
  assign n32776 = ( n8125 & ~n27696 ) | ( n8125 & n32775 ) | ( ~n27696 & n32775 ) ;
  assign n32777 = n32774 | n32776 ;
  assign n32778 = x5 | n32774 ;
  assign n32779 = n32776 | n32778 ;
  assign n32780 = ~x5 & n32778 ;
  assign n32781 = ( ~x5 & n32776 ) | ( ~x5 & n32780 ) | ( n32776 & n32780 ) ;
  assign n32782 = ( ~n32777 & n32779 ) | ( ~n32777 & n32781 ) | ( n32779 & n32781 ) ;
  assign n32783 = n32766 & n32782 ;
  assign n32784 = n32766 | n32782 ;
  assign n32785 = ~n32783 & n32784 ;
  assign n32786 = n31955 & n31957 ;
  assign n32787 = n31955 | n31957 ;
  assign n32788 = ~n32786 & n32787 ;
  assign n32789 = n8115 & n26017 ;
  assign n32790 = n8118 & ~n26270 ;
  assign n32791 = ~n26263 & n32790 ;
  assign n32792 = n32789 | n32791 ;
  assign n32793 = n8122 & ~n26526 ;
  assign n32794 = ~n26520 & n32793 ;
  assign n32796 = n8125 | n32794 ;
  assign n32797 = n32792 | n32796 ;
  assign n32795 = n32792 | n32794 ;
  assign n32798 = n32795 & n32797 ;
  assign n32799 = ( ~n26555 & n32797 ) | ( ~n26555 & n32798 ) | ( n32797 & n32798 ) ;
  assign n32800 = ( n26528 & n32797 ) | ( n26528 & n32798 ) | ( n32797 & n32798 ) ;
  assign n32801 = ( ~n26543 & n32799 ) | ( ~n26543 & n32800 ) | ( n32799 & n32800 ) ;
  assign n32802 = ~x5 & n32801 ;
  assign n32803 = x5 | n32801 ;
  assign n32804 = ( ~n32801 & n32802 ) | ( ~n32801 & n32803 ) | ( n32802 & n32803 ) ;
  assign n32805 = n32788 & n32804 ;
  assign n32806 = n31720 | n31953 ;
  assign n32807 = ~n31954 & n32806 ;
  assign n32808 = n8115 & ~n25728 ;
  assign n32809 = n8118 & n26017 ;
  assign n32810 = n32808 | n32809 ;
  assign n32811 = n8122 & ~n26270 ;
  assign n32812 = ~n26263 & n32811 ;
  assign n32814 = n8125 | n32812 ;
  assign n32815 = n32810 | n32814 ;
  assign n32813 = n32810 | n32812 ;
  assign n32816 = n32813 & n32815 ;
  assign n32817 = ( n26571 & n32815 ) | ( n26571 & n32816 ) | ( n32815 & n32816 ) ;
  assign n32818 = x5 & n32816 ;
  assign n32819 = x5 & n32815 ;
  assign n32820 = ( n26571 & n32818 ) | ( n26571 & n32819 ) | ( n32818 & n32819 ) ;
  assign n32821 = x5 & ~n32818 ;
  assign n32822 = x5 & ~n32819 ;
  assign n32823 = ( ~n26571 & n32821 ) | ( ~n26571 & n32822 ) | ( n32821 & n32822 ) ;
  assign n32824 = ( n32817 & ~n32820 ) | ( n32817 & n32823 ) | ( ~n32820 & n32823 ) ;
  assign n32825 = n32807 & n32824 ;
  assign n32826 = n32807 & ~n32825 ;
  assign n32827 = ~n32807 & n32824 ;
  assign n32828 = n32826 | n32827 ;
  assign n32829 = n31741 & n31951 ;
  assign n32830 = n31741 | n31951 ;
  assign n32831 = ~n32829 & n32830 ;
  assign n32832 = n8122 & n26017 ;
  assign n32833 = n8115 & ~n25046 ;
  assign n32834 = n8118 & ~n25728 ;
  assign n32835 = n32833 | n32834 ;
  assign n32836 = n32832 | n32835 ;
  assign n32837 = n8125 | n32832 ;
  assign n32838 = n32835 | n32837 ;
  assign n32839 = ( n26613 & n32836 ) | ( n26613 & n32838 ) | ( n32836 & n32838 ) ;
  assign n32840 = n32836 | n32838 ;
  assign n32841 = ( n26605 & n32839 ) | ( n26605 & n32840 ) | ( n32839 & n32840 ) ;
  assign n32842 = x5 & n32841 ;
  assign n32843 = x5 & ~n32841 ;
  assign n32844 = ( n32841 & ~n32842 ) | ( n32841 & n32843 ) | ( ~n32842 & n32843 ) ;
  assign n32845 = n32831 & n32844 ;
  assign n32846 = n32831 & ~n32845 ;
  assign n32847 = ~n32831 & n32844 ;
  assign n32848 = n32846 | n32847 ;
  assign n32849 = ( n31777 & n31778 ) | ( n31777 & n31949 ) | ( n31778 & n31949 ) ;
  assign n32850 = n31756 | n31777 ;
  assign n32851 = n31949 | n32850 ;
  assign n32852 = ~n32849 & n32851 ;
  assign n32853 = n8122 & ~n25728 ;
  assign n32854 = n8115 & n24770 ;
  assign n32855 = n8118 & ~n25046 ;
  assign n32856 = n32854 | n32855 ;
  assign n32857 = n32853 | n32856 ;
  assign n32858 = n8125 & n25740 ;
  assign n32859 = n8125 & n25731 ;
  assign n32860 = ( ~n25441 & n32858 ) | ( ~n25441 & n32859 ) | ( n32858 & n32859 ) ;
  assign n32861 = n32857 | n32860 ;
  assign n32862 = n8125 | n32857 ;
  assign n32863 = ( n25733 & n32861 ) | ( n25733 & n32862 ) | ( n32861 & n32862 ) ;
  assign n32864 = x5 | n32863 ;
  assign n32865 = ~x5 & n32863 ;
  assign n32866 = ( ~n32863 & n32864 ) | ( ~n32863 & n32865 ) | ( n32864 & n32865 ) ;
  assign n32867 = n32852 & n32866 ;
  assign n32868 = n31946 & ~n31949 ;
  assign n32871 = n8122 & ~n25046 ;
  assign n32872 = n8115 & ~n25054 ;
  assign n32873 = n8118 & n24770 ;
  assign n32874 = n32872 | n32873 ;
  assign n32875 = n32871 | n32874 ;
  assign n32876 = n8125 | n32871 ;
  assign n32877 = n32874 | n32876 ;
  assign n32878 = ( ~n25069 & n32875 ) | ( ~n25069 & n32877 ) | ( n32875 & n32877 ) ;
  assign n32879 = ~x5 & n32877 ;
  assign n32880 = ~x5 & n32875 ;
  assign n32881 = ( ~n25069 & n32879 ) | ( ~n25069 & n32880 ) | ( n32879 & n32880 ) ;
  assign n32882 = x5 | n32880 ;
  assign n32883 = x5 | n32879 ;
  assign n32884 = ( ~n25069 & n32882 ) | ( ~n25069 & n32883 ) | ( n32882 & n32883 ) ;
  assign n32885 = ( ~n32878 & n32881 ) | ( ~n32878 & n32884 ) | ( n32881 & n32884 ) ;
  assign n32869 = ~n31946 & n31948 ;
  assign n32886 = n32869 & n32885 ;
  assign n32887 = ( n32868 & n32885 ) | ( n32868 & n32886 ) | ( n32885 & n32886 ) ;
  assign n32870 = n32868 | n32869 ;
  assign n32888 = n32870 & ~n32887 ;
  assign n32889 = ~n32869 & n32885 ;
  assign n32890 = ~n32868 & n32889 ;
  assign n32891 = n32888 | n32890 ;
  assign n32892 = n31944 & ~n31945 ;
  assign n32893 = n31801 & ~n31945 ;
  assign n32894 = n32892 | n32893 ;
  assign n32895 = n8122 & n24770 ;
  assign n32896 = n8115 & n24167 ;
  assign n32897 = n8118 & ~n25054 ;
  assign n32898 = n32896 | n32897 ;
  assign n32899 = n32895 | n32898 ;
  assign n32900 = n8125 | n32899 ;
  assign n32901 = ( ~n25095 & n32899 ) | ( ~n25095 & n32900 ) | ( n32899 & n32900 ) ;
  assign n32902 = ~x5 & n32900 ;
  assign n32903 = ~x5 & n32899 ;
  assign n32904 = ( ~n25095 & n32902 ) | ( ~n25095 & n32903 ) | ( n32902 & n32903 ) ;
  assign n32905 = x5 | n32902 ;
  assign n32906 = x5 | n32903 ;
  assign n32907 = ( ~n25095 & n32905 ) | ( ~n25095 & n32906 ) | ( n32905 & n32906 ) ;
  assign n32908 = ( ~n32901 & n32904 ) | ( ~n32901 & n32907 ) | ( n32904 & n32907 ) ;
  assign n32909 = n32894 & n32908 ;
  assign n32910 = n32894 & ~n32909 ;
  assign n32911 = ~n32894 & n32908 ;
  assign n32912 = n32910 | n32911 ;
  assign n32913 = n31823 | n31917 ;
  assign n32914 = ~n31918 & n32913 ;
  assign n32915 = n8122 & n24167 ;
  assign n32916 = n8115 & n23316 ;
  assign n32917 = n8118 & n23614 ;
  assign n32918 = n32916 | n32917 ;
  assign n32919 = n32915 | n32918 ;
  assign n32920 = n8125 | n32919 ;
  assign n32921 = ( n24182 & n32919 ) | ( n24182 & n32920 ) | ( n32919 & n32920 ) ;
  assign n32922 = n32919 | n32920 ;
  assign n32923 = ( n24175 & n32921 ) | ( n24175 & n32922 ) | ( n32921 & n32922 ) ;
  assign n32924 = x5 & n32923 ;
  assign n32925 = x5 & ~n32923 ;
  assign n32926 = ( n32923 & ~n32924 ) | ( n32923 & n32925 ) | ( ~n32924 & n32925 ) ;
  assign n32927 = n32914 & n32926 ;
  assign n32928 = n31919 & n31942 ;
  assign n32929 = n31919 | n31942 ;
  assign n32930 = ~n32928 & n32929 ;
  assign n32931 = n8122 & ~n25054 ;
  assign n32932 = n8115 & n23614 ;
  assign n32933 = n8118 & n24167 ;
  assign n32934 = n32932 | n32933 ;
  assign n32935 = n32931 | n32934 ;
  assign n32936 = n8125 | n32931 ;
  assign n32937 = n32934 | n32936 ;
  assign n32938 = ( ~n25122 & n32935 ) | ( ~n25122 & n32937 ) | ( n32935 & n32937 ) ;
  assign n32939 = ~x5 & n32937 ;
  assign n32940 = ~x5 & n32935 ;
  assign n32941 = ( ~n25122 & n32939 ) | ( ~n25122 & n32940 ) | ( n32939 & n32940 ) ;
  assign n32942 = x5 | n32940 ;
  assign n32943 = x5 | n32939 ;
  assign n32944 = ( ~n25122 & n32942 ) | ( ~n25122 & n32943 ) | ( n32942 & n32943 ) ;
  assign n32945 = ( ~n32938 & n32941 ) | ( ~n32938 & n32944 ) | ( n32941 & n32944 ) ;
  assign n32946 = n32930 & n32945 ;
  assign n32947 = n32930 | n32945 ;
  assign n32948 = ~n32946 & n32947 ;
  assign n32949 = n32927 & n32948 ;
  assign n32950 = n32946 | n32948 ;
  assign n32951 = n31842 | n31915 ;
  assign n32952 = ~n31916 & n32951 ;
  assign n32953 = n8122 & n23614 ;
  assign n32954 = n8115 & n23620 ;
  assign n32955 = ( n8118 & n8446 ) | ( n8118 & n23620 ) | ( n8446 & n23620 ) ;
  assign n32956 = ( n23316 & n32954 ) | ( n23316 & n32955 ) | ( n32954 & n32955 ) ;
  assign n32958 = n8125 | n32956 ;
  assign n32959 = n32953 | n32958 ;
  assign n32957 = n32953 | n32956 ;
  assign n32960 = n32957 & n32959 ;
  assign n32961 = ( n23634 & n32959 ) | ( n23634 & n32960 ) | ( n32959 & n32960 ) ;
  assign n32962 = x5 & n32960 ;
  assign n32963 = x5 & n32959 ;
  assign n32964 = ( n23634 & n32962 ) | ( n23634 & n32963 ) | ( n32962 & n32963 ) ;
  assign n32965 = x5 & ~n32962 ;
  assign n32966 = x5 & ~n32963 ;
  assign n32967 = ( ~n23634 & n32965 ) | ( ~n23634 & n32966 ) | ( n32965 & n32966 ) ;
  assign n32968 = ( n32961 & ~n32964 ) | ( n32961 & n32967 ) | ( ~n32964 & n32967 ) ;
  assign n32969 = n32952 & n32968 ;
  assign n32970 = n32952 & ~n32969 ;
  assign n32971 = ~n32952 & n32968 ;
  assign n32972 = n32970 | n32971 ;
  assign n32973 = n31895 & n31909 ;
  assign n32974 = n31895 & ~n32973 ;
  assign n32975 = n8115 & ~n22385 ;
  assign n32976 = ( n8118 & n8446 ) | ( n8118 & ~n22385 ) | ( n8446 & ~n22385 ) ;
  assign n32977 = ( n22381 & n32975 ) | ( n22381 & n32976 ) | ( n32975 & n32976 ) ;
  assign n32978 = n8122 | n32977 ;
  assign n32979 = ( n23620 & n32977 ) | ( n23620 & n32978 ) | ( n32977 & n32978 ) ;
  assign n32980 = n8125 | n32979 ;
  assign n32981 = ( ~n23686 & n32979 ) | ( ~n23686 & n32980 ) | ( n32979 & n32980 ) ;
  assign n32982 = ~x5 & n32980 ;
  assign n32983 = ~x5 & n32979 ;
  assign n32984 = ( ~n23686 & n32982 ) | ( ~n23686 & n32983 ) | ( n32982 & n32983 ) ;
  assign n32985 = x5 | n32982 ;
  assign n32986 = x5 | n32983 ;
  assign n32987 = ( ~n23686 & n32985 ) | ( ~n23686 & n32986 ) | ( n32985 & n32986 ) ;
  assign n32988 = ( ~n32981 & n32984 ) | ( ~n32981 & n32987 ) | ( n32984 & n32987 ) ;
  assign n32989 = ~n31895 & n31909 ;
  assign n32990 = n32988 & n32989 ;
  assign n32991 = ( n32974 & n32988 ) | ( n32974 & n32990 ) | ( n32988 & n32990 ) ;
  assign n32992 = n32988 | n32989 ;
  assign n32993 = n32974 | n32992 ;
  assign n32994 = ~n32991 & n32993 ;
  assign n32995 = n31874 & n31892 ;
  assign n32996 = n31874 | n31892 ;
  assign n32997 = ~n32995 & n32996 ;
  assign n32998 = n8122 & n22381 ;
  assign n32999 = n8115 & ~n22398 ;
  assign n33000 = n8118 & ~n22385 ;
  assign n33001 = n32999 | n33000 ;
  assign n33002 = n32998 | n33001 ;
  assign n33003 = n8125 | n33002 ;
  assign n33004 = x5 & n33003 ;
  assign n33005 = x5 & n33002 ;
  assign n33006 = ( n22422 & n33004 ) | ( n22422 & n33005 ) | ( n33004 & n33005 ) ;
  assign n33007 = x5 | n33003 ;
  assign n33008 = x5 | n33002 ;
  assign n33009 = ( n22422 & n33007 ) | ( n22422 & n33008 ) | ( n33007 & n33008 ) ;
  assign n33010 = ~n33006 & n33009 ;
  assign n33011 = n32997 & n33010 ;
  assign n33012 = ~n32997 & n33010 ;
  assign n33013 = ( n32997 & ~n33011 ) | ( n32997 & n33012 ) | ( ~n33011 & n33012 ) ;
  assign n33014 = n31868 | n31870 ;
  assign n33015 = ~n31870 & n31872 ;
  assign n33016 = ( n31869 & n33014 ) | ( n31869 & ~n33015 ) | ( n33014 & ~n33015 ) ;
  assign n33017 = ~n31874 & n33016 ;
  assign n33018 = n8122 & ~n22385 ;
  assign n33019 = n8115 & n22393 ;
  assign n33020 = n8118 & ~n22398 ;
  assign n33021 = n33019 | n33020 ;
  assign n33022 = n33018 | n33021 ;
  assign n33023 = n8125 | n33018 ;
  assign n33024 = n33021 | n33023 ;
  assign n33025 = ( ~n22545 & n33022 ) | ( ~n22545 & n33024 ) | ( n33022 & n33024 ) ;
  assign n33026 = ~x5 & n33024 ;
  assign n33027 = ~x5 & n33022 ;
  assign n33028 = ( ~n22545 & n33026 ) | ( ~n22545 & n33027 ) | ( n33026 & n33027 ) ;
  assign n33029 = x5 | n33027 ;
  assign n33030 = x5 | n33026 ;
  assign n33031 = ( ~n22545 & n33029 ) | ( ~n22545 & n33030 ) | ( n33029 & n33030 ) ;
  assign n33032 = ( ~n33025 & n33028 ) | ( ~n33025 & n33031 ) | ( n33028 & n33031 ) ;
  assign n33033 = n33017 & n33032 ;
  assign n33034 = n8125 & n22474 ;
  assign n33035 = n8118 & ~n22409 ;
  assign n33036 = n8122 & ~n22406 ;
  assign n33037 = n33035 | n33036 ;
  assign n33038 = x5 | n33037 ;
  assign n33039 = n33034 | n33038 ;
  assign n33040 = ~x5 & n33039 ;
  assign n33041 = ( x5 & n21296 ) | ( x5 & n22409 ) | ( n21296 & n22409 ) ;
  assign n33042 = n33039 & n33041 ;
  assign n33043 = n33034 | n33037 ;
  assign n33044 = n33041 & ~n33043 ;
  assign n33045 = ( n33040 & n33042 ) | ( n33040 & n33044 ) | ( n33042 & n33044 ) ;
  assign n33046 = n8122 & n22393 ;
  assign n33047 = n8115 & ~n22409 ;
  assign n33048 = n8118 & ~n22406 ;
  assign n33049 = n33047 | n33048 ;
  assign n33050 = n33046 | n33049 ;
  assign n33051 = n22439 | n33050 ;
  assign n33052 = n8125 | n33046 ;
  assign n33053 = n33049 | n33052 ;
  assign n33054 = ~x5 & n33053 ;
  assign n33055 = n33051 & n33054 ;
  assign n33056 = x5 | n33055 ;
  assign n33057 = n7067 & ~n22409 ;
  assign n33058 = n33055 & n33057 ;
  assign n33059 = n33051 & n33053 ;
  assign n33060 = n33057 & ~n33059 ;
  assign n33061 = ( n33056 & n33058 ) | ( n33056 & n33060 ) | ( n33058 & n33060 ) ;
  assign n33062 = n33045 & n33061 ;
  assign n33063 = ( n33055 & n33056 ) | ( n33055 & ~n33059 ) | ( n33056 & ~n33059 ) ;
  assign n33064 = n33045 | n33057 ;
  assign n33065 = ( n33057 & n33063 ) | ( n33057 & n33064 ) | ( n33063 & n33064 ) ;
  assign n33066 = ~n33062 & n33065 ;
  assign n33067 = n8115 & ~n22406 ;
  assign n33068 = n8118 & n22393 ;
  assign n33069 = n33067 | n33068 ;
  assign n33070 = n8122 & ~n22398 ;
  assign n33071 = n8125 | n33070 ;
  assign n33072 = n33069 | n33071 ;
  assign n33073 = x5 & n33072 ;
  assign n33074 = n33069 | n33070 ;
  assign n33075 = x5 & n33074 ;
  assign n33076 = ( n22608 & n33073 ) | ( n22608 & n33075 ) | ( n33073 & n33075 ) ;
  assign n33077 = x5 | n33072 ;
  assign n33078 = x5 | n33074 ;
  assign n33079 = ( n22608 & n33077 ) | ( n22608 & n33078 ) | ( n33077 & n33078 ) ;
  assign n33080 = ~n33076 & n33079 ;
  assign n33081 = n33062 | n33080 ;
  assign n33082 = ( n33062 & n33066 ) | ( n33062 & n33081 ) | ( n33066 & n33081 ) ;
  assign n33083 = n33017 | n33032 ;
  assign n33084 = ~n33033 & n33083 ;
  assign n33085 = n33033 | n33084 ;
  assign n33086 = ( n33033 & n33082 ) | ( n33033 & n33085 ) | ( n33082 & n33085 ) ;
  assign n33087 = n33013 & n33086 ;
  assign n33088 = n33011 | n33087 ;
  assign n33089 = n32994 & n33088 ;
  assign n33090 = n32991 | n33089 ;
  assign n33091 = n8115 & n22381 ;
  assign n33092 = ( n8118 & n8446 ) | ( n8118 & n22381 ) | ( n8446 & n22381 ) ;
  assign n33093 = ( n23620 & n33091 ) | ( n23620 & n33092 ) | ( n33091 & n33092 ) ;
  assign n33094 = n8122 | n33092 ;
  assign n33095 = n8122 | n33091 ;
  assign n33096 = ( n23620 & n33094 ) | ( n23620 & n33095 ) | ( n33094 & n33095 ) ;
  assign n33097 = ( n23316 & n33093 ) | ( n23316 & n33096 ) | ( n33093 & n33096 ) ;
  assign n33098 = n8125 | n33097 ;
  assign n33099 = ~x5 & n33098 ;
  assign n33100 = ~x5 & n33097 ;
  assign n33101 = ( n23661 & n33099 ) | ( n23661 & n33100 ) | ( n33099 & n33100 ) ;
  assign n33102 = ( x5 & n21256 ) | ( x5 & n33097 ) | ( n21256 & n33097 ) ;
  assign n33103 = x5 & ~n33102 ;
  assign n33104 = x5 & n33097 ;
  assign n33105 = x5 & ~n33104 ;
  assign n33106 = ( ~n23661 & n33103 ) | ( ~n23661 & n33105 ) | ( n33103 & n33105 ) ;
  assign n33107 = n33101 | n33106 ;
  assign n33108 = n31911 & n31913 ;
  assign n33109 = n31911 | n31913 ;
  assign n33110 = ~n33108 & n33109 ;
  assign n33111 = n33107 & n33110 ;
  assign n33112 = n33107 | n33110 ;
  assign n33113 = ~n33111 & n33112 ;
  assign n33114 = n33111 | n33113 ;
  assign n33115 = ( n33090 & n33111 ) | ( n33090 & n33114 ) | ( n33111 & n33114 ) ;
  assign n33116 = n32972 & n33115 ;
  assign n33117 = n32969 | n33116 ;
  assign n33118 = ~n32914 & n32926 ;
  assign n33119 = ( n32914 & ~n32927 ) | ( n32914 & n33118 ) | ( ~n32927 & n33118 ) ;
  assign n33120 = n33117 & n33119 ;
  assign n33121 = n32946 | n33120 ;
  assign n33122 = ( n32949 & n32950 ) | ( n32949 & n33121 ) | ( n32950 & n33121 ) ;
  assign n33123 = n32909 | n33122 ;
  assign n33124 = ( n32909 & n32912 ) | ( n32909 & n33123 ) | ( n32912 & n33123 ) ;
  assign n33125 = n32891 & n33124 ;
  assign n33126 = n32887 | n33125 ;
  assign n33127 = ~n32852 & n32866 ;
  assign n33128 = ( n32852 & ~n32867 ) | ( n32852 & n33127 ) | ( ~n32867 & n33127 ) ;
  assign n33129 = n32867 | n33128 ;
  assign n33130 = ( n32867 & n33126 ) | ( n32867 & n33129 ) | ( n33126 & n33129 ) ;
  assign n33131 = n32845 | n33130 ;
  assign n33132 = ( n32845 & n32848 ) | ( n32845 & n33131 ) | ( n32848 & n33131 ) ;
  assign n33133 = n32828 & n33132 ;
  assign n33134 = n32825 | n33133 ;
  assign n33135 = n32788 | n32804 ;
  assign n33136 = ~n32805 & n33135 ;
  assign n33137 = n32805 | n33136 ;
  assign n33138 = ( n32805 & n33134 ) | ( n32805 & n33137 ) | ( n33134 & n33137 ) ;
  assign n33139 = n32785 & n33138 ;
  assign n33140 = n32783 | n33139 ;
  assign n33141 = n32744 | n32762 ;
  assign n33142 = ~n32763 & n33141 ;
  assign n33143 = n32763 | n33142 ;
  assign n33144 = ( n32763 & n33140 ) | ( n32763 & n33143 ) | ( n33140 & n33143 ) ;
  assign n33145 = n32741 & n33144 ;
  assign n33146 = n32739 | n33145 ;
  assign n33147 = n32699 & ~n32718 ;
  assign n33148 = ~n32699 & n32717 ;
  assign n33149 = n33147 | n33148 ;
  assign n33150 = n33146 & n33149 ;
  assign n33151 = n32718 | n33150 ;
  assign n33152 = n31969 & n31971 ;
  assign n33153 = n31969 | n31971 ;
  assign n33154 = ~n33152 & n33153 ;
  assign n33155 = n8122 & n28492 ;
  assign n33156 = n8115 & ~n27606 ;
  assign n33157 = ~n27597 & n33156 ;
  assign n33158 = n8118 & ~n28503 ;
  assign n33159 = n28498 & n33158 ;
  assign n33160 = n33157 | n33159 ;
  assign n33161 = n33155 | n33160 ;
  assign n33162 = n8125 | n33161 ;
  assign n33163 = n33161 & n33162 ;
  assign n33164 = ( ~n28749 & n33162 ) | ( ~n28749 & n33163 ) | ( n33162 & n33163 ) ;
  assign n33165 = ~x5 & n33163 ;
  assign n33166 = ~x5 & n33162 ;
  assign n33167 = ( ~n28749 & n33165 ) | ( ~n28749 & n33166 ) | ( n33165 & n33166 ) ;
  assign n33168 = x5 | n33165 ;
  assign n33169 = x5 | n33166 ;
  assign n33170 = ( ~n28749 & n33168 ) | ( ~n28749 & n33169 ) | ( n33168 & n33169 ) ;
  assign n33171 = ( ~n33164 & n33167 ) | ( ~n33164 & n33170 ) | ( n33167 & n33170 ) ;
  assign n33172 = n33154 & n33171 ;
  assign n33173 = n33154 & ~n33172 ;
  assign n33174 = ~n33154 & n33171 ;
  assign n33175 = n33173 | n33174 ;
  assign n33176 = n33151 & n33175 ;
  assign n33177 = n32681 | n32696 ;
  assign n33178 = ~n32697 & n33177 ;
  assign n33179 = n33172 & n33178 ;
  assign n33180 = ( n33176 & n33178 ) | ( n33176 & n33179 ) | ( n33178 & n33179 ) ;
  assign n33181 = n32697 | n33180 ;
  assign n33182 = n32676 | n33181 ;
  assign n33183 = ( n32676 & n32679 ) | ( n32676 & n33182 ) | ( n32679 & n33182 ) ;
  assign n33184 = n32656 | n33183 ;
  assign n33185 = ( n32656 & n32659 ) | ( n32656 & n33184 ) | ( n32659 & n33184 ) ;
  assign n33186 = ~n32623 & n32636 ;
  assign n33187 = ( n32623 & ~n32637 ) | ( n32623 & n33186 ) | ( ~n32637 & n33186 ) ;
  assign n33188 = n32637 | n33187 ;
  assign n33189 = ( n32637 & n33185 ) | ( n32637 & n33188 ) | ( n33185 & n33188 ) ;
  assign n33190 = n32617 | n33189 ;
  assign n33191 = ( n32617 & n32620 ) | ( n32617 & n33190 ) | ( n32620 & n33190 ) ;
  assign n33192 = n32580 | n32596 ;
  assign n33193 = ~n32597 & n33192 ;
  assign n33194 = n32597 | n33193 ;
  assign n33195 = ( n32597 & n33191 ) | ( n32597 & n33194 ) | ( n33191 & n33194 ) ;
  assign n33196 = ~n32577 & n33195 ;
  assign n33197 = n32575 | n33196 ;
  assign n33198 = n32541 & ~n32556 ;
  assign n33199 = n32557 | n33198 ;
  assign n33200 = ~n32557 & n33199 ;
  assign n33201 = ( n32557 & n33197 ) | ( n32557 & ~n33200 ) | ( n33197 & ~n33200 ) ;
  assign n33202 = n32538 & n33201 ;
  assign n33203 = n32536 | n33202 ;
  assign n33204 = n32506 | n33203 ;
  assign n33205 = ( n32506 & ~n32508 ) | ( n32506 & n33204 ) | ( ~n32508 & n33204 ) ;
  assign n33206 = n32476 & ~n33205 ;
  assign n33207 = ~n32476 & n33205 ;
  assign n33208 = n33206 | n33207 ;
  assign n33209 = n1062 & ~n21570 ;
  assign n33210 = n22270 & n33209 ;
  assign n33211 = ( n1062 & n22304 ) | ( n1062 & n33210 ) | ( n22304 & n33210 ) ;
  assign n33212 = n110 | n255 ;
  assign n33213 = n262 | n33212 ;
  assign n33214 = n8012 | n33213 ;
  assign n33215 = n8999 | n33214 ;
  assign n33216 = n170 | n33215 ;
  assign n33217 = n8995 | n33216 ;
  assign n33218 = n401 | n33217 ;
  assign n33219 = n1002 | n7998 ;
  assign n33220 = n7996 | n33219 ;
  assign n33221 = n33218 | n33220 ;
  assign n33222 = n7947 & ~n33221 ;
  assign n33223 = n32348 & n33222 ;
  assign n33224 = n32348 | n33222 ;
  assign n33225 = ~n33223 & n33224 ;
  assign n33226 = n2308 | n2315 ;
  assign n33227 = n2312 | n33226 ;
  assign n33228 = n2306 | n33227 ;
  assign n33229 = ~n23229 & n33228 ;
  assign n33230 = ( n23154 & n33228 ) | ( n23154 & n33229 ) | ( n33228 & n33229 ) ;
  assign n33231 = ~n23232 & n33228 ;
  assign n33232 = ~n23231 & n33228 ;
  assign n33233 = ( n9072 & n33231 ) | ( n9072 & n33232 ) | ( n33231 & n33232 ) ;
  assign n33234 = ( ~n21543 & n33230 ) | ( ~n21543 & n33233 ) | ( n33230 & n33233 ) ;
  assign n33235 = ( ~n21545 & n33230 ) | ( ~n21545 & n33233 ) | ( n33230 & n33233 ) ;
  assign n33236 = ( ~n15882 & n33234 ) | ( ~n15882 & n33235 ) | ( n33234 & n33235 ) ;
  assign n33237 = ~x26 & n33234 ;
  assign n33238 = ~x26 & n33235 ;
  assign n33239 = ( ~n15882 & n33237 ) | ( ~n15882 & n33238 ) | ( n33237 & n33238 ) ;
  assign n33240 = x26 | n33237 ;
  assign n33241 = x26 | n33238 ;
  assign n33242 = ( ~n15882 & n33240 ) | ( ~n15882 & n33241 ) | ( n33240 & n33241 ) ;
  assign n33243 = ( ~n33236 & n33239 ) | ( ~n33236 & n33242 ) | ( n33239 & n33242 ) ;
  assign n33244 = n33225 & ~n33243 ;
  assign n33245 = ~n33225 & n33243 ;
  assign n33246 = n33244 | n33245 ;
  assign n33247 = n4247 | n5948 ;
  assign n33248 = n7888 | n33247 ;
  assign n33249 = n7988 | n33248 ;
  assign n33250 = n7871 | n33249 ;
  assign n33251 = n2853 | n20360 ;
  assign n33252 = n8004 | n33251 ;
  assign n33253 = n796 | n33252 ;
  assign n33254 = n33250 | n33253 ;
  assign n33255 = n262 | n406 ;
  assign n33256 = n447 | n33255 ;
  assign n33257 = n401 | n8026 ;
  assign n33258 = n33256 | n33257 ;
  assign n33259 = n7863 | n33258 ;
  assign n33260 = n33254 | n33259 ;
  assign n33261 = n32348 & n33260 ;
  assign n33262 = n1060 & ~n20618 ;
  assign n33263 = n1065 & n20609 ;
  assign n33264 = n33262 | n33263 ;
  assign n33265 = n1057 & ~n21563 ;
  assign n33266 = ~n33261 & n33265 ;
  assign n33267 = ( ~n33261 & n33264 ) | ( ~n33261 & n33266 ) | ( n33264 & n33266 ) ;
  assign n33268 = n32348 | n33260 ;
  assign n33269 = n33261 | n33268 ;
  assign n33270 = ( n33261 & n33267 ) | ( n33261 & n33269 ) | ( n33267 & n33269 ) ;
  assign n33271 = ~n33246 & n33270 ;
  assign n33272 = ~n33261 & n33268 ;
  assign n33273 = n33261 | n33272 ;
  assign n33274 = ~n33246 & n33273 ;
  assign n33275 = ( n33211 & n33271 ) | ( n33211 & n33274 ) | ( n33271 & n33274 ) ;
  assign n33276 = n33246 & ~n33270 ;
  assign n33277 = n33246 & ~n33273 ;
  assign n33278 = ( ~n33211 & n33276 ) | ( ~n33211 & n33277 ) | ( n33276 & n33277 ) ;
  assign n33279 = n33275 | n33278 ;
  assign n33280 = n1057 & ~n21517 ;
  assign n33281 = n1060 & n20609 ;
  assign n33282 = n1065 & ~n21563 ;
  assign n33283 = n33281 | n33282 ;
  assign n33284 = n33280 | n33283 ;
  assign n33285 = n1062 | n33280 ;
  assign n33286 = n33283 | n33285 ;
  assign n33287 = ( ~n22283 & n33284 ) | ( ~n22283 & n33286 ) | ( n33284 & n33286 ) ;
  assign n33288 = n33284 & n33286 ;
  assign n33289 = ( ~n22271 & n33287 ) | ( ~n22271 & n33288 ) | ( n33287 & n33288 ) ;
  assign n33290 = n33279 & n33289 ;
  assign n33291 = n33279 | n33289 ;
  assign n33292 = ~n33290 & n33291 ;
  assign n33293 = n1829 & ~n23240 ;
  assign n33294 = n1826 & ~n21551 ;
  assign n33295 = n1823 & n23227 ;
  assign n33296 = ( n1823 & n23217 ) | ( n1823 & n33295 ) | ( n23217 & n33295 ) ;
  assign n33297 = n33294 | n33296 ;
  assign n33298 = n33293 | n33297 ;
  assign n33299 = n1821 | n33293 ;
  assign n33300 = n33297 | n33299 ;
  assign n33301 = ( n23260 & n33298 ) | ( n23260 & n33300 ) | ( n33298 & n33300 ) ;
  assign n33302 = x29 & n33300 ;
  assign n33303 = x29 & n33298 ;
  assign n33304 = ( n23260 & n33302 ) | ( n23260 & n33303 ) | ( n33302 & n33303 ) ;
  assign n33305 = x29 & ~n33303 ;
  assign n33306 = x29 & ~n33302 ;
  assign n33307 = ( ~n23260 & n33305 ) | ( ~n23260 & n33306 ) | ( n33305 & n33306 ) ;
  assign n33308 = ( n33301 & ~n33304 ) | ( n33301 & n33307 ) | ( ~n33304 & n33307 ) ;
  assign n33309 = ~n33292 & n33308 ;
  assign n33310 = n33292 & ~n33308 ;
  assign n33311 = n33309 | n33310 ;
  assign n33312 = n32351 | n32372 ;
  assign n33313 = n33268 & ~n33269 ;
  assign n33314 = ( ~n33267 & n33272 ) | ( ~n33267 & n33313 ) | ( n33272 & n33313 ) ;
  assign n33315 = ~n33211 & n33314 ;
  assign n33316 = n33312 & n33315 ;
  assign n33317 = n33264 | n33265 ;
  assign n33318 = ~n33272 & n33317 ;
  assign n33319 = ( n33211 & ~n33272 ) | ( n33211 & n33318 ) | ( ~n33272 & n33318 ) ;
  assign n33320 = ( n33312 & n33316 ) | ( n33312 & n33319 ) | ( n33316 & n33319 ) ;
  assign n33321 = n32376 | n32392 ;
  assign n33322 = ( n32376 & ~n32377 ) | ( n32376 & n33321 ) | ( ~n32377 & n33321 ) ;
  assign n33323 = n33312 | n33315 ;
  assign n33324 = n33319 | n33323 ;
  assign n33325 = ~n33320 & n33324 ;
  assign n33326 = n33320 | n33325 ;
  assign n33327 = ( n33320 & n33322 ) | ( n33320 & n33326 ) | ( n33322 & n33326 ) ;
  assign n33328 = n33311 & ~n33327 ;
  assign n33329 = ~n33311 & n33327 ;
  assign n33330 = n33328 | n33329 ;
  assign n33331 = n33322 & n33325 ;
  assign n33332 = n33322 | n33325 ;
  assign n33333 = ~n33331 & n33332 ;
  assign n33334 = ~n23234 & n33226 ;
  assign n33335 = ~n23235 & n33226 ;
  assign n33336 = ( ~n15882 & n33334 ) | ( ~n15882 & n33335 ) | ( n33334 & n33335 ) ;
  assign n33337 = n2312 | n33334 ;
  assign n33338 = n2312 | n33335 ;
  assign n33339 = ( ~n15882 & n33337 ) | ( ~n15882 & n33338 ) | ( n33337 & n33338 ) ;
  assign n33340 = ( ~n23240 & n33336 ) | ( ~n23240 & n33339 ) | ( n33336 & n33339 ) ;
  assign n33341 = n2306 & ~n24135 ;
  assign n33342 = n2306 & ~n23240 ;
  assign n33343 = ( ~n23575 & n33341 ) | ( ~n23575 & n33342 ) | ( n33341 & n33342 ) ;
  assign n33344 = ( ~n23577 & n33341 ) | ( ~n23577 & n33342 ) | ( n33341 & n33342 ) ;
  assign n33345 = n33343 & n33344 ;
  assign n33346 = n33340 | n33345 ;
  assign n33347 = ( n21554 & n33343 ) | ( n21554 & n33344 ) | ( n33343 & n33344 ) ;
  assign n33348 = n33340 | n33347 ;
  assign n33349 = ( ~n21584 & n33346 ) | ( ~n21584 & n33348 ) | ( n33346 & n33348 ) ;
  assign n33350 = x26 & n33348 ;
  assign n33351 = x26 & n33346 ;
  assign n33352 = ( ~n21584 & n33350 ) | ( ~n21584 & n33351 ) | ( n33350 & n33351 ) ;
  assign n33353 = n33349 & ~n33352 ;
  assign n33354 = x26 & ~n33348 ;
  assign n33355 = x26 & ~n33346 ;
  assign n33356 = ( n21584 & n33354 ) | ( n21584 & n33355 ) | ( n33354 & n33355 ) ;
  assign n33357 = n33353 | n33356 ;
  assign n33358 = n1826 & ~n21517 ;
  assign n33359 = n1823 & ~n21551 ;
  assign n33360 = n33358 | n33359 ;
  assign n33361 = n1829 & n23227 ;
  assign n33362 = ( n1829 & n23217 ) | ( n1829 & n33361 ) | ( n23217 & n33361 ) ;
  assign n33363 = n33360 | n33362 ;
  assign n33364 = n1821 & n23299 ;
  assign n33365 = n1821 & n23298 ;
  assign n33366 = ( n21584 & n33364 ) | ( n21584 & n33365 ) | ( n33364 & n33365 ) ;
  assign n33367 = n33363 | n33366 ;
  assign n33368 = n1821 | n33363 ;
  assign n33369 = ( n23289 & n33367 ) | ( n23289 & n33368 ) | ( n33367 & n33368 ) ;
  assign n33370 = ~x29 & n33369 ;
  assign n33371 = x29 & n33362 ;
  assign n33372 = ( x29 & n33360 ) | ( x29 & n33371 ) | ( n33360 & n33371 ) ;
  assign n33373 = x29 & ~n33372 ;
  assign n33374 = ~n33366 & n33373 ;
  assign n33375 = ~n1821 & n33373 ;
  assign n33376 = ( ~n23289 & n33374 ) | ( ~n23289 & n33375 ) | ( n33374 & n33375 ) ;
  assign n33377 = n33357 & n33376 ;
  assign n33378 = ( n33357 & n33370 ) | ( n33357 & n33377 ) | ( n33370 & n33377 ) ;
  assign n33379 = n33357 | n33376 ;
  assign n33380 = n33370 | n33379 ;
  assign n33381 = ~n33378 & n33380 ;
  assign n33382 = n33378 | n33381 ;
  assign n33383 = ( n33333 & n33378 ) | ( n33333 & n33382 ) | ( n33378 & n33382 ) ;
  assign n33384 = ~n33330 & n33383 ;
  assign n33385 = n33330 & ~n33383 ;
  assign n33386 = n33384 | n33385 ;
  assign n33387 = n33333 & n33381 ;
  assign n33388 = n33333 | n33381 ;
  assign n33389 = ~n33387 & n33388 ;
  assign n33390 = n32397 | n32417 ;
  assign n33391 = ( n32397 & ~n32399 ) | ( n32397 & n33390 ) | ( ~n32399 & n33390 ) ;
  assign n33392 = n33389 & n33391 ;
  assign n33393 = n33389 | n33391 ;
  assign n33394 = ~n33392 & n33393 ;
  assign n33395 = n32421 | n32425 ;
  assign n33396 = n33394 & n33395 ;
  assign n33397 = n33392 | n33396 ;
  assign n33398 = ~n33386 & n33397 ;
  assign n33399 = ~n32421 & n32424 ;
  assign n33400 = n33394 & ~n33399 ;
  assign n33401 = n33392 | n33400 ;
  assign n33402 = ~n33386 & n33401 ;
  assign n33403 = ( n32274 & n33398 ) | ( n32274 & n33402 ) | ( n33398 & n33402 ) ;
  assign n33404 = n32421 | n32428 ;
  assign n33405 = n33394 & n33404 ;
  assign n33406 = n33392 | n33405 ;
  assign n33407 = ~n33386 & n33406 ;
  assign n33408 = n32421 | n32430 ;
  assign n33409 = n33394 & n33408 ;
  assign n33410 = n33392 | n33409 ;
  assign n33411 = ~n33386 & n33410 ;
  assign n33412 = ( n31274 & n33407 ) | ( n31274 & n33411 ) | ( n33407 & n33411 ) ;
  assign n33413 = ( n28465 & n33403 ) | ( n28465 & n33412 ) | ( n33403 & n33412 ) ;
  assign n33414 = n33403 & n33412 ;
  assign n33415 = ( n28489 & n33413 ) | ( n28489 & n33414 ) | ( n33413 & n33414 ) ;
  assign n33416 = ( n32274 & n33397 ) | ( n32274 & n33401 ) | ( n33397 & n33401 ) ;
  assign n33417 = ( n31274 & n33406 ) | ( n31274 & n33410 ) | ( n33406 & n33410 ) ;
  assign n33418 = n33416 & n33417 ;
  assign n33419 = n33386 & ~n33418 ;
  assign n33420 = ( n28465 & n33416 ) | ( n28465 & n33417 ) | ( n33416 & n33417 ) ;
  assign n33421 = n33386 & ~n33420 ;
  assign n33422 = ( ~n28489 & n33419 ) | ( ~n28489 & n33421 ) | ( n33419 & n33421 ) ;
  assign n33423 = n33415 | n33422 ;
  assign n33424 = ( n32274 & n33396 ) | ( n32274 & n33400 ) | ( n33396 & n33400 ) ;
  assign n33425 = ( n31274 & n33405 ) | ( n31274 & n33409 ) | ( n33405 & n33409 ) ;
  assign n33426 = ( n28465 & n33424 ) | ( n28465 & n33425 ) | ( n33424 & n33425 ) ;
  assign n33427 = n33424 & n33425 ;
  assign n33428 = ( n28489 & n33426 ) | ( n28489 & n33427 ) | ( n33426 & n33427 ) ;
  assign n33429 = ( n32274 & n33395 ) | ( n32274 & ~n33399 ) | ( n33395 & ~n33399 ) ;
  assign n33430 = ( n31274 & n33404 ) | ( n31274 & n33408 ) | ( n33404 & n33408 ) ;
  assign n33431 = n33429 & n33430 ;
  assign n33432 = n33394 | n33431 ;
  assign n33433 = ( n28465 & n33429 ) | ( n28465 & n33430 ) | ( n33429 & n33430 ) ;
  assign n33434 = n33394 | n33433 ;
  assign n33435 = ( n28489 & n33432 ) | ( n28489 & n33434 ) | ( n33432 & n33434 ) ;
  assign n33436 = ~n33428 & n33435 ;
  assign n33437 = ~n33423 & n33436 ;
  assign n33438 = n33423 & ~n33436 ;
  assign n33439 = ~n32442 & n33436 ;
  assign n33440 = n32442 & ~n33436 ;
  assign n33441 = n33439 | n33440 ;
  assign n33442 = ~n33438 & n33439 ;
  assign n33443 = ( n33438 & n33441 ) | ( n33438 & ~n33442 ) | ( n33441 & ~n33442 ) ;
  assign n33444 = ~n33437 & n33443 ;
  assign n33445 = n33437 | n33442 ;
  assign n33446 = ( n32456 & ~n33444 ) | ( n32456 & n33445 ) | ( ~n33444 & n33445 ) ;
  assign n33447 = n1057 & ~n21551 ;
  assign n33448 = n1060 & ~n21563 ;
  assign n33449 = n1065 & ~n21517 ;
  assign n33450 = n33448 | n33449 ;
  assign n33451 = n33447 | n33450 ;
  assign n33452 = n1062 | n33447 ;
  assign n33453 = n33450 | n33452 ;
  assign n33454 = ( ~n21587 & n33451 ) | ( ~n21587 & n33453 ) | ( n33451 & n33453 ) ;
  assign n33455 = n8995 | n33215 ;
  assign n33456 = n9044 | n9045 ;
  assign n33457 = n9040 | n33456 ;
  assign n33458 = n33455 | n33457 ;
  assign n33459 = n7980 | n33458 ;
  assign n33460 = n170 | n33459 ;
  assign n33461 = ( n33224 & ~n33225 ) | ( n33224 & n33460 ) | ( ~n33225 & n33460 ) ;
  assign n33462 = n33224 | n33460 ;
  assign n33463 = ( n33243 & n33461 ) | ( n33243 & n33462 ) | ( n33461 & n33462 ) ;
  assign n33464 = n33224 & ~n33225 ;
  assign n33465 = n33460 & n33464 ;
  assign n33466 = n33224 & n33460 ;
  assign n33467 = ( n33243 & n33465 ) | ( n33243 & n33466 ) | ( n33465 & n33466 ) ;
  assign n33468 = n33463 & ~n33467 ;
  assign n33469 = n33453 & n33468 ;
  assign n33470 = n33451 & n33468 ;
  assign n33471 = ( ~n21587 & n33469 ) | ( ~n21587 & n33470 ) | ( n33469 & n33470 ) ;
  assign n33472 = n33468 & ~n33470 ;
  assign n33473 = n33468 & ~n33469 ;
  assign n33474 = ( n21587 & n33472 ) | ( n21587 & n33473 ) | ( n33472 & n33473 ) ;
  assign n33475 = ( n33454 & ~n33471 ) | ( n33454 & n33474 ) | ( ~n33471 & n33474 ) ;
  assign n33476 = n33275 | n33289 ;
  assign n33477 = ( n33275 & ~n33279 ) | ( n33275 & n33476 ) | ( ~n33279 & n33476 ) ;
  assign n33478 = n33475 | n33477 ;
  assign n33479 = n33475 & n33477 ;
  assign n33480 = n33478 & ~n33479 ;
  assign n33481 = n1823 & ~n23240 ;
  assign n33482 = n1826 & n23227 ;
  assign n33483 = ( n1826 & n23217 ) | ( n1826 & n33482 ) | ( n23217 & n33482 ) ;
  assign n33484 = n33481 | n33483 ;
  assign n33485 = n1829 & ~n23234 ;
  assign n33486 = n1829 & ~n23235 ;
  assign n33487 = ( ~n15882 & n33485 ) | ( ~n15882 & n33486 ) | ( n33485 & n33486 ) ;
  assign n33489 = n1821 | n33487 ;
  assign n33490 = n33484 | n33489 ;
  assign n33488 = n33484 | n33487 ;
  assign n33491 = n33488 & n33490 ;
  assign n33492 = ( ~n23587 & n33490 ) | ( ~n23587 & n33491 ) | ( n33490 & n33491 ) ;
  assign n33493 = ~x29 & n33491 ;
  assign n33494 = ~x29 & n33490 ;
  assign n33495 = ( ~n23587 & n33493 ) | ( ~n23587 & n33494 ) | ( n33493 & n33494 ) ;
  assign n33496 = x29 | n33493 ;
  assign n33497 = x29 | n33494 ;
  assign n33498 = ( ~n23587 & n33496 ) | ( ~n23587 & n33497 ) | ( n33496 & n33497 ) ;
  assign n33499 = ( ~n33492 & n33495 ) | ( ~n33492 & n33498 ) | ( n33495 & n33498 ) ;
  assign n33500 = n33480 & n33499 ;
  assign n33501 = n33480 | n33499 ;
  assign n33502 = ~n33500 & n33501 ;
  assign n33503 = ~n33309 & n33311 ;
  assign n33504 = ( n33309 & n33327 ) | ( n33309 & ~n33503 ) | ( n33327 & ~n33503 ) ;
  assign n33505 = n33502 & n33504 ;
  assign n33506 = n33502 | n33504 ;
  assign n33507 = ~n33505 & n33506 ;
  assign n33508 = n33384 | n33407 ;
  assign n33509 = n33384 | n33411 ;
  assign n33510 = ( n31274 & n33508 ) | ( n31274 & n33509 ) | ( n33508 & n33509 ) ;
  assign n33511 = n33507 & n33510 ;
  assign n33512 = n33384 | n33398 ;
  assign n33513 = n33507 & n33512 ;
  assign n33514 = n33384 | n33402 ;
  assign n33515 = n33507 & n33514 ;
  assign n33516 = ( n32274 & n33513 ) | ( n32274 & n33515 ) | ( n33513 & n33515 ) ;
  assign n33517 = ( n28465 & n33511 ) | ( n28465 & n33516 ) | ( n33511 & n33516 ) ;
  assign n33518 = n33511 & n33516 ;
  assign n33519 = ( n28489 & n33517 ) | ( n28489 & n33518 ) | ( n33517 & n33518 ) ;
  assign n33520 = ( n32274 & n33512 ) | ( n32274 & n33514 ) | ( n33512 & n33514 ) ;
  assign n33521 = n33510 & n33520 ;
  assign n33522 = n33507 | n33521 ;
  assign n33523 = ( n28465 & n33510 ) | ( n28465 & n33520 ) | ( n33510 & n33520 ) ;
  assign n33524 = n33507 | n33523 ;
  assign n33525 = ( n28489 & n33522 ) | ( n28489 & n33524 ) | ( n33522 & n33524 ) ;
  assign n33526 = ~n33519 & n33525 ;
  assign n33527 = ~n33423 & n33526 ;
  assign n33528 = n33423 & ~n33526 ;
  assign n33529 = n33437 & ~n33528 ;
  assign n33530 = ( n33442 & ~n33528 ) | ( n33442 & n33529 ) | ( ~n33528 & n33529 ) ;
  assign n33531 = ~n33527 & n33530 ;
  assign n33532 = ~n33527 & n33529 ;
  assign n33533 = n33527 | n33528 ;
  assign n33534 = ( n33443 & ~n33532 ) | ( n33443 & n33533 ) | ( ~n33532 & n33533 ) ;
  assign n33535 = ( n32456 & n33531 ) | ( n32456 & ~n33534 ) | ( n33531 & ~n33534 ) ;
  assign n33536 = n33446 & ~n33535 ;
  assign n33537 = n9021 & n33436 ;
  assign n33538 = n9024 & ~n33423 ;
  assign n33539 = n33537 | n33538 ;
  assign n33540 = n9475 & n33526 ;
  assign n33541 = n8970 | n33540 ;
  assign n33542 = n33539 | n33541 ;
  assign n33543 = n33539 | n33540 ;
  assign n33544 = ~n33527 & n33534 ;
  assign n33545 = ~n33528 & n33544 ;
  assign n33546 = n33543 | n33545 ;
  assign n33547 = n33527 | n33530 ;
  assign n33548 = n33528 | n33547 ;
  assign n33549 = ~n33543 & n33548 ;
  assign n33550 = ( n32456 & ~n33546 ) | ( n32456 & n33549 ) | ( ~n33546 & n33549 ) ;
  assign n33551 = n33542 & ~n33550 ;
  assign n33552 = ( n33536 & n33542 ) | ( n33536 & n33551 ) | ( n33542 & n33551 ) ;
  assign n33553 = x2 & n33552 ;
  assign n33554 = x2 & ~n33552 ;
  assign n33555 = ( n33552 & ~n33553 ) | ( n33552 & n33554 ) | ( ~n33553 & n33554 ) ;
  assign n33556 = ~n33208 & n33555 ;
  assign n33557 = n33208 & ~n33555 ;
  assign n33558 = n33556 | n33557 ;
  assign n33559 = ~n32508 & n33203 ;
  assign n33560 = n32508 & ~n33203 ;
  assign n33561 = n33559 | n33560 ;
  assign n33562 = ~n33439 & n33441 ;
  assign n33563 = ( n32456 & n33439 ) | ( n32456 & ~n33562 ) | ( n33439 & ~n33562 ) ;
  assign n33564 = n33437 | n33443 ;
  assign n33565 = ~n33437 & n33442 ;
  assign n33566 = ( n32456 & ~n33564 ) | ( n32456 & n33565 ) | ( ~n33564 & n33565 ) ;
  assign n33567 = n33563 & ~n33566 ;
  assign n33568 = n9021 & ~n32442 ;
  assign n33569 = n9024 & n33436 ;
  assign n33570 = n33568 | n33569 ;
  assign n33571 = n9475 & ~n33423 ;
  assign n33572 = n8970 | n33571 ;
  assign n33573 = n33570 | n33572 ;
  assign n33574 = n33570 | n33571 ;
  assign n33575 = ~n33438 & n33444 ;
  assign n33576 = n33574 | n33575 ;
  assign n33577 = n33438 | n33445 ;
  assign n33578 = ~n33574 & n33577 ;
  assign n33579 = ( n32456 & ~n33576 ) | ( n32456 & n33578 ) | ( ~n33576 & n33578 ) ;
  assign n33580 = n33573 & ~n33579 ;
  assign n33581 = ( n33567 & n33573 ) | ( n33567 & n33580 ) | ( n33573 & n33580 ) ;
  assign n33582 = x2 & n33581 ;
  assign n33583 = x2 & ~n33581 ;
  assign n33584 = ( n33581 & ~n33582 ) | ( n33581 & n33583 ) | ( ~n33582 & n33583 ) ;
  assign n33585 = ~n33561 & n33584 ;
  assign n33586 = ~n33558 & n33585 ;
  assign n33587 = n33561 | n33585 ;
  assign n33588 = n33561 & n33584 ;
  assign n33589 = n33587 & ~n33588 ;
  assign n33590 = n32538 & ~n33201 ;
  assign n33592 = n9021 & n32306 ;
  assign n33593 = n9024 & n32293 ;
  assign n33594 = n33592 | n33593 ;
  assign n33591 = n9475 & ~n32442 ;
  assign n33596 = n8970 | n33591 ;
  assign n33597 = n33594 | n33596 ;
  assign n33595 = n33591 | n33594 ;
  assign n33598 = n33595 & n33597 ;
  assign n33599 = ( ~n32458 & n33597 ) | ( ~n32458 & n33598 ) | ( n33597 & n33598 ) ;
  assign n33600 = ~x2 & n33598 ;
  assign n33601 = ~x2 & n33597 ;
  assign n33602 = ( ~n32458 & n33600 ) | ( ~n32458 & n33601 ) | ( n33600 & n33601 ) ;
  assign n33603 = x2 | n33600 ;
  assign n33604 = x2 | n33601 ;
  assign n33605 = ( ~n32458 & n33603 ) | ( ~n32458 & n33604 ) | ( n33603 & n33604 ) ;
  assign n33606 = ( ~n33599 & n33602 ) | ( ~n33599 & n33605 ) | ( n33602 & n33605 ) ;
  assign n33607 = n9021 & ~n30186 ;
  assign n33608 = n9024 & ~n31309 ;
  assign n33609 = n33607 | n33608 ;
  assign n33610 = n9475 & ~n31323 ;
  assign n33611 = n8970 | n33610 ;
  assign n33612 = n33609 | n33611 ;
  assign n33613 = n33609 | n33610 ;
  assign n33614 = n31384 | n33613 ;
  assign n33615 = n31386 | n33613 ;
  assign n33616 = ( ~n30232 & n33614 ) | ( ~n30232 & n33615 ) | ( n33614 & n33615 ) ;
  assign n33617 = n33612 & n33616 ;
  assign n33618 = ( ~n31376 & n33612 ) | ( ~n31376 & n33617 ) | ( n33612 & n33617 ) ;
  assign n33619 = x2 & n33618 ;
  assign n33620 = x2 & ~n33618 ;
  assign n33621 = ( n33618 & ~n33619 ) | ( n33618 & n33620 ) | ( ~n33619 & n33620 ) ;
  assign n33623 = n9021 & n30212 ;
  assign n33624 = n9024 & ~n30186 ;
  assign n33625 = n33623 | n33624 ;
  assign n33622 = n9475 & ~n31309 ;
  assign n33627 = n8970 | n33622 ;
  assign n33628 = n33625 | n33627 ;
  assign n33626 = n33622 | n33625 ;
  assign n33629 = n33626 & n33628 ;
  assign n33630 = ( n31404 & n33628 ) | ( n31404 & n33629 ) | ( n33628 & n33629 ) ;
  assign n33631 = x2 & n33629 ;
  assign n33632 = x2 & n33628 ;
  assign n33633 = ( n31404 & n33631 ) | ( n31404 & n33632 ) | ( n33631 & n33632 ) ;
  assign n33634 = x2 & ~n33631 ;
  assign n33635 = x2 & ~n33632 ;
  assign n33636 = ( ~n31404 & n33634 ) | ( ~n31404 & n33635 ) | ( n33634 & n33635 ) ;
  assign n33637 = ( n33630 & ~n33633 ) | ( n33630 & n33636 ) | ( ~n33633 & n33636 ) ;
  assign n33639 = n9021 & ~n30199 ;
  assign n33640 = n9024 & n30212 ;
  assign n33641 = n33639 | n33640 ;
  assign n33638 = n9475 & ~n30186 ;
  assign n33643 = n8970 | n33638 ;
  assign n33644 = n33641 | n33643 ;
  assign n33642 = n33638 | n33641 ;
  assign n33645 = n33642 & n33644 ;
  assign n33646 = ( ~n30241 & n33644 ) | ( ~n30241 & n33645 ) | ( n33644 & n33645 ) ;
  assign n33647 = ~x2 & n33645 ;
  assign n33648 = ~x2 & n33644 ;
  assign n33649 = ( ~n30241 & n33647 ) | ( ~n30241 & n33648 ) | ( n33647 & n33648 ) ;
  assign n33650 = x2 | n33647 ;
  assign n33651 = x2 | n33648 ;
  assign n33652 = ( ~n30241 & n33650 ) | ( ~n30241 & n33651 ) | ( n33650 & n33651 ) ;
  assign n33653 = ( ~n33646 & n33649 ) | ( ~n33646 & n33652 ) | ( n33649 & n33652 ) ;
  assign n33654 = n32741 | n33144 ;
  assign n33655 = ~n33145 & n33654 ;
  assign n33656 = n9475 & n28492 ;
  assign n33657 = n9021 & ~n27606 ;
  assign n33658 = ~n27597 & n33657 ;
  assign n33659 = n9024 & ~n28503 ;
  assign n33660 = n28498 & n33659 ;
  assign n33661 = n33658 | n33660 ;
  assign n33662 = n33656 | n33661 ;
  assign n33663 = n8970 | n33662 ;
  assign n33664 = n33662 & n33663 ;
  assign n33665 = ( ~n28749 & n33663 ) | ( ~n28749 & n33664 ) | ( n33663 & n33664 ) ;
  assign n33666 = ~x2 & n33664 ;
  assign n33667 = ~x2 & n33663 ;
  assign n33668 = ( ~n28749 & n33666 ) | ( ~n28749 & n33667 ) | ( n33666 & n33667 ) ;
  assign n33669 = x2 | n33666 ;
  assign n33670 = x2 | n33667 ;
  assign n33671 = ( ~n28749 & n33669 ) | ( ~n28749 & n33670 ) | ( n33669 & n33670 ) ;
  assign n33672 = ( ~n33665 & n33668 ) | ( ~n33665 & n33671 ) | ( n33668 & n33671 ) ;
  assign n33673 = n9021 & ~n27371 ;
  assign n33674 = ~n27363 & n33673 ;
  assign n33675 = n9024 & ~n27606 ;
  assign n33676 = ~n27597 & n33675 ;
  assign n33677 = n33674 | n33676 ;
  assign n33678 = n9475 & ~n28503 ;
  assign n33679 = n28498 & n33678 ;
  assign n33680 = n33677 | n33679 ;
  assign n33681 = n28794 | n33680 ;
  assign n33682 = n28783 | n33681 ;
  assign n33683 = n8970 | n33679 ;
  assign n33684 = n33677 | n33683 ;
  assign n33685 = n33682 & n33684 ;
  assign n33686 = ~x2 & n33684 ;
  assign n33687 = n33682 & n33686 ;
  assign n33688 = x2 | n33686 ;
  assign n33689 = ( x2 & n33682 ) | ( x2 & n33688 ) | ( n33682 & n33688 ) ;
  assign n33690 = ( ~n33685 & n33687 ) | ( ~n33685 & n33689 ) | ( n33687 & n33689 ) ;
  assign n33691 = n32848 | n33130 ;
  assign n33692 = n32848 & ~n33130 ;
  assign n33693 = ( ~n32848 & n33691 ) | ( ~n32848 & n33692 ) | ( n33691 & n33692 ) ;
  assign n33694 = n9021 & n26017 ;
  assign n33695 = n9024 & ~n26270 ;
  assign n33696 = ~n26263 & n33695 ;
  assign n33697 = n33694 | n33696 ;
  assign n33698 = n9475 & ~n26526 ;
  assign n33699 = ~n26520 & n33698 ;
  assign n33701 = n8970 | n33699 ;
  assign n33702 = n33697 | n33701 ;
  assign n33700 = n33697 | n33699 ;
  assign n33703 = n33700 & n33702 ;
  assign n33704 = ( ~n26555 & n33702 ) | ( ~n26555 & n33703 ) | ( n33702 & n33703 ) ;
  assign n33705 = ( n26528 & n33702 ) | ( n26528 & n33703 ) | ( n33702 & n33703 ) ;
  assign n33706 = ( ~n26543 & n33704 ) | ( ~n26543 & n33705 ) | ( n33704 & n33705 ) ;
  assign n33707 = ~x2 & n33706 ;
  assign n33708 = x2 | n33706 ;
  assign n33709 = ( ~n33706 & n33707 ) | ( ~n33706 & n33708 ) | ( n33707 & n33708 ) ;
  assign n33710 = n9021 & ~n25728 ;
  assign n33711 = n9024 & n26017 ;
  assign n33712 = n33710 | n33711 ;
  assign n33713 = n9475 & ~n26270 ;
  assign n33714 = ~n26263 & n33713 ;
  assign n33716 = n8970 | n33714 ;
  assign n33717 = n33712 | n33716 ;
  assign n33715 = n33712 | n33714 ;
  assign n33718 = n33715 & n33717 ;
  assign n33719 = ( n26571 & n33717 ) | ( n26571 & n33718 ) | ( n33717 & n33718 ) ;
  assign n33720 = x2 & n33718 ;
  assign n33721 = x2 & n33717 ;
  assign n33722 = ( n26571 & n33720 ) | ( n26571 & n33721 ) | ( n33720 & n33721 ) ;
  assign n33723 = x2 & ~n33720 ;
  assign n33724 = x2 & ~n33721 ;
  assign n33725 = ( ~n26571 & n33723 ) | ( ~n26571 & n33724 ) | ( n33723 & n33724 ) ;
  assign n33726 = ( n33719 & ~n33722 ) | ( n33719 & n33725 ) | ( ~n33722 & n33725 ) ;
  assign n33727 = n9475 & n26017 ;
  assign n33728 = n9021 & ~n25046 ;
  assign n33729 = n9024 & ~n25728 ;
  assign n33730 = n33728 | n33729 ;
  assign n33731 = n33727 | n33730 ;
  assign n33732 = n8970 | n33727 ;
  assign n33733 = n33730 | n33732 ;
  assign n33734 = ( n26613 & n33731 ) | ( n26613 & n33733 ) | ( n33731 & n33733 ) ;
  assign n33735 = n33731 | n33733 ;
  assign n33736 = ( n26605 & n33734 ) | ( n26605 & n33735 ) | ( n33734 & n33735 ) ;
  assign n33737 = x2 & n33736 ;
  assign n33738 = x2 & ~n33736 ;
  assign n33739 = ( n33736 & ~n33737 ) | ( n33736 & n33738 ) | ( ~n33737 & n33738 ) ;
  assign n33740 = n32972 | n33115 ;
  assign n33741 = ~n33116 & n33740 ;
  assign n33742 = n32994 | n33088 ;
  assign n33743 = ~n33089 & n33742 ;
  assign n33744 = n33082 & n33084 ;
  assign n33745 = n33082 | n33084 ;
  assign n33746 = ~n33744 & n33745 ;
  assign n33747 = n9021 & ~n22385 ;
  assign n33748 = ( n9024 & n9994 ) | ( n9024 & ~n22385 ) | ( n9994 & ~n22385 ) ;
  assign n33749 = ( n22381 & n33747 ) | ( n22381 & n33748 ) | ( n33747 & n33748 ) ;
  assign n33750 = n9475 | n33749 ;
  assign n33751 = ( n23620 & n33749 ) | ( n23620 & n33750 ) | ( n33749 & n33750 ) ;
  assign n33752 = n8970 | n33751 ;
  assign n33753 = ( ~n23686 & n33751 ) | ( ~n23686 & n33752 ) | ( n33751 & n33752 ) ;
  assign n33754 = ~x2 & n33752 ;
  assign n33755 = ~x2 & n33751 ;
  assign n33756 = ( ~n23686 & n33754 ) | ( ~n23686 & n33755 ) | ( n33754 & n33755 ) ;
  assign n33757 = x2 | n33754 ;
  assign n33758 = x2 | n33755 ;
  assign n33759 = ( ~n23686 & n33757 ) | ( ~n23686 & n33758 ) | ( n33757 & n33758 ) ;
  assign n33760 = ( ~n33753 & n33756 ) | ( ~n33753 & n33759 ) | ( n33756 & n33759 ) ;
  assign n33761 = n33045 & n33063 ;
  assign n33762 = n33045 | n33063 ;
  assign n33763 = ~n33761 & n33762 ;
  assign n33764 = n8113 & ~n22409 ;
  assign n33765 = n9633 & n22474 ;
  assign n33766 = n9644 & ~n22409 ;
  assign n33767 = ( x2 & n9640 ) | ( x2 & n22406 ) | ( n9640 & n22406 ) ;
  assign n33768 = ~n33766 & n33767 ;
  assign n33769 = ~n33765 & n33768 ;
  assign n33770 = n9021 & ~n22409 ;
  assign n33771 = n9024 & ~n22406 ;
  assign n33772 = n33770 | n33771 ;
  assign n33773 = n21756 & n22393 ;
  assign n33774 = ( x2 & n33772 ) | ( x2 & n33773 ) | ( n33772 & n33773 ) ;
  assign n33775 = n33769 & ~n33774 ;
  assign n33776 = n9660 & ~n22409 ;
  assign n33777 = n9633 | n33776 ;
  assign n33778 = ( n22439 & n33776 ) | ( n22439 & n33777 ) | ( n33776 & n33777 ) ;
  assign n33779 = n33775 & ~n33778 ;
  assign n33780 = n9475 & ~n22398 ;
  assign n33781 = n9021 & ~n22406 ;
  assign n33782 = n9024 & n22393 ;
  assign n33783 = n33781 | n33782 ;
  assign n33784 = n33780 | n33783 ;
  assign n33785 = n8970 | n33780 ;
  assign n33786 = n33783 | n33785 ;
  assign n33787 = ( n22608 & n33784 ) | ( n22608 & n33786 ) | ( n33784 & n33786 ) ;
  assign n33788 = x2 & n33786 ;
  assign n33789 = x2 & n33784 ;
  assign n33790 = ( n22608 & n33788 ) | ( n22608 & n33789 ) | ( n33788 & n33789 ) ;
  assign n33791 = x2 & ~n33790 ;
  assign n33792 = ( n33787 & ~n33790 ) | ( n33787 & n33791 ) | ( ~n33790 & n33791 ) ;
  assign n33793 = ( n33764 & n33779 ) | ( n33764 & n33792 ) | ( n33779 & n33792 ) ;
  assign n33794 = n9475 & ~n22385 ;
  assign n33795 = n9021 & n22393 ;
  assign n33796 = n9024 & ~n22398 ;
  assign n33797 = n33795 | n33796 ;
  assign n33798 = n33794 | n33797 ;
  assign n33799 = n8970 | n33794 ;
  assign n33800 = n33797 | n33799 ;
  assign n33801 = ( ~n22545 & n33798 ) | ( ~n22545 & n33800 ) | ( n33798 & n33800 ) ;
  assign n33802 = ~x2 & n33800 ;
  assign n33803 = ~x2 & n33798 ;
  assign n33804 = ( ~n22545 & n33802 ) | ( ~n22545 & n33803 ) | ( n33802 & n33803 ) ;
  assign n33805 = x2 | n33803 ;
  assign n33806 = x2 | n33802 ;
  assign n33807 = ( ~n22545 & n33805 ) | ( ~n22545 & n33806 ) | ( n33805 & n33806 ) ;
  assign n33808 = ( ~n33801 & n33804 ) | ( ~n33801 & n33807 ) | ( n33804 & n33807 ) ;
  assign n33809 = n33793 & n33808 ;
  assign n33810 = n33763 & n33809 ;
  assign n33811 = n33039 | n33041 ;
  assign n33812 = ~n33041 & n33043 ;
  assign n33813 = ( n33040 & n33811 ) | ( n33040 & ~n33812 ) | ( n33811 & ~n33812 ) ;
  assign n33814 = ~n33045 & n33813 ;
  assign n33815 = n33808 & n33814 ;
  assign n33816 = ( n33793 & n33814 ) | ( n33793 & n33815 ) | ( n33814 & n33815 ) ;
  assign n33817 = ( n33763 & n33810 ) | ( n33763 & n33816 ) | ( n33810 & n33816 ) ;
  assign n33818 = n33760 & n33817 ;
  assign n33819 = n33763 | n33809 ;
  assign n33820 = n9475 & n22381 ;
  assign n33821 = n9021 & ~n22398 ;
  assign n33822 = n9024 & ~n22385 ;
  assign n33823 = n33821 | n33822 ;
  assign n33824 = n33820 | n33823 ;
  assign n33825 = n8970 | n33824 ;
  assign n33826 = ( n22422 & n33824 ) | ( n22422 & n33825 ) | ( n33824 & n33825 ) ;
  assign n33827 = x2 & n33825 ;
  assign n33828 = x2 & n33824 ;
  assign n33829 = ( n22422 & n33827 ) | ( n22422 & n33828 ) | ( n33827 & n33828 ) ;
  assign n33830 = x2 & ~n33827 ;
  assign n33831 = x2 & ~n33828 ;
  assign n33832 = ( ~n22422 & n33830 ) | ( ~n22422 & n33831 ) | ( n33830 & n33831 ) ;
  assign n33833 = ( n33826 & ~n33829 ) | ( n33826 & n33832 ) | ( ~n33829 & n33832 ) ;
  assign n33834 = n33816 & n33833 ;
  assign n33835 = ( n33819 & n33833 ) | ( n33819 & n33834 ) | ( n33833 & n33834 ) ;
  assign n33836 = ( n33760 & n33818 ) | ( n33760 & n33835 ) | ( n33818 & n33835 ) ;
  assign n33837 = n33746 | n33836 ;
  assign n33838 = n33066 & ~n33080 ;
  assign n33839 = n33760 | n33817 ;
  assign n33840 = ( n33080 & n33835 ) | ( n33080 & n33838 ) | ( n33835 & n33838 ) ;
  assign n33841 = n33080 | n33838 ;
  assign n33842 = ( n33839 & n33840 ) | ( n33839 & n33841 ) | ( n33840 & n33841 ) ;
  assign n33843 = ( ~n33066 & n33838 ) | ( ~n33066 & n33842 ) | ( n33838 & n33842 ) ;
  assign n33844 = n33837 | n33843 ;
  assign n33845 = n9021 & n22381 ;
  assign n33846 = ( n9024 & n9994 ) | ( n9024 & n22381 ) | ( n9994 & n22381 ) ;
  assign n33847 = ( n23620 & n33845 ) | ( n23620 & n33846 ) | ( n33845 & n33846 ) ;
  assign n33848 = n9475 | n33846 ;
  assign n33849 = n9475 | n33845 ;
  assign n33850 = ( n23620 & n33848 ) | ( n23620 & n33849 ) | ( n33848 & n33849 ) ;
  assign n33851 = ( n23316 & n33847 ) | ( n23316 & n33850 ) | ( n33847 & n33850 ) ;
  assign n33852 = n8970 | n33851 ;
  assign n33853 = ( n23661 & n33851 ) | ( n23661 & n33852 ) | ( n33851 & n33852 ) ;
  assign n33854 = x2 & n33852 ;
  assign n33855 = x2 & n33851 ;
  assign n33856 = ( n23661 & n33854 ) | ( n23661 & n33855 ) | ( n33854 & n33855 ) ;
  assign n33857 = x2 & ~n33854 ;
  assign n33858 = x2 & ~n33855 ;
  assign n33859 = ( ~n23661 & n33857 ) | ( ~n23661 & n33858 ) | ( n33857 & n33858 ) ;
  assign n33860 = ( n33853 & ~n33856 ) | ( n33853 & n33859 ) | ( ~n33856 & n33859 ) ;
  assign n33861 = n33844 & n33860 ;
  assign n33862 = n9475 & n23614 ;
  assign n33863 = n9021 & n23620 ;
  assign n33864 = ( n9024 & n9994 ) | ( n9024 & n23620 ) | ( n9994 & n23620 ) ;
  assign n33865 = ( n23316 & n33863 ) | ( n23316 & n33864 ) | ( n33863 & n33864 ) ;
  assign n33867 = n8970 | n33865 ;
  assign n33868 = n33862 | n33867 ;
  assign n33866 = n33862 | n33865 ;
  assign n33869 = n33866 & n33868 ;
  assign n33870 = ( n23634 & n33868 ) | ( n23634 & n33869 ) | ( n33868 & n33869 ) ;
  assign n33871 = x2 & n33869 ;
  assign n33872 = x2 & n33868 ;
  assign n33873 = ( n23634 & n33871 ) | ( n23634 & n33872 ) | ( n33871 & n33872 ) ;
  assign n33874 = x2 & ~n33871 ;
  assign n33875 = x2 & ~n33872 ;
  assign n33876 = ( ~n23634 & n33874 ) | ( ~n23634 & n33875 ) | ( n33874 & n33875 ) ;
  assign n33877 = ( n33870 & ~n33873 ) | ( n33870 & n33876 ) | ( ~n33873 & n33876 ) ;
  assign n33878 = n33746 & n33836 ;
  assign n33879 = ( n33746 & n33843 ) | ( n33746 & n33878 ) | ( n33843 & n33878 ) ;
  assign n33880 = n33877 & n33879 ;
  assign n33881 = ( n33861 & n33877 ) | ( n33861 & n33880 ) | ( n33877 & n33880 ) ;
  assign n33882 = n9475 & n24167 ;
  assign n33883 = n9021 & n23316 ;
  assign n33884 = n9024 & n23614 ;
  assign n33885 = n33883 | n33884 ;
  assign n33886 = n33882 | n33885 ;
  assign n33887 = n8970 | n33886 ;
  assign n33888 = ( n24182 & n33886 ) | ( n24182 & n33887 ) | ( n33886 & n33887 ) ;
  assign n33889 = n33886 | n33887 ;
  assign n33890 = ( n24175 & n33888 ) | ( n24175 & n33889 ) | ( n33888 & n33889 ) ;
  assign n33891 = x2 & n33890 ;
  assign n33892 = x2 & ~n33890 ;
  assign n33893 = ( n33890 & ~n33891 ) | ( n33890 & n33892 ) | ( ~n33891 & n33892 ) ;
  assign n33894 = n33881 | n33893 ;
  assign n33895 = n33013 & ~n33086 ;
  assign n33896 = n33877 | n33879 ;
  assign n33897 = n33861 | n33896 ;
  assign n33898 = ( ~n33013 & n33086 ) | ( ~n33013 & n33895 ) | ( n33086 & n33895 ) ;
  assign n33899 = ( n33895 & n33897 ) | ( n33895 & n33898 ) | ( n33897 & n33898 ) ;
  assign n33900 = n33894 | n33899 ;
  assign n33901 = n33743 & n33900 ;
  assign n33902 = n9475 & ~n25054 ;
  assign n33903 = n9021 & n23614 ;
  assign n33904 = n9024 & n24167 ;
  assign n33905 = n33903 | n33904 ;
  assign n33906 = n33902 | n33905 ;
  assign n33907 = n8970 | n33902 ;
  assign n33908 = n33905 | n33907 ;
  assign n33909 = ( ~n25122 & n33906 ) | ( ~n25122 & n33908 ) | ( n33906 & n33908 ) ;
  assign n33910 = ~x2 & n33908 ;
  assign n33911 = ~x2 & n33906 ;
  assign n33912 = ( ~n25122 & n33910 ) | ( ~n25122 & n33911 ) | ( n33910 & n33911 ) ;
  assign n33913 = x2 | n33911 ;
  assign n33914 = x2 | n33910 ;
  assign n33915 = ( ~n25122 & n33913 ) | ( ~n25122 & n33914 ) | ( n33913 & n33914 ) ;
  assign n33916 = ( ~n33909 & n33912 ) | ( ~n33909 & n33915 ) | ( n33912 & n33915 ) ;
  assign n33917 = n33881 & n33893 ;
  assign n33918 = ( n33893 & n33899 ) | ( n33893 & n33917 ) | ( n33899 & n33917 ) ;
  assign n33919 = n33916 & n33918 ;
  assign n33920 = ( n33901 & n33916 ) | ( n33901 & n33919 ) | ( n33916 & n33919 ) ;
  assign n33921 = n33741 | n33920 ;
  assign n33922 = n33916 | n33918 ;
  assign n33923 = n33901 | n33922 ;
  assign n33924 = n33090 & n33113 ;
  assign n33925 = n33090 & ~n33924 ;
  assign n33926 = n33113 & ~n33924 ;
  assign n33927 = ( n33923 & n33925 ) | ( n33923 & n33926 ) | ( n33925 & n33926 ) ;
  assign n33928 = n33921 | n33927 ;
  assign n33929 = n9475 & n24770 ;
  assign n33930 = n9021 & n24167 ;
  assign n33931 = n9024 & ~n25054 ;
  assign n33932 = n33930 | n33931 ;
  assign n33933 = n33929 | n33932 ;
  assign n33934 = n8970 | n33933 ;
  assign n33935 = ( ~n25095 & n33933 ) | ( ~n25095 & n33934 ) | ( n33933 & n33934 ) ;
  assign n33936 = ~x2 & n33934 ;
  assign n33937 = ~x2 & n33933 ;
  assign n33938 = ( ~n25095 & n33936 ) | ( ~n25095 & n33937 ) | ( n33936 & n33937 ) ;
  assign n33939 = x2 | n33936 ;
  assign n33940 = x2 | n33937 ;
  assign n33941 = ( ~n25095 & n33939 ) | ( ~n25095 & n33940 ) | ( n33939 & n33940 ) ;
  assign n33942 = ( ~n33935 & n33938 ) | ( ~n33935 & n33941 ) | ( n33938 & n33941 ) ;
  assign n33943 = n33928 & n33942 ;
  assign n33944 = n33117 | n33119 ;
  assign n33945 = ~n33120 & n33944 ;
  assign n33946 = n33741 & n33920 ;
  assign n33947 = ( n33741 & n33927 ) | ( n33741 & n33946 ) | ( n33927 & n33946 ) ;
  assign n33948 = n33945 | n33947 ;
  assign n33949 = n33943 | n33948 ;
  assign n33950 = n9475 & ~n25046 ;
  assign n33951 = n9021 & ~n25054 ;
  assign n33952 = n9024 & n24770 ;
  assign n33953 = n33951 | n33952 ;
  assign n33954 = n33950 | n33953 ;
  assign n33955 = n8970 | n33950 ;
  assign n33956 = n33953 | n33955 ;
  assign n33957 = ( ~n25069 & n33954 ) | ( ~n25069 & n33956 ) | ( n33954 & n33956 ) ;
  assign n33958 = ~x2 & n33956 ;
  assign n33959 = ~x2 & n33954 ;
  assign n33960 = ( ~n25069 & n33958 ) | ( ~n25069 & n33959 ) | ( n33958 & n33959 ) ;
  assign n33961 = x2 | n33959 ;
  assign n33962 = x2 | n33958 ;
  assign n33963 = ( ~n25069 & n33961 ) | ( ~n25069 & n33962 ) | ( n33961 & n33962 ) ;
  assign n33964 = ( ~n33957 & n33960 ) | ( ~n33957 & n33963 ) | ( n33960 & n33963 ) ;
  assign n33965 = n33949 & n33964 ;
  assign n33966 = ( n32948 & n32949 ) | ( n32948 & n33120 ) | ( n32949 & n33120 ) ;
  assign n33967 = n32927 | n32948 ;
  assign n33968 = n33120 | n33967 ;
  assign n33969 = ~n33966 & n33968 ;
  assign n33970 = n33945 & n33947 ;
  assign n33971 = ( n33943 & n33945 ) | ( n33943 & n33970 ) | ( n33945 & n33970 ) ;
  assign n33972 = n33969 & n33971 ;
  assign n33973 = ( n33965 & n33969 ) | ( n33965 & n33972 ) | ( n33969 & n33972 ) ;
  assign n33974 = n33739 & n33973 ;
  assign n33975 = n33969 | n33971 ;
  assign n33976 = n33965 | n33975 ;
  assign n33977 = n9475 & ~n25728 ;
  assign n33978 = n9021 & n24770 ;
  assign n33979 = n9024 & ~n25046 ;
  assign n33980 = n33978 | n33979 ;
  assign n33981 = n33977 | n33980 ;
  assign n33982 = n8970 & n25740 ;
  assign n33983 = n8970 & n25731 ;
  assign n33984 = ( ~n25441 & n33982 ) | ( ~n25441 & n33983 ) | ( n33982 & n33983 ) ;
  assign n33985 = n33981 | n33984 ;
  assign n33986 = n8970 | n33981 ;
  assign n33987 = ( n25733 & n33985 ) | ( n25733 & n33986 ) | ( n33985 & n33986 ) ;
  assign n33988 = x2 & n33987 ;
  assign n33989 = n33987 & ~n33988 ;
  assign n33990 = x2 & ~n33988 ;
  assign n33991 = ( n33976 & n33989 ) | ( n33976 & n33990 ) | ( n33989 & n33990 ) ;
  assign n33992 = ( n33739 & n33974 ) | ( n33739 & n33991 ) | ( n33974 & n33991 ) ;
  assign n33993 = n33726 & n33992 ;
  assign n33994 = n32912 & ~n33122 ;
  assign n33995 = n33739 | n33973 ;
  assign n33996 = n33991 | n33995 ;
  assign n33997 = ( ~n32912 & n33122 ) | ( ~n32912 & n33994 ) | ( n33122 & n33994 ) ;
  assign n33998 = ( n33994 & n33996 ) | ( n33994 & n33997 ) | ( n33996 & n33997 ) ;
  assign n33999 = ( n33726 & n33993 ) | ( n33726 & n33998 ) | ( n33993 & n33998 ) ;
  assign n34000 = n33709 & n33999 ;
  assign n34001 = n32891 & ~n33124 ;
  assign n34002 = n33726 | n33992 ;
  assign n34003 = n33998 | n34002 ;
  assign n34004 = ( ~n32891 & n33124 ) | ( ~n32891 & n34001 ) | ( n33124 & n34001 ) ;
  assign n34005 = ( n34001 & n34003 ) | ( n34001 & n34004 ) | ( n34003 & n34004 ) ;
  assign n34006 = ( n33709 & n34000 ) | ( n33709 & n34005 ) | ( n34000 & n34005 ) ;
  assign n34007 = n33693 & n34006 ;
  assign n34008 = n33126 & ~n33128 ;
  assign n34009 = n33709 | n33999 ;
  assign n34010 = n34005 | n34009 ;
  assign n34011 = ( ~n33126 & n33128 ) | ( ~n33126 & n34008 ) | ( n33128 & n34008 ) ;
  assign n34012 = ( n34008 & n34010 ) | ( n34008 & n34011 ) | ( n34010 & n34011 ) ;
  assign n34013 = ( n33693 & n34007 ) | ( n33693 & n34012 ) | ( n34007 & n34012 ) ;
  assign n34014 = n32828 | n33132 ;
  assign n34015 = ~n33132 & n34014 ;
  assign n34016 = ( ~n32828 & n34014 ) | ( ~n32828 & n34015 ) | ( n34014 & n34015 ) ;
  assign n34017 = n34013 | n34016 ;
  assign n34018 = n33693 | n34006 ;
  assign n34019 = n34012 | n34018 ;
  assign n34020 = n8970 & n27699 ;
  assign n34021 = ( n8970 & ~n27696 ) | ( n8970 & n34020 ) | ( ~n27696 & n34020 ) ;
  assign n34022 = n9021 & ~n26270 ;
  assign n34023 = ~n26263 & n34022 ;
  assign n34024 = n9024 & ~n26526 ;
  assign n34025 = ~n26520 & n34024 ;
  assign n34026 = n34023 | n34025 ;
  assign n34027 = n9475 & ~n27133 ;
  assign n34028 = ~n27125 & n34027 ;
  assign n34029 = n34026 | n34028 ;
  assign n34030 = n34021 | n34029 ;
  assign n34031 = x2 & n34029 ;
  assign n34032 = ( x2 & n34021 ) | ( x2 & n34031 ) | ( n34021 & n34031 ) ;
  assign n34033 = n34030 & ~n34032 ;
  assign n34034 = x2 & ~n34032 ;
  assign n34035 = ( n34019 & n34033 ) | ( n34019 & n34034 ) | ( n34033 & n34034 ) ;
  assign n34036 = n34017 | n34035 ;
  assign n34037 = n9021 & ~n26526 ;
  assign n34038 = ~n26520 & n34037 ;
  assign n34039 = n9024 & ~n27133 ;
  assign n34040 = ~n27125 & n34039 ;
  assign n34041 = n34038 | n34040 ;
  assign n34042 = n9475 & ~n27371 ;
  assign n34043 = ~n27363 & n34042 ;
  assign n34044 = n34041 | n34043 ;
  assign n34045 = n8970 | n34043 ;
  assign n34046 = n34041 | n34045 ;
  assign n34047 = ( ~n27654 & n34044 ) | ( ~n27654 & n34046 ) | ( n34044 & n34046 ) ;
  assign n34048 = ~x2 & n34046 ;
  assign n34049 = ~x2 & n34044 ;
  assign n34050 = ( ~n27654 & n34048 ) | ( ~n27654 & n34049 ) | ( n34048 & n34049 ) ;
  assign n34051 = x2 | n34049 ;
  assign n34052 = x2 | n34048 ;
  assign n34053 = ( ~n27654 & n34051 ) | ( ~n27654 & n34052 ) | ( n34051 & n34052 ) ;
  assign n34054 = ( ~n34047 & n34050 ) | ( ~n34047 & n34053 ) | ( n34050 & n34053 ) ;
  assign n34055 = n34036 & n34054 ;
  assign n34056 = n33134 & n33136 ;
  assign n34057 = n33134 | n33136 ;
  assign n34058 = ~n34056 & n34057 ;
  assign n34059 = n34013 & n34016 ;
  assign n34060 = ( n34016 & n34035 ) | ( n34016 & n34059 ) | ( n34035 & n34059 ) ;
  assign n34061 = n34058 & n34060 ;
  assign n34062 = ( n34055 & n34058 ) | ( n34055 & n34061 ) | ( n34058 & n34061 ) ;
  assign n34063 = n33690 & n34062 ;
  assign n34064 = n34058 | n34060 ;
  assign n34065 = n34055 | n34064 ;
  assign n34066 = n8970 & n27630 ;
  assign n34067 = ~n27625 & n34066 ;
  assign n34068 = ( n8970 & ~n27634 ) | ( n8970 & n34067 ) | ( ~n27634 & n34067 ) ;
  assign n34069 = n9021 & ~n27133 ;
  assign n34070 = ~n27125 & n34069 ;
  assign n34071 = n9024 & ~n27371 ;
  assign n34072 = ~n27363 & n34071 ;
  assign n34073 = n34070 | n34072 ;
  assign n34074 = n9475 & ~n27606 ;
  assign n34075 = ~n27597 & n34074 ;
  assign n34076 = n34073 | n34075 ;
  assign n34077 = n34068 | n34076 ;
  assign n34078 = x2 & n34076 ;
  assign n34079 = ( x2 & n34068 ) | ( x2 & n34078 ) | ( n34068 & n34078 ) ;
  assign n34080 = n34077 & ~n34079 ;
  assign n34081 = x2 & ~n34079 ;
  assign n34082 = ( n34065 & n34080 ) | ( n34065 & n34081 ) | ( n34080 & n34081 ) ;
  assign n34083 = ( n33690 & n34063 ) | ( n33690 & n34082 ) | ( n34063 & n34082 ) ;
  assign n34084 = n33672 & n34083 ;
  assign n34085 = n32785 & ~n33138 ;
  assign n34086 = n33690 | n34062 ;
  assign n34087 = n34082 | n34086 ;
  assign n34088 = ( ~n32785 & n33138 ) | ( ~n32785 & n34085 ) | ( n33138 & n34085 ) ;
  assign n34089 = ( n34085 & n34087 ) | ( n34085 & n34088 ) | ( n34087 & n34088 ) ;
  assign n34090 = ( n33672 & n34084 ) | ( n33672 & n34089 ) | ( n34084 & n34089 ) ;
  assign n34091 = n9024 & n28492 ;
  assign n34092 = n9021 & ~n28503 ;
  assign n34093 = n28498 & n34092 ;
  assign n34094 = n34091 | n34093 ;
  assign n34095 = n9475 & ~n28714 ;
  assign n34096 = n8970 | n34095 ;
  assign n34097 = n34094 | n34096 ;
  assign n34098 = n34094 | n34095 ;
  assign n34099 = n28731 & ~n34098 ;
  assign n34100 = ( n28518 & ~n34098 ) | ( n28518 & n34099 ) | ( ~n34098 & n34099 ) ;
  assign n34101 = n34097 & ~n34100 ;
  assign n34102 = ( n28720 & n34097 ) | ( n28720 & n34101 ) | ( n34097 & n34101 ) ;
  assign n34103 = x2 & n34102 ;
  assign n34104 = x2 & ~n34102 ;
  assign n34105 = ( n34102 & ~n34103 ) | ( n34102 & n34104 ) | ( ~n34103 & n34104 ) ;
  assign n34106 = n34090 | n34105 ;
  assign n34107 = ~n33140 & n33142 ;
  assign n34108 = n33672 | n34083 ;
  assign n34109 = n34089 | n34108 ;
  assign n34110 = ( n33140 & ~n33142 ) | ( n33140 & n34107 ) | ( ~n33142 & n34107 ) ;
  assign n34111 = ( n34107 & n34109 ) | ( n34107 & n34110 ) | ( n34109 & n34110 ) ;
  assign n34112 = n34106 | n34111 ;
  assign n34113 = n33655 & n34112 ;
  assign n34114 = ( ~n33146 & n33147 ) | ( ~n33146 & n33148 ) | ( n33147 & n33148 ) ;
  assign n34115 = n33146 | n34114 ;
  assign n34116 = ~n33150 & n34115 ;
  assign n34117 = n34090 & n34105 ;
  assign n34118 = ( n34105 & n34111 ) | ( n34105 & n34117 ) | ( n34111 & n34117 ) ;
  assign n34119 = n34116 | n34118 ;
  assign n34120 = n34113 | n34119 ;
  assign n34121 = n9475 & n29620 ;
  assign n34122 = n9021 & n28492 ;
  assign n34123 = n9024 & ~n28714 ;
  assign n34124 = n34122 | n34123 ;
  assign n34125 = n34121 | n34124 ;
  assign n34126 = n8970 | n34121 ;
  assign n34127 = n34124 | n34126 ;
  assign n34128 = ( ~n29642 & n34125 ) | ( ~n29642 & n34127 ) | ( n34125 & n34127 ) ;
  assign n34129 = n34125 | n34127 ;
  assign n34130 = ( n29629 & n34128 ) | ( n29629 & n34129 ) | ( n34128 & n34129 ) ;
  assign n34131 = ~x2 & n34130 ;
  assign n34132 = x2 | n34130 ;
  assign n34133 = ( ~n34130 & n34131 ) | ( ~n34130 & n34132 ) | ( n34131 & n34132 ) ;
  assign n34134 = n34120 & n34133 ;
  assign n34135 = ( ~n33151 & n33173 ) | ( ~n33151 & n33174 ) | ( n33173 & n33174 ) ;
  assign n34136 = n33151 | n34135 ;
  assign n34137 = ~n33176 & n34136 ;
  assign n34138 = n34116 & n34118 ;
  assign n34139 = ( n34113 & n34116 ) | ( n34113 & n34138 ) | ( n34116 & n34138 ) ;
  assign n34140 = n34137 | n34139 ;
  assign n34141 = n34134 | n34140 ;
  assign n34142 = n9475 & ~n30199 ;
  assign n34143 = n9021 & ~n28714 ;
  assign n34144 = n9024 & n29620 ;
  assign n34145 = n34143 | n34144 ;
  assign n34146 = n34142 | n34145 ;
  assign n34147 = n8970 | n34142 ;
  assign n34148 = n34145 | n34147 ;
  assign n34149 = ( ~n30299 & n34146 ) | ( ~n30299 & n34148 ) | ( n34146 & n34148 ) ;
  assign n34150 = ~x2 & n34148 ;
  assign n34151 = ~x2 & n34146 ;
  assign n34152 = ( ~n30299 & n34150 ) | ( ~n30299 & n34151 ) | ( n34150 & n34151 ) ;
  assign n34153 = x2 | n34151 ;
  assign n34154 = x2 | n34150 ;
  assign n34155 = ( ~n30299 & n34153 ) | ( ~n30299 & n34154 ) | ( n34153 & n34154 ) ;
  assign n34156 = ( ~n34149 & n34152 ) | ( ~n34149 & n34155 ) | ( n34152 & n34155 ) ;
  assign n34157 = n34141 & n34156 ;
  assign n34158 = n33172 | n33178 ;
  assign n34159 = n33176 | n34158 ;
  assign n34160 = ~n33180 & n34159 ;
  assign n34161 = n34137 & n34139 ;
  assign n34162 = ( n34134 & n34137 ) | ( n34134 & n34161 ) | ( n34137 & n34161 ) ;
  assign n34163 = n34160 & n34162 ;
  assign n34164 = ( n34157 & n34160 ) | ( n34157 & n34163 ) | ( n34160 & n34163 ) ;
  assign n34165 = n33653 & n34164 ;
  assign n34166 = n34160 | n34162 ;
  assign n34167 = n34157 | n34166 ;
  assign n34168 = n8970 & ~n30266 ;
  assign n34169 = ( n8970 & n30276 ) | ( n8970 & n34168 ) | ( n30276 & n34168 ) ;
  assign n34170 = n9475 & n30212 ;
  assign n34171 = n9021 & n29620 ;
  assign n34172 = n9024 & ~n30199 ;
  assign n34173 = n34171 | n34172 ;
  assign n34174 = n34170 | n34173 ;
  assign n34175 = n34169 | n34174 ;
  assign n34176 = x2 & n34174 ;
  assign n34177 = ( x2 & n34169 ) | ( x2 & n34176 ) | ( n34169 & n34176 ) ;
  assign n34178 = n34175 & ~n34177 ;
  assign n34179 = x2 & ~n34177 ;
  assign n34180 = ( n34167 & n34178 ) | ( n34167 & n34179 ) | ( n34178 & n34179 ) ;
  assign n34181 = ( n33653 & n34165 ) | ( n33653 & n34180 ) | ( n34165 & n34180 ) ;
  assign n34182 = n33637 & n34181 ;
  assign n34183 = n32679 & ~n33181 ;
  assign n34184 = n33653 | n34164 ;
  assign n34185 = n34180 | n34184 ;
  assign n34186 = ( ~n32679 & n33181 ) | ( ~n32679 & n34183 ) | ( n33181 & n34183 ) ;
  assign n34187 = ( n34183 & n34185 ) | ( n34183 & n34186 ) | ( n34185 & n34186 ) ;
  assign n34188 = ( n33637 & n34182 ) | ( n33637 & n34187 ) | ( n34182 & n34187 ) ;
  assign n34189 = n33621 & n34188 ;
  assign n34190 = n32659 & ~n33183 ;
  assign n34191 = n33637 | n34181 ;
  assign n34192 = n34187 | n34191 ;
  assign n34193 = ( ~n32659 & n33183 ) | ( ~n32659 & n34190 ) | ( n33183 & n34190 ) ;
  assign n34194 = ( n34190 & n34192 ) | ( n34190 & n34193 ) | ( n34192 & n34193 ) ;
  assign n34195 = ( n33621 & n34189 ) | ( n33621 & n34194 ) | ( n34189 & n34194 ) ;
  assign n34196 = n32620 | n33189 ;
  assign n34197 = n32620 & ~n33189 ;
  assign n34198 = ( ~n32620 & n34196 ) | ( ~n32620 & n34197 ) | ( n34196 & n34197 ) ;
  assign n34199 = n34195 | n34198 ;
  assign n34200 = n33185 & ~n33187 ;
  assign n34201 = n33621 | n34188 ;
  assign n34202 = n34194 | n34201 ;
  assign n34203 = ( ~n33185 & n33187 ) | ( ~n33185 & n34200 ) | ( n33187 & n34200 ) ;
  assign n34204 = ( n34200 & n34202 ) | ( n34200 & n34203 ) | ( n34202 & n34203 ) ;
  assign n34205 = n34199 | n34204 ;
  assign n34206 = n9475 & n31295 ;
  assign n34207 = n9021 & ~n31309 ;
  assign n34208 = n9024 & ~n31323 ;
  assign n34209 = n34207 | n34208 ;
  assign n34210 = n34206 | n34209 ;
  assign n34211 = n8970 | n34206 ;
  assign n34212 = n34209 | n34211 ;
  assign n34213 = ( n31355 & n34210 ) | ( n31355 & n34212 ) | ( n34210 & n34212 ) ;
  assign n34214 = x2 & n34212 ;
  assign n34215 = x2 & n34210 ;
  assign n34216 = ( n31355 & n34214 ) | ( n31355 & n34215 ) | ( n34214 & n34215 ) ;
  assign n34217 = x2 & ~n34215 ;
  assign n34218 = x2 & ~n34214 ;
  assign n34219 = ( ~n31355 & n34217 ) | ( ~n31355 & n34218 ) | ( n34217 & n34218 ) ;
  assign n34220 = ( n34213 & ~n34216 ) | ( n34213 & n34219 ) | ( ~n34216 & n34219 ) ;
  assign n34221 = n34205 & n34220 ;
  assign n34222 = n33191 & n33193 ;
  assign n34223 = n33191 | n33193 ;
  assign n34224 = ~n34222 & n34223 ;
  assign n34225 = n34195 & n34198 ;
  assign n34226 = ( n34198 & n34204 ) | ( n34198 & n34225 ) | ( n34204 & n34225 ) ;
  assign n34227 = n34224 | n34226 ;
  assign n34228 = n34221 | n34227 ;
  assign n34229 = n9475 & n32306 ;
  assign n34230 = n9021 & ~n31323 ;
  assign n34231 = n9024 & n31295 ;
  assign n34232 = n34230 | n34231 ;
  assign n34233 = n34229 | n34232 ;
  assign n34234 = n8970 | n34229 ;
  assign n34235 = n34232 | n34234 ;
  assign n34236 = ( ~n32525 & n34233 ) | ( ~n32525 & n34235 ) | ( n34233 & n34235 ) ;
  assign n34237 = ~x2 & n34235 ;
  assign n34238 = ~x2 & n34233 ;
  assign n34239 = ( ~n32525 & n34237 ) | ( ~n32525 & n34238 ) | ( n34237 & n34238 ) ;
  assign n34240 = x2 | n34238 ;
  assign n34241 = x2 | n34237 ;
  assign n34242 = ( ~n32525 & n34240 ) | ( ~n32525 & n34241 ) | ( n34240 & n34241 ) ;
  assign n34243 = ( ~n34236 & n34239 ) | ( ~n34236 & n34242 ) | ( n34239 & n34242 ) ;
  assign n34244 = n34228 & n34243 ;
  assign n34245 = n9475 & n32293 ;
  assign n34246 = n9021 & n31295 ;
  assign n34247 = n9024 & n32306 ;
  assign n34248 = n34246 | n34247 ;
  assign n34249 = n34245 | n34248 ;
  assign n34250 = n32497 | n34249 ;
  assign n34251 = n32494 | n34250 ;
  assign n34252 = n8970 | n34245 ;
  assign n34253 = n34248 | n34252 ;
  assign n34254 = n34251 & n34253 ;
  assign n34255 = ~x2 & n34253 ;
  assign n34256 = n34251 & n34255 ;
  assign n34257 = x2 | n34255 ;
  assign n34258 = ( x2 & n34251 ) | ( x2 & n34257 ) | ( n34251 & n34257 ) ;
  assign n34259 = ( ~n34254 & n34256 ) | ( ~n34254 & n34258 ) | ( n34256 & n34258 ) ;
  assign n34260 = n34224 & n34226 ;
  assign n34261 = ( n34221 & n34224 ) | ( n34221 & n34260 ) | ( n34224 & n34260 ) ;
  assign n34262 = n34259 & n34261 ;
  assign n34263 = ( n34244 & n34259 ) | ( n34244 & n34262 ) | ( n34259 & n34262 ) ;
  assign n34264 = n33606 & n34263 ;
  assign n34265 = n32577 | n33195 ;
  assign n34266 = n34259 | n34261 ;
  assign n34267 = n34244 | n34266 ;
  assign n34268 = ( n32577 & n33195 ) | ( n32577 & ~n34265 ) | ( n33195 & ~n34265 ) ;
  assign n34269 = ( ~n34265 & n34267 ) | ( ~n34265 & n34268 ) | ( n34267 & n34268 ) ;
  assign n34270 = ( n33606 & n34264 ) | ( n33606 & n34269 ) | ( n34264 & n34269 ) ;
  assign n34271 = n32456 & n33441 ;
  assign n34272 = n9475 & n33436 ;
  assign n34273 = n9021 & n32293 ;
  assign n34274 = n9024 & ~n32442 ;
  assign n34275 = n34273 | n34274 ;
  assign n34276 = n34272 | n34275 ;
  assign n34277 = n33441 & ~n34276 ;
  assign n34278 = ( n32456 & ~n34276 ) | ( n32456 & n34277 ) | ( ~n34276 & n34277 ) ;
  assign n34279 = ~n34271 & n34278 ;
  assign n34280 = n8970 | n34272 ;
  assign n34281 = n34275 | n34280 ;
  assign n34282 = ~n34279 & n34281 ;
  assign n34283 = x2 & n34281 ;
  assign n34284 = ~n34279 & n34283 ;
  assign n34285 = x2 & ~n34283 ;
  assign n34286 = ( x2 & n34279 ) | ( x2 & n34285 ) | ( n34279 & n34285 ) ;
  assign n34287 = ( n34282 & ~n34284 ) | ( n34282 & n34286 ) | ( ~n34284 & n34286 ) ;
  assign n34288 = n34270 | n34287 ;
  assign n34289 = n33197 | n33199 ;
  assign n34290 = n33606 | n34263 ;
  assign n34291 = n34269 | n34290 ;
  assign n34292 = ( n33197 & n33199 ) | ( n33197 & ~n34289 ) | ( n33199 & ~n34289 ) ;
  assign n34293 = ( ~n34289 & n34291 ) | ( ~n34289 & n34292 ) | ( n34291 & n34292 ) ;
  assign n34294 = n34288 | n34293 ;
  assign n34295 = ( ~n32538 & n33201 ) | ( ~n32538 & n33590 ) | ( n33201 & n33590 ) ;
  assign n34296 = ( n33590 & n34294 ) | ( n33590 & n34295 ) | ( n34294 & n34295 ) ;
  assign n34297 = n34270 & n34287 ;
  assign n34298 = ( n34287 & n34293 ) | ( n34287 & n34297 ) | ( n34293 & n34297 ) ;
  assign n34299 = ~n33589 & n34298 ;
  assign n34300 = ( ~n33589 & n34296 ) | ( ~n33589 & n34299 ) | ( n34296 & n34299 ) ;
  assign n34301 = ( ~n33558 & n33586 ) | ( ~n33558 & n34300 ) | ( n33586 & n34300 ) ;
  assign n34302 = n33558 & ~n33585 ;
  assign n34303 = ~n34300 & n34302 ;
  assign n34304 = n34301 | n34303 ;
  assign n34305 = n33589 & ~n34298 ;
  assign n34306 = ~n34296 & n34305 ;
  assign n34307 = n34300 | n34306 ;
  assign n34308 = n34304 | n34307 ;
  assign n34309 = ~n34307 & n34308 ;
  assign n34310 = ( ~n34304 & n34308 ) | ( ~n34304 & n34309 ) | ( n34308 & n34309 ) ;
  assign n34311 = n29649 | n29653 ;
  assign n34312 = n29404 | n29408 ;
  assign n34396 = ~n29353 & n29356 ;
  assign n34397 = ( n29353 & n29358 ) | ( n29353 & ~n34396 ) | ( n29358 & ~n34396 ) ;
  assign n34313 = n29331 | n29337 ;
  assign n34352 = ~n29321 & n29326 ;
  assign n34353 = ( n29267 & n29321 ) | ( n29267 & ~n34352 ) | ( n29321 & ~n34352 ) ;
  assign n34314 = n1057 & n23620 ;
  assign n34315 = n1065 & n22381 ;
  assign n34316 = n1060 & ~n22385 ;
  assign n34317 = n34315 | n34316 ;
  assign n34318 = n34314 | n34317 ;
  assign n34319 = n1062 | n34316 ;
  assign n34320 = n34315 | n34319 ;
  assign n34321 = n34314 | n34320 ;
  assign n34322 = ( ~n23686 & n34318 ) | ( ~n23686 & n34321 ) | ( n34318 & n34321 ) ;
  assign n34323 = n168 | n202 ;
  assign n34324 = n3330 | n34323 ;
  assign n34325 = n143 & ~n262 ;
  assign n34326 = ~n39 & n34325 ;
  assign n34327 = ~n34324 & n34326 ;
  assign n34328 = ~n245 & n34327 ;
  assign n34329 = n2841 | n6973 ;
  assign n34330 = n397 | n34329 ;
  assign n34331 = n1122 | n34330 ;
  assign n34332 = n1512 | n34331 ;
  assign n34333 = n25775 | n34332 ;
  assign n34334 = n3495 | n6932 ;
  assign n34335 = n575 | n967 ;
  assign n34336 = n34334 | n34335 ;
  assign n34337 = n431 | n34336 ;
  assign n34338 = n474 | n34337 ;
  assign n34339 = n6028 | n34338 ;
  assign n34340 = n34333 | n34339 ;
  assign n34341 = n34328 & ~n34340 ;
  assign n34342 = n34320 & ~n34341 ;
  assign n34343 = ( n34314 & ~n34341 ) | ( n34314 & n34342 ) | ( ~n34341 & n34342 ) ;
  assign n34344 = n34317 & ~n34341 ;
  assign n34345 = ( n34314 & ~n34341 ) | ( n34314 & n34344 ) | ( ~n34341 & n34344 ) ;
  assign n34346 = ( ~n23686 & n34343 ) | ( ~n23686 & n34345 ) | ( n34343 & n34345 ) ;
  assign n34347 = n34322 & ~n34346 ;
  assign n34348 = n34321 | n34341 ;
  assign n34349 = n34318 | n34341 ;
  assign n34350 = ( ~n23686 & n34348 ) | ( ~n23686 & n34349 ) | ( n34348 & n34349 ) ;
  assign n34351 = ~n34347 & n34350 ;
  assign n34354 = ~n34351 & n34353 ;
  assign n34355 = n34353 & ~n34354 ;
  assign n34356 = n34351 | n34354 ;
  assign n34357 = ~n34355 & n34356 ;
  assign n34358 = n1829 & n24167 ;
  assign n34359 = n1826 & n23316 ;
  assign n34360 = n1823 & n23614 ;
  assign n34361 = n34359 | n34360 ;
  assign n34362 = n34358 | n34361 ;
  assign n34363 = n1821 | n34362 ;
  assign n34364 = ( n24182 & n34362 ) | ( n24182 & n34363 ) | ( n34362 & n34363 ) ;
  assign n34365 = n34362 | n34363 ;
  assign n34366 = ( n24175 & n34364 ) | ( n24175 & n34365 ) | ( n34364 & n34365 ) ;
  assign n34367 = x29 & n34366 ;
  assign n34368 = x29 & ~n34366 ;
  assign n34369 = ( n34366 & ~n34367 ) | ( n34366 & n34368 ) | ( ~n34367 & n34368 ) ;
  assign n34370 = ~n34357 & n34369 ;
  assign n34371 = n34357 & ~n34369 ;
  assign n34372 = n34370 | n34371 ;
  assign n34373 = n34313 & ~n34372 ;
  assign n34374 = ~n34313 & n34372 ;
  assign n34375 = n34373 | n34374 ;
  assign n34377 = n2312 & ~n25054 ;
  assign n34378 = n2308 & n24770 ;
  assign n34379 = n34377 | n34378 ;
  assign n34376 = n2315 & ~n25046 ;
  assign n34381 = n2306 | n34376 ;
  assign n34382 = n34379 | n34381 ;
  assign n34380 = n34376 | n34379 ;
  assign n34383 = n34380 & n34382 ;
  assign n34384 = ( ~n25069 & n34382 ) | ( ~n25069 & n34383 ) | ( n34382 & n34383 ) ;
  assign n34385 = ~x26 & n34383 ;
  assign n34386 = ~x26 & n34382 ;
  assign n34387 = ( ~n25069 & n34385 ) | ( ~n25069 & n34386 ) | ( n34385 & n34386 ) ;
  assign n34388 = x26 | n34385 ;
  assign n34389 = x26 | n34386 ;
  assign n34390 = ( ~n25069 & n34388 ) | ( ~n25069 & n34389 ) | ( n34388 & n34389 ) ;
  assign n34391 = ( ~n34384 & n34387 ) | ( ~n34384 & n34390 ) | ( n34387 & n34390 ) ;
  assign n34392 = ~n34375 & n34391 ;
  assign n34393 = n34375 | n34392 ;
  assign n34394 = n34375 & n34391 ;
  assign n34395 = n34393 & ~n34394 ;
  assign n34398 = ~n34395 & n34397 ;
  assign n34399 = n34397 & ~n34398 ;
  assign n34400 = n34395 | n34398 ;
  assign n34401 = ~n34399 & n34400 ;
  assign n34402 = n2925 & ~n25728 ;
  assign n34403 = n2928 & n26017 ;
  assign n34404 = n34402 | n34403 ;
  assign n34405 = n2932 & ~n26270 ;
  assign n34406 = ~n26263 & n34405 ;
  assign n34407 = n34404 | n34406 ;
  assign n34408 = n2936 | n34406 ;
  assign n34409 = n34404 | n34408 ;
  assign n34410 = ( n26571 & n34407 ) | ( n26571 & n34409 ) | ( n34407 & n34409 ) ;
  assign n34411 = x23 & n34409 ;
  assign n34412 = x23 & n34407 ;
  assign n34413 = ( n26571 & n34411 ) | ( n26571 & n34412 ) | ( n34411 & n34412 ) ;
  assign n34414 = x23 & ~n34412 ;
  assign n34415 = x23 & ~n34411 ;
  assign n34416 = ( ~n26571 & n34414 ) | ( ~n26571 & n34415 ) | ( n34414 & n34415 ) ;
  assign n34417 = ( n34410 & ~n34413 ) | ( n34410 & n34416 ) | ( ~n34413 & n34416 ) ;
  assign n34418 = ~n34401 & n34417 ;
  assign n34419 = n34401 | n34418 ;
  assign n34420 = n34401 & n34417 ;
  assign n34421 = n34419 & ~n34420 ;
  assign n34422 = ~n29377 & n29381 ;
  assign n34423 = ( n29377 & n29382 ) | ( n29377 & ~n34422 ) | ( n29382 & ~n34422 ) ;
  assign n34424 = n34421 & ~n34423 ;
  assign n34425 = ~n34421 & n34423 ;
  assign n34426 = n34424 | n34425 ;
  assign n34427 = n3544 & ~n26526 ;
  assign n34428 = ~n26520 & n34427 ;
  assign n34429 = n3541 & ~n27133 ;
  assign n34430 = ~n27125 & n34429 ;
  assign n34431 = n34428 | n34430 ;
  assign n34432 = n3547 & ~n27371 ;
  assign n34433 = ~n27363 & n34432 ;
  assign n34435 = n3537 | n34433 ;
  assign n34436 = n34431 | n34435 ;
  assign n34434 = n34431 | n34433 ;
  assign n34437 = n34434 & n34436 ;
  assign n34438 = ( ~n27654 & n34436 ) | ( ~n27654 & n34437 ) | ( n34436 & n34437 ) ;
  assign n34439 = ~x20 & n34437 ;
  assign n34440 = ~x20 & n34436 ;
  assign n34441 = ( ~n27654 & n34439 ) | ( ~n27654 & n34440 ) | ( n34439 & n34440 ) ;
  assign n34442 = x20 | n34439 ;
  assign n34443 = x20 | n34440 ;
  assign n34444 = ( ~n27654 & n34442 ) | ( ~n27654 & n34443 ) | ( n34442 & n34443 ) ;
  assign n34445 = ( ~n34438 & n34441 ) | ( ~n34438 & n34444 ) | ( n34441 & n34444 ) ;
  assign n34446 = ~n34426 & n34445 ;
  assign n34447 = n34426 | n34446 ;
  assign n34448 = n34426 & n34445 ;
  assign n34449 = n34447 & ~n34448 ;
  assign n34450 = n34312 & ~n34449 ;
  assign n34451 = n34312 & ~n34450 ;
  assign n34452 = n34312 | n34449 ;
  assign n34453 = ~n34451 & n34452 ;
  assign n34454 = n4471 & n28492 ;
  assign n34455 = n4466 & ~n27606 ;
  assign n34456 = ~n27597 & n34455 ;
  assign n34457 = n4468 & ~n28503 ;
  assign n34458 = n28498 & n34457 ;
  assign n34459 = n34456 | n34458 ;
  assign n34460 = n34454 | n34459 ;
  assign n34461 = n4475 | n34460 ;
  assign n34462 = ( ~n28749 & n34460 ) | ( ~n28749 & n34461 ) | ( n34460 & n34461 ) ;
  assign n34463 = ~x17 & n34461 ;
  assign n34464 = ~x17 & n34460 ;
  assign n34465 = ( ~n28749 & n34463 ) | ( ~n28749 & n34464 ) | ( n34463 & n34464 ) ;
  assign n34466 = x17 | n34463 ;
  assign n34467 = x17 | n34464 ;
  assign n34468 = ( ~n28749 & n34466 ) | ( ~n28749 & n34467 ) | ( n34466 & n34467 ) ;
  assign n34469 = ( ~n34462 & n34465 ) | ( ~n34462 & n34468 ) | ( n34465 & n34468 ) ;
  assign n34470 = ~n34452 & n34469 ;
  assign n34471 = ( n34451 & n34469 ) | ( n34451 & n34470 ) | ( n34469 & n34470 ) ;
  assign n34472 = n34453 | n34471 ;
  assign n34473 = n34452 & n34469 ;
  assign n34474 = ~n34451 & n34473 ;
  assign n34475 = n34472 & ~n34474 ;
  assign n34476 = n29428 | n29436 ;
  assign n34477 = n34475 & ~n34476 ;
  assign n34478 = ~n34475 & n34476 ;
  assign n34479 = n34477 | n34478 ;
  assign n34481 = n5237 & ~n28714 ;
  assign n34482 = n5231 & n29620 ;
  assign n34483 = n34481 | n34482 ;
  assign n34480 = n5234 & ~n30199 ;
  assign n34485 = n5227 | n34480 ;
  assign n34486 = n34483 | n34485 ;
  assign n34484 = n34480 | n34483 ;
  assign n34487 = n34484 & n34486 ;
  assign n34488 = ( ~n30299 & n34486 ) | ( ~n30299 & n34487 ) | ( n34486 & n34487 ) ;
  assign n34489 = ~x14 & n34487 ;
  assign n34490 = ~x14 & n34486 ;
  assign n34491 = ( ~n30299 & n34489 ) | ( ~n30299 & n34490 ) | ( n34489 & n34490 ) ;
  assign n34492 = x14 | n34489 ;
  assign n34493 = x14 | n34490 ;
  assign n34494 = ( ~n30299 & n34492 ) | ( ~n30299 & n34493 ) | ( n34492 & n34493 ) ;
  assign n34495 = ( ~n34488 & n34491 ) | ( ~n34488 & n34494 ) | ( n34491 & n34494 ) ;
  assign n34496 = ~n34479 & n34495 ;
  assign n34497 = n34479 | n34496 ;
  assign n34498 = n34479 & n34495 ;
  assign n34499 = n34497 & ~n34498 ;
  assign n34500 = n34311 & ~n34499 ;
  assign n34501 = n34311 & ~n34500 ;
  assign n34502 = n34499 | n34500 ;
  assign n34503 = ~n34501 & n34502 ;
  assign n34504 = n6122 & ~n31309 ;
  assign n34505 = n6125 & n30212 ;
  assign n34506 = n6119 & ~n30186 ;
  assign n34507 = n34505 | n34506 ;
  assign n34508 = n34504 | n34507 ;
  assign n34509 = n6115 | n34504 ;
  assign n34510 = n34507 | n34509 ;
  assign n34511 = ( n31404 & n34508 ) | ( n31404 & n34510 ) | ( n34508 & n34510 ) ;
  assign n34512 = x11 & n34510 ;
  assign n34513 = x11 & n34508 ;
  assign n34514 = ( n31404 & n34512 ) | ( n31404 & n34513 ) | ( n34512 & n34513 ) ;
  assign n34515 = x11 & ~n34513 ;
  assign n34516 = x11 & ~n34512 ;
  assign n34517 = ( ~n31404 & n34515 ) | ( ~n31404 & n34516 ) | ( n34515 & n34516 ) ;
  assign n34518 = ( n34511 & ~n34514 ) | ( n34511 & n34517 ) | ( ~n34514 & n34517 ) ;
  assign n34519 = ~n34503 & n34518 ;
  assign n34520 = n34503 | n34519 ;
  assign n34521 = n34503 & n34518 ;
  assign n34522 = n34520 & ~n34521 ;
  assign n34523 = n30252 | n30843 ;
  assign n34524 = ( n30252 & ~n30255 ) | ( n30252 & n34523 ) | ( ~n30255 & n34523 ) ;
  assign n34525 = n34522 & ~n34524 ;
  assign n34526 = ~n34522 & n34524 ;
  assign n34527 = n34525 | n34526 ;
  assign n34529 = n7074 & ~n31323 ;
  assign n34530 = n7068 & n31295 ;
  assign n34531 = n34529 | n34530 ;
  assign n34528 = n7079 & n32306 ;
  assign n34533 = n7078 | n34528 ;
  assign n34534 = n34531 | n34533 ;
  assign n34532 = n34528 | n34531 ;
  assign n34535 = n34532 & n34534 ;
  assign n34536 = ( ~n32525 & n34534 ) | ( ~n32525 & n34535 ) | ( n34534 & n34535 ) ;
  assign n34537 = ~x8 & n34535 ;
  assign n34538 = ~x8 & n34534 ;
  assign n34539 = ( ~n32525 & n34537 ) | ( ~n32525 & n34538 ) | ( n34537 & n34538 ) ;
  assign n34540 = x8 | n34537 ;
  assign n34541 = x8 | n34538 ;
  assign n34542 = ( ~n32525 & n34540 ) | ( ~n32525 & n34541 ) | ( n34540 & n34541 ) ;
  assign n34543 = ( ~n34536 & n34539 ) | ( ~n34536 & n34542 ) | ( n34539 & n34542 ) ;
  assign n34544 = ~n34527 & n34543 ;
  assign n34545 = n34527 | n34544 ;
  assign n34546 = n34527 & n34543 ;
  assign n34547 = n34545 & ~n34546 ;
  assign n34548 = n31364 | n32024 ;
  assign n34549 = ( n31364 & ~n31367 ) | ( n31364 & n34548 ) | ( ~n31367 & n34548 ) ;
  assign n34550 = n34547 & n34549 ;
  assign n34551 = n34547 | n34549 ;
  assign n34552 = ~n34550 & n34551 ;
  assign n34553 = n8122 & n33436 ;
  assign n34554 = n8115 & n32293 ;
  assign n34555 = n8118 & ~n32442 ;
  assign n34556 = n34554 | n34555 ;
  assign n34557 = n34553 | n34556 ;
  assign n34558 = n8125 & ~n33441 ;
  assign n34559 = ~n32456 & n34558 ;
  assign n34560 = ( n8125 & n34271 ) | ( n8125 & n34559 ) | ( n34271 & n34559 ) ;
  assign n34561 = n34557 | n34560 ;
  assign n34562 = x5 | n34557 ;
  assign n34563 = n34560 | n34562 ;
  assign n34564 = ~x5 & n34562 ;
  assign n34565 = ( ~x5 & n34560 ) | ( ~x5 & n34564 ) | ( n34560 & n34564 ) ;
  assign n34566 = ( ~n34561 & n34563 ) | ( ~n34561 & n34565 ) | ( n34563 & n34565 ) ;
  assign n34567 = ~n34552 & n34566 ;
  assign n34568 = n34552 & ~n34566 ;
  assign n34569 = n34567 | n34568 ;
  assign n34570 = n32474 | n33205 ;
  assign n34571 = ( n32474 & ~n32476 ) | ( n32474 & n34570 ) | ( ~n32476 & n34570 ) ;
  assign n34572 = n34569 & ~n34571 ;
  assign n34573 = ~n34569 & n34571 ;
  assign n34574 = n34572 | n34573 ;
  assign n34575 = n33463 & ~n33468 ;
  assign n34576 = ( ~n33453 & n33463 ) | ( ~n33453 & n34575 ) | ( n33463 & n34575 ) ;
  assign n34577 = ( ~n33451 & n33463 ) | ( ~n33451 & n34575 ) | ( n33463 & n34575 ) ;
  assign n34578 = ( n21587 & n34576 ) | ( n21587 & n34577 ) | ( n34576 & n34577 ) ;
  assign n34579 = n9018 | n9051 ;
  assign n34580 = ~n33460 & n34579 ;
  assign n34581 = n33460 & ~n34579 ;
  assign n34582 = n34580 | n34581 ;
  assign n34583 = n34576 | n34582 ;
  assign n34584 = n34577 | n34582 ;
  assign n34585 = ( n21587 & n34583 ) | ( n21587 & n34584 ) | ( n34583 & n34584 ) ;
  assign n34586 = ~n34578 & n34585 ;
  assign n34587 = ~n34581 & n34582 ;
  assign n34588 = ( n34577 & ~n34581 ) | ( n34577 & n34587 ) | ( ~n34581 & n34587 ) ;
  assign n34589 = ~n34580 & n34588 ;
  assign n34590 = ( n34576 & ~n34581 ) | ( n34576 & n34587 ) | ( ~n34581 & n34587 ) ;
  assign n34591 = ~n34580 & n34590 ;
  assign n34592 = ( n21587 & n34589 ) | ( n21587 & n34591 ) | ( n34589 & n34591 ) ;
  assign n34593 = n34586 | n34592 ;
  assign n34594 = n1823 | n1829 ;
  assign n34595 = ~n23234 & n34594 ;
  assign n34596 = ~n23235 & n34594 ;
  assign n34597 = ( ~n15882 & n34595 ) | ( ~n15882 & n34596 ) | ( n34595 & n34596 ) ;
  assign n34598 = n1826 | n34595 ;
  assign n34599 = n1826 | n34596 ;
  assign n34600 = ( ~n15882 & n34598 ) | ( ~n15882 & n34599 ) | ( n34598 & n34599 ) ;
  assign n34601 = ( ~n23240 & n34597 ) | ( ~n23240 & n34600 ) | ( n34597 & n34600 ) ;
  assign n34602 = n1821 & ~n24135 ;
  assign n34603 = n1821 & ~n23240 ;
  assign n34604 = ( ~n23575 & n34602 ) | ( ~n23575 & n34603 ) | ( n34602 & n34603 ) ;
  assign n34605 = ( ~n23577 & n34602 ) | ( ~n23577 & n34603 ) | ( n34602 & n34603 ) ;
  assign n34606 = n34604 & n34605 ;
  assign n34607 = n34601 | n34606 ;
  assign n34608 = ( n21554 & n34604 ) | ( n21554 & n34605 ) | ( n34604 & n34605 ) ;
  assign n34609 = n34601 | n34608 ;
  assign n34610 = ( ~n21584 & n34607 ) | ( ~n21584 & n34609 ) | ( n34607 & n34609 ) ;
  assign n34611 = x29 & n34609 ;
  assign n34612 = x29 & n34607 ;
  assign n34613 = ( ~n21584 & n34611 ) | ( ~n21584 & n34612 ) | ( n34611 & n34612 ) ;
  assign n34614 = n34610 & ~n34613 ;
  assign n34615 = x29 & ~n34609 ;
  assign n34616 = x29 & ~n34607 ;
  assign n34617 = ( n21584 & n34615 ) | ( n21584 & n34616 ) | ( n34615 & n34616 ) ;
  assign n34618 = n34614 | n34617 ;
  assign n34619 = n1060 & ~n21517 ;
  assign n34620 = n1065 & ~n21551 ;
  assign n34621 = n34619 | n34620 ;
  assign n34622 = n1057 & n23227 ;
  assign n34623 = ( n1057 & n23217 ) | ( n1057 & n34622 ) | ( n23217 & n34622 ) ;
  assign n34624 = n34621 | n34623 ;
  assign n34625 = n1062 & n23299 ;
  assign n34626 = n1062 & n23298 ;
  assign n34627 = ( n21584 & n34625 ) | ( n21584 & n34626 ) | ( n34625 & n34626 ) ;
  assign n34628 = n34624 | n34627 ;
  assign n34629 = n1062 | n34624 ;
  assign n34630 = ( n23289 & n34628 ) | ( n23289 & n34629 ) | ( n34628 & n34629 ) ;
  assign n34631 = n34618 & n34630 ;
  assign n34632 = n34618 & ~n34631 ;
  assign n34633 = n34630 & ~n34631 ;
  assign n34634 = n34632 | n34633 ;
  assign n34635 = n34593 & ~n34634 ;
  assign n34636 = ~n34593 & n34634 ;
  assign n34637 = n34635 | n34636 ;
  assign n34638 = n33479 | n33499 ;
  assign n34639 = ( n33479 & n33480 ) | ( n33479 & n34638 ) | ( n33480 & n34638 ) ;
  assign n34640 = n34637 & n34639 ;
  assign n34641 = n34637 | n34639 ;
  assign n34642 = ~n34640 & n34641 ;
  assign n34643 = n33505 | n33513 ;
  assign n34644 = n33505 | n33515 ;
  assign n34645 = ( n32274 & n34643 ) | ( n32274 & n34644 ) | ( n34643 & n34644 ) ;
  assign n34646 = n33505 | n33507 ;
  assign n34647 = ( n33505 & n33510 ) | ( n33505 & n34646 ) | ( n33510 & n34646 ) ;
  assign n34648 = n34645 & n34647 ;
  assign n34649 = n34642 & n34648 ;
  assign n34650 = ( n28465 & n34645 ) | ( n28465 & n34647 ) | ( n34645 & n34647 ) ;
  assign n34651 = n34642 & n34650 ;
  assign n34652 = ( n28489 & n34649 ) | ( n28489 & n34651 ) | ( n34649 & n34651 ) ;
  assign n34653 = n34642 | n34648 ;
  assign n34654 = n34642 | n34650 ;
  assign n34655 = ( n28489 & n34653 ) | ( n28489 & n34654 ) | ( n34653 & n34654 ) ;
  assign n34656 = ~n34652 & n34655 ;
  assign n34657 = n33526 | n34656 ;
  assign n34658 = n33526 & n34656 ;
  assign n34659 = n34657 & ~n34658 ;
  assign n34660 = n33527 & n34659 ;
  assign n34661 = ( ~n33534 & n34659 ) | ( ~n33534 & n34660 ) | ( n34659 & n34660 ) ;
  assign n34662 = ( n33530 & n34659 ) | ( n33530 & n34660 ) | ( n34659 & n34660 ) ;
  assign n34663 = ( n32456 & n34661 ) | ( n32456 & n34662 ) | ( n34661 & n34662 ) ;
  assign n34664 = n33544 & ~n34659 ;
  assign n34665 = n33547 | n34659 ;
  assign n34666 = ( n32456 & ~n34664 ) | ( n32456 & n34665 ) | ( ~n34664 & n34665 ) ;
  assign n34667 = ~n34663 & n34666 ;
  assign n34669 = n9021 & ~n33423 ;
  assign n34670 = n9024 & n33526 ;
  assign n34671 = n34669 | n34670 ;
  assign n34668 = n9475 & n34656 ;
  assign n34673 = n8970 | n34668 ;
  assign n34674 = n34671 | n34673 ;
  assign n34672 = n34668 | n34671 ;
  assign n34675 = n34672 & n34674 ;
  assign n34676 = ( n34667 & n34674 ) | ( n34667 & n34675 ) | ( n34674 & n34675 ) ;
  assign n34677 = x2 & n34675 ;
  assign n34678 = x2 & n34674 ;
  assign n34679 = ( n34667 & n34677 ) | ( n34667 & n34678 ) | ( n34677 & n34678 ) ;
  assign n34680 = x2 & ~n34677 ;
  assign n34681 = x2 & ~n34678 ;
  assign n34682 = ( ~n34667 & n34680 ) | ( ~n34667 & n34681 ) | ( n34680 & n34681 ) ;
  assign n34683 = ( n34676 & ~n34679 ) | ( n34676 & n34682 ) | ( ~n34679 & n34682 ) ;
  assign n34684 = ~n34574 & n34683 ;
  assign n34685 = n34574 & ~n34683 ;
  assign n34686 = n34684 | n34685 ;
  assign n34687 = n33556 | n33585 ;
  assign n34688 = ( n33556 & ~n33558 ) | ( n33556 & n34687 ) | ( ~n33558 & n34687 ) ;
  assign n34689 = ~n34686 & n34688 ;
  assign n34690 = ~n33556 & n33558 ;
  assign n34691 = n34686 | n34690 ;
  assign n34692 = ( n34300 & n34689 ) | ( n34300 & ~n34691 ) | ( n34689 & ~n34691 ) ;
  assign n34693 = n34686 & ~n34688 ;
  assign n34694 = n34686 & n34690 ;
  assign n34695 = ( ~n34300 & n34693 ) | ( ~n34300 & n34694 ) | ( n34693 & n34694 ) ;
  assign n34696 = n34692 | n34695 ;
  assign n34697 = n34308 | n34696 ;
  assign n34698 = n34308 & n34696 ;
  assign n34699 = n34697 & ~n34698 ;
  assign n34700 = n34496 | n34500 ;
  assign n34837 = ~n34446 & n34449 ;
  assign n34838 = ( n34312 & n34446 ) | ( n34312 & ~n34837 ) | ( n34446 & ~n34837 ) ;
  assign n34701 = n34392 | n34398 ;
  assign n34702 = n34346 | n34354 ;
  assign n34703 = n1057 & n23316 ;
  assign n34704 = n1060 & n22381 ;
  assign n34705 = n1065 | n34704 ;
  assign n34706 = ( n23620 & n34704 ) | ( n23620 & n34705 ) | ( n34704 & n34705 ) ;
  assign n34707 = n34703 | n34706 ;
  assign n34708 = n1062 | n34706 ;
  assign n34709 = n34703 | n34708 ;
  assign n34710 = ( n23661 & n34707 ) | ( n23661 & n34709 ) | ( n34707 & n34709 ) ;
  assign n34711 = n17922 | n17924 ;
  assign n34712 = n160 | n26285 ;
  assign n34713 = n24262 | n34712 ;
  assign n34714 = n129 | n1382 ;
  assign n34715 = n34713 | n34714 ;
  assign n34716 = n5091 | n17928 ;
  assign n34717 = n34715 | n34716 ;
  assign n34718 = n10868 | n34717 ;
  assign n34719 = n34711 | n34718 ;
  assign n34720 = n2060 | n34719 ;
  assign n34721 = n240 | n3376 ;
  assign n34722 = n979 | n34721 ;
  assign n34723 = n2747 | n34722 ;
  assign n34724 = n2856 | n3430 ;
  assign n34725 = n643 | n34724 ;
  assign n34726 = n34723 | n34725 ;
  assign n34727 = n237 | n356 ;
  assign n34728 = n103 | n555 ;
  assign n34729 = n34727 | n34728 ;
  assign n34730 = n34726 | n34729 ;
  assign n34731 = n34720 | n34730 ;
  assign n34732 = n34709 & n34731 ;
  assign n34733 = n34706 & n34731 ;
  assign n34734 = ( n34703 & n34731 ) | ( n34703 & n34733 ) | ( n34731 & n34733 ) ;
  assign n34735 = ( n23661 & n34732 ) | ( n23661 & n34734 ) | ( n34732 & n34734 ) ;
  assign n34736 = n34710 & ~n34735 ;
  assign n34737 = ~n34709 & n34731 ;
  assign n34738 = ~n34707 & n34731 ;
  assign n34739 = ( ~n23661 & n34737 ) | ( ~n23661 & n34738 ) | ( n34737 & n34738 ) ;
  assign n34740 = n34736 | n34739 ;
  assign n34741 = n34702 & n34740 ;
  assign n34742 = n34702 & ~n34741 ;
  assign n34743 = n1829 & ~n25054 ;
  assign n34744 = n1826 & n23614 ;
  assign n34745 = n1823 & n24167 ;
  assign n34746 = n34744 | n34745 ;
  assign n34747 = n34743 | n34746 ;
  assign n34748 = n1821 | n34743 ;
  assign n34749 = n34746 | n34748 ;
  assign n34750 = ( ~n25122 & n34747 ) | ( ~n25122 & n34749 ) | ( n34747 & n34749 ) ;
  assign n34751 = ~x29 & n34749 ;
  assign n34752 = ~x29 & n34747 ;
  assign n34753 = ( ~n25122 & n34751 ) | ( ~n25122 & n34752 ) | ( n34751 & n34752 ) ;
  assign n34754 = x29 | n34752 ;
  assign n34755 = x29 | n34751 ;
  assign n34756 = ( ~n25122 & n34754 ) | ( ~n25122 & n34755 ) | ( n34754 & n34755 ) ;
  assign n34757 = ( ~n34750 & n34753 ) | ( ~n34750 & n34756 ) | ( n34753 & n34756 ) ;
  assign n34758 = ~n34702 & n34740 ;
  assign n34759 = n34757 & n34758 ;
  assign n34760 = ( n34742 & n34757 ) | ( n34742 & n34759 ) | ( n34757 & n34759 ) ;
  assign n34761 = n34757 | n34758 ;
  assign n34762 = n34742 | n34761 ;
  assign n34763 = ~n34760 & n34762 ;
  assign n34764 = ~n34370 & n34372 ;
  assign n34765 = ( n34313 & n34370 ) | ( n34313 & ~n34764 ) | ( n34370 & ~n34764 ) ;
  assign n34766 = n34763 & n34765 ;
  assign n34767 = n34763 | n34765 ;
  assign n34768 = ~n34766 & n34767 ;
  assign n34769 = n2312 & n24770 ;
  assign n34770 = n2308 & ~n25046 ;
  assign n34771 = n34769 | n34770 ;
  assign n34772 = n2315 & ~n25728 ;
  assign n34773 = n2306 | n34772 ;
  assign n34774 = n34771 | n34773 ;
  assign n34775 = n34771 | n34772 ;
  assign n34776 = n25740 | n34775 ;
  assign n34777 = n25731 | n34775 ;
  assign n34778 = ( ~n25441 & n34776 ) | ( ~n25441 & n34777 ) | ( n34776 & n34777 ) ;
  assign n34779 = n34774 & n34778 ;
  assign n34780 = ( n25733 & n34774 ) | ( n25733 & n34779 ) | ( n34774 & n34779 ) ;
  assign n34781 = ~x26 & n34780 ;
  assign n34782 = x26 | n34780 ;
  assign n34783 = ( ~n34780 & n34781 ) | ( ~n34780 & n34782 ) | ( n34781 & n34782 ) ;
  assign n34784 = n34768 & n34783 ;
  assign n34785 = n34768 & ~n34784 ;
  assign n34786 = ~n34768 & n34783 ;
  assign n34787 = n34785 | n34786 ;
  assign n34788 = ~n34701 & n34787 ;
  assign n34789 = n34701 & ~n34787 ;
  assign n34790 = n34788 | n34789 ;
  assign n34791 = n2925 & n26017 ;
  assign n34792 = n2928 & ~n26270 ;
  assign n34793 = ~n26263 & n34792 ;
  assign n34794 = n34791 | n34793 ;
  assign n34795 = n2932 & ~n26526 ;
  assign n34796 = ~n26520 & n34795 ;
  assign n34797 = n34794 | n34796 ;
  assign n34798 = n2936 | n34796 ;
  assign n34799 = n34794 | n34798 ;
  assign n34800 = ( ~n26555 & n34797 ) | ( ~n26555 & n34799 ) | ( n34797 & n34799 ) ;
  assign n34801 = ( n26528 & n34797 ) | ( n26528 & n34799 ) | ( n34797 & n34799 ) ;
  assign n34802 = ( ~n26543 & n34800 ) | ( ~n26543 & n34801 ) | ( n34800 & n34801 ) ;
  assign n34803 = ~x23 & n34802 ;
  assign n34804 = x23 | n34802 ;
  assign n34805 = ( ~n34802 & n34803 ) | ( ~n34802 & n34804 ) | ( n34803 & n34804 ) ;
  assign n34806 = n34790 & n34805 ;
  assign n34807 = n34790 | n34805 ;
  assign n34808 = ~n34806 & n34807 ;
  assign n34809 = n34418 | n34808 ;
  assign n34810 = n34425 | n34809 ;
  assign n34811 = n34418 & n34808 ;
  assign n34812 = ( n34425 & n34808 ) | ( n34425 & n34811 ) | ( n34808 & n34811 ) ;
  assign n34813 = n34810 & ~n34812 ;
  assign n34814 = n3544 & ~n27133 ;
  assign n34815 = ~n27125 & n34814 ;
  assign n34816 = n3541 & ~n27371 ;
  assign n34817 = ~n27363 & n34816 ;
  assign n34818 = n34815 | n34817 ;
  assign n34819 = n3547 & ~n27606 ;
  assign n34820 = ~n27597 & n34819 ;
  assign n34821 = n34818 | n34820 ;
  assign n34822 = n27630 | n34821 ;
  assign n34823 = ( ~n27625 & n34821 ) | ( ~n27625 & n34822 ) | ( n34821 & n34822 ) ;
  assign n34824 = n27634 & ~n34823 ;
  assign n34825 = n3537 | n34820 ;
  assign n34826 = n34818 | n34825 ;
  assign n34827 = ~n34824 & n34826 ;
  assign n34828 = x20 & n34826 ;
  assign n34829 = ~n34824 & n34828 ;
  assign n34830 = x20 & ~n34828 ;
  assign n34831 = ( x20 & n34824 ) | ( x20 & n34830 ) | ( n34824 & n34830 ) ;
  assign n34832 = ( n34827 & ~n34829 ) | ( n34827 & n34831 ) | ( ~n34829 & n34831 ) ;
  assign n34833 = n34813 & n34832 ;
  assign n34834 = n34813 & ~n34833 ;
  assign n34835 = ~n34813 & n34832 ;
  assign n34836 = n34834 | n34835 ;
  assign n34839 = n34836 & n34838 ;
  assign n34840 = n34838 & ~n34839 ;
  assign n34841 = n34836 & ~n34838 ;
  assign n34842 = n34840 | n34841 ;
  assign n34843 = n4471 & ~n28714 ;
  assign n34844 = n4468 & n28492 ;
  assign n34845 = n4466 & ~n28503 ;
  assign n34846 = n28498 & n34845 ;
  assign n34847 = n34844 | n34846 ;
  assign n34848 = n34843 | n34847 ;
  assign n34849 = n4475 & ~n28731 ;
  assign n34850 = ~n28518 & n34849 ;
  assign n34851 = n34848 | n34850 ;
  assign n34852 = n4475 | n34848 ;
  assign n34853 = ( n28720 & n34851 ) | ( n28720 & n34852 ) | ( n34851 & n34852 ) ;
  assign n34854 = x17 | n34853 ;
  assign n34855 = ~x17 & n34853 ;
  assign n34856 = ( ~n34853 & n34854 ) | ( ~n34853 & n34855 ) | ( n34854 & n34855 ) ;
  assign n34857 = n34841 & n34856 ;
  assign n34858 = ( n34840 & n34856 ) | ( n34840 & n34857 ) | ( n34856 & n34857 ) ;
  assign n34859 = n34842 & ~n34858 ;
  assign n34860 = ~n34841 & n34856 ;
  assign n34861 = ~n34840 & n34860 ;
  assign n34862 = n34859 | n34861 ;
  assign n34863 = n34471 | n34478 ;
  assign n34864 = n34862 | n34863 ;
  assign n34865 = n34862 & n34863 ;
  assign n34866 = n34864 & ~n34865 ;
  assign n34867 = n5234 & n30212 ;
  assign n34868 = n5237 & n29620 ;
  assign n34869 = n5231 & ~n30199 ;
  assign n34870 = n34868 | n34869 ;
  assign n34871 = n34867 | n34870 ;
  assign n34872 = n30266 & ~n34871 ;
  assign n34873 = ~n30276 & n34872 ;
  assign n34874 = n5227 | n34867 ;
  assign n34875 = n34870 | n34874 ;
  assign n34876 = ~n34873 & n34875 ;
  assign n34877 = x14 & n34875 ;
  assign n34878 = ~n34873 & n34877 ;
  assign n34879 = x14 & ~n34877 ;
  assign n34880 = ( x14 & n34873 ) | ( x14 & n34879 ) | ( n34873 & n34879 ) ;
  assign n34881 = ( n34876 & ~n34878 ) | ( n34876 & n34880 ) | ( ~n34878 & n34880 ) ;
  assign n34882 = n34866 & n34881 ;
  assign n34883 = n34866 & ~n34882 ;
  assign n34884 = ~n34866 & n34881 ;
  assign n34885 = n34883 | n34884 ;
  assign n34886 = n34700 & n34885 ;
  assign n34887 = n34700 & ~n34886 ;
  assign n34888 = n34885 & ~n34886 ;
  assign n34889 = n34887 | n34888 ;
  assign n34890 = n6122 & ~n31323 ;
  assign n34891 = n6125 & ~n30186 ;
  assign n34892 = n6119 & ~n31309 ;
  assign n34893 = n34891 | n34892 ;
  assign n34894 = n34890 | n34893 ;
  assign n34895 = n6115 & n31384 ;
  assign n34896 = n6115 & n31386 ;
  assign n34897 = ( ~n30232 & n34895 ) | ( ~n30232 & n34896 ) | ( n34895 & n34896 ) ;
  assign n34898 = n34894 | n34897 ;
  assign n34899 = n6115 | n34894 ;
  assign n34900 = ( ~n31376 & n34898 ) | ( ~n31376 & n34899 ) | ( n34898 & n34899 ) ;
  assign n34901 = x11 | n34900 ;
  assign n34902 = ~x11 & n34900 ;
  assign n34903 = ( ~n34900 & n34901 ) | ( ~n34900 & n34902 ) | ( n34901 & n34902 ) ;
  assign n34904 = n34889 & n34903 ;
  assign n34905 = n34889 & ~n34904 ;
  assign n34906 = ~n34889 & n34903 ;
  assign n34907 = n34905 | n34906 ;
  assign n34908 = n34519 | n34524 ;
  assign n34909 = ( n34519 & ~n34522 ) | ( n34519 & n34908 ) | ( ~n34522 & n34908 ) ;
  assign n34910 = n34907 | n34909 ;
  assign n34911 = n34907 & n34909 ;
  assign n34912 = n34910 & ~n34911 ;
  assign n34913 = n7079 & n32293 ;
  assign n34914 = n7074 & n31295 ;
  assign n34915 = n7068 & n32306 ;
  assign n34916 = n34914 | n34915 ;
  assign n34917 = n34913 | n34916 ;
  assign n34918 = n32497 | n34917 ;
  assign n34919 = n32494 | n34918 ;
  assign n34920 = n7078 | n34913 ;
  assign n34921 = n34916 | n34920 ;
  assign n34922 = n34919 & n34921 ;
  assign n34923 = ~x8 & n34921 ;
  assign n34924 = n34919 & n34923 ;
  assign n34925 = x8 | n34923 ;
  assign n34926 = ( x8 & n34919 ) | ( x8 & n34925 ) | ( n34919 & n34925 ) ;
  assign n34927 = ( ~n34922 & n34924 ) | ( ~n34922 & n34926 ) | ( n34924 & n34926 ) ;
  assign n34928 = n34912 & n34927 ;
  assign n34929 = n34912 & ~n34928 ;
  assign n34930 = ~n34912 & n34927 ;
  assign n34931 = n34929 | n34930 ;
  assign n34932 = n34544 | n34549 ;
  assign n34933 = ( n34544 & ~n34547 ) | ( n34544 & n34932 ) | ( ~n34547 & n34932 ) ;
  assign n34934 = ~n34931 & n34933 ;
  assign n34935 = n34931 & ~n34933 ;
  assign n34936 = n34934 | n34935 ;
  assign n34937 = n8122 & ~n33423 ;
  assign n34938 = n8115 & ~n32442 ;
  assign n34939 = n8118 & n33436 ;
  assign n34940 = n34938 | n34939 ;
  assign n34941 = n34937 | n34940 ;
  assign n34942 = n8125 & n33575 ;
  assign n34943 = n8125 & ~n33577 ;
  assign n34944 = ( ~n32456 & n34942 ) | ( ~n32456 & n34943 ) | ( n34942 & n34943 ) ;
  assign n34945 = n34941 | n34944 ;
  assign n34946 = n8125 | n34941 ;
  assign n34947 = ( n33567 & n34945 ) | ( n33567 & n34946 ) | ( n34945 & n34946 ) ;
  assign n34948 = x5 | n34947 ;
  assign n34949 = ~x5 & n34947 ;
  assign n34950 = ( ~n34947 & n34948 ) | ( ~n34947 & n34949 ) | ( n34948 & n34949 ) ;
  assign n34951 = n34936 & n34950 ;
  assign n34952 = n34936 | n34950 ;
  assign n34953 = ~n34951 & n34952 ;
  assign n34954 = n34567 | n34571 ;
  assign n34955 = ( n34567 & ~n34569 ) | ( n34567 & n34954 ) | ( ~n34569 & n34954 ) ;
  assign n34956 = n34953 | n34955 ;
  assign n34957 = n34953 & n34955 ;
  assign n34958 = n34956 & ~n34957 ;
  assign n34959 = ( n21587 & n34588 ) | ( n21587 & n34590 ) | ( n34588 & n34590 ) ;
  assign n34960 = n1057 & ~n23240 ;
  assign n34961 = n1060 & ~n21551 ;
  assign n34962 = n1065 & n23227 ;
  assign n34963 = ( n1065 & n23217 ) | ( n1065 & n34962 ) | ( n23217 & n34962 ) ;
  assign n34964 = n34961 | n34963 ;
  assign n34965 = n34960 | n34964 ;
  assign n34966 = n1062 | n34960 ;
  assign n34967 = n34964 | n34966 ;
  assign n34968 = ( n23260 & n34965 ) | ( n23260 & n34967 ) | ( n34965 & n34967 ) ;
  assign n34969 = n9051 & n23199 ;
  assign n34970 = ( n9018 & n23199 ) | ( n9018 & n34969 ) | ( n23199 & n34969 ) ;
  assign n34971 = ( n23192 & n34579 ) | ( n23192 & n34970 ) | ( n34579 & n34970 ) ;
  assign n34972 = n9051 | n23199 ;
  assign n34973 = n9018 | n34972 ;
  assign n34974 = n23192 | n34973 ;
  assign n34975 = ~n34971 & n34974 ;
  assign n34976 = n1820 | n1823 ;
  assign n34977 = n1826 | n34976 ;
  assign n34978 = ~n23229 & n34977 ;
  assign n34979 = ( n23154 & n34977 ) | ( n23154 & n34978 ) | ( n34977 & n34978 ) ;
  assign n34980 = ~n23232 & n34977 ;
  assign n34981 = ~n23231 & n34977 ;
  assign n34982 = ( n9072 & n34980 ) | ( n9072 & n34981 ) | ( n34980 & n34981 ) ;
  assign n34983 = ( ~n21543 & n34979 ) | ( ~n21543 & n34982 ) | ( n34979 & n34982 ) ;
  assign n34984 = ( ~n21545 & n34979 ) | ( ~n21545 & n34982 ) | ( n34979 & n34982 ) ;
  assign n34985 = ( ~n15882 & n34983 ) | ( ~n15882 & n34984 ) | ( n34983 & n34984 ) ;
  assign n34986 = ~x29 & n34983 ;
  assign n34987 = ~x29 & n34984 ;
  assign n34988 = ( ~n15882 & n34986 ) | ( ~n15882 & n34987 ) | ( n34986 & n34987 ) ;
  assign n34989 = x29 | n34986 ;
  assign n34990 = x29 | n34987 ;
  assign n34991 = ( ~n15882 & n34989 ) | ( ~n15882 & n34990 ) | ( n34989 & n34990 ) ;
  assign n34992 = ( ~n34985 & n34988 ) | ( ~n34985 & n34991 ) | ( n34988 & n34991 ) ;
  assign n34993 = n34975 & ~n34992 ;
  assign n34994 = ~n34975 & n34992 ;
  assign n34995 = n34993 | n34994 ;
  assign n34996 = n34967 & ~n34995 ;
  assign n34997 = n34965 & ~n34995 ;
  assign n34998 = ( n23260 & n34996 ) | ( n23260 & n34997 ) | ( n34996 & n34997 ) ;
  assign n34999 = n34968 & ~n34998 ;
  assign n35000 = n34967 | n34995 ;
  assign n35001 = n34965 | n34995 ;
  assign n35002 = ( n23260 & n35000 ) | ( n23260 & n35001 ) | ( n35000 & n35001 ) ;
  assign n35003 = n34959 | n35002 ;
  assign n35004 = ( n34959 & ~n34999 ) | ( n34959 & n35003 ) | ( ~n34999 & n35003 ) ;
  assign n35005 = n34959 & n35002 ;
  assign n35006 = ~n34999 & n35005 ;
  assign n35007 = n35004 & ~n35006 ;
  assign n35008 = n34593 | n34631 ;
  assign n35009 = ( n34631 & n34634 ) | ( n34631 & n35008 ) | ( n34634 & n35008 ) ;
  assign n35010 = n35007 & n35009 ;
  assign n35011 = n35007 | n35009 ;
  assign n35012 = ~n35010 & n35011 ;
  assign n35013 = n34640 & n35012 ;
  assign n35014 = ( n34651 & n35012 ) | ( n34651 & n35013 ) | ( n35012 & n35013 ) ;
  assign n35015 = ( n34649 & n35012 ) | ( n34649 & n35013 ) | ( n35012 & n35013 ) ;
  assign n35016 = ( n28489 & n35014 ) | ( n28489 & n35015 ) | ( n35014 & n35015 ) ;
  assign n35017 = n34640 | n35012 ;
  assign n35018 = n34651 | n35017 ;
  assign n35019 = n34649 | n35017 ;
  assign n35020 = ( n28489 & n35018 ) | ( n28489 & n35019 ) | ( n35018 & n35019 ) ;
  assign n35021 = ~n35016 & n35020 ;
  assign n35022 = n34656 | n35021 ;
  assign n35023 = n34656 & n35021 ;
  assign n35024 = n35022 & ~n35023 ;
  assign n35025 = n34658 | n34661 ;
  assign n35026 = n35024 & n35025 ;
  assign n35027 = n34658 | n34662 ;
  assign n35028 = n35024 & n35027 ;
  assign n35029 = ( n32456 & n35026 ) | ( n32456 & n35028 ) | ( n35026 & n35028 ) ;
  assign n35030 = n35024 | n35025 ;
  assign n35031 = n35024 | n35027 ;
  assign n35032 = ( n32456 & n35030 ) | ( n32456 & n35031 ) | ( n35030 & n35031 ) ;
  assign n35033 = ~n35029 & n35032 ;
  assign n35034 = n9475 & n35021 ;
  assign n35035 = n9021 & n33526 ;
  assign n35036 = n9024 & n34656 ;
  assign n35037 = n35035 | n35036 ;
  assign n35038 = n35034 | n35037 ;
  assign n35039 = n8970 | n35034 ;
  assign n35040 = n35037 | n35039 ;
  assign n35041 = ( n35033 & n35038 ) | ( n35033 & n35040 ) | ( n35038 & n35040 ) ;
  assign n35042 = x2 & n35040 ;
  assign n35043 = x2 & n35038 ;
  assign n35044 = ( n35033 & n35042 ) | ( n35033 & n35043 ) | ( n35042 & n35043 ) ;
  assign n35045 = x2 & ~n35043 ;
  assign n35046 = x2 & ~n35042 ;
  assign n35047 = ( ~n35033 & n35045 ) | ( ~n35033 & n35046 ) | ( n35045 & n35046 ) ;
  assign n35048 = ( n35041 & ~n35044 ) | ( n35041 & n35047 ) | ( ~n35044 & n35047 ) ;
  assign n35049 = n34958 & n35048 ;
  assign n35050 = n34958 | n35048 ;
  assign n35051 = ~n35049 & n35050 ;
  assign n35052 = n34684 | n34689 ;
  assign n35053 = n35051 & n35052 ;
  assign n35054 = ~n34684 & n34691 ;
  assign n35055 = n35051 & ~n35054 ;
  assign n35056 = ( n34300 & n35053 ) | ( n34300 & n35055 ) | ( n35053 & n35055 ) ;
  assign n35057 = n35051 | n35052 ;
  assign n35058 = ~n35051 & n35054 ;
  assign n35059 = ( n34300 & n35057 ) | ( n34300 & ~n35058 ) | ( n35057 & ~n35058 ) ;
  assign n35060 = ~n35056 & n35059 ;
  assign n35061 = n34697 & ~n35060 ;
  assign n35062 = ~n34696 & n35060 ;
  assign n35063 = ~n34308 & n35062 ;
  assign n35064 = n35061 | n35063 ;
  assign n35065 = n34882 | n34886 ;
  assign n35147 = n34784 | n34787 ;
  assign n35148 = ( n34701 & n34784 ) | ( n34701 & n35147 ) | ( n34784 & n35147 ) ;
  assign n35101 = n34735 | n34740 ;
  assign n35102 = ( n34702 & n34735 ) | ( n34702 & n35101 ) | ( n34735 & n35101 ) ;
  assign n35066 = n1057 & n23614 ;
  assign n35067 = n1065 & n23316 ;
  assign n35068 = n1060 & n23620 ;
  assign n35069 = n35067 | n35068 ;
  assign n35070 = n35066 | n35069 ;
  assign n35071 = n1062 | n35068 ;
  assign n35072 = n35067 | n35071 ;
  assign n35073 = n35066 | n35072 ;
  assign n35074 = ( n23634 & n35070 ) | ( n23634 & n35073 ) | ( n35070 & n35073 ) ;
  assign n35075 = n758 | n23898 ;
  assign n35076 = n54 | n319 ;
  assign n35077 = n6029 | n35076 ;
  assign n35078 = n2843 | n2865 ;
  assign n35079 = n35077 | n35078 ;
  assign n35080 = n129 | n15233 ;
  assign n35081 = n35079 | n35080 ;
  assign n35082 = ( ~n1379 & n35075 ) | ( ~n1379 & n35081 ) | ( n35075 & n35081 ) ;
  assign n35083 = n35075 & n35081 ;
  assign n35084 = ( n1410 & n35082 ) | ( n1410 & n35083 ) | ( n35082 & n35083 ) ;
  assign n35085 = n1411 & ~n35084 ;
  assign n35086 = n1231 | n18485 ;
  assign n35087 = n1521 | n2748 ;
  assign n35088 = n309 | n710 ;
  assign n35089 = n35087 | n35088 ;
  assign n35090 = n151 | n35089 ;
  assign n35091 = n35086 | n35090 ;
  assign n35092 = n35085 & ~n35091 ;
  assign n35093 = n35073 & ~n35092 ;
  assign n35094 = n35070 & ~n35092 ;
  assign n35095 = ( n23634 & n35093 ) | ( n23634 & n35094 ) | ( n35093 & n35094 ) ;
  assign n35096 = n35074 & ~n35095 ;
  assign n35097 = n35073 | n35092 ;
  assign n35098 = n35070 | n35092 ;
  assign n35099 = ( n23634 & n35097 ) | ( n23634 & n35098 ) | ( n35097 & n35098 ) ;
  assign n35100 = ~n35096 & n35099 ;
  assign n35103 = ~n35100 & n35102 ;
  assign n35104 = n35102 & ~n35103 ;
  assign n35105 = n1829 & n24770 ;
  assign n35106 = n1826 & n24167 ;
  assign n35107 = n1823 & ~n25054 ;
  assign n35108 = n35106 | n35107 ;
  assign n35109 = n35105 | n35108 ;
  assign n35110 = n1821 | n35109 ;
  assign n35111 = ( ~n25095 & n35109 ) | ( ~n25095 & n35110 ) | ( n35109 & n35110 ) ;
  assign n35112 = ~x29 & n35110 ;
  assign n35113 = ~x29 & n35109 ;
  assign n35114 = ( ~n25095 & n35112 ) | ( ~n25095 & n35113 ) | ( n35112 & n35113 ) ;
  assign n35115 = x29 | n35112 ;
  assign n35116 = x29 | n35113 ;
  assign n35117 = ( ~n25095 & n35115 ) | ( ~n25095 & n35116 ) | ( n35115 & n35116 ) ;
  assign n35118 = ( ~n35111 & n35114 ) | ( ~n35111 & n35117 ) | ( n35114 & n35117 ) ;
  assign n35119 = n35100 | n35102 ;
  assign n35120 = n35118 & ~n35119 ;
  assign n35121 = ( n35104 & n35118 ) | ( n35104 & n35120 ) | ( n35118 & n35120 ) ;
  assign n35122 = ~n35118 & n35119 ;
  assign n35123 = ~n35104 & n35122 ;
  assign n35124 = n35121 | n35123 ;
  assign n35125 = n34760 | n34763 ;
  assign n35126 = ( n34760 & n34765 ) | ( n34760 & n35125 ) | ( n34765 & n35125 ) ;
  assign n35127 = ~n35124 & n35126 ;
  assign n35128 = n35124 & ~n35126 ;
  assign n35129 = n35127 | n35128 ;
  assign n35130 = n2315 & n26017 ;
  assign n35131 = n2312 & ~n25046 ;
  assign n35132 = n2308 & ~n25728 ;
  assign n35133 = n35131 | n35132 ;
  assign n35134 = n35130 | n35133 ;
  assign n35135 = n2306 | n35130 ;
  assign n35136 = n35133 | n35135 ;
  assign n35137 = ( n26613 & n35134 ) | ( n26613 & n35136 ) | ( n35134 & n35136 ) ;
  assign n35138 = n35134 | n35136 ;
  assign n35139 = ( n26605 & n35137 ) | ( n26605 & n35138 ) | ( n35137 & n35138 ) ;
  assign n35140 = x26 & n35139 ;
  assign n35141 = x26 & ~n35139 ;
  assign n35142 = ( n35139 & ~n35140 ) | ( n35139 & n35141 ) | ( ~n35140 & n35141 ) ;
  assign n35143 = ~n35129 & n35142 ;
  assign n35144 = n35129 | n35143 ;
  assign n35145 = n35129 & n35142 ;
  assign n35146 = n35144 & ~n35145 ;
  assign n35149 = ~n35146 & n35148 ;
  assign n35150 = n35148 & ~n35149 ;
  assign n35151 = n2925 & ~n26270 ;
  assign n35152 = ~n26263 & n35151 ;
  assign n35153 = n2928 & ~n26526 ;
  assign n35154 = ~n26520 & n35153 ;
  assign n35155 = n35152 | n35154 ;
  assign n35156 = n2932 & ~n27133 ;
  assign n35157 = ~n27125 & n35156 ;
  assign n35158 = n35155 | n35157 ;
  assign n35159 = n2936 & n27699 ;
  assign n35160 = ( n2936 & ~n27696 ) | ( n2936 & n35159 ) | ( ~n27696 & n35159 ) ;
  assign n35161 = n35158 | n35160 ;
  assign n35162 = x23 | n35158 ;
  assign n35163 = n35160 | n35162 ;
  assign n35164 = ~x23 & n35162 ;
  assign n35165 = ( ~x23 & n35160 ) | ( ~x23 & n35164 ) | ( n35160 & n35164 ) ;
  assign n35166 = ( ~n35161 & n35163 ) | ( ~n35161 & n35165 ) | ( n35163 & n35165 ) ;
  assign n35167 = n35146 | n35148 ;
  assign n35168 = n35166 & ~n35167 ;
  assign n35169 = ( n35150 & n35166 ) | ( n35150 & n35168 ) | ( n35166 & n35168 ) ;
  assign n35170 = ~n35166 & n35167 ;
  assign n35171 = ~n35150 & n35170 ;
  assign n35172 = n35169 | n35171 ;
  assign n35173 = ~n34806 & n35172 ;
  assign n35174 = ~n34812 & n35173 ;
  assign n35175 = n34806 & ~n35172 ;
  assign n35176 = ( n34812 & ~n35172 ) | ( n34812 & n35175 ) | ( ~n35172 & n35175 ) ;
  assign n35177 = n35174 | n35176 ;
  assign n35178 = n3544 & ~n27371 ;
  assign n35179 = ~n27363 & n35178 ;
  assign n35180 = n3541 & ~n27606 ;
  assign n35181 = ~n27597 & n35180 ;
  assign n35182 = n35179 | n35181 ;
  assign n35183 = n3547 & ~n28503 ;
  assign n35184 = n28498 & n35183 ;
  assign n35185 = n35182 | n35184 ;
  assign n35186 = n28794 | n35185 ;
  assign n35187 = n28783 | n35186 ;
  assign n35188 = n3537 | n35184 ;
  assign n35189 = n35182 | n35188 ;
  assign n35190 = n35187 & n35189 ;
  assign n35191 = ~x20 & n35189 ;
  assign n35192 = n35187 & n35191 ;
  assign n35193 = x20 | n35191 ;
  assign n35194 = ( x20 & n35187 ) | ( x20 & n35193 ) | ( n35187 & n35193 ) ;
  assign n35195 = ( ~n35190 & n35192 ) | ( ~n35190 & n35194 ) | ( n35192 & n35194 ) ;
  assign n35196 = ~n35177 & n35195 ;
  assign n35197 = n35177 | n35196 ;
  assign n35198 = n35177 & n35195 ;
  assign n35199 = n35197 & ~n35198 ;
  assign n35200 = n34833 | n34836 ;
  assign n35201 = ( n34833 & n34838 ) | ( n34833 & n35200 ) | ( n34838 & n35200 ) ;
  assign n35202 = n35199 | n35201 ;
  assign n35203 = n35199 & n35201 ;
  assign n35204 = n35202 & ~n35203 ;
  assign n35205 = n4471 & n29620 ;
  assign n35206 = n4466 & n28492 ;
  assign n35207 = n4468 & ~n28714 ;
  assign n35208 = n35206 | n35207 ;
  assign n35209 = n35205 | n35208 ;
  assign n35210 = n4475 | n35205 ;
  assign n35211 = n35208 | n35210 ;
  assign n35212 = ( ~n29642 & n35209 ) | ( ~n29642 & n35211 ) | ( n35209 & n35211 ) ;
  assign n35213 = n35209 | n35211 ;
  assign n35214 = ( n29629 & n35212 ) | ( n29629 & n35213 ) | ( n35212 & n35213 ) ;
  assign n35215 = ~x17 & n35214 ;
  assign n35216 = x17 | n35214 ;
  assign n35217 = ( ~n35214 & n35215 ) | ( ~n35214 & n35216 ) | ( n35215 & n35216 ) ;
  assign n35218 = ~n35204 & n35217 ;
  assign n35219 = n35204 & ~n35217 ;
  assign n35220 = n35218 | n35219 ;
  assign n35221 = n34858 | n34862 ;
  assign n35222 = ( n34858 & n34863 ) | ( n34858 & n35221 ) | ( n34863 & n35221 ) ;
  assign n35223 = n35220 & ~n35222 ;
  assign n35224 = ~n35220 & n35222 ;
  assign n35225 = n35223 | n35224 ;
  assign n35227 = n5237 & ~n30199 ;
  assign n35228 = n5231 & n30212 ;
  assign n35229 = n35227 | n35228 ;
  assign n35226 = n5234 & ~n30186 ;
  assign n35231 = n5227 | n35226 ;
  assign n35232 = n35229 | n35231 ;
  assign n35230 = n35226 | n35229 ;
  assign n35233 = n35230 & n35232 ;
  assign n35234 = ( ~n30241 & n35232 ) | ( ~n30241 & n35233 ) | ( n35232 & n35233 ) ;
  assign n35235 = ~x14 & n35233 ;
  assign n35236 = ~x14 & n35232 ;
  assign n35237 = ( ~n30241 & n35235 ) | ( ~n30241 & n35236 ) | ( n35235 & n35236 ) ;
  assign n35238 = x14 | n35235 ;
  assign n35239 = x14 | n35236 ;
  assign n35240 = ( ~n30241 & n35238 ) | ( ~n30241 & n35239 ) | ( n35238 & n35239 ) ;
  assign n35241 = ( ~n35234 & n35237 ) | ( ~n35234 & n35240 ) | ( n35237 & n35240 ) ;
  assign n35242 = ~n35225 & n35241 ;
  assign n35243 = n35225 | n35242 ;
  assign n35244 = n35225 & n35241 ;
  assign n35245 = n35243 & ~n35244 ;
  assign n35246 = n35065 & ~n35245 ;
  assign n35247 = n35065 & ~n35246 ;
  assign n35248 = n35065 | n35245 ;
  assign n35249 = ~n35247 & n35248 ;
  assign n35250 = n6122 & n31295 ;
  assign n35251 = n6125 & ~n31309 ;
  assign n35252 = n6119 & ~n31323 ;
  assign n35253 = n35251 | n35252 ;
  assign n35254 = n35250 | n35253 ;
  assign n35255 = n6115 | n35250 ;
  assign n35256 = n35253 | n35255 ;
  assign n35257 = ( n31355 & n35254 ) | ( n31355 & n35256 ) | ( n35254 & n35256 ) ;
  assign n35258 = x11 & n35256 ;
  assign n35259 = x11 & n35254 ;
  assign n35260 = ( n31355 & n35258 ) | ( n31355 & n35259 ) | ( n35258 & n35259 ) ;
  assign n35261 = x11 & ~n35259 ;
  assign n35262 = x11 & ~n35258 ;
  assign n35263 = ( ~n31355 & n35261 ) | ( ~n31355 & n35262 ) | ( n35261 & n35262 ) ;
  assign n35264 = ( n35257 & ~n35260 ) | ( n35257 & n35263 ) | ( ~n35260 & n35263 ) ;
  assign n35265 = ~n35248 & n35264 ;
  assign n35266 = ( n35247 & n35264 ) | ( n35247 & n35265 ) | ( n35264 & n35265 ) ;
  assign n35267 = n35249 | n35266 ;
  assign n35268 = n35248 & n35264 ;
  assign n35269 = ~n35247 & n35268 ;
  assign n35270 = n35267 & ~n35269 ;
  assign n35271 = n34904 | n34909 ;
  assign n35272 = ( n34904 & n34907 ) | ( n34904 & n35271 ) | ( n34907 & n35271 ) ;
  assign n35273 = n35270 & ~n35272 ;
  assign n35274 = ~n35270 & n35272 ;
  assign n35275 = n35273 | n35274 ;
  assign n35277 = n7074 & n32306 ;
  assign n35278 = n7068 & n32293 ;
  assign n35279 = n35277 | n35278 ;
  assign n35276 = n7079 & ~n32442 ;
  assign n35281 = n7078 | n35276 ;
  assign n35282 = n35279 | n35281 ;
  assign n35280 = n35276 | n35279 ;
  assign n35283 = n35280 & n35282 ;
  assign n35284 = ( ~n32458 & n35282 ) | ( ~n32458 & n35283 ) | ( n35282 & n35283 ) ;
  assign n35285 = ~x8 & n35283 ;
  assign n35286 = ~x8 & n35282 ;
  assign n35287 = ( ~n32458 & n35285 ) | ( ~n32458 & n35286 ) | ( n35285 & n35286 ) ;
  assign n35288 = x8 | n35285 ;
  assign n35289 = x8 | n35286 ;
  assign n35290 = ( ~n32458 & n35288 ) | ( ~n32458 & n35289 ) | ( n35288 & n35289 ) ;
  assign n35291 = ( ~n35284 & n35287 ) | ( ~n35284 & n35290 ) | ( n35287 & n35290 ) ;
  assign n35292 = ~n35275 & n35291 ;
  assign n35293 = n35275 | n35292 ;
  assign n35294 = n35275 & n35291 ;
  assign n35295 = n35293 & ~n35294 ;
  assign n35296 = n34928 | n34933 ;
  assign n35297 = ( n34928 & n34931 ) | ( n34928 & n35296 ) | ( n34931 & n35296 ) ;
  assign n35298 = n35295 & n35297 ;
  assign n35299 = n35295 | n35297 ;
  assign n35300 = ~n35298 & n35299 ;
  assign n35301 = n8122 & n33526 ;
  assign n35302 = n8115 & n33436 ;
  assign n35303 = n8118 & ~n33423 ;
  assign n35304 = n35302 | n35303 ;
  assign n35305 = n35301 | n35304 ;
  assign n35306 = n8125 & n33545 ;
  assign n35307 = n8125 & ~n33548 ;
  assign n35308 = ( ~n32456 & n35306 ) | ( ~n32456 & n35307 ) | ( n35306 & n35307 ) ;
  assign n35309 = n35305 | n35308 ;
  assign n35310 = n8125 | n35305 ;
  assign n35311 = ( n33536 & n35309 ) | ( n33536 & n35310 ) | ( n35309 & n35310 ) ;
  assign n35312 = x5 | n35311 ;
  assign n35313 = ~x5 & n35311 ;
  assign n35314 = ( ~n35311 & n35312 ) | ( ~n35311 & n35313 ) | ( n35312 & n35313 ) ;
  assign n35315 = ~n35300 & n35314 ;
  assign n35316 = n35300 & ~n35314 ;
  assign n35317 = n35315 | n35316 ;
  assign n35318 = n34951 | n34955 ;
  assign n35319 = ( n34951 & n34953 ) | ( n34951 & n35318 ) | ( n34953 & n35318 ) ;
  assign n35320 = n35317 & ~n35319 ;
  assign n35321 = ~n35317 & n35319 ;
  assign n35322 = n35320 | n35321 ;
  assign n35323 = n35023 | n35024 ;
  assign n35324 = ( n35023 & n35025 ) | ( n35023 & n35323 ) | ( n35025 & n35323 ) ;
  assign n35325 = ( n35023 & n35027 ) | ( n35023 & n35323 ) | ( n35027 & n35323 ) ;
  assign n35326 = ( n32456 & n35324 ) | ( n32456 & n35325 ) | ( n35324 & n35325 ) ;
  assign n35327 = n1065 & ~n23240 ;
  assign n35328 = n1060 & n23227 ;
  assign n35329 = ( n1060 & n23217 ) | ( n1060 & n35328 ) | ( n23217 & n35328 ) ;
  assign n35330 = n35327 | n35329 ;
  assign n35331 = n1057 & ~n23234 ;
  assign n35332 = n1057 & ~n23235 ;
  assign n35333 = ( ~n15882 & n35331 ) | ( ~n15882 & n35332 ) | ( n35331 & n35332 ) ;
  assign n35334 = n35330 | n35333 ;
  assign n35335 = n1062 | n35333 ;
  assign n35336 = n35330 | n35335 ;
  assign n35337 = ( ~n23587 & n35334 ) | ( ~n23587 & n35336 ) | ( n35334 & n35336 ) ;
  assign n35338 = ( n8982 & n34971 ) | ( n8982 & n34975 ) | ( n34971 & n34975 ) ;
  assign n35339 = n8982 & n34971 ;
  assign n35340 = ( ~n34992 & n35338 ) | ( ~n34992 & n35339 ) | ( n35338 & n35339 ) ;
  assign n35341 = n34971 | n34975 ;
  assign n35342 = n8982 | n35341 ;
  assign n35343 = n8982 | n34971 ;
  assign n35344 = ( ~n34992 & n35342 ) | ( ~n34992 & n35343 ) | ( n35342 & n35343 ) ;
  assign n35345 = ~n35340 & n35344 ;
  assign n35346 = n35336 & n35345 ;
  assign n35347 = n35334 & n35345 ;
  assign n35348 = ( ~n23587 & n35346 ) | ( ~n23587 & n35347 ) | ( n35346 & n35347 ) ;
  assign n35349 = n35345 & ~n35347 ;
  assign n35350 = n35345 & ~n35346 ;
  assign n35351 = ( n23587 & n35349 ) | ( n23587 & n35350 ) | ( n35349 & n35350 ) ;
  assign n35352 = ( n35337 & ~n35348 ) | ( n35337 & n35351 ) | ( ~n35348 & n35351 ) ;
  assign n35353 = n34998 | n35352 ;
  assign n35354 = n35004 & ~n35353 ;
  assign n35355 = n34998 & n35352 ;
  assign n35356 = ( ~n35004 & n35352 ) | ( ~n35004 & n35355 ) | ( n35352 & n35355 ) ;
  assign n35357 = n35354 | n35356 ;
  assign n35358 = n35010 & ~n35357 ;
  assign n35359 = ( n35013 & ~n35357 ) | ( n35013 & n35358 ) | ( ~n35357 & n35358 ) ;
  assign n35360 = ( n35012 & ~n35357 ) | ( n35012 & n35358 ) | ( ~n35357 & n35358 ) ;
  assign n35361 = ( n34651 & n35359 ) | ( n34651 & n35360 ) | ( n35359 & n35360 ) ;
  assign n35362 = ( n34649 & n35359 ) | ( n34649 & n35360 ) | ( n35359 & n35360 ) ;
  assign n35363 = ( n28489 & n35361 ) | ( n28489 & n35362 ) | ( n35361 & n35362 ) ;
  assign n35364 = n35010 | n35013 ;
  assign n35365 = n35010 | n35012 ;
  assign n35366 = ( n34649 & n35364 ) | ( n34649 & n35365 ) | ( n35364 & n35365 ) ;
  assign n35367 = n35357 & ~n35366 ;
  assign n35368 = ( n34651 & n35364 ) | ( n34651 & n35365 ) | ( n35364 & n35365 ) ;
  assign n35369 = n35357 & ~n35368 ;
  assign n35370 = ( ~n28489 & n35367 ) | ( ~n28489 & n35369 ) | ( n35367 & n35369 ) ;
  assign n35371 = n35363 | n35370 ;
  assign n35372 = n35021 & ~n35371 ;
  assign n35373 = ~n35021 & n35371 ;
  assign n35374 = n35023 & ~n35373 ;
  assign n35375 = ( n35024 & ~n35373 ) | ( n35024 & n35374 ) | ( ~n35373 & n35374 ) ;
  assign n35376 = ~n35372 & n35375 ;
  assign n35377 = ~n35372 & n35374 ;
  assign n35378 = ( n35025 & n35376 ) | ( n35025 & n35377 ) | ( n35376 & n35377 ) ;
  assign n35379 = ( n35027 & n35376 ) | ( n35027 & n35377 ) | ( n35376 & n35377 ) ;
  assign n35380 = ( n32456 & n35378 ) | ( n32456 & n35379 ) | ( n35378 & n35379 ) ;
  assign n35381 = n35326 & ~n35380 ;
  assign n35382 = n9021 & n34656 ;
  assign n35383 = n9024 & n35021 ;
  assign n35384 = n35382 | n35383 ;
  assign n35385 = n9475 & ~n35371 ;
  assign n35386 = n8970 | n35385 ;
  assign n35387 = n35384 | n35386 ;
  assign n35388 = n35384 | n35385 ;
  assign n35389 = n35372 | n35375 ;
  assign n35390 = n35372 | n35374 ;
  assign n35391 = ( n35025 & n35389 ) | ( n35025 & n35390 ) | ( n35389 & n35390 ) ;
  assign n35392 = n35373 | n35391 ;
  assign n35393 = ~n35388 & n35392 ;
  assign n35394 = ( n35027 & n35389 ) | ( n35027 & n35390 ) | ( n35389 & n35390 ) ;
  assign n35395 = n35373 | n35394 ;
  assign n35396 = ~n35388 & n35395 ;
  assign n35397 = ( n32456 & n35393 ) | ( n32456 & n35396 ) | ( n35393 & n35396 ) ;
  assign n35398 = n35387 & ~n35397 ;
  assign n35399 = ( n35381 & n35387 ) | ( n35381 & n35398 ) | ( n35387 & n35398 ) ;
  assign n35400 = x2 & n35399 ;
  assign n35401 = x2 & ~n35399 ;
  assign n35402 = ( n35399 & ~n35400 ) | ( n35399 & n35401 ) | ( ~n35400 & n35401 ) ;
  assign n35403 = ~n35322 & n35402 ;
  assign n35404 = n35322 & ~n35402 ;
  assign n35405 = n35403 | n35404 ;
  assign n35406 = n35049 | n35053 ;
  assign n35407 = ~n35405 & n35406 ;
  assign n35408 = n35049 | n35055 ;
  assign n35409 = ~n35405 & n35408 ;
  assign n35410 = ( n34300 & n35407 ) | ( n34300 & n35409 ) | ( n35407 & n35409 ) ;
  assign n35411 = n35405 & ~n35406 ;
  assign n35412 = n35405 & ~n35408 ;
  assign n35413 = ( ~n34300 & n35411 ) | ( ~n34300 & n35412 ) | ( n35411 & n35412 ) ;
  assign n35414 = n35410 | n35413 ;
  assign n35415 = n35063 & ~n35414 ;
  assign n35416 = ~n35063 & n35414 ;
  assign n35417 = n35415 | n35416 ;
  assign n35418 = ~n35295 & n35297 ;
  assign n35419 = n35292 | n35418 ;
  assign n35572 = ~n35196 & n35199 ;
  assign n35573 = ( n35196 & n35201 ) | ( n35196 & ~n35572 ) | ( n35201 & ~n35572 ) ;
  assign n35518 = ~n35143 & n35146 ;
  assign n35519 = ( n35143 & n35148 ) | ( n35143 & ~n35518 ) | ( n35148 & ~n35518 ) ;
  assign n35466 = ~n35095 & n35100 ;
  assign n35467 = ( n35095 & n35102 ) | ( n35095 & ~n35466 ) | ( n35102 & ~n35466 ) ;
  assign n35420 = n1057 & n24167 ;
  assign n35421 = n1065 & n23614 ;
  assign n35422 = n1060 & n23316 ;
  assign n35423 = n35421 | n35422 ;
  assign n35424 = n35420 | n35423 ;
  assign n35425 = n1062 | n35422 ;
  assign n35426 = n35421 | n35425 ;
  assign n35427 = n35420 | n35426 ;
  assign n35428 = ( n24182 & n35424 ) | ( n24182 & n35427 ) | ( n35424 & n35427 ) ;
  assign n35429 = n35424 | n35427 ;
  assign n35430 = ( n24175 & n35428 ) | ( n24175 & n35429 ) | ( n35428 & n35429 ) ;
  assign n35431 = n1445 | n4305 ;
  assign n35432 = n2795 | n4153 ;
  assign n35433 = n35431 | n35432 ;
  assign n35434 = n1636 | n7880 ;
  assign n35435 = n929 | n35434 ;
  assign n35436 = ( ~n16784 & n35433 ) | ( ~n16784 & n35435 ) | ( n35433 & n35435 ) ;
  assign n35437 = n2033 & ~n16784 ;
  assign n35438 = ~n35436 & n35437 ;
  assign n35439 = n1221 | n3412 ;
  assign n35440 = n34334 | n35439 ;
  assign n35441 = n246 | n841 ;
  assign n35442 = n193 | n340 ;
  assign n35443 = n35441 | n35442 ;
  assign n35444 = n237 | n435 ;
  assign n35445 = n349 | n413 ;
  assign n35446 = n35444 | n35445 ;
  assign n35447 = n35443 | n35446 ;
  assign n35448 = n35440 | n35447 ;
  assign n35449 = n1304 | n2050 ;
  assign n35450 = n4249 | n35449 ;
  assign n35451 = n168 | n35450 ;
  assign n35452 = n35448 | n35451 ;
  assign n35453 = n11734 | n35452 ;
  assign n35454 = n35438 & ~n35453 ;
  assign n35455 = n354 | n555 ;
  assign n35456 = n5082 | n35455 ;
  assign n35457 = n35454 & ~n35456 ;
  assign n35458 = n35427 & ~n35457 ;
  assign n35459 = n35424 & ~n35457 ;
  assign n35460 = ( n24182 & n35458 ) | ( n24182 & n35459 ) | ( n35458 & n35459 ) ;
  assign n35461 = n35458 | n35459 ;
  assign n35462 = ( n24175 & n35460 ) | ( n24175 & n35461 ) | ( n35460 & n35461 ) ;
  assign n35463 = n35430 & ~n35462 ;
  assign n35464 = n35430 | n35457 ;
  assign n35465 = ~n35463 & n35464 ;
  assign n35468 = ~n35465 & n35467 ;
  assign n35469 = n35467 & ~n35468 ;
  assign n35471 = n1826 & ~n25054 ;
  assign n35472 = n1823 & n24770 ;
  assign n35473 = n35471 | n35472 ;
  assign n35470 = n1829 & ~n25046 ;
  assign n35475 = n1821 | n35470 ;
  assign n35476 = n35473 | n35475 ;
  assign n35474 = n35470 | n35473 ;
  assign n35477 = n35474 & n35476 ;
  assign n35478 = ( ~n25069 & n35476 ) | ( ~n25069 & n35477 ) | ( n35476 & n35477 ) ;
  assign n35479 = ~x29 & n35477 ;
  assign n35480 = ~x29 & n35476 ;
  assign n35481 = ( ~n25069 & n35479 ) | ( ~n25069 & n35480 ) | ( n35479 & n35480 ) ;
  assign n35482 = x29 | n35479 ;
  assign n35483 = x29 | n35480 ;
  assign n35484 = ( ~n25069 & n35482 ) | ( ~n25069 & n35483 ) | ( n35482 & n35483 ) ;
  assign n35485 = ( ~n35478 & n35481 ) | ( ~n35478 & n35484 ) | ( n35481 & n35484 ) ;
  assign n35486 = n35465 | n35467 ;
  assign n35487 = n35485 & ~n35486 ;
  assign n35488 = ( n35469 & n35485 ) | ( n35469 & n35487 ) | ( n35485 & n35487 ) ;
  assign n35489 = ~n35485 & n35486 ;
  assign n35490 = ~n35469 & n35489 ;
  assign n35491 = n35488 | n35490 ;
  assign n35492 = ~n35121 & n35124 ;
  assign n35493 = ( n35121 & n35126 ) | ( n35121 & ~n35492 ) | ( n35126 & ~n35492 ) ;
  assign n35494 = ~n35491 & n35493 ;
  assign n35495 = n35491 & ~n35493 ;
  assign n35496 = n35494 | n35495 ;
  assign n35497 = n2312 & ~n25728 ;
  assign n35498 = n2308 & n26017 ;
  assign n35499 = n35497 | n35498 ;
  assign n35500 = n2315 & ~n26270 ;
  assign n35501 = ~n26263 & n35500 ;
  assign n35503 = n2306 | n35501 ;
  assign n35504 = n35499 | n35503 ;
  assign n35502 = n35499 | n35501 ;
  assign n35505 = n35502 & n35504 ;
  assign n35506 = ( n26571 & n35504 ) | ( n26571 & n35505 ) | ( n35504 & n35505 ) ;
  assign n35507 = x26 & n35505 ;
  assign n35508 = x26 & n35504 ;
  assign n35509 = ( n26571 & n35507 ) | ( n26571 & n35508 ) | ( n35507 & n35508 ) ;
  assign n35510 = x26 & ~n35507 ;
  assign n35511 = x26 & ~n35508 ;
  assign n35512 = ( ~n26571 & n35510 ) | ( ~n26571 & n35511 ) | ( n35510 & n35511 ) ;
  assign n35513 = ( n35506 & ~n35509 ) | ( n35506 & n35512 ) | ( ~n35509 & n35512 ) ;
  assign n35514 = ~n35496 & n35513 ;
  assign n35515 = n35496 | n35514 ;
  assign n35516 = n35496 & n35513 ;
  assign n35517 = n35515 & ~n35516 ;
  assign n35520 = ~n35517 & n35519 ;
  assign n35521 = n35519 & ~n35520 ;
  assign n35522 = n2925 & ~n26526 ;
  assign n35523 = ~n26520 & n35522 ;
  assign n35524 = n2928 & ~n27133 ;
  assign n35525 = ~n27125 & n35524 ;
  assign n35526 = n35523 | n35525 ;
  assign n35527 = n2932 & ~n27371 ;
  assign n35528 = ~n27363 & n35527 ;
  assign n35529 = n35526 | n35528 ;
  assign n35530 = n2936 | n35528 ;
  assign n35531 = n35526 | n35530 ;
  assign n35532 = ( ~n27654 & n35529 ) | ( ~n27654 & n35531 ) | ( n35529 & n35531 ) ;
  assign n35533 = ~x23 & n35531 ;
  assign n35534 = ~x23 & n35529 ;
  assign n35535 = ( ~n27654 & n35533 ) | ( ~n27654 & n35534 ) | ( n35533 & n35534 ) ;
  assign n35536 = x23 | n35534 ;
  assign n35537 = x23 | n35533 ;
  assign n35538 = ( ~n27654 & n35536 ) | ( ~n27654 & n35537 ) | ( n35536 & n35537 ) ;
  assign n35539 = ( ~n35532 & n35535 ) | ( ~n35532 & n35538 ) | ( n35535 & n35538 ) ;
  assign n35540 = n35517 | n35519 ;
  assign n35541 = n35539 & ~n35540 ;
  assign n35542 = ( n35521 & n35539 ) | ( n35521 & n35541 ) | ( n35539 & n35541 ) ;
  assign n35543 = ~n35539 & n35540 ;
  assign n35544 = ~n35521 & n35543 ;
  assign n35545 = n35542 | n35544 ;
  assign n35546 = ~n35169 & n35545 ;
  assign n35547 = ~n35176 & n35546 ;
  assign n35548 = n35169 & ~n35545 ;
  assign n35549 = ( n35176 & ~n35545 ) | ( n35176 & n35548 ) | ( ~n35545 & n35548 ) ;
  assign n35550 = n35547 | n35549 ;
  assign n35551 = n3547 & n28492 ;
  assign n35552 = n3544 & ~n27606 ;
  assign n35553 = ~n27597 & n35552 ;
  assign n35554 = n3541 & ~n28503 ;
  assign n35555 = n28498 & n35554 ;
  assign n35556 = n35553 | n35555 ;
  assign n35557 = n35551 | n35556 ;
  assign n35558 = n3537 | n35557 ;
  assign n35559 = n35557 & n35558 ;
  assign n35560 = ( ~n28749 & n35558 ) | ( ~n28749 & n35559 ) | ( n35558 & n35559 ) ;
  assign n35561 = ~x20 & n35559 ;
  assign n35562 = ~x20 & n35558 ;
  assign n35563 = ( ~n28749 & n35561 ) | ( ~n28749 & n35562 ) | ( n35561 & n35562 ) ;
  assign n35564 = x20 | n35561 ;
  assign n35565 = x20 | n35562 ;
  assign n35566 = ( ~n28749 & n35564 ) | ( ~n28749 & n35565 ) | ( n35564 & n35565 ) ;
  assign n35567 = ( ~n35560 & n35563 ) | ( ~n35560 & n35566 ) | ( n35563 & n35566 ) ;
  assign n35568 = ~n35550 & n35567 ;
  assign n35569 = n35550 | n35568 ;
  assign n35570 = n35550 & n35567 ;
  assign n35571 = n35569 & ~n35570 ;
  assign n35574 = ~n35571 & n35573 ;
  assign n35575 = n35573 & ~n35574 ;
  assign n35576 = n4471 & ~n30199 ;
  assign n35577 = n4466 & ~n28714 ;
  assign n35578 = n4468 & n29620 ;
  assign n35579 = n35577 | n35578 ;
  assign n35580 = n35576 | n35579 ;
  assign n35581 = n4475 | n35576 ;
  assign n35582 = n35579 | n35581 ;
  assign n35583 = ( ~n30299 & n35580 ) | ( ~n30299 & n35582 ) | ( n35580 & n35582 ) ;
  assign n35584 = ~x17 & n35582 ;
  assign n35585 = ~x17 & n35580 ;
  assign n35586 = ( ~n30299 & n35584 ) | ( ~n30299 & n35585 ) | ( n35584 & n35585 ) ;
  assign n35587 = x17 | n35585 ;
  assign n35588 = x17 | n35584 ;
  assign n35589 = ( ~n30299 & n35587 ) | ( ~n30299 & n35588 ) | ( n35587 & n35588 ) ;
  assign n35590 = ( ~n35583 & n35586 ) | ( ~n35583 & n35589 ) | ( n35586 & n35589 ) ;
  assign n35591 = n35571 | n35573 ;
  assign n35592 = n35590 & ~n35591 ;
  assign n35593 = ( n35575 & n35590 ) | ( n35575 & n35592 ) | ( n35590 & n35592 ) ;
  assign n35594 = ~n35590 & n35591 ;
  assign n35595 = ~n35575 & n35594 ;
  assign n35596 = n35593 | n35595 ;
  assign n35597 = ~n35218 & n35220 ;
  assign n35598 = n35596 & n35597 ;
  assign n35599 = ~n35218 & n35596 ;
  assign n35600 = ( ~n35222 & n35598 ) | ( ~n35222 & n35599 ) | ( n35598 & n35599 ) ;
  assign n35601 = n35596 | n35597 ;
  assign n35602 = n35218 & ~n35596 ;
  assign n35603 = ( n35222 & ~n35601 ) | ( n35222 & n35602 ) | ( ~n35601 & n35602 ) ;
  assign n35604 = n35600 | n35603 ;
  assign n35606 = n5237 & n30212 ;
  assign n35607 = n5231 & ~n30186 ;
  assign n35608 = n35606 | n35607 ;
  assign n35605 = n5234 & ~n31309 ;
  assign n35610 = n5227 | n35605 ;
  assign n35611 = n35608 | n35610 ;
  assign n35609 = n35605 | n35608 ;
  assign n35612 = n35609 & n35611 ;
  assign n35613 = ( n31404 & n35611 ) | ( n31404 & n35612 ) | ( n35611 & n35612 ) ;
  assign n35614 = x14 & n35612 ;
  assign n35615 = x14 & n35611 ;
  assign n35616 = ( n31404 & n35614 ) | ( n31404 & n35615 ) | ( n35614 & n35615 ) ;
  assign n35617 = x14 & ~n35614 ;
  assign n35618 = x14 & ~n35615 ;
  assign n35619 = ( ~n31404 & n35617 ) | ( ~n31404 & n35618 ) | ( n35617 & n35618 ) ;
  assign n35620 = ( n35613 & ~n35616 ) | ( n35613 & n35619 ) | ( ~n35616 & n35619 ) ;
  assign n35621 = ~n35604 & n35620 ;
  assign n35622 = n35604 | n35621 ;
  assign n35623 = n35604 & n35620 ;
  assign n35624 = n35622 & ~n35623 ;
  assign n35625 = ~n35242 & n35245 ;
  assign n35626 = ( n35065 & n35242 ) | ( n35065 & ~n35625 ) | ( n35242 & ~n35625 ) ;
  assign n35627 = n35624 | n35626 ;
  assign n35628 = n35624 & n35626 ;
  assign n35629 = n35627 & ~n35628 ;
  assign n35630 = n6122 & n32306 ;
  assign n35631 = n6125 & ~n31323 ;
  assign n35632 = n6119 & n31295 ;
  assign n35633 = n35631 | n35632 ;
  assign n35634 = n35630 | n35633 ;
  assign n35635 = n6115 | n35630 ;
  assign n35636 = n35633 | n35635 ;
  assign n35637 = ( ~n32525 & n35634 ) | ( ~n32525 & n35636 ) | ( n35634 & n35636 ) ;
  assign n35638 = ~x11 & n35636 ;
  assign n35639 = ~x11 & n35634 ;
  assign n35640 = ( ~n32525 & n35638 ) | ( ~n32525 & n35639 ) | ( n35638 & n35639 ) ;
  assign n35641 = x11 | n35639 ;
  assign n35642 = x11 | n35638 ;
  assign n35643 = ( ~n32525 & n35641 ) | ( ~n32525 & n35642 ) | ( n35641 & n35642 ) ;
  assign n35644 = ( ~n35637 & n35640 ) | ( ~n35637 & n35643 ) | ( n35640 & n35643 ) ;
  assign n35645 = ~n35629 & n35644 ;
  assign n35646 = n35629 & ~n35644 ;
  assign n35647 = n35645 | n35646 ;
  assign n35648 = ~n35266 & n35647 ;
  assign n35649 = ~n35274 & n35648 ;
  assign n35650 = n35266 & ~n35647 ;
  assign n35651 = ( n35274 & ~n35647 ) | ( n35274 & n35650 ) | ( ~n35647 & n35650 ) ;
  assign n35652 = n35649 | n35651 ;
  assign n35653 = n7079 & n33436 ;
  assign n35654 = n7074 & n32293 ;
  assign n35655 = n7068 & ~n32442 ;
  assign n35656 = n35654 | n35655 ;
  assign n35657 = n35653 | n35656 ;
  assign n35658 = n33441 & ~n35657 ;
  assign n35659 = ( n32456 & ~n35657 ) | ( n32456 & n35658 ) | ( ~n35657 & n35658 ) ;
  assign n35660 = ~n34271 & n35659 ;
  assign n35661 = n7078 | n35653 ;
  assign n35662 = n35656 | n35661 ;
  assign n35663 = ~n35660 & n35662 ;
  assign n35664 = x8 & n35662 ;
  assign n35665 = ~n35660 & n35664 ;
  assign n35666 = x8 & ~n35664 ;
  assign n35667 = ( x8 & n35660 ) | ( x8 & n35666 ) | ( n35660 & n35666 ) ;
  assign n35668 = ( n35663 & ~n35665 ) | ( n35663 & n35667 ) | ( ~n35665 & n35667 ) ;
  assign n35669 = ~n35652 & n35668 ;
  assign n35670 = n35652 | n35669 ;
  assign n35671 = n35652 & n35668 ;
  assign n35672 = n35670 & ~n35671 ;
  assign n35673 = n35419 & ~n35672 ;
  assign n35674 = n35419 & ~n35673 ;
  assign n35675 = n35419 | n35672 ;
  assign n35676 = ~n35674 & n35675 ;
  assign n35677 = n8122 & n34656 ;
  assign n35678 = n8115 & ~n33423 ;
  assign n35679 = n8118 & n33526 ;
  assign n35680 = n35678 | n35679 ;
  assign n35681 = n35677 | n35680 ;
  assign n35682 = n8125 | n35677 ;
  assign n35683 = n35680 | n35682 ;
  assign n35684 = ( n34667 & n35681 ) | ( n34667 & n35683 ) | ( n35681 & n35683 ) ;
  assign n35685 = x5 & n35683 ;
  assign n35686 = x5 & n35681 ;
  assign n35687 = ( n34667 & n35685 ) | ( n34667 & n35686 ) | ( n35685 & n35686 ) ;
  assign n35688 = x5 & ~n35686 ;
  assign n35689 = x5 & ~n35685 ;
  assign n35690 = ( ~n34667 & n35688 ) | ( ~n34667 & n35689 ) | ( n35688 & n35689 ) ;
  assign n35691 = ( n35684 & ~n35687 ) | ( n35684 & n35690 ) | ( ~n35687 & n35690 ) ;
  assign n35692 = ~n35675 & n35691 ;
  assign n35693 = ( n35674 & n35691 ) | ( n35674 & n35692 ) | ( n35691 & n35692 ) ;
  assign n35694 = n35676 | n35693 ;
  assign n35695 = n35675 & n35691 ;
  assign n35696 = ~n35674 & n35695 ;
  assign n35697 = n35694 & ~n35696 ;
  assign n35698 = n35315 | n35321 ;
  assign n35699 = n35697 & ~n35698 ;
  assign n35700 = ~n35697 & n35698 ;
  assign n35701 = n35699 | n35700 ;
  assign n35702 = n1057 | n1065 ;
  assign n35703 = ~n23234 & n35702 ;
  assign n35704 = ~n23235 & n35702 ;
  assign n35705 = ( ~n15882 & n35703 ) | ( ~n15882 & n35704 ) | ( n35703 & n35704 ) ;
  assign n35706 = n1060 | n35703 ;
  assign n35707 = n1060 | n35704 ;
  assign n35708 = ( ~n15882 & n35706 ) | ( ~n15882 & n35707 ) | ( n35706 & n35707 ) ;
  assign n35709 = ( ~n23240 & n35705 ) | ( ~n23240 & n35708 ) | ( n35705 & n35708 ) ;
  assign n35710 = n1062 & ~n24135 ;
  assign n35711 = n1062 & ~n23240 ;
  assign n35712 = ( ~n23575 & n35710 ) | ( ~n23575 & n35711 ) | ( n35710 & n35711 ) ;
  assign n35713 = ( ~n23577 & n35710 ) | ( ~n23577 & n35711 ) | ( n35710 & n35711 ) ;
  assign n35714 = ( n21554 & n35712 ) | ( n21554 & n35713 ) | ( n35712 & n35713 ) ;
  assign n35715 = n35709 | n35714 ;
  assign n35716 = n8982 & ~n35715 ;
  assign n35717 = n35712 & n35713 ;
  assign n35718 = n35709 | n35717 ;
  assign n35719 = n8982 & ~n35718 ;
  assign n35720 = ( n21584 & n35716 ) | ( n21584 & n35719 ) | ( n35716 & n35719 ) ;
  assign n35721 = ~n8982 & n35715 ;
  assign n35722 = ~n8982 & n35718 ;
  assign n35723 = ( ~n21584 & n35721 ) | ( ~n21584 & n35722 ) | ( n35721 & n35722 ) ;
  assign n35724 = n35720 | n35723 ;
  assign n35725 = n35340 | n35347 ;
  assign n35726 = n35340 | n35346 ;
  assign n35727 = ( ~n23587 & n35725 ) | ( ~n23587 & n35726 ) | ( n35725 & n35726 ) ;
  assign n35728 = n35724 | n35727 ;
  assign n35729 = n35724 & n35727 ;
  assign n35730 = n35728 & ~n35729 ;
  assign n35731 = n35356 | n35358 ;
  assign n35732 = ~n35356 & n35357 ;
  assign n35733 = ( n35013 & n35731 ) | ( n35013 & ~n35732 ) | ( n35731 & ~n35732 ) ;
  assign n35734 = n35730 & n35733 ;
  assign n35735 = n35356 & n35730 ;
  assign n35736 = ( n35360 & n35730 ) | ( n35360 & n35735 ) | ( n35730 & n35735 ) ;
  assign n35737 = ( n34651 & n35734 ) | ( n34651 & n35736 ) | ( n35734 & n35736 ) ;
  assign n35738 = ( n34649 & n35734 ) | ( n34649 & n35736 ) | ( n35734 & n35736 ) ;
  assign n35739 = ( n28489 & n35737 ) | ( n28489 & n35738 ) | ( n35737 & n35738 ) ;
  assign n35740 = n35356 | n35360 ;
  assign n35741 = ( n34649 & n35733 ) | ( n34649 & n35740 ) | ( n35733 & n35740 ) ;
  assign n35742 = n35730 | n35741 ;
  assign n35743 = ( n34651 & n35733 ) | ( n34651 & n35740 ) | ( n35733 & n35740 ) ;
  assign n35744 = n35730 | n35743 ;
  assign n35745 = ( n28489 & n35742 ) | ( n28489 & n35744 ) | ( n35742 & n35744 ) ;
  assign n35746 = ~n35739 & n35745 ;
  assign n35747 = n35371 & ~n35746 ;
  assign n35748 = ~n35371 & n35746 ;
  assign n35749 = n35747 | n35748 ;
  assign n35750 = n35390 & ~n35749 ;
  assign n35751 = n35372 & ~n35749 ;
  assign n35752 = ( n35375 & ~n35749 ) | ( n35375 & n35751 ) | ( ~n35749 & n35751 ) ;
  assign n35753 = ( n35025 & n35750 ) | ( n35025 & n35752 ) | ( n35750 & n35752 ) ;
  assign n35754 = ( n35027 & n35750 ) | ( n35027 & n35752 ) | ( n35750 & n35752 ) ;
  assign n35755 = ( n32456 & n35753 ) | ( n32456 & n35754 ) | ( n35753 & n35754 ) ;
  assign n35756 = ~n35391 & n35749 ;
  assign n35757 = ~n35394 & n35749 ;
  assign n35758 = ( ~n32456 & n35756 ) | ( ~n32456 & n35757 ) | ( n35756 & n35757 ) ;
  assign n35759 = n35755 | n35758 ;
  assign n35761 = n9021 & n35021 ;
  assign n35762 = n9024 & ~n35371 ;
  assign n35763 = n35761 | n35762 ;
  assign n35760 = n9475 & n35746 ;
  assign n35765 = n8970 | n35760 ;
  assign n35766 = n35763 | n35765 ;
  assign n35764 = n35760 | n35763 ;
  assign n35767 = n35764 & n35766 ;
  assign n35768 = ( ~n35759 & n35766 ) | ( ~n35759 & n35767 ) | ( n35766 & n35767 ) ;
  assign n35769 = ~x2 & n35767 ;
  assign n35770 = ~x2 & n35766 ;
  assign n35771 = ( ~n35759 & n35769 ) | ( ~n35759 & n35770 ) | ( n35769 & n35770 ) ;
  assign n35772 = x2 | n35769 ;
  assign n35773 = x2 | n35770 ;
  assign n35774 = ( ~n35759 & n35772 ) | ( ~n35759 & n35773 ) | ( n35772 & n35773 ) ;
  assign n35775 = ( ~n35768 & n35771 ) | ( ~n35768 & n35774 ) | ( n35771 & n35774 ) ;
  assign n35776 = ~n35701 & n35775 ;
  assign n35777 = n35701 & ~n35775 ;
  assign n35778 = n35776 | n35777 ;
  assign n35779 = n35403 | n35409 ;
  assign n35780 = n35403 | n35407 ;
  assign n35781 = ( n34300 & n35779 ) | ( n34300 & n35780 ) | ( n35779 & n35780 ) ;
  assign n35782 = ~n35778 & n35781 ;
  assign n35783 = n35778 & ~n35781 ;
  assign n35784 = n35782 | n35783 ;
  assign n35785 = ~n35415 & n35784 ;
  assign n35786 = n35414 | n35784 ;
  assign n35787 = n35063 & ~n35786 ;
  assign n35788 = n35785 | n35787 ;
  assign n36025 = ~n35669 & n35672 ;
  assign n36026 = ( n35419 & n35669 ) | ( n35419 & ~n36025 ) | ( n35669 & ~n36025 ) ;
  assign n35789 = ~n35621 & n35624 ;
  assign n35790 = ( n35621 & n35626 ) | ( n35621 & ~n35789 ) | ( n35626 & ~n35789 ) ;
  assign n35929 = ~n35568 & n35571 ;
  assign n35930 = ( n35568 & n35573 ) | ( n35568 & ~n35929 ) | ( n35573 & ~n35929 ) ;
  assign n35877 = ~n35514 & n35517 ;
  assign n35878 = ( n35514 & n35519 ) | ( n35514 & ~n35877 ) | ( n35519 & ~n35877 ) ;
  assign n35791 = n1057 & ~n25054 ;
  assign n35792 = n1065 & n24167 ;
  assign n35793 = n1060 & n23614 ;
  assign n35794 = n35792 | n35793 ;
  assign n35795 = n35791 | n35794 ;
  assign n35796 = n1062 | n35793 ;
  assign n35797 = n35792 | n35796 ;
  assign n35798 = n35791 | n35797 ;
  assign n35799 = ( ~n25122 & n35795 ) | ( ~n25122 & n35798 ) | ( n35795 & n35798 ) ;
  assign n35800 = n13023 | n13027 ;
  assign n35801 = n1771 | n5072 ;
  assign n35802 = n6914 | n35801 ;
  assign n35803 = n12291 | n18464 ;
  assign n35804 = n35802 | n35803 ;
  assign n35805 = n18233 | n35804 ;
  assign n35806 = n12286 & ~n35805 ;
  assign n35807 = ~n35800 & n35806 ;
  assign n35808 = n273 | n333 ;
  assign n35809 = n390 | n35808 ;
  assign n35810 = n138 | n246 ;
  assign n35811 = n4246 | n35810 ;
  assign n35812 = n112 | n458 ;
  assign n35813 = n401 | n35812 ;
  assign n35814 = n35811 | n35813 ;
  assign n35815 = n277 | n600 ;
  assign n35816 = n198 | n35815 ;
  assign n35817 = n35814 | n35816 ;
  assign n35818 = n35809 | n35817 ;
  assign n35819 = n35807 & ~n35818 ;
  assign n35820 = n35791 & ~n35819 ;
  assign n35821 = ( n35797 & ~n35819 ) | ( n35797 & n35820 ) | ( ~n35819 & n35820 ) ;
  assign n35822 = ( n35794 & ~n35819 ) | ( n35794 & n35820 ) | ( ~n35819 & n35820 ) ;
  assign n35823 = ( ~n25122 & n35821 ) | ( ~n25122 & n35822 ) | ( n35821 & n35822 ) ;
  assign n35824 = n35799 & ~n35823 ;
  assign n35825 = n35798 | n35819 ;
  assign n35826 = n35795 | n35819 ;
  assign n35827 = ( ~n25122 & n35825 ) | ( ~n25122 & n35826 ) | ( n35825 & n35826 ) ;
  assign n35828 = ~n35824 & n35827 ;
  assign n35829 = ~n35462 & n35465 ;
  assign n35830 = ( n35462 & n35467 ) | ( n35462 & ~n35829 ) | ( n35467 & ~n35829 ) ;
  assign n35831 = ~n35828 & n35830 ;
  assign n35832 = n35828 & ~n35830 ;
  assign n35833 = n35831 | n35832 ;
  assign n35834 = n1826 & n24770 ;
  assign n35835 = n1823 & ~n25046 ;
  assign n35836 = n35834 | n35835 ;
  assign n35837 = n1829 & ~n25728 ;
  assign n35838 = n1821 | n35837 ;
  assign n35839 = n35836 | n35838 ;
  assign n35840 = n35836 | n35837 ;
  assign n35841 = n25740 | n35840 ;
  assign n35842 = n25731 | n35840 ;
  assign n35843 = ( ~n25441 & n35841 ) | ( ~n25441 & n35842 ) | ( n35841 & n35842 ) ;
  assign n35844 = n35839 & n35843 ;
  assign n35845 = ( n25733 & n35839 ) | ( n25733 & n35844 ) | ( n35839 & n35844 ) ;
  assign n35846 = ~x29 & n35845 ;
  assign n35847 = x29 | n35845 ;
  assign n35848 = ( ~n35845 & n35846 ) | ( ~n35845 & n35847 ) | ( n35846 & n35847 ) ;
  assign n35849 = ~n35833 & n35848 ;
  assign n35850 = n35833 & ~n35848 ;
  assign n35851 = n35849 | n35850 ;
  assign n35852 = ~n35488 & n35491 ;
  assign n35853 = ( n35488 & n35493 ) | ( n35488 & ~n35852 ) | ( n35493 & ~n35852 ) ;
  assign n35854 = ~n35851 & n35853 ;
  assign n35855 = n35851 & ~n35853 ;
  assign n35856 = n35854 | n35855 ;
  assign n35857 = n2312 & n26017 ;
  assign n35858 = n2308 & ~n26270 ;
  assign n35859 = ~n26263 & n35858 ;
  assign n35860 = n35857 | n35859 ;
  assign n35861 = n2315 & ~n26526 ;
  assign n35862 = ~n26520 & n35861 ;
  assign n35864 = n2306 | n35862 ;
  assign n35865 = n35860 | n35864 ;
  assign n35863 = n35860 | n35862 ;
  assign n35866 = n35863 & n35865 ;
  assign n35867 = ( ~n26555 & n35865 ) | ( ~n26555 & n35866 ) | ( n35865 & n35866 ) ;
  assign n35868 = ( n26528 & n35865 ) | ( n26528 & n35866 ) | ( n35865 & n35866 ) ;
  assign n35869 = ( ~n26543 & n35867 ) | ( ~n26543 & n35868 ) | ( n35867 & n35868 ) ;
  assign n35870 = ~x26 & n35869 ;
  assign n35871 = x26 | n35869 ;
  assign n35872 = ( ~n35869 & n35870 ) | ( ~n35869 & n35871 ) | ( n35870 & n35871 ) ;
  assign n35873 = ~n35856 & n35872 ;
  assign n35874 = n35856 | n35873 ;
  assign n35875 = n35856 & n35872 ;
  assign n35876 = n35874 & ~n35875 ;
  assign n35879 = ~n35876 & n35878 ;
  assign n35880 = n35878 & ~n35879 ;
  assign n35881 = n35876 | n35878 ;
  assign n35882 = ~n35880 & n35881 ;
  assign n35883 = n2925 & ~n27133 ;
  assign n35884 = ~n27125 & n35883 ;
  assign n35885 = n2928 & ~n27371 ;
  assign n35886 = ~n27363 & n35885 ;
  assign n35887 = n35884 | n35886 ;
  assign n35888 = n2932 & ~n27606 ;
  assign n35889 = ~n27597 & n35888 ;
  assign n35890 = n35887 | n35889 ;
  assign n35891 = n2936 & n27630 ;
  assign n35892 = ~n27625 & n35891 ;
  assign n35893 = ( n2936 & ~n27634 ) | ( n2936 & n35892 ) | ( ~n27634 & n35892 ) ;
  assign n35894 = n35890 | n35893 ;
  assign n35895 = x23 | n35890 ;
  assign n35896 = n35893 | n35895 ;
  assign n35897 = ~x23 & n35895 ;
  assign n35898 = ( ~x23 & n35893 ) | ( ~x23 & n35897 ) | ( n35893 & n35897 ) ;
  assign n35899 = ( ~n35894 & n35896 ) | ( ~n35894 & n35898 ) | ( n35896 & n35898 ) ;
  assign n35900 = ~n35881 & n35899 ;
  assign n35901 = ( n35880 & n35899 ) | ( n35880 & n35900 ) | ( n35899 & n35900 ) ;
  assign n35902 = n35882 | n35901 ;
  assign n35903 = n35881 & n35899 ;
  assign n35904 = ~n35880 & n35903 ;
  assign n35905 = n35902 & ~n35904 ;
  assign n35906 = n35542 | n35549 ;
  assign n35907 = n35905 & ~n35906 ;
  assign n35908 = ~n35905 & n35906 ;
  assign n35909 = n35907 | n35908 ;
  assign n35910 = n3541 & n28492 ;
  assign n35911 = n3544 & ~n28503 ;
  assign n35912 = n28498 & n35911 ;
  assign n35913 = n35910 | n35912 ;
  assign n35914 = n3547 & ~n28714 ;
  assign n35915 = n3537 | n35914 ;
  assign n35916 = n35913 | n35915 ;
  assign n35917 = n35913 | n35914 ;
  assign n35918 = n28731 & ~n35917 ;
  assign n35919 = ( n28518 & ~n35917 ) | ( n28518 & n35918 ) | ( ~n35917 & n35918 ) ;
  assign n35920 = n35916 & ~n35919 ;
  assign n35921 = ( n28720 & n35916 ) | ( n28720 & n35920 ) | ( n35916 & n35920 ) ;
  assign n35922 = x20 & n35921 ;
  assign n35923 = x20 & ~n35921 ;
  assign n35924 = ( n35921 & ~n35922 ) | ( n35921 & n35923 ) | ( ~n35922 & n35923 ) ;
  assign n35925 = ~n35909 & n35924 ;
  assign n35926 = n35909 | n35925 ;
  assign n35927 = n35909 & n35924 ;
  assign n35928 = n35926 & ~n35927 ;
  assign n35931 = ~n35928 & n35930 ;
  assign n35932 = n35930 & ~n35931 ;
  assign n35933 = n4471 & n30212 ;
  assign n35934 = n4466 & n29620 ;
  assign n35935 = n4468 & ~n30199 ;
  assign n35936 = n35934 | n35935 ;
  assign n35937 = n35933 | n35936 ;
  assign n35938 = n4475 & ~n30266 ;
  assign n35939 = ( n4475 & n30276 ) | ( n4475 & n35938 ) | ( n30276 & n35938 ) ;
  assign n35940 = n35937 | n35939 ;
  assign n35941 = x17 | n35937 ;
  assign n35942 = n35939 | n35941 ;
  assign n35943 = ~x17 & n35941 ;
  assign n35944 = ( ~x17 & n35939 ) | ( ~x17 & n35943 ) | ( n35939 & n35943 ) ;
  assign n35945 = ( ~n35940 & n35942 ) | ( ~n35940 & n35944 ) | ( n35942 & n35944 ) ;
  assign n35946 = n35928 | n35930 ;
  assign n35947 = n35945 & ~n35946 ;
  assign n35948 = ( n35932 & n35945 ) | ( n35932 & n35947 ) | ( n35945 & n35947 ) ;
  assign n35949 = ~n35945 & n35946 ;
  assign n35950 = ~n35932 & n35949 ;
  assign n35951 = n35948 | n35950 ;
  assign n35952 = ~n35593 & n35951 ;
  assign n35953 = ~n35603 & n35952 ;
  assign n35954 = n35593 & ~n35951 ;
  assign n35955 = ( n35603 & ~n35951 ) | ( n35603 & n35954 ) | ( ~n35951 & n35954 ) ;
  assign n35956 = n35953 | n35955 ;
  assign n35957 = n5237 & ~n30186 ;
  assign n35958 = n5231 & ~n31309 ;
  assign n35959 = n35957 | n35958 ;
  assign n35960 = n5234 & ~n31323 ;
  assign n35961 = n5227 | n35960 ;
  assign n35962 = n35959 | n35961 ;
  assign n35963 = n35959 | n35960 ;
  assign n35964 = n31384 | n35963 ;
  assign n35965 = n31386 | n35963 ;
  assign n35966 = ( ~n30232 & n35964 ) | ( ~n30232 & n35965 ) | ( n35964 & n35965 ) ;
  assign n35967 = n35962 & n35966 ;
  assign n35968 = ( ~n31376 & n35962 ) | ( ~n31376 & n35967 ) | ( n35962 & n35967 ) ;
  assign n35969 = x14 & n35968 ;
  assign n35970 = x14 & ~n35968 ;
  assign n35971 = ( n35968 & ~n35969 ) | ( n35968 & n35970 ) | ( ~n35969 & n35970 ) ;
  assign n35972 = ~n35956 & n35971 ;
  assign n35973 = n35956 | n35972 ;
  assign n35974 = n35956 & n35971 ;
  assign n35975 = n35973 & ~n35974 ;
  assign n35976 = n35789 | n35975 ;
  assign n35977 = n35621 & ~n35975 ;
  assign n35978 = ( n35626 & ~n35976 ) | ( n35626 & n35977 ) | ( ~n35976 & n35977 ) ;
  assign n35979 = n35790 & ~n35978 ;
  assign n35980 = n6122 & n32293 ;
  assign n35981 = n6125 & n31295 ;
  assign n35982 = n6119 & n32306 ;
  assign n35983 = n35981 | n35982 ;
  assign n35984 = n35980 | n35983 ;
  assign n35985 = n6115 & n32497 ;
  assign n35986 = ( n6115 & n32494 ) | ( n6115 & n35985 ) | ( n32494 & n35985 ) ;
  assign n35987 = n35984 | n35986 ;
  assign n35988 = x11 | n35984 ;
  assign n35989 = n35986 | n35988 ;
  assign n35990 = ~x11 & n35988 ;
  assign n35991 = ( ~x11 & n35986 ) | ( ~x11 & n35990 ) | ( n35986 & n35990 ) ;
  assign n35992 = ( ~n35987 & n35989 ) | ( ~n35987 & n35991 ) | ( n35989 & n35991 ) ;
  assign n35993 = n35789 & ~n35975 ;
  assign n35994 = n35621 | n35975 ;
  assign n35995 = ( n35626 & ~n35993 ) | ( n35626 & n35994 ) | ( ~n35993 & n35994 ) ;
  assign n35996 = n35992 & ~n35995 ;
  assign n35997 = ( n35979 & n35992 ) | ( n35979 & n35996 ) | ( n35992 & n35996 ) ;
  assign n35998 = ~n35992 & n35995 ;
  assign n35999 = ~n35979 & n35998 ;
  assign n36000 = n35997 | n35999 ;
  assign n36001 = ~n35645 & n36000 ;
  assign n36002 = ~n35651 & n36001 ;
  assign n36003 = n35645 & ~n36000 ;
  assign n36004 = ( n35651 & ~n36000 ) | ( n35651 & n36003 ) | ( ~n36000 & n36003 ) ;
  assign n36005 = n36002 | n36004 ;
  assign n36006 = n7074 & ~n32442 ;
  assign n36007 = n7068 & n33436 ;
  assign n36008 = n36006 | n36007 ;
  assign n36009 = n7079 & ~n33423 ;
  assign n36010 = n7078 | n36009 ;
  assign n36011 = n36008 | n36010 ;
  assign n36012 = n36008 | n36009 ;
  assign n36013 = n33575 | n36012 ;
  assign n36014 = n33577 & ~n36012 ;
  assign n36015 = ( n32456 & ~n36013 ) | ( n32456 & n36014 ) | ( ~n36013 & n36014 ) ;
  assign n36016 = n36011 & ~n36015 ;
  assign n36017 = ( n33567 & n36011 ) | ( n33567 & n36016 ) | ( n36011 & n36016 ) ;
  assign n36018 = x8 & n36017 ;
  assign n36019 = x8 & ~n36017 ;
  assign n36020 = ( n36017 & ~n36018 ) | ( n36017 & n36019 ) | ( ~n36018 & n36019 ) ;
  assign n36021 = ~n36005 & n36020 ;
  assign n36022 = n36005 | n36021 ;
  assign n36023 = n36005 & n36020 ;
  assign n36024 = n36022 & ~n36023 ;
  assign n36027 = ~n36024 & n36026 ;
  assign n36028 = n36026 & ~n36027 ;
  assign n36029 = n36024 | n36026 ;
  assign n36030 = ~n36028 & n36029 ;
  assign n36031 = n8122 & n35021 ;
  assign n36032 = n8115 & n33526 ;
  assign n36033 = n8118 & n34656 ;
  assign n36034 = n36032 | n36033 ;
  assign n36035 = n36031 | n36034 ;
  assign n36036 = n8125 | n36031 ;
  assign n36037 = n36034 | n36036 ;
  assign n36038 = ( n35033 & n36035 ) | ( n35033 & n36037 ) | ( n36035 & n36037 ) ;
  assign n36039 = x5 & n36037 ;
  assign n36040 = x5 & n36035 ;
  assign n36041 = ( n35033 & n36039 ) | ( n35033 & n36040 ) | ( n36039 & n36040 ) ;
  assign n36042 = x5 & ~n36040 ;
  assign n36043 = x5 & ~n36039 ;
  assign n36044 = ( ~n35033 & n36042 ) | ( ~n35033 & n36043 ) | ( n36042 & n36043 ) ;
  assign n36045 = ( n36038 & ~n36041 ) | ( n36038 & n36044 ) | ( ~n36041 & n36044 ) ;
  assign n36046 = ~n36029 & n36045 ;
  assign n36047 = ( n36028 & n36045 ) | ( n36028 & n36046 ) | ( n36045 & n36046 ) ;
  assign n36048 = n36030 | n36047 ;
  assign n36049 = n36029 & n36045 ;
  assign n36050 = ~n36028 & n36049 ;
  assign n36051 = n36048 & ~n36050 ;
  assign n36052 = n35693 | n35698 ;
  assign n36053 = ( n35693 & ~n35697 ) | ( n35693 & n36052 ) | ( ~n35697 & n36052 ) ;
  assign n36054 = n36051 & ~n36053 ;
  assign n36055 = ~n36051 & n36053 ;
  assign n36056 = n36054 | n36055 ;
  assign n36057 = n35748 | n35752 ;
  assign n36058 = ~n35748 & n35749 ;
  assign n36059 = ( n35390 & n35748 ) | ( n35390 & ~n36058 ) | ( n35748 & ~n36058 ) ;
  assign n36060 = ( n35025 & n36057 ) | ( n35025 & n36059 ) | ( n36057 & n36059 ) ;
  assign n36061 = ( n35027 & n36057 ) | ( n35027 & n36059 ) | ( n36057 & n36059 ) ;
  assign n36062 = ( n32456 & n36060 ) | ( n32456 & n36061 ) | ( n36060 & n36061 ) ;
  assign n36063 = n35729 | n35730 ;
  assign n36064 = ( n35729 & n35733 ) | ( n35729 & n36063 ) | ( n35733 & n36063 ) ;
  assign n36065 = n35729 | n35735 ;
  assign n36066 = ( n35360 & n36063 ) | ( n35360 & n36065 ) | ( n36063 & n36065 ) ;
  assign n36067 = ( n34651 & n36064 ) | ( n34651 & n36066 ) | ( n36064 & n36066 ) ;
  assign n36068 = ( n34649 & n36064 ) | ( n34649 & n36066 ) | ( n36064 & n36066 ) ;
  assign n36069 = ( n28489 & n36067 ) | ( n28489 & n36068 ) | ( n36067 & n36068 ) ;
  assign n36070 = x31 | n33 ;
  assign n36071 = ~n23234 & n36070 ;
  assign n36072 = ~n23235 & n36070 ;
  assign n36073 = ( ~n15882 & n36071 ) | ( ~n15882 & n36072 ) | ( n36071 & n36072 ) ;
  assign n36074 = n35720 & ~n36073 ;
  assign n36075 = n35720 | n36073 ;
  assign n36076 = ( ~n35720 & n36074 ) | ( ~n35720 & n36075 ) | ( n36074 & n36075 ) ;
  assign n36077 = n36068 & n36076 ;
  assign n36078 = n36067 & n36076 ;
  assign n36079 = ( n28489 & n36077 ) | ( n28489 & n36078 ) | ( n36077 & n36078 ) ;
  assign n36080 = n36076 & ~n36078 ;
  assign n36081 = n36076 & ~n36077 ;
  assign n36082 = ( ~n28489 & n36080 ) | ( ~n28489 & n36081 ) | ( n36080 & n36081 ) ;
  assign n36083 = ( n36069 & ~n36079 ) | ( n36069 & n36082 ) | ( ~n36079 & n36082 ) ;
  assign n36084 = n35746 & n36083 ;
  assign n36085 = n35746 | n36083 ;
  assign n36086 = n35748 & n36085 ;
  assign n36087 = ~n36084 & n36086 ;
  assign n36088 = ~n36084 & n36085 ;
  assign n36089 = ( n35752 & n36087 ) | ( n35752 & n36088 ) | ( n36087 & n36088 ) ;
  assign n36090 = n36059 & n36088 ;
  assign n36091 = ( n35025 & n36089 ) | ( n35025 & n36090 ) | ( n36089 & n36090 ) ;
  assign n36092 = ( n35027 & n36089 ) | ( n35027 & n36090 ) | ( n36089 & n36090 ) ;
  assign n36093 = ( n32456 & n36091 ) | ( n32456 & n36092 ) | ( n36091 & n36092 ) ;
  assign n36094 = n36062 & ~n36093 ;
  assign n36096 = n9021 & ~n35371 ;
  assign n36097 = n9024 & n35746 ;
  assign n36098 = n36096 | n36097 ;
  assign n36095 = n9475 & n36083 ;
  assign n36100 = n8970 | n36095 ;
  assign n36101 = n36098 | n36100 ;
  assign n36099 = n36095 | n36098 ;
  assign n36102 = n36099 & n36101 ;
  assign n36103 = n36084 | n36091 ;
  assign n36104 = n36085 & ~n36103 ;
  assign n36105 = n36084 | n36092 ;
  assign n36106 = n36085 & ~n36105 ;
  assign n36107 = ( ~n32456 & n36104 ) | ( ~n32456 & n36106 ) | ( n36104 & n36106 ) ;
  assign n36108 = ( n36101 & n36102 ) | ( n36101 & n36107 ) | ( n36102 & n36107 ) ;
  assign n36109 = n36101 | n36102 ;
  assign n36110 = ( n36094 & n36108 ) | ( n36094 & n36109 ) | ( n36108 & n36109 ) ;
  assign n36111 = x2 & n36110 ;
  assign n36112 = x2 & ~n36110 ;
  assign n36113 = ( n36110 & ~n36111 ) | ( n36110 & n36112 ) | ( ~n36111 & n36112 ) ;
  assign n36114 = ~n36056 & n36113 ;
  assign n36115 = n36056 & ~n36113 ;
  assign n36116 = n36114 | n36115 ;
  assign n36117 = ~n35776 & n35778 ;
  assign n36118 = ( n35776 & n35781 ) | ( n35776 & ~n36117 ) | ( n35781 & ~n36117 ) ;
  assign n36119 = ~n36116 & n36118 ;
  assign n36120 = n36116 & ~n36118 ;
  assign n36121 = n36119 | n36120 ;
  assign n36122 = n35787 & ~n36121 ;
  assign n36123 = ~n35787 & n36121 ;
  assign n36124 = n36122 | n36123 ;
  assign n36125 = n1057 & n24770 ;
  assign n36126 = n1065 & ~n25054 ;
  assign n36127 = n1060 & n24167 ;
  assign n36128 = n36126 | n36127 ;
  assign n36129 = n36125 | n36128 ;
  assign n36130 = n1062 | n36128 ;
  assign n36131 = n36125 | n36130 ;
  assign n36132 = ( ~n25095 & n36129 ) | ( ~n25095 & n36131 ) | ( n36129 & n36131 ) ;
  assign n36133 = n184 | n381 ;
  assign n36134 = n333 | n36133 ;
  assign n36135 = n1678 | n2787 ;
  assign n36136 = n399 | n595 ;
  assign n36137 = n36135 | n36136 ;
  assign n36138 = n36134 | n36137 ;
  assign n36139 = n1742 | n7880 ;
  assign n36140 = n2066 | n6029 ;
  assign n36141 = n35076 | n36140 ;
  assign n36142 = n36139 | n36141 ;
  assign n36143 = n36138 | n36142 ;
  assign n36144 = n26290 | n36143 ;
  assign n36145 = n13321 | n36144 ;
  assign n36146 = n1016 | n24282 ;
  assign n36147 = n431 | n4276 ;
  assign n36148 = n474 | n36147 ;
  assign n36149 = n36146 | n36148 ;
  assign n36150 = n36145 | n36149 ;
  assign n36151 = n477 | n762 ;
  assign n36152 = n1251 | n36151 ;
  assign n36153 = n143 & ~n197 ;
  assign n36154 = ~n363 & n36153 ;
  assign n36155 = ~n36152 & n36154 ;
  assign n36156 = n405 | n413 ;
  assign n36157 = n375 | n36156 ;
  assign n36158 = n36155 & ~n36157 ;
  assign n36159 = ~n36150 & n36158 ;
  assign n36160 = n36129 & ~n36159 ;
  assign n36161 = n36125 & ~n36159 ;
  assign n36162 = ( n36130 & ~n36159 ) | ( n36130 & n36161 ) | ( ~n36159 & n36161 ) ;
  assign n36163 = ( ~n25095 & n36160 ) | ( ~n25095 & n36162 ) | ( n36160 & n36162 ) ;
  assign n36164 = n36132 & ~n36163 ;
  assign n36165 = n36131 | n36159 ;
  assign n36166 = n36129 | n36159 ;
  assign n36167 = ( ~n25095 & n36165 ) | ( ~n25095 & n36166 ) | ( n36165 & n36166 ) ;
  assign n36168 = ~n36164 & n36167 ;
  assign n36169 = ~n35823 & n35828 ;
  assign n36170 = ( n35823 & n35830 ) | ( n35823 & ~n36169 ) | ( n35830 & ~n36169 ) ;
  assign n36171 = ~n36168 & n36170 ;
  assign n36172 = n36168 & ~n36170 ;
  assign n36173 = n36171 | n36172 ;
  assign n36174 = n1829 & n26017 ;
  assign n36175 = n1826 & ~n25046 ;
  assign n36176 = n1823 & ~n25728 ;
  assign n36177 = n36175 | n36176 ;
  assign n36178 = n36174 | n36177 ;
  assign n36179 = n1821 | n36174 ;
  assign n36180 = n36177 | n36179 ;
  assign n36181 = ( n26613 & n36178 ) | ( n26613 & n36180 ) | ( n36178 & n36180 ) ;
  assign n36182 = n36178 | n36180 ;
  assign n36183 = ( n26605 & n36181 ) | ( n26605 & n36182 ) | ( n36181 & n36182 ) ;
  assign n36184 = x29 & n36183 ;
  assign n36185 = x29 & ~n36183 ;
  assign n36186 = ( n36183 & ~n36184 ) | ( n36183 & n36185 ) | ( ~n36184 & n36185 ) ;
  assign n36187 = ~n36173 & n36186 ;
  assign n36188 = n36173 & ~n36186 ;
  assign n36189 = n36187 | n36188 ;
  assign n36190 = ~n35849 & n35851 ;
  assign n36191 = ( n35849 & n35853 ) | ( n35849 & ~n36190 ) | ( n35853 & ~n36190 ) ;
  assign n36192 = ~n36189 & n36191 ;
  assign n36193 = n36189 & ~n36191 ;
  assign n36194 = n36192 | n36193 ;
  assign n36195 = n2312 & ~n26270 ;
  assign n36196 = ~n26263 & n36195 ;
  assign n36197 = n2308 & ~n26526 ;
  assign n36198 = ~n26520 & n36197 ;
  assign n36199 = n36196 | n36198 ;
  assign n36200 = n2315 & ~n27133 ;
  assign n36201 = ~n27125 & n36200 ;
  assign n36202 = n36199 | n36201 ;
  assign n36203 = n27699 | n36202 ;
  assign n36204 = n27696 & ~n36203 ;
  assign n36205 = n2306 | n36201 ;
  assign n36206 = n36199 | n36205 ;
  assign n36207 = ~n36204 & n36206 ;
  assign n36208 = x26 & n36206 ;
  assign n36209 = ~n36204 & n36208 ;
  assign n36210 = x26 & ~n36208 ;
  assign n36211 = ( x26 & n36204 ) | ( x26 & n36210 ) | ( n36204 & n36210 ) ;
  assign n36212 = ( n36207 & ~n36209 ) | ( n36207 & n36211 ) | ( ~n36209 & n36211 ) ;
  assign n36213 = ~n36194 & n36212 ;
  assign n36214 = n36194 & ~n36212 ;
  assign n36215 = n36213 | n36214 ;
  assign n36216 = n35873 & ~n36215 ;
  assign n36217 = ( n35879 & ~n36215 ) | ( n35879 & n36216 ) | ( ~n36215 & n36216 ) ;
  assign n36218 = ~n35873 & n36215 ;
  assign n36219 = ~n35879 & n36218 ;
  assign n36220 = n36217 | n36219 ;
  assign n36221 = n2925 & ~n27371 ;
  assign n36222 = ~n27363 & n36221 ;
  assign n36223 = n2928 & ~n27606 ;
  assign n36224 = ~n27597 & n36223 ;
  assign n36225 = n36222 | n36224 ;
  assign n36226 = n2932 & ~n28503 ;
  assign n36227 = n28498 & n36226 ;
  assign n36228 = n36225 | n36227 ;
  assign n36229 = n2936 & n28794 ;
  assign n36230 = ( n2936 & n28783 ) | ( n2936 & n36229 ) | ( n28783 & n36229 ) ;
  assign n36231 = n36228 | n36230 ;
  assign n36232 = x23 | n36228 ;
  assign n36233 = n36230 | n36232 ;
  assign n36234 = ~x23 & n36232 ;
  assign n36235 = ( ~x23 & n36230 ) | ( ~x23 & n36234 ) | ( n36230 & n36234 ) ;
  assign n36236 = ( ~n36231 & n36233 ) | ( ~n36231 & n36235 ) | ( n36233 & n36235 ) ;
  assign n36237 = ~n36220 & n36236 ;
  assign n36238 = n36220 | n36237 ;
  assign n36239 = n36220 & n36236 ;
  assign n36240 = n36238 & ~n36239 ;
  assign n36241 = n35901 & n36239 ;
  assign n36242 = ( n35901 & ~n36238 ) | ( n35901 & n36241 ) | ( ~n36238 & n36241 ) ;
  assign n36243 = ( n35908 & ~n36240 ) | ( n35908 & n36242 ) | ( ~n36240 & n36242 ) ;
  assign n36244 = n35901 | n36239 ;
  assign n36245 = n36238 & ~n36244 ;
  assign n36246 = ~n35908 & n36245 ;
  assign n36247 = n36243 | n36246 ;
  assign n36249 = n3544 & n28492 ;
  assign n36250 = n3541 & ~n28714 ;
  assign n36251 = n36249 | n36250 ;
  assign n36248 = n3547 & n29620 ;
  assign n36253 = n3537 | n36248 ;
  assign n36254 = n36251 | n36253 ;
  assign n36252 = n36248 | n36251 ;
  assign n36255 = n36252 & n36254 ;
  assign n36256 = ( ~n29642 & n36254 ) | ( ~n29642 & n36255 ) | ( n36254 & n36255 ) ;
  assign n36257 = n36254 | n36255 ;
  assign n36258 = ( n29629 & n36256 ) | ( n29629 & n36257 ) | ( n36256 & n36257 ) ;
  assign n36259 = ~x20 & n36258 ;
  assign n36260 = x20 | n36258 ;
  assign n36261 = ( ~n36258 & n36259 ) | ( ~n36258 & n36260 ) | ( n36259 & n36260 ) ;
  assign n36262 = ~n36247 & n36261 ;
  assign n36263 = n36247 & ~n36261 ;
  assign n36264 = n36262 | n36263 ;
  assign n36265 = n35925 & ~n36264 ;
  assign n36266 = ( n35931 & ~n36264 ) | ( n35931 & n36265 ) | ( ~n36264 & n36265 ) ;
  assign n36267 = ~n35925 & n36264 ;
  assign n36268 = ~n35931 & n36267 ;
  assign n36269 = n36266 | n36268 ;
  assign n36270 = n4471 & ~n30186 ;
  assign n36271 = n4466 & ~n30199 ;
  assign n36272 = n4468 & n30212 ;
  assign n36273 = n36271 | n36272 ;
  assign n36274 = n36270 | n36273 ;
  assign n36275 = n4475 | n36270 ;
  assign n36276 = n36273 | n36275 ;
  assign n36277 = ( ~n30241 & n36274 ) | ( ~n30241 & n36276 ) | ( n36274 & n36276 ) ;
  assign n36278 = ~x17 & n36276 ;
  assign n36279 = ~x17 & n36274 ;
  assign n36280 = ( ~n30241 & n36278 ) | ( ~n30241 & n36279 ) | ( n36278 & n36279 ) ;
  assign n36281 = x17 | n36279 ;
  assign n36282 = x17 | n36278 ;
  assign n36283 = ( ~n30241 & n36281 ) | ( ~n30241 & n36282 ) | ( n36281 & n36282 ) ;
  assign n36284 = ( ~n36277 & n36280 ) | ( ~n36277 & n36283 ) | ( n36280 & n36283 ) ;
  assign n36285 = ~n36269 & n36284 ;
  assign n36286 = n36269 | n36285 ;
  assign n36287 = n36269 & n36284 ;
  assign n36288 = n36286 & ~n36287 ;
  assign n36289 = n35948 | n35955 ;
  assign n36290 = n36288 & ~n36289 ;
  assign n36291 = ~n36288 & n36289 ;
  assign n36292 = n36290 | n36291 ;
  assign n36294 = n5237 & ~n31309 ;
  assign n36295 = n5231 & ~n31323 ;
  assign n36296 = n36294 | n36295 ;
  assign n36293 = n5234 & n31295 ;
  assign n36298 = n5227 | n36293 ;
  assign n36299 = n36296 | n36298 ;
  assign n36297 = n36293 | n36296 ;
  assign n36300 = n36297 & n36299 ;
  assign n36301 = ( n31355 & n36299 ) | ( n31355 & n36300 ) | ( n36299 & n36300 ) ;
  assign n36302 = x14 & n36300 ;
  assign n36303 = x14 & n36299 ;
  assign n36304 = ( n31355 & n36302 ) | ( n31355 & n36303 ) | ( n36302 & n36303 ) ;
  assign n36305 = x14 & ~n36302 ;
  assign n36306 = x14 & ~n36303 ;
  assign n36307 = ( ~n31355 & n36305 ) | ( ~n31355 & n36306 ) | ( n36305 & n36306 ) ;
  assign n36308 = ( n36301 & ~n36304 ) | ( n36301 & n36307 ) | ( ~n36304 & n36307 ) ;
  assign n36309 = ~n36292 & n36308 ;
  assign n36310 = n36292 & ~n36308 ;
  assign n36311 = n36309 | n36310 ;
  assign n36312 = n35972 & ~n36311 ;
  assign n36313 = ( n35978 & ~n36311 ) | ( n35978 & n36312 ) | ( ~n36311 & n36312 ) ;
  assign n36314 = ~n35972 & n36311 ;
  assign n36315 = ~n35978 & n36314 ;
  assign n36316 = n36313 | n36315 ;
  assign n36317 = n6122 & ~n32442 ;
  assign n36318 = n6125 & n32306 ;
  assign n36319 = n6119 & n32293 ;
  assign n36320 = n36318 | n36319 ;
  assign n36321 = n36317 | n36320 ;
  assign n36322 = n6115 | n36317 ;
  assign n36323 = n36320 | n36322 ;
  assign n36324 = ( ~n32458 & n36321 ) | ( ~n32458 & n36323 ) | ( n36321 & n36323 ) ;
  assign n36325 = ~x11 & n36323 ;
  assign n36326 = ~x11 & n36321 ;
  assign n36327 = ( ~n32458 & n36325 ) | ( ~n32458 & n36326 ) | ( n36325 & n36326 ) ;
  assign n36328 = x11 | n36326 ;
  assign n36329 = x11 | n36325 ;
  assign n36330 = ( ~n32458 & n36328 ) | ( ~n32458 & n36329 ) | ( n36328 & n36329 ) ;
  assign n36331 = ( ~n36324 & n36327 ) | ( ~n36324 & n36330 ) | ( n36327 & n36330 ) ;
  assign n36332 = ~n36316 & n36331 ;
  assign n36333 = n36316 | n36332 ;
  assign n36334 = n36316 & n36331 ;
  assign n36335 = n36333 & ~n36334 ;
  assign n36336 = n35997 | n36003 ;
  assign n36337 = ~n35997 & n36000 ;
  assign n36338 = ( n35651 & n36336 ) | ( n35651 & ~n36337 ) | ( n36336 & ~n36337 ) ;
  assign n36339 = n36335 & ~n36338 ;
  assign n36340 = ~n36335 & n36338 ;
  assign n36341 = n36339 | n36340 ;
  assign n36342 = n7074 & n33436 ;
  assign n36343 = n7068 & ~n33423 ;
  assign n36344 = n36342 | n36343 ;
  assign n36345 = n7079 & n33526 ;
  assign n36346 = n7078 | n36345 ;
  assign n36347 = n36344 | n36346 ;
  assign n36348 = n36344 | n36345 ;
  assign n36349 = n33545 | n36348 ;
  assign n36350 = n33548 & ~n36348 ;
  assign n36351 = ( n32456 & ~n36349 ) | ( n32456 & n36350 ) | ( ~n36349 & n36350 ) ;
  assign n36352 = n36347 & ~n36351 ;
  assign n36353 = ( n33536 & n36347 ) | ( n33536 & n36352 ) | ( n36347 & n36352 ) ;
  assign n36354 = x8 & n36353 ;
  assign n36355 = x8 & ~n36353 ;
  assign n36356 = ( n36353 & ~n36354 ) | ( n36353 & n36355 ) | ( ~n36354 & n36355 ) ;
  assign n36357 = ~n36341 & n36356 ;
  assign n36358 = n36341 & ~n36356 ;
  assign n36359 = n36357 | n36358 ;
  assign n36360 = n36021 & ~n36359 ;
  assign n36361 = ( n36027 & ~n36359 ) | ( n36027 & n36360 ) | ( ~n36359 & n36360 ) ;
  assign n36362 = ~n36021 & n36359 ;
  assign n36363 = ~n36027 & n36362 ;
  assign n36364 = n36361 | n36363 ;
  assign n36365 = n8122 & ~n35371 ;
  assign n36366 = n8115 & n34656 ;
  assign n36367 = n8118 & n35021 ;
  assign n36368 = n36366 | n36367 ;
  assign n36369 = n36365 | n36368 ;
  assign n36370 = n8125 & ~n35392 ;
  assign n36371 = n8125 & ~n35395 ;
  assign n36372 = ( ~n32456 & n36370 ) | ( ~n32456 & n36371 ) | ( n36370 & n36371 ) ;
  assign n36373 = n36369 | n36372 ;
  assign n36374 = n8125 | n36369 ;
  assign n36375 = ( n35381 & n36373 ) | ( n35381 & n36374 ) | ( n36373 & n36374 ) ;
  assign n36376 = x5 | n36375 ;
  assign n36377 = ~x5 & n36375 ;
  assign n36378 = ( ~n36375 & n36376 ) | ( ~n36375 & n36377 ) | ( n36376 & n36377 ) ;
  assign n36379 = ~n36364 & n36378 ;
  assign n36380 = n36364 | n36379 ;
  assign n36381 = n24127 & n36083 ;
  assign n36382 = n9021 & n35746 ;
  assign n36383 = n36381 | n36382 ;
  assign n36384 = n8970 | n36383 ;
  assign n36385 = ( n36103 & n36383 ) | ( n36103 & n36384 ) | ( n36383 & n36384 ) ;
  assign n36386 = ( n36105 & n36383 ) | ( n36105 & n36384 ) | ( n36383 & n36384 ) ;
  assign n36387 = ( n32456 & n36385 ) | ( n32456 & n36386 ) | ( n36385 & n36386 ) ;
  assign n36388 = x2 & n36387 ;
  assign n36389 = x2 & ~n36387 ;
  assign n36390 = ( n36387 & ~n36388 ) | ( n36387 & n36389 ) | ( ~n36388 & n36389 ) ;
  assign n36391 = n36364 & n36378 ;
  assign n36392 = n36390 & n36391 ;
  assign n36393 = ( ~n36380 & n36390 ) | ( ~n36380 & n36392 ) | ( n36390 & n36392 ) ;
  assign n36394 = n36390 | n36391 ;
  assign n36395 = n36380 & ~n36394 ;
  assign n36396 = n36393 | n36395 ;
  assign n36397 = n36047 | n36055 ;
  assign n36398 = n36396 & ~n36397 ;
  assign n36399 = ~n36396 & n36397 ;
  assign n36400 = n36398 | n36399 ;
  assign n36401 = ~n36114 & n36400 ;
  assign n36402 = ~n36119 & n36401 ;
  assign n36403 = ( ~n36114 & n36116 ) | ( ~n36114 & n36400 ) | ( n36116 & n36400 ) ;
  assign n36404 = n36114 & ~n36400 ;
  assign n36405 = ( n36118 & ~n36403 ) | ( n36118 & n36404 ) | ( ~n36403 & n36404 ) ;
  assign n36406 = n36402 | n36405 ;
  assign n36407 = n36122 & ~n36406 ;
  assign n36408 = ~n36122 & n36406 ;
  assign n36409 = n36407 | n36408 ;
  assign n36410 = n1057 & ~n25046 ;
  assign n36411 = n1060 & ~n25054 ;
  assign n36412 = n1065 & n24770 ;
  assign n36413 = n36411 | n36412 ;
  assign n36414 = n36410 | n36413 ;
  assign n36415 = n1062 | n36410 ;
  assign n36416 = n36413 | n36415 ;
  assign n36417 = ( ~n25069 & n36414 ) | ( ~n25069 & n36416 ) | ( n36414 & n36416 ) ;
  assign n36418 = x2 | n9020 ;
  assign n36419 = n8969 | n36418 ;
  assign n36420 = ( x2 & n36083 ) | ( x2 & ~n36419 ) | ( n36083 & ~n36419 ) ;
  assign n36421 = x2 & n36419 ;
  assign n36422 = ~n36083 & n36421 ;
  assign n36423 = ( n36083 & ~n36420 ) | ( n36083 & n36422 ) | ( ~n36420 & n36422 ) ;
  assign n36424 = n76 | n2217 ;
  assign n36425 = n1372 | n29749 ;
  assign n36426 = n36424 | n36425 ;
  assign n36427 = n407 | n36426 ;
  assign n36428 = n448 | n1028 ;
  assign n36429 = n29920 & ~n36428 ;
  assign n36430 = ~n2683 & n36429 ;
  assign n36431 = ~n36427 & n36430 ;
  assign n36432 = ~n2192 & n36431 ;
  assign n36433 = ~n7863 & n36432 ;
  assign n36434 = n334 | n8004 ;
  assign n36435 = n329 | n36434 ;
  assign n36436 = n821 | n36435 ;
  assign n36437 = n401 | n469 ;
  assign n36438 = n24228 | n36437 ;
  assign n36439 = n234 | n514 ;
  assign n36440 = n36438 | n36439 ;
  assign n36441 = n36436 | n36440 ;
  assign n36442 = n36433 & ~n36441 ;
  assign n36443 = n36423 & ~n36442 ;
  assign n36444 = ~n36423 & n36442 ;
  assign n36445 = n36443 | n36444 ;
  assign n36446 = n36416 & ~n36445 ;
  assign n36447 = n36414 & ~n36445 ;
  assign n36448 = ( ~n25069 & n36446 ) | ( ~n25069 & n36447 ) | ( n36446 & n36447 ) ;
  assign n36449 = n36417 & ~n36448 ;
  assign n36450 = n36445 | n36448 ;
  assign n36451 = ~n36449 & n36450 ;
  assign n36452 = ~n36163 & n36168 ;
  assign n36453 = n36451 & n36452 ;
  assign n36454 = ~n36163 & n36451 ;
  assign n36455 = ( ~n36170 & n36453 ) | ( ~n36170 & n36454 ) | ( n36453 & n36454 ) ;
  assign n36456 = n36451 | n36452 ;
  assign n36457 = n36163 & ~n36451 ;
  assign n36458 = ( n36170 & ~n36456 ) | ( n36170 & n36457 ) | ( ~n36456 & n36457 ) ;
  assign n36459 = n36455 | n36458 ;
  assign n36460 = n1826 & ~n25728 ;
  assign n36461 = n1823 & n26017 ;
  assign n36462 = n36460 | n36461 ;
  assign n36463 = n1829 & ~n26270 ;
  assign n36464 = ~n26263 & n36463 ;
  assign n36466 = n1821 | n36464 ;
  assign n36467 = n36462 | n36466 ;
  assign n36465 = n36462 | n36464 ;
  assign n36468 = n36465 & n36467 ;
  assign n36469 = ( n26571 & n36467 ) | ( n26571 & n36468 ) | ( n36467 & n36468 ) ;
  assign n36470 = x29 & n36468 ;
  assign n36471 = x29 & n36467 ;
  assign n36472 = ( n26571 & n36470 ) | ( n26571 & n36471 ) | ( n36470 & n36471 ) ;
  assign n36473 = x29 & ~n36470 ;
  assign n36474 = x29 & ~n36471 ;
  assign n36475 = ( ~n26571 & n36473 ) | ( ~n26571 & n36474 ) | ( n36473 & n36474 ) ;
  assign n36476 = ( n36469 & ~n36472 ) | ( n36469 & n36475 ) | ( ~n36472 & n36475 ) ;
  assign n36477 = ~n36459 & n36476 ;
  assign n36478 = n36459 & ~n36476 ;
  assign n36479 = n36477 | n36478 ;
  assign n36480 = ~n36187 & n36189 ;
  assign n36481 = ( n36187 & n36191 ) | ( n36187 & ~n36480 ) | ( n36191 & ~n36480 ) ;
  assign n36482 = ~n36479 & n36481 ;
  assign n36483 = n36479 & ~n36481 ;
  assign n36484 = n36482 | n36483 ;
  assign n36485 = n2312 & ~n26526 ;
  assign n36486 = ~n26520 & n36485 ;
  assign n36487 = n2308 & ~n27133 ;
  assign n36488 = ~n27125 & n36487 ;
  assign n36489 = n36486 | n36488 ;
  assign n36490 = n2315 & ~n27371 ;
  assign n36491 = ~n27363 & n36490 ;
  assign n36492 = n36489 | n36491 ;
  assign n36493 = n2306 | n36491 ;
  assign n36494 = n36489 | n36493 ;
  assign n36495 = ( ~n27654 & n36492 ) | ( ~n27654 & n36494 ) | ( n36492 & n36494 ) ;
  assign n36496 = ~x26 & n36494 ;
  assign n36497 = ~x26 & n36492 ;
  assign n36498 = ( ~n27654 & n36496 ) | ( ~n27654 & n36497 ) | ( n36496 & n36497 ) ;
  assign n36499 = x26 | n36497 ;
  assign n36500 = x26 | n36496 ;
  assign n36501 = ( ~n27654 & n36499 ) | ( ~n27654 & n36500 ) | ( n36499 & n36500 ) ;
  assign n36502 = ( ~n36495 & n36498 ) | ( ~n36495 & n36501 ) | ( n36498 & n36501 ) ;
  assign n36503 = n36484 | n36502 ;
  assign n36504 = n36484 & ~n36502 ;
  assign n36505 = ( ~n36484 & n36503 ) | ( ~n36484 & n36504 ) | ( n36503 & n36504 ) ;
  assign n36506 = n36213 | n36216 ;
  assign n36507 = ~n36213 & n36215 ;
  assign n36508 = ( n35879 & n36506 ) | ( n35879 & ~n36507 ) | ( n36506 & ~n36507 ) ;
  assign n36509 = n36505 & ~n36508 ;
  assign n36510 = ~n36505 & n36508 ;
  assign n36511 = n36509 | n36510 ;
  assign n36512 = n2932 & n28492 ;
  assign n36513 = n2925 & ~n27606 ;
  assign n36514 = ~n27597 & n36513 ;
  assign n36515 = n2928 & ~n28503 ;
  assign n36516 = n28498 & n36515 ;
  assign n36517 = n36514 | n36516 ;
  assign n36518 = n36512 | n36517 ;
  assign n36519 = n2936 | n36518 ;
  assign n36520 = ( ~n28749 & n36518 ) | ( ~n28749 & n36519 ) | ( n36518 & n36519 ) ;
  assign n36521 = ~x23 & n36519 ;
  assign n36522 = ~x23 & n36518 ;
  assign n36523 = ( ~n28749 & n36521 ) | ( ~n28749 & n36522 ) | ( n36521 & n36522 ) ;
  assign n36524 = x23 | n36521 ;
  assign n36525 = x23 | n36522 ;
  assign n36526 = ( ~n28749 & n36524 ) | ( ~n28749 & n36525 ) | ( n36524 & n36525 ) ;
  assign n36527 = ( ~n36520 & n36523 ) | ( ~n36520 & n36526 ) | ( n36523 & n36526 ) ;
  assign n36528 = n36511 & n36527 ;
  assign n36529 = n36505 & ~n36527 ;
  assign n36530 = ( n36508 & n36527 ) | ( n36508 & ~n36529 ) | ( n36527 & ~n36529 ) ;
  assign n36531 = n36509 | n36530 ;
  assign n36532 = ~n36528 & n36531 ;
  assign n36533 = n36237 | n36242 ;
  assign n36534 = ~n36237 & n36240 ;
  assign n36535 = ( n35908 & n36533 ) | ( n35908 & ~n36534 ) | ( n36533 & ~n36534 ) ;
  assign n36536 = n36532 & ~n36535 ;
  assign n36537 = ~n36532 & n36535 ;
  assign n36538 = n36536 | n36537 ;
  assign n36539 = n3547 & ~n30199 ;
  assign n36540 = n3544 & ~n28714 ;
  assign n36541 = n3541 & n29620 ;
  assign n36542 = n36540 | n36541 ;
  assign n36543 = n36539 | n36542 ;
  assign n36544 = n3537 | n36539 ;
  assign n36545 = n36542 | n36544 ;
  assign n36546 = ( ~n30299 & n36543 ) | ( ~n30299 & n36545 ) | ( n36543 & n36545 ) ;
  assign n36547 = ~x20 & n36545 ;
  assign n36548 = ~x20 & n36543 ;
  assign n36549 = ( ~n30299 & n36547 ) | ( ~n30299 & n36548 ) | ( n36547 & n36548 ) ;
  assign n36550 = x20 | n36548 ;
  assign n36551 = x20 | n36547 ;
  assign n36552 = ( ~n30299 & n36550 ) | ( ~n30299 & n36551 ) | ( n36550 & n36551 ) ;
  assign n36553 = ( ~n36546 & n36549 ) | ( ~n36546 & n36552 ) | ( n36549 & n36552 ) ;
  assign n36554 = n36538 & n36553 ;
  assign n36555 = n36532 & ~n36553 ;
  assign n36556 = ( n36535 & n36553 ) | ( n36535 & ~n36555 ) | ( n36553 & ~n36555 ) ;
  assign n36557 = n36536 | n36556 ;
  assign n36558 = ~n36554 & n36557 ;
  assign n36559 = ~n36262 & n36558 ;
  assign n36560 = ~n36266 & n36559 ;
  assign n36561 = n36262 & ~n36558 ;
  assign n36562 = ( n36266 & ~n36558 ) | ( n36266 & n36561 ) | ( ~n36558 & n36561 ) ;
  assign n36563 = n36560 | n36562 ;
  assign n36564 = n4471 & ~n31309 ;
  assign n36565 = n4466 & n30212 ;
  assign n36566 = n4468 & ~n30186 ;
  assign n36567 = n36565 | n36566 ;
  assign n36568 = n36564 | n36567 ;
  assign n36569 = n4475 | n36564 ;
  assign n36570 = n36567 | n36569 ;
  assign n36571 = ( n31404 & n36568 ) | ( n31404 & n36570 ) | ( n36568 & n36570 ) ;
  assign n36572 = x17 & n36570 ;
  assign n36573 = x17 & n36568 ;
  assign n36574 = ( n31404 & n36572 ) | ( n31404 & n36573 ) | ( n36572 & n36573 ) ;
  assign n36575 = x17 & ~n36573 ;
  assign n36576 = x17 & ~n36572 ;
  assign n36577 = ( ~n31404 & n36575 ) | ( ~n31404 & n36576 ) | ( n36575 & n36576 ) ;
  assign n36578 = ( n36571 & ~n36574 ) | ( n36571 & n36577 ) | ( ~n36574 & n36577 ) ;
  assign n36579 = n36563 & n36578 ;
  assign n36580 = n36562 | n36578 ;
  assign n36581 = n36560 | n36580 ;
  assign n36582 = ~n36579 & n36581 ;
  assign n36583 = ~n36285 & n36288 ;
  assign n36584 = ( n36285 & n36289 ) | ( n36285 & ~n36583 ) | ( n36289 & ~n36583 ) ;
  assign n36585 = n36582 & ~n36584 ;
  assign n36586 = ~n36582 & n36584 ;
  assign n36587 = n36585 | n36586 ;
  assign n36588 = n5234 & n32306 ;
  assign n36589 = n5237 & ~n31323 ;
  assign n36590 = n5231 & n31295 ;
  assign n36591 = n36589 | n36590 ;
  assign n36592 = n36588 | n36591 ;
  assign n36593 = n5227 | n36588 ;
  assign n36594 = n36591 | n36593 ;
  assign n36595 = ( ~n32525 & n36592 ) | ( ~n32525 & n36594 ) | ( n36592 & n36594 ) ;
  assign n36596 = ~x14 & n36594 ;
  assign n36597 = ~x14 & n36592 ;
  assign n36598 = ( ~n32525 & n36596 ) | ( ~n32525 & n36597 ) | ( n36596 & n36597 ) ;
  assign n36599 = x14 | n36597 ;
  assign n36600 = x14 | n36596 ;
  assign n36601 = ( ~n32525 & n36599 ) | ( ~n32525 & n36600 ) | ( n36599 & n36600 ) ;
  assign n36602 = ( ~n36595 & n36598 ) | ( ~n36595 & n36601 ) | ( n36598 & n36601 ) ;
  assign n36603 = n36587 & n36602 ;
  assign n36604 = n36582 & ~n36602 ;
  assign n36605 = ( n36584 & n36602 ) | ( n36584 & ~n36604 ) | ( n36602 & ~n36604 ) ;
  assign n36606 = n36585 | n36605 ;
  assign n36607 = ~n36603 & n36606 ;
  assign n36608 = ~n36309 & n36607 ;
  assign n36609 = ~n36313 & n36608 ;
  assign n36610 = n36309 & ~n36607 ;
  assign n36611 = ( n36313 & ~n36607 ) | ( n36313 & n36610 ) | ( ~n36607 & n36610 ) ;
  assign n36612 = n36609 | n36611 ;
  assign n36613 = n6122 & n33436 ;
  assign n36614 = n6125 & n32293 ;
  assign n36615 = n6119 & ~n32442 ;
  assign n36616 = n36614 | n36615 ;
  assign n36617 = n36613 | n36616 ;
  assign n36618 = n6115 & ~n33441 ;
  assign n36619 = ~n32456 & n36618 ;
  assign n36620 = ( n6115 & n34271 ) | ( n6115 & n36619 ) | ( n34271 & n36619 ) ;
  assign n36621 = n36617 | n36620 ;
  assign n36622 = x11 | n36617 ;
  assign n36623 = n36620 | n36622 ;
  assign n36624 = ~x11 & n36622 ;
  assign n36625 = ( ~x11 & n36620 ) | ( ~x11 & n36624 ) | ( n36620 & n36624 ) ;
  assign n36626 = ( ~n36621 & n36623 ) | ( ~n36621 & n36625 ) | ( n36623 & n36625 ) ;
  assign n36627 = n36612 & n36626 ;
  assign n36628 = n36611 | n36626 ;
  assign n36629 = n36609 | n36628 ;
  assign n36630 = ~n36627 & n36629 ;
  assign n36631 = ~n36332 & n36335 ;
  assign n36632 = ( n36332 & n36338 ) | ( n36332 & ~n36631 ) | ( n36338 & ~n36631 ) ;
  assign n36633 = n36630 & ~n36632 ;
  assign n36634 = ~n36630 & n36632 ;
  assign n36635 = n36633 | n36634 ;
  assign n36636 = n7079 & n34656 ;
  assign n36637 = n7074 & ~n33423 ;
  assign n36638 = n7068 & n33526 ;
  assign n36639 = n36637 | n36638 ;
  assign n36640 = n36636 | n36639 ;
  assign n36641 = n7078 | n36636 ;
  assign n36642 = n36639 | n36641 ;
  assign n36643 = ( n34667 & n36640 ) | ( n34667 & n36642 ) | ( n36640 & n36642 ) ;
  assign n36644 = x8 & n36642 ;
  assign n36645 = x8 & n36640 ;
  assign n36646 = ( n34667 & n36644 ) | ( n34667 & n36645 ) | ( n36644 & n36645 ) ;
  assign n36647 = x8 & ~n36645 ;
  assign n36648 = x8 & ~n36644 ;
  assign n36649 = ( ~n34667 & n36647 ) | ( ~n34667 & n36648 ) | ( n36647 & n36648 ) ;
  assign n36650 = ( n36643 & ~n36646 ) | ( n36643 & n36649 ) | ( ~n36646 & n36649 ) ;
  assign n36651 = n36635 & n36650 ;
  assign n36652 = n36630 & ~n36650 ;
  assign n36653 = ( n36632 & n36650 ) | ( n36632 & ~n36652 ) | ( n36650 & ~n36652 ) ;
  assign n36654 = n36633 | n36653 ;
  assign n36655 = ~n36651 & n36654 ;
  assign n36656 = n36357 | n36360 ;
  assign n36657 = ~n36357 & n36359 ;
  assign n36658 = ( n36027 & n36656 ) | ( n36027 & ~n36657 ) | ( n36656 & ~n36657 ) ;
  assign n36659 = n36655 & ~n36658 ;
  assign n36660 = ~n36655 & n36658 ;
  assign n36661 = n36659 | n36660 ;
  assign n36662 = n8122 & n35746 ;
  assign n36663 = n8115 & n35021 ;
  assign n36664 = n8118 & ~n35371 ;
  assign n36665 = n36663 | n36664 ;
  assign n36666 = n36662 | n36665 ;
  assign n36667 = n8125 | n36662 ;
  assign n36668 = n36665 | n36667 ;
  assign n36669 = ( ~n35759 & n36666 ) | ( ~n35759 & n36668 ) | ( n36666 & n36668 ) ;
  assign n36670 = ~x5 & n36668 ;
  assign n36671 = ~x5 & n36666 ;
  assign n36672 = ( ~n35759 & n36670 ) | ( ~n35759 & n36671 ) | ( n36670 & n36671 ) ;
  assign n36673 = x5 | n36671 ;
  assign n36674 = x5 | n36670 ;
  assign n36675 = ( ~n35759 & n36673 ) | ( ~n35759 & n36674 ) | ( n36673 & n36674 ) ;
  assign n36676 = ( ~n36669 & n36672 ) | ( ~n36669 & n36675 ) | ( n36672 & n36675 ) ;
  assign n36677 = n36661 & n36676 ;
  assign n36678 = n36655 & ~n36676 ;
  assign n36679 = ( n36658 & n36676 ) | ( n36658 & ~n36678 ) | ( n36676 & ~n36678 ) ;
  assign n36680 = n36659 | n36679 ;
  assign n36681 = ~n36677 & n36680 ;
  assign n36682 = n36379 | n36393 ;
  assign n36683 = n36681 & ~n36682 ;
  assign n36684 = ~n36681 & n36682 ;
  assign n36685 = n36683 | n36684 ;
  assign n36686 = n36399 & ~n36685 ;
  assign n36687 = ( n36405 & ~n36685 ) | ( n36405 & n36686 ) | ( ~n36685 & n36686 ) ;
  assign n36688 = ~n36399 & n36685 ;
  assign n36689 = ~n36405 & n36688 ;
  assign n36690 = n36687 | n36689 ;
  assign n36691 = ~n36407 & n36690 ;
  assign n36692 = n36406 | n36690 ;
  assign n36693 = n36122 & ~n36692 ;
  assign n36694 = n36691 | n36693 ;
  assign n36695 = n10811 | n10816 ;
  assign n36696 = n1149 | n4145 ;
  assign n36697 = n22449 | n36696 ;
  assign n36698 = n129 | n36697 ;
  assign n36699 = n274 | n364 ;
  assign n36700 = n10737 | n36699 ;
  assign n36701 = n413 | n775 ;
  assign n36702 = n36700 | n36701 ;
  assign n36703 = n36698 | n36702 ;
  assign n36704 = n758 | n2644 ;
  assign n36705 = n857 | n36704 ;
  assign n36706 = n36703 | n36705 ;
  assign n36707 = n36695 | n36706 ;
  assign n36708 = ( n504 & ~n894 ) | ( n504 & n1523 ) | ( ~n894 & n1523 ) ;
  assign n36709 = n894 | n36708 ;
  assign n36710 = n2265 | n36709 ;
  assign n36711 = n1166 | n12387 ;
  assign n36712 = n249 | n325 ;
  assign n36713 = n517 | n36712 ;
  assign n36714 = n36711 | n36713 ;
  assign n36715 = n229 | n36714 ;
  assign n36716 = n36710 | n36715 ;
  assign n36717 = n36707 | n36716 ;
  assign n36718 = n36423 & n36717 ;
  assign n36719 = n36423 | n36717 ;
  assign n36720 = ~n36718 & n36719 ;
  assign n36721 = n36443 & n36720 ;
  assign n36722 = ( n36448 & n36720 ) | ( n36448 & n36721 ) | ( n36720 & n36721 ) ;
  assign n36723 = ( n36443 & n36448 ) | ( n36443 & ~n36722 ) | ( n36448 & ~n36722 ) ;
  assign n36724 = n36720 & ~n36721 ;
  assign n36725 = ~n36448 & n36724 ;
  assign n36726 = n36723 | n36725 ;
  assign n36727 = n1057 & ~n25728 ;
  assign n36728 = n1060 & n24770 ;
  assign n36729 = n1065 & ~n25046 ;
  assign n36730 = n36728 | n36729 ;
  assign n36731 = n36727 | n36730 ;
  assign n36732 = n1062 & n25740 ;
  assign n36733 = n1062 & n25731 ;
  assign n36734 = ( ~n25441 & n36732 ) | ( ~n25441 & n36733 ) | ( n36732 & n36733 ) ;
  assign n36735 = n36731 | n36734 ;
  assign n36736 = n1062 | n36731 ;
  assign n36737 = ( n25733 & n36735 ) | ( n25733 & n36736 ) | ( n36735 & n36736 ) ;
  assign n36738 = n36725 & n36737 ;
  assign n36739 = ( n36723 & n36737 ) | ( n36723 & n36738 ) | ( n36737 & n36738 ) ;
  assign n36740 = n36726 & ~n36739 ;
  assign n36741 = ~n36725 & n36737 ;
  assign n36742 = ~n36723 & n36741 ;
  assign n36743 = n36740 | n36742 ;
  assign n36744 = n36458 | n36476 ;
  assign n36745 = ( n36458 & ~n36459 ) | ( n36458 & n36744 ) | ( ~n36459 & n36744 ) ;
  assign n36746 = n36743 | n36745 ;
  assign n36747 = n36743 & n36745 ;
  assign n36748 = n36746 & ~n36747 ;
  assign n36749 = n1826 & n26017 ;
  assign n36750 = n1823 & ~n26270 ;
  assign n36751 = ~n26263 & n36750 ;
  assign n36752 = n36749 | n36751 ;
  assign n36753 = n1829 & ~n26526 ;
  assign n36754 = ~n26520 & n36753 ;
  assign n36755 = n36752 | n36754 ;
  assign n36756 = n1821 | n36754 ;
  assign n36757 = n36752 | n36756 ;
  assign n36758 = ( ~n26555 & n36755 ) | ( ~n26555 & n36757 ) | ( n36755 & n36757 ) ;
  assign n36759 = ( n26528 & n36755 ) | ( n26528 & n36757 ) | ( n36755 & n36757 ) ;
  assign n36760 = ( ~n26543 & n36758 ) | ( ~n26543 & n36759 ) | ( n36758 & n36759 ) ;
  assign n36761 = ~x29 & n36760 ;
  assign n36762 = x29 | n36760 ;
  assign n36763 = ( ~n36760 & n36761 ) | ( ~n36760 & n36762 ) | ( n36761 & n36762 ) ;
  assign n36764 = n36748 & n36763 ;
  assign n36765 = n36748 & ~n36764 ;
  assign n36766 = n2312 & ~n27133 ;
  assign n36767 = ~n27125 & n36766 ;
  assign n36768 = n2308 & ~n27371 ;
  assign n36769 = ~n27363 & n36768 ;
  assign n36770 = n36767 | n36769 ;
  assign n36771 = n2315 & ~n27606 ;
  assign n36772 = ~n27597 & n36771 ;
  assign n36773 = n36770 | n36772 ;
  assign n36774 = n2306 & n27630 ;
  assign n36775 = ~n27625 & n36774 ;
  assign n36776 = ( n2306 & ~n27634 ) | ( n2306 & n36775 ) | ( ~n27634 & n36775 ) ;
  assign n36777 = n36773 | n36776 ;
  assign n36778 = x26 | n36773 ;
  assign n36779 = n36776 | n36778 ;
  assign n36780 = ~x26 & n36778 ;
  assign n36781 = ( ~x26 & n36776 ) | ( ~x26 & n36780 ) | ( n36776 & n36780 ) ;
  assign n36782 = ( ~n36777 & n36779 ) | ( ~n36777 & n36781 ) | ( n36779 & n36781 ) ;
  assign n36783 = ~n36748 & n36763 ;
  assign n36784 = n36782 & n36783 ;
  assign n36785 = ( n36765 & n36782 ) | ( n36765 & n36784 ) | ( n36782 & n36784 ) ;
  assign n36786 = n36782 | n36783 ;
  assign n36787 = n36765 | n36786 ;
  assign n36788 = ~n36785 & n36787 ;
  assign n36789 = n36482 | n36502 ;
  assign n36790 = ( n36482 & ~n36484 ) | ( n36482 & n36789 ) | ( ~n36484 & n36789 ) ;
  assign n36791 = n36788 | n36790 ;
  assign n36792 = n36788 & n36790 ;
  assign n36793 = n36791 & ~n36792 ;
  assign n36794 = n2932 & ~n28714 ;
  assign n36795 = n2928 & n28492 ;
  assign n36796 = n2925 & ~n28503 ;
  assign n36797 = n28498 & n36796 ;
  assign n36798 = n36795 | n36797 ;
  assign n36799 = n36794 | n36798 ;
  assign n36800 = n2936 & ~n28731 ;
  assign n36801 = ~n28518 & n36800 ;
  assign n36802 = n36799 | n36801 ;
  assign n36803 = n2936 | n36799 ;
  assign n36804 = ( n28720 & n36802 ) | ( n28720 & n36803 ) | ( n36802 & n36803 ) ;
  assign n36805 = x23 | n36804 ;
  assign n36806 = ~x23 & n36804 ;
  assign n36807 = ( ~n36804 & n36805 ) | ( ~n36804 & n36806 ) | ( n36805 & n36806 ) ;
  assign n36808 = ~n36793 & n36807 ;
  assign n36809 = n36792 | n36807 ;
  assign n36810 = n36791 & ~n36809 ;
  assign n36811 = n36808 | n36810 ;
  assign n36812 = n36510 | n36527 ;
  assign n36813 = ( n36510 & ~n36511 ) | ( n36510 & n36812 ) | ( ~n36511 & n36812 ) ;
  assign n36814 = n36811 | n36813 ;
  assign n36815 = n36811 & n36813 ;
  assign n36816 = n36814 & ~n36815 ;
  assign n36817 = n3547 & n30212 ;
  assign n36818 = n3544 & n29620 ;
  assign n36819 = n3541 & ~n30199 ;
  assign n36820 = n36818 | n36819 ;
  assign n36821 = n36817 | n36820 ;
  assign n36822 = n3537 & ~n30266 ;
  assign n36823 = ( n3537 & n30276 ) | ( n3537 & n36822 ) | ( n30276 & n36822 ) ;
  assign n36824 = n36821 | n36823 ;
  assign n36825 = x20 | n36821 ;
  assign n36826 = n36823 | n36825 ;
  assign n36827 = ~x20 & n36825 ;
  assign n36828 = ( ~x20 & n36823 ) | ( ~x20 & n36827 ) | ( n36823 & n36827 ) ;
  assign n36829 = ( ~n36824 & n36826 ) | ( ~n36824 & n36828 ) | ( n36826 & n36828 ) ;
  assign n36830 = ~n36816 & n36829 ;
  assign n36831 = n36811 | n36829 ;
  assign n36832 = ( n36813 & n36829 ) | ( n36813 & n36831 ) | ( n36829 & n36831 ) ;
  assign n36833 = n36814 & ~n36832 ;
  assign n36834 = n36830 | n36833 ;
  assign n36835 = n36537 | n36553 ;
  assign n36836 = ( n36537 & ~n36538 ) | ( n36537 & n36835 ) | ( ~n36538 & n36835 ) ;
  assign n36837 = n36834 | n36836 ;
  assign n36838 = n36834 & n36836 ;
  assign n36839 = n36837 & ~n36838 ;
  assign n36840 = n4471 & ~n31323 ;
  assign n36841 = n4466 & ~n30186 ;
  assign n36842 = n4468 & ~n31309 ;
  assign n36843 = n36841 | n36842 ;
  assign n36844 = n36840 | n36843 ;
  assign n36845 = n4475 & n31384 ;
  assign n36846 = n4475 & n31386 ;
  assign n36847 = ( ~n30232 & n36845 ) | ( ~n30232 & n36846 ) | ( n36845 & n36846 ) ;
  assign n36848 = n36844 | n36847 ;
  assign n36849 = n4475 | n36844 ;
  assign n36850 = ( ~n31376 & n36848 ) | ( ~n31376 & n36849 ) | ( n36848 & n36849 ) ;
  assign n36851 = x17 | n36850 ;
  assign n36852 = ~x17 & n36850 ;
  assign n36853 = ( ~n36850 & n36851 ) | ( ~n36850 & n36852 ) | ( n36851 & n36852 ) ;
  assign n36854 = ~n36839 & n36853 ;
  assign n36855 = n36834 | n36853 ;
  assign n36856 = ( n36836 & n36853 ) | ( n36836 & n36855 ) | ( n36853 & n36855 ) ;
  assign n36857 = n36837 & ~n36856 ;
  assign n36858 = n36854 | n36857 ;
  assign n36859 = ( n36562 & ~n36563 ) | ( n36562 & n36580 ) | ( ~n36563 & n36580 ) ;
  assign n36860 = n36858 | n36859 ;
  assign n36861 = n36858 & n36859 ;
  assign n36862 = n36860 & ~n36861 ;
  assign n36863 = n5234 & n32293 ;
  assign n36864 = n5237 & n31295 ;
  assign n36865 = n5231 & n32306 ;
  assign n36866 = n36864 | n36865 ;
  assign n36867 = n36863 | n36866 ;
  assign n36868 = n5227 & n32497 ;
  assign n36869 = ( n5227 & n32494 ) | ( n5227 & n36868 ) | ( n32494 & n36868 ) ;
  assign n36870 = n36867 | n36869 ;
  assign n36871 = x14 | n36867 ;
  assign n36872 = n36869 | n36871 ;
  assign n36873 = ~x14 & n36871 ;
  assign n36874 = ( ~x14 & n36869 ) | ( ~x14 & n36873 ) | ( n36869 & n36873 ) ;
  assign n36875 = ( ~n36870 & n36872 ) | ( ~n36870 & n36874 ) | ( n36872 & n36874 ) ;
  assign n36876 = ~n36862 & n36875 ;
  assign n36877 = n36858 | n36875 ;
  assign n36878 = ( n36859 & n36875 ) | ( n36859 & n36877 ) | ( n36875 & n36877 ) ;
  assign n36879 = n36860 & ~n36878 ;
  assign n36880 = n36876 | n36879 ;
  assign n36881 = n36586 | n36602 ;
  assign n36882 = ( n36586 & ~n36587 ) | ( n36586 & n36881 ) | ( ~n36587 & n36881 ) ;
  assign n36883 = n36880 | n36882 ;
  assign n36884 = n36880 & n36882 ;
  assign n36885 = n36883 & ~n36884 ;
  assign n36886 = n6122 & ~n33423 ;
  assign n36887 = n6125 & ~n32442 ;
  assign n36888 = n6119 & n33436 ;
  assign n36889 = n36887 | n36888 ;
  assign n36890 = n36886 | n36889 ;
  assign n36891 = n6115 & n33575 ;
  assign n36892 = n6115 & ~n33577 ;
  assign n36893 = ( ~n32456 & n36891 ) | ( ~n32456 & n36892 ) | ( n36891 & n36892 ) ;
  assign n36894 = n36890 | n36893 ;
  assign n36895 = n6115 | n36890 ;
  assign n36896 = ( n33567 & n36894 ) | ( n33567 & n36895 ) | ( n36894 & n36895 ) ;
  assign n36897 = x11 | n36896 ;
  assign n36898 = ~x11 & n36896 ;
  assign n36899 = ( ~n36896 & n36897 ) | ( ~n36896 & n36898 ) | ( n36897 & n36898 ) ;
  assign n36900 = ~n36885 & n36899 ;
  assign n36901 = n36880 | n36899 ;
  assign n36902 = ( n36882 & n36899 ) | ( n36882 & n36901 ) | ( n36899 & n36901 ) ;
  assign n36903 = n36883 & ~n36902 ;
  assign n36904 = n36900 | n36903 ;
  assign n36905 = ( n36611 & ~n36612 ) | ( n36611 & n36628 ) | ( ~n36612 & n36628 ) ;
  assign n36906 = n36904 | n36905 ;
  assign n36907 = n36904 & n36905 ;
  assign n36908 = n36906 & ~n36907 ;
  assign n36909 = n7079 & n35021 ;
  assign n36910 = n7074 & n33526 ;
  assign n36911 = n7068 & n34656 ;
  assign n36912 = n36910 | n36911 ;
  assign n36913 = n36909 | n36912 ;
  assign n36914 = n7078 | n36909 ;
  assign n36915 = n36912 | n36914 ;
  assign n36916 = ( n35033 & n36913 ) | ( n35033 & n36915 ) | ( n36913 & n36915 ) ;
  assign n36917 = x8 & n36915 ;
  assign n36918 = x8 & n36913 ;
  assign n36919 = ( n35033 & n36917 ) | ( n35033 & n36918 ) | ( n36917 & n36918 ) ;
  assign n36920 = x8 & ~n36918 ;
  assign n36921 = x8 & ~n36917 ;
  assign n36922 = ( ~n35033 & n36920 ) | ( ~n35033 & n36921 ) | ( n36920 & n36921 ) ;
  assign n36923 = ( n36916 & ~n36919 ) | ( n36916 & n36922 ) | ( ~n36919 & n36922 ) ;
  assign n36924 = ~n36908 & n36923 ;
  assign n36925 = n36904 | n36923 ;
  assign n36926 = ( n36905 & n36923 ) | ( n36905 & n36925 ) | ( n36923 & n36925 ) ;
  assign n36927 = n36906 & ~n36926 ;
  assign n36928 = n36924 | n36927 ;
  assign n36929 = n36634 | n36650 ;
  assign n36930 = ( n36634 & ~n36635 ) | ( n36634 & n36929 ) | ( ~n36635 & n36929 ) ;
  assign n36931 = n36928 | n36930 ;
  assign n36932 = n36928 & n36930 ;
  assign n36933 = n36931 & ~n36932 ;
  assign n36934 = n8122 & n36083 ;
  assign n36935 = n8115 & ~n35371 ;
  assign n36936 = n8118 & n35746 ;
  assign n36937 = n36935 | n36936 ;
  assign n36938 = n36934 | n36937 ;
  assign n36939 = n8125 | n36934 ;
  assign n36940 = n36937 | n36939 ;
  assign n36941 = ( n36107 & n36938 ) | ( n36107 & n36940 ) | ( n36938 & n36940 ) ;
  assign n36942 = n36938 | n36940 ;
  assign n36943 = ( n36094 & n36941 ) | ( n36094 & n36942 ) | ( n36941 & n36942 ) ;
  assign n36944 = x5 & n36943 ;
  assign n36945 = x5 & ~n36943 ;
  assign n36946 = ( n36943 & ~n36944 ) | ( n36943 & n36945 ) | ( ~n36944 & n36945 ) ;
  assign n36947 = ~n36933 & n36946 ;
  assign n36948 = n36928 | n36946 ;
  assign n36949 = ( n36930 & n36946 ) | ( n36930 & n36948 ) | ( n36946 & n36948 ) ;
  assign n36950 = n36931 & ~n36949 ;
  assign n36951 = n36947 | n36950 ;
  assign n36952 = n36660 | n36676 ;
  assign n36953 = ( n36660 & ~n36661 ) | ( n36660 & n36952 ) | ( ~n36661 & n36952 ) ;
  assign n36954 = n36951 | n36953 ;
  assign n36955 = n36951 & n36953 ;
  assign n36956 = n36954 & ~n36955 ;
  assign n36957 = n36684 | n36686 ;
  assign n36958 = ~n36684 & n36685 ;
  assign n36959 = ( n36405 & n36957 ) | ( n36405 & ~n36958 ) | ( n36957 & ~n36958 ) ;
  assign n36960 = n36956 | n36959 ;
  assign n36961 = n36956 & n36959 ;
  assign n36962 = n36960 & ~n36961 ;
  assign n36963 = n36693 & n36962 ;
  assign n36964 = n36693 | n36962 ;
  assign n36965 = ~n36963 & n36964 ;
  assign n36966 = n24771 & n36083 ;
  assign n36967 = n8115 & n35746 ;
  assign n36968 = n36966 | n36967 ;
  assign n36969 = n8125 | n36968 ;
  assign n36970 = ( n36103 & n36968 ) | ( n36103 & n36969 ) | ( n36968 & n36969 ) ;
  assign n36971 = ( n36105 & n36968 ) | ( n36105 & n36969 ) | ( n36968 & n36969 ) ;
  assign n36972 = ( n32456 & n36970 ) | ( n32456 & n36971 ) | ( n36970 & n36971 ) ;
  assign n36973 = x5 & n36972 ;
  assign n36974 = x5 & ~n36972 ;
  assign n36975 = ( n36972 & ~n36973 ) | ( n36972 & n36974 ) | ( ~n36973 & n36974 ) ;
  assign n36976 = n36907 | n36923 ;
  assign n36977 = ( n36907 & n36908 ) | ( n36907 & n36976 ) | ( n36908 & n36976 ) ;
  assign n36978 = n36975 & n36977 ;
  assign n36979 = n36975 | n36977 ;
  assign n36980 = ~n36978 & n36979 ;
  assign n36981 = n36764 | n36785 ;
  assign n37018 = n1057 & n26017 ;
  assign n37019 = n1060 & ~n25046 ;
  assign n37020 = n1065 & ~n25728 ;
  assign n37021 = n37019 | n37020 ;
  assign n37022 = n37018 | n37021 ;
  assign n37023 = n1062 | n37018 ;
  assign n37024 = n37021 | n37023 ;
  assign n37025 = ( n26613 & n37022 ) | ( n26613 & n37024 ) | ( n37022 & n37024 ) ;
  assign n37026 = n37022 | n37024 ;
  assign n37027 = ( n26605 & n37025 ) | ( n26605 & n37026 ) | ( n37025 & n37026 ) ;
  assign n36982 = n36718 | n36721 ;
  assign n36983 = n36718 | n36720 ;
  assign n36984 = ( n36448 & n36982 ) | ( n36448 & n36983 ) | ( n36982 & n36983 ) ;
  assign n36985 = n80 | n170 ;
  assign n36986 = n24284 | n36985 ;
  assign n36987 = n836 | n4184 ;
  assign n36988 = n36986 | n36987 ;
  assign n36989 = n18248 | n36988 ;
  assign n36990 = n1094 | n36989 ;
  assign n36991 = ( ~n5004 & n5993 ) | ( ~n5004 & n36990 ) | ( n5993 & n36990 ) ;
  assign n36992 = n5993 & n36990 ;
  assign n36993 = ( ~n5025 & n36991 ) | ( ~n5025 & n36992 ) | ( n36991 & n36992 ) ;
  assign n36994 = n5026 | n36993 ;
  assign n36995 = n702 | n710 ;
  assign n36996 = n12280 | n36995 ;
  assign n36997 = n126 | n36996 ;
  assign n36998 = n938 | n36997 ;
  assign n36999 = n1597 | n36998 ;
  assign n37000 = n318 | n839 ;
  assign n37001 = n348 | n418 ;
  assign n37002 = n37000 | n37001 ;
  assign n37003 = n36999 | n37002 ;
  assign n37004 = n36994 | n37003 ;
  assign n37005 = n36423 & n37004 ;
  assign n37006 = n36423 | n37004 ;
  assign n37007 = n36718 & n37006 ;
  assign n37008 = ~n37005 & n37007 ;
  assign n37009 = ~n37005 & n37006 ;
  assign n37010 = ( n36721 & n37008 ) | ( n36721 & n37009 ) | ( n37008 & n37009 ) ;
  assign n37011 = ( n36720 & n37008 ) | ( n36720 & n37009 ) | ( n37008 & n37009 ) ;
  assign n37012 = ( n36448 & n37010 ) | ( n36448 & n37011 ) | ( n37010 & n37011 ) ;
  assign n37013 = n36984 & ~n37012 ;
  assign n37014 = ~n36423 & n37006 ;
  assign n37015 = ~n37004 & n37006 ;
  assign n37016 = ( ~n36984 & n37014 ) | ( ~n36984 & n37015 ) | ( n37014 & n37015 ) ;
  assign n37017 = n37013 | n37016 ;
  assign n37028 = n37017 & n37027 ;
  assign n37029 = n37017 & ~n37028 ;
  assign n37030 = ( n37027 & ~n37028 ) | ( n37027 & n37029 ) | ( ~n37028 & n37029 ) ;
  assign n37031 = n36739 | n36743 ;
  assign n37032 = ( n36739 & n36745 ) | ( n36739 & n37031 ) | ( n36745 & n37031 ) ;
  assign n37033 = n37030 | n37032 ;
  assign n37034 = n37030 & n37032 ;
  assign n37035 = n37033 & ~n37034 ;
  assign n37036 = n1826 & ~n26270 ;
  assign n37037 = ~n26263 & n37036 ;
  assign n37038 = n1823 & ~n26526 ;
  assign n37039 = ~n26520 & n37038 ;
  assign n37040 = n37037 | n37039 ;
  assign n37041 = n1829 & ~n27133 ;
  assign n37042 = ~n27125 & n37041 ;
  assign n37043 = n37040 | n37042 ;
  assign n37044 = n1821 & n27699 ;
  assign n37045 = ( n1821 & ~n27696 ) | ( n1821 & n37044 ) | ( ~n27696 & n37044 ) ;
  assign n37046 = n37043 | n37045 ;
  assign n37047 = x29 | n37043 ;
  assign n37048 = n37045 | n37047 ;
  assign n37049 = ~x29 & n37047 ;
  assign n37050 = ( ~x29 & n37045 ) | ( ~x29 & n37049 ) | ( n37045 & n37049 ) ;
  assign n37051 = ( ~n37046 & n37048 ) | ( ~n37046 & n37050 ) | ( n37048 & n37050 ) ;
  assign n37052 = n37035 & n37051 ;
  assign n37053 = n37035 & ~n37052 ;
  assign n37054 = n2312 & ~n27371 ;
  assign n37055 = ~n27363 & n37054 ;
  assign n37056 = n2308 & ~n27606 ;
  assign n37057 = ~n27597 & n37056 ;
  assign n37058 = n37055 | n37057 ;
  assign n37059 = n2315 & ~n28503 ;
  assign n37060 = n28498 & n37059 ;
  assign n37061 = n37058 | n37060 ;
  assign n37062 = n2306 & n28794 ;
  assign n37063 = ( n2306 & n28783 ) | ( n2306 & n37062 ) | ( n28783 & n37062 ) ;
  assign n37064 = n37061 | n37063 ;
  assign n37065 = x26 | n37061 ;
  assign n37066 = n37063 | n37065 ;
  assign n37067 = ~x26 & n37065 ;
  assign n37068 = ( ~x26 & n37063 ) | ( ~x26 & n37067 ) | ( n37063 & n37067 ) ;
  assign n37069 = ( ~n37064 & n37066 ) | ( ~n37064 & n37068 ) | ( n37066 & n37068 ) ;
  assign n37070 = ~n37035 & n37051 ;
  assign n37071 = n37069 & n37070 ;
  assign n37072 = ( n37053 & n37069 ) | ( n37053 & n37071 ) | ( n37069 & n37071 ) ;
  assign n37073 = n37069 | n37070 ;
  assign n37074 = n37053 | n37073 ;
  assign n37075 = ~n37072 & n37074 ;
  assign n37076 = n36981 | n37075 ;
  assign n37077 = n36981 & n37075 ;
  assign n37078 = n37076 & ~n37077 ;
  assign n37079 = n2932 & n29620 ;
  assign n37080 = n2925 & n28492 ;
  assign n37081 = n2928 & ~n28714 ;
  assign n37082 = n37080 | n37081 ;
  assign n37083 = n37079 | n37082 ;
  assign n37084 = n2936 | n37079 ;
  assign n37085 = n37082 | n37084 ;
  assign n37086 = ( ~n29642 & n37083 ) | ( ~n29642 & n37085 ) | ( n37083 & n37085 ) ;
  assign n37087 = n37083 | n37085 ;
  assign n37088 = ( n29629 & n37086 ) | ( n29629 & n37087 ) | ( n37086 & n37087 ) ;
  assign n37089 = ~x23 & n37088 ;
  assign n37090 = x23 | n37088 ;
  assign n37091 = ( ~n37088 & n37089 ) | ( ~n37088 & n37090 ) | ( n37089 & n37090 ) ;
  assign n37092 = ~n37078 & n37091 ;
  assign n37093 = ( n36792 & n36793 ) | ( n36792 & n36809 ) | ( n36793 & n36809 ) ;
  assign n37094 = n36981 | n37091 ;
  assign n37095 = ( n37075 & n37091 ) | ( n37075 & n37094 ) | ( n37091 & n37094 ) ;
  assign n37096 = n37076 & ~n37095 ;
  assign n37097 = n37093 & n37096 ;
  assign n37098 = ( n37092 & n37093 ) | ( n37092 & n37097 ) | ( n37093 & n37097 ) ;
  assign n37099 = n37093 | n37096 ;
  assign n37100 = n37092 | n37099 ;
  assign n37101 = ~n37098 & n37100 ;
  assign n37102 = n3547 & ~n30186 ;
  assign n37103 = n3544 & ~n30199 ;
  assign n37104 = n3541 & n30212 ;
  assign n37105 = n37103 | n37104 ;
  assign n37106 = n37102 | n37105 ;
  assign n37107 = n3537 | n37102 ;
  assign n37108 = n37105 | n37107 ;
  assign n37109 = ( ~n30241 & n37106 ) | ( ~n30241 & n37108 ) | ( n37106 & n37108 ) ;
  assign n37110 = ~x20 & n37108 ;
  assign n37111 = ~x20 & n37106 ;
  assign n37112 = ( ~n30241 & n37110 ) | ( ~n30241 & n37111 ) | ( n37110 & n37111 ) ;
  assign n37113 = x20 | n37111 ;
  assign n37114 = x20 | n37110 ;
  assign n37115 = ( ~n30241 & n37113 ) | ( ~n30241 & n37114 ) | ( n37113 & n37114 ) ;
  assign n37116 = ( ~n37109 & n37112 ) | ( ~n37109 & n37115 ) | ( n37112 & n37115 ) ;
  assign n37117 = n37101 & n37116 ;
  assign n37118 = n37101 & ~n37117 ;
  assign n37120 = n36815 | n36829 ;
  assign n37121 = ( n36815 & n36816 ) | ( n36815 & n37120 ) | ( n36816 & n37120 ) ;
  assign n37119 = ~n37101 & n37116 ;
  assign n37122 = n37119 & n37121 ;
  assign n37123 = ( n37118 & n37121 ) | ( n37118 & n37122 ) | ( n37121 & n37122 ) ;
  assign n37124 = n37118 | n37119 ;
  assign n37125 = n37121 | n37124 ;
  assign n37126 = ~n37123 & n37125 ;
  assign n37127 = n4471 & n31295 ;
  assign n37128 = n4466 & ~n31309 ;
  assign n37129 = n4468 & ~n31323 ;
  assign n37130 = n37128 | n37129 ;
  assign n37131 = n37127 | n37130 ;
  assign n37132 = n4475 | n37127 ;
  assign n37133 = n37130 | n37132 ;
  assign n37134 = ( n31355 & n37131 ) | ( n31355 & n37133 ) | ( n37131 & n37133 ) ;
  assign n37135 = x17 & n37133 ;
  assign n37136 = x17 & n37131 ;
  assign n37137 = ( n31355 & n37135 ) | ( n31355 & n37136 ) | ( n37135 & n37136 ) ;
  assign n37138 = x17 & ~n37136 ;
  assign n37139 = x17 & ~n37135 ;
  assign n37140 = ( ~n31355 & n37138 ) | ( ~n31355 & n37139 ) | ( n37138 & n37139 ) ;
  assign n37141 = ( n37134 & ~n37137 ) | ( n37134 & n37140 ) | ( ~n37137 & n37140 ) ;
  assign n37142 = n37125 & n37141 ;
  assign n37143 = ~n37123 & n37142 ;
  assign n37144 = n37126 & ~n37143 ;
  assign n37145 = n36838 | n36853 ;
  assign n37146 = ( n36838 & n36839 ) | ( n36838 & n37145 ) | ( n36839 & n37145 ) ;
  assign n37147 = ~n37125 & n37141 ;
  assign n37148 = ( n37123 & n37141 ) | ( n37123 & n37147 ) | ( n37141 & n37147 ) ;
  assign n37149 = n37146 & n37148 ;
  assign n37150 = ( n37144 & n37146 ) | ( n37144 & n37149 ) | ( n37146 & n37149 ) ;
  assign n37151 = n37144 | n37148 ;
  assign n37152 = n37146 | n37151 ;
  assign n37153 = ~n37150 & n37152 ;
  assign n37154 = n5234 & ~n32442 ;
  assign n37155 = n5237 & n32306 ;
  assign n37156 = n5231 & n32293 ;
  assign n37157 = n37155 | n37156 ;
  assign n37158 = n37154 | n37157 ;
  assign n37159 = n5227 | n37154 ;
  assign n37160 = n37157 | n37159 ;
  assign n37161 = ( ~n32458 & n37158 ) | ( ~n32458 & n37160 ) | ( n37158 & n37160 ) ;
  assign n37162 = ~x14 & n37160 ;
  assign n37163 = ~x14 & n37158 ;
  assign n37164 = ( ~n32458 & n37162 ) | ( ~n32458 & n37163 ) | ( n37162 & n37163 ) ;
  assign n37165 = x14 | n37163 ;
  assign n37166 = x14 | n37162 ;
  assign n37167 = ( ~n32458 & n37165 ) | ( ~n32458 & n37166 ) | ( n37165 & n37166 ) ;
  assign n37168 = ( ~n37161 & n37164 ) | ( ~n37161 & n37167 ) | ( n37164 & n37167 ) ;
  assign n37169 = n37152 & ~n37168 ;
  assign n37170 = ~n37150 & n37169 ;
  assign n37171 = n37168 | n37170 ;
  assign n37172 = ( ~n37153 & n37170 ) | ( ~n37153 & n37171 ) | ( n37170 & n37171 ) ;
  assign n37173 = n36861 | n36875 ;
  assign n37174 = ( n36861 & n36862 ) | ( n36861 & n37173 ) | ( n36862 & n37173 ) ;
  assign n37175 = n37172 | n37174 ;
  assign n37176 = n37172 & n37174 ;
  assign n37177 = n37175 & ~n37176 ;
  assign n37178 = n6122 & n33526 ;
  assign n37179 = n6125 & n33436 ;
  assign n37180 = n6119 & ~n33423 ;
  assign n37181 = n37179 | n37180 ;
  assign n37182 = n37178 | n37181 ;
  assign n37183 = n6115 & n33545 ;
  assign n37184 = n6115 & ~n33548 ;
  assign n37185 = ( ~n32456 & n37183 ) | ( ~n32456 & n37184 ) | ( n37183 & n37184 ) ;
  assign n37186 = n37182 | n37185 ;
  assign n37187 = n6115 | n37182 ;
  assign n37188 = ( n33536 & n37186 ) | ( n33536 & n37187 ) | ( n37186 & n37187 ) ;
  assign n37189 = x11 | n37188 ;
  assign n37190 = ~x11 & n37188 ;
  assign n37191 = ( ~n37188 & n37189 ) | ( ~n37188 & n37190 ) | ( n37189 & n37190 ) ;
  assign n37192 = ~n37177 & n37191 ;
  assign n37193 = n37176 | n37191 ;
  assign n37194 = n37175 & ~n37193 ;
  assign n37195 = n37192 | n37194 ;
  assign n37196 = n36884 | n36899 ;
  assign n37197 = ( n36884 & n36885 ) | ( n36884 & n37196 ) | ( n36885 & n37196 ) ;
  assign n37198 = n37195 | n37197 ;
  assign n37199 = n37195 & n37197 ;
  assign n37200 = n37198 & ~n37199 ;
  assign n37201 = n7079 & ~n35371 ;
  assign n37202 = n7074 & n34656 ;
  assign n37203 = n7068 & n35021 ;
  assign n37204 = n37202 | n37203 ;
  assign n37205 = n37201 | n37204 ;
  assign n37206 = n7078 & ~n35392 ;
  assign n37207 = n7078 & ~n35395 ;
  assign n37208 = ( ~n32456 & n37206 ) | ( ~n32456 & n37207 ) | ( n37206 & n37207 ) ;
  assign n37209 = n37205 | n37208 ;
  assign n37210 = n7078 | n37205 ;
  assign n37211 = ( n35381 & n37209 ) | ( n35381 & n37210 ) | ( n37209 & n37210 ) ;
  assign n37212 = x8 | n37211 ;
  assign n37213 = ~x8 & n37211 ;
  assign n37214 = ( ~n37211 & n37212 ) | ( ~n37211 & n37213 ) | ( n37212 & n37213 ) ;
  assign n37215 = ~n37200 & n37214 ;
  assign n37216 = n37195 | n37214 ;
  assign n37217 = ( n37197 & n37214 ) | ( n37197 & n37216 ) | ( n37214 & n37216 ) ;
  assign n37218 = n37198 & ~n37217 ;
  assign n37219 = n37215 | n37218 ;
  assign n37220 = n36980 & ~n37219 ;
  assign n37221 = n36980 | n37219 ;
  assign n37222 = ( ~n36980 & n37220 ) | ( ~n36980 & n37221 ) | ( n37220 & n37221 ) ;
  assign n37223 = n36932 | n36946 ;
  assign n37224 = ( n36932 & n36933 ) | ( n36932 & n37223 ) | ( n36933 & n37223 ) ;
  assign n37225 = n37222 | n37224 ;
  assign n37226 = n37222 & n37224 ;
  assign n37227 = n37225 & ~n37226 ;
  assign n37228 = n36951 & n37227 ;
  assign n37229 = n36953 & n37228 ;
  assign n37230 = ( n36956 & n37227 ) | ( n36956 & n37229 ) | ( n37227 & n37229 ) ;
  assign n37231 = ( n36959 & n37229 ) | ( n36959 & n37230 ) | ( n37229 & n37230 ) ;
  assign n37232 = n36953 | n37227 ;
  assign n37233 = n36951 | n37227 ;
  assign n37234 = ( n36959 & n37232 ) | ( n36959 & n37233 ) | ( n37232 & n37233 ) ;
  assign n37235 = ~n37231 & n37234 ;
  assign n37236 = n36963 & n37235 ;
  assign n37237 = n36963 | n37235 ;
  assign n37238 = ~n37236 & n37237 ;
  assign n37239 = n37052 | n37072 ;
  assign n37240 = ( n36423 & n36984 ) | ( n36423 & n37004 ) | ( n36984 & n37004 ) ;
  assign n37241 = ~x5 & n8125 ;
  assign n37242 = ( ~x5 & n25463 ) | ( ~x5 & n37241 ) | ( n25463 & n37241 ) ;
  assign n37243 = n36083 & n37242 ;
  assign n37244 = x5 & ~n8125 ;
  assign n37245 = ~n25463 & n37244 ;
  assign n37246 = ( x5 & ~n36083 ) | ( x5 & n37245 ) | ( ~n36083 & n37245 ) ;
  assign n37247 = n37243 | n37246 ;
  assign n37248 = n1473 | n9151 ;
  assign n37249 = n1636 | n3282 ;
  assign n37250 = n37248 | n37249 ;
  assign n37251 = n28524 | n37250 ;
  assign n37252 = n18122 | n37251 ;
  assign n37253 = n2759 | n11388 ;
  assign n37254 = n2765 | n37253 ;
  assign n37255 = n2751 | n37254 ;
  assign n37256 = n314 | n1398 ;
  assign n37257 = n433 | n37256 ;
  assign n37258 = n22501 | n37257 ;
  assign n37259 = n22497 | n37258 ;
  assign n37260 = n176 | n406 ;
  assign n37261 = n75 | n37260 ;
  assign n37262 = n37259 | n37261 ;
  assign n37263 = n37255 | n37262 ;
  assign n37264 = n37252 | n37263 ;
  assign n37265 = n443 | n37264 ;
  assign n37266 = n36423 | n37265 ;
  assign n37267 = n36423 & n37265 ;
  assign n37268 = n37266 & ~n37267 ;
  assign n37269 = n37247 | n37268 ;
  assign n37270 = ~n37268 & n37269 ;
  assign n37271 = ( ~n37247 & n37269 ) | ( ~n37247 & n37270 ) | ( n37269 & n37270 ) ;
  assign n37272 = n37240 & ~n37271 ;
  assign n37273 = ~n37240 & n37271 ;
  assign n37274 = n37272 | n37273 ;
  assign n37275 = n1060 & ~n25728 ;
  assign n37276 = n1065 & n26017 ;
  assign n37277 = n37275 | n37276 ;
  assign n37278 = n1057 & ~n26270 ;
  assign n37279 = ~n26263 & n37278 ;
  assign n37280 = n37277 | n37279 ;
  assign n37281 = n1062 | n37279 ;
  assign n37282 = n37277 | n37281 ;
  assign n37283 = ( n26571 & n37280 ) | ( n26571 & n37282 ) | ( n37280 & n37282 ) ;
  assign n37284 = n37274 & n37283 ;
  assign n37285 = n37274 | n37283 ;
  assign n37286 = ~n37284 & n37285 ;
  assign n37287 = n37028 | n37030 ;
  assign n37288 = ( n37028 & n37032 ) | ( n37028 & n37287 ) | ( n37032 & n37287 ) ;
  assign n37289 = n37286 | n37288 ;
  assign n37290 = n37286 & n37288 ;
  assign n37291 = n37289 & ~n37290 ;
  assign n37292 = n1826 & ~n26526 ;
  assign n37293 = ~n26520 & n37292 ;
  assign n37294 = n1823 & ~n27133 ;
  assign n37295 = ~n27125 & n37294 ;
  assign n37296 = n37293 | n37295 ;
  assign n37297 = n1829 & ~n27371 ;
  assign n37298 = ~n27363 & n37297 ;
  assign n37299 = n37296 | n37298 ;
  assign n37300 = n1821 | n37298 ;
  assign n37301 = n37296 | n37300 ;
  assign n37302 = ( ~n27654 & n37299 ) | ( ~n27654 & n37301 ) | ( n37299 & n37301 ) ;
  assign n37303 = ~x29 & n37301 ;
  assign n37304 = ~x29 & n37299 ;
  assign n37305 = ( ~n27654 & n37303 ) | ( ~n27654 & n37304 ) | ( n37303 & n37304 ) ;
  assign n37306 = x29 | n37304 ;
  assign n37307 = x29 | n37303 ;
  assign n37308 = ( ~n27654 & n37306 ) | ( ~n27654 & n37307 ) | ( n37306 & n37307 ) ;
  assign n37309 = ( ~n37302 & n37305 ) | ( ~n37302 & n37308 ) | ( n37305 & n37308 ) ;
  assign n37310 = ~n37291 & n37309 ;
  assign n37311 = n2315 & n28492 ;
  assign n37312 = n2312 & ~n27606 ;
  assign n37313 = ~n27597 & n37312 ;
  assign n37314 = n2308 & ~n28503 ;
  assign n37315 = n28498 & n37314 ;
  assign n37316 = n37313 | n37315 ;
  assign n37317 = n37311 | n37316 ;
  assign n37318 = n2306 | n37317 ;
  assign n37319 = ( ~n28749 & n37317 ) | ( ~n28749 & n37318 ) | ( n37317 & n37318 ) ;
  assign n37320 = ~x26 & n37318 ;
  assign n37321 = ~x26 & n37317 ;
  assign n37322 = ( ~n28749 & n37320 ) | ( ~n28749 & n37321 ) | ( n37320 & n37321 ) ;
  assign n37323 = x26 | n37320 ;
  assign n37324 = x26 | n37321 ;
  assign n37325 = ( ~n28749 & n37323 ) | ( ~n28749 & n37324 ) | ( n37323 & n37324 ) ;
  assign n37326 = ( ~n37319 & n37322 ) | ( ~n37319 & n37325 ) | ( n37322 & n37325 ) ;
  assign n37327 = n37286 | n37309 ;
  assign n37328 = ( n37288 & n37309 ) | ( n37288 & n37327 ) | ( n37309 & n37327 ) ;
  assign n37329 = n37289 & ~n37328 ;
  assign n37330 = n37326 & n37329 ;
  assign n37331 = ( n37310 & n37326 ) | ( n37310 & n37330 ) | ( n37326 & n37330 ) ;
  assign n37332 = n37326 | n37329 ;
  assign n37333 = n37310 | n37332 ;
  assign n37334 = ~n37331 & n37333 ;
  assign n37335 = n37239 | n37334 ;
  assign n37336 = n37239 & n37334 ;
  assign n37337 = n37335 & ~n37336 ;
  assign n37338 = n2932 & ~n30199 ;
  assign n37339 = n2925 & ~n28714 ;
  assign n37340 = n2928 & n29620 ;
  assign n37341 = n37339 | n37340 ;
  assign n37342 = n37338 | n37341 ;
  assign n37343 = n2936 | n37338 ;
  assign n37344 = n37341 | n37343 ;
  assign n37345 = ( ~n30299 & n37342 ) | ( ~n30299 & n37344 ) | ( n37342 & n37344 ) ;
  assign n37346 = ~x23 & n37344 ;
  assign n37347 = ~x23 & n37342 ;
  assign n37348 = ( ~n30299 & n37346 ) | ( ~n30299 & n37347 ) | ( n37346 & n37347 ) ;
  assign n37349 = x23 | n37347 ;
  assign n37350 = x23 | n37346 ;
  assign n37351 = ( ~n30299 & n37349 ) | ( ~n30299 & n37350 ) | ( n37349 & n37350 ) ;
  assign n37352 = ( ~n37345 & n37348 ) | ( ~n37345 & n37351 ) | ( n37348 & n37351 ) ;
  assign n37353 = n37337 & n37352 ;
  assign n37354 = n37337 & ~n37353 ;
  assign n37356 = n37077 | n37091 ;
  assign n37357 = ( n37077 & n37078 ) | ( n37077 & n37356 ) | ( n37078 & n37356 ) ;
  assign n37355 = ~n37337 & n37352 ;
  assign n37358 = n37355 & n37357 ;
  assign n37359 = ( n37354 & n37357 ) | ( n37354 & n37358 ) | ( n37357 & n37358 ) ;
  assign n37360 = n37355 | n37357 ;
  assign n37361 = n37354 | n37360 ;
  assign n37362 = ~n37359 & n37361 ;
  assign n37363 = n3547 & ~n31309 ;
  assign n37364 = n3544 & n30212 ;
  assign n37365 = n3541 & ~n30186 ;
  assign n37366 = n37364 | n37365 ;
  assign n37367 = n37363 | n37366 ;
  assign n37368 = n3537 | n37363 ;
  assign n37369 = n37366 | n37368 ;
  assign n37370 = ( n31404 & n37367 ) | ( n31404 & n37369 ) | ( n37367 & n37369 ) ;
  assign n37371 = x20 & n37369 ;
  assign n37372 = x20 & n37367 ;
  assign n37373 = ( n31404 & n37371 ) | ( n31404 & n37372 ) | ( n37371 & n37372 ) ;
  assign n37374 = x20 & ~n37372 ;
  assign n37375 = x20 & ~n37371 ;
  assign n37376 = ( ~n31404 & n37374 ) | ( ~n31404 & n37375 ) | ( n37374 & n37375 ) ;
  assign n37377 = ( n37370 & ~n37373 ) | ( n37370 & n37376 ) | ( ~n37373 & n37376 ) ;
  assign n37378 = n37362 & n37377 ;
  assign n37379 = n37362 & ~n37378 ;
  assign n37381 = n37098 | n37116 ;
  assign n37382 = ( n37098 & n37101 ) | ( n37098 & n37381 ) | ( n37101 & n37381 ) ;
  assign n37380 = ~n37362 & n37377 ;
  assign n37383 = n37380 & n37382 ;
  assign n37384 = ( n37379 & n37382 ) | ( n37379 & n37383 ) | ( n37382 & n37383 ) ;
  assign n37385 = n37380 | n37382 ;
  assign n37386 = n37379 | n37385 ;
  assign n37387 = ~n37384 & n37386 ;
  assign n37388 = n4471 & n32306 ;
  assign n37389 = n4466 & ~n31323 ;
  assign n37390 = n4468 & n31295 ;
  assign n37391 = n37389 | n37390 ;
  assign n37392 = n37388 | n37391 ;
  assign n37393 = n4475 | n37388 ;
  assign n37394 = n37391 | n37393 ;
  assign n37395 = ( ~n32525 & n37392 ) | ( ~n32525 & n37394 ) | ( n37392 & n37394 ) ;
  assign n37396 = ~x17 & n37394 ;
  assign n37397 = ~x17 & n37392 ;
  assign n37398 = ( ~n32525 & n37396 ) | ( ~n32525 & n37397 ) | ( n37396 & n37397 ) ;
  assign n37399 = x17 | n37397 ;
  assign n37400 = x17 | n37396 ;
  assign n37401 = ( ~n32525 & n37399 ) | ( ~n32525 & n37400 ) | ( n37399 & n37400 ) ;
  assign n37402 = ( ~n37395 & n37398 ) | ( ~n37395 & n37401 ) | ( n37398 & n37401 ) ;
  assign n37403 = n37387 & n37402 ;
  assign n37404 = n37387 & ~n37403 ;
  assign n37405 = n37123 | n37143 ;
  assign n37406 = ~n37387 & n37402 ;
  assign n37407 = n37405 & n37406 ;
  assign n37408 = ( n37404 & n37405 ) | ( n37404 & n37407 ) | ( n37405 & n37407 ) ;
  assign n37409 = n37405 | n37406 ;
  assign n37410 = n37404 | n37409 ;
  assign n37411 = ~n37408 & n37410 ;
  assign n37412 = n37152 & n37168 ;
  assign n37413 = ~n37150 & n37412 ;
  assign n37414 = n37150 | n37413 ;
  assign n37415 = n5234 & n33436 ;
  assign n37416 = n5237 & n32293 ;
  assign n37417 = n5231 & ~n32442 ;
  assign n37418 = n37416 | n37417 ;
  assign n37419 = n37415 | n37418 ;
  assign n37420 = n5227 & ~n33441 ;
  assign n37421 = ~n32456 & n37420 ;
  assign n37422 = ( n5227 & n34271 ) | ( n5227 & n37421 ) | ( n34271 & n37421 ) ;
  assign n37423 = n37419 | n37422 ;
  assign n37424 = x14 | n37419 ;
  assign n37425 = n37422 | n37424 ;
  assign n37426 = ~x14 & n37424 ;
  assign n37427 = ( ~x14 & n37422 ) | ( ~x14 & n37426 ) | ( n37422 & n37426 ) ;
  assign n37428 = ( ~n37423 & n37425 ) | ( ~n37423 & n37427 ) | ( n37425 & n37427 ) ;
  assign n37429 = n37150 & n37428 ;
  assign n37430 = ( n37413 & n37428 ) | ( n37413 & n37429 ) | ( n37428 & n37429 ) ;
  assign n37431 = n37414 & ~n37430 ;
  assign n37432 = ~n37150 & n37428 ;
  assign n37433 = ~n37413 & n37432 ;
  assign n37434 = n37411 & n37433 ;
  assign n37435 = ( n37411 & n37431 ) | ( n37411 & n37434 ) | ( n37431 & n37434 ) ;
  assign n37436 = n37411 | n37433 ;
  assign n37437 = n37431 | n37436 ;
  assign n37438 = ~n37435 & n37437 ;
  assign n37439 = n6122 & n34656 ;
  assign n37440 = n6125 & ~n33423 ;
  assign n37441 = n6119 & n33526 ;
  assign n37442 = n37440 | n37441 ;
  assign n37443 = n37439 | n37442 ;
  assign n37444 = n6115 | n37439 ;
  assign n37445 = n37442 | n37444 ;
  assign n37446 = ( n34667 & n37443 ) | ( n34667 & n37445 ) | ( n37443 & n37445 ) ;
  assign n37447 = x11 & n37445 ;
  assign n37448 = x11 & n37443 ;
  assign n37449 = ( n34667 & n37447 ) | ( n34667 & n37448 ) | ( n37447 & n37448 ) ;
  assign n37450 = x11 & ~n37448 ;
  assign n37451 = x11 & ~n37447 ;
  assign n37452 = ( ~n34667 & n37450 ) | ( ~n34667 & n37451 ) | ( n37450 & n37451 ) ;
  assign n37453 = ( n37446 & ~n37449 ) | ( n37446 & n37452 ) | ( ~n37449 & n37452 ) ;
  assign n37454 = n37438 & n37453 ;
  assign n37455 = n37438 & ~n37454 ;
  assign n37457 = ( n37176 & n37177 ) | ( n37176 & n37193 ) | ( n37177 & n37193 ) ;
  assign n37456 = ~n37438 & n37453 ;
  assign n37458 = n37456 & n37457 ;
  assign n37459 = ( n37455 & n37457 ) | ( n37455 & n37458 ) | ( n37457 & n37458 ) ;
  assign n37460 = n37456 | n37457 ;
  assign n37461 = n37455 | n37460 ;
  assign n37462 = ~n37459 & n37461 ;
  assign n37478 = n37199 | n37214 ;
  assign n37479 = ( n37199 & n37200 ) | ( n37199 & n37478 ) | ( n37200 & n37478 ) ;
  assign n37463 = n7079 & n35746 ;
  assign n37464 = n7074 & n35021 ;
  assign n37465 = n7068 & ~n35371 ;
  assign n37466 = n37464 | n37465 ;
  assign n37467 = n37463 | n37466 ;
  assign n37468 = n7078 | n37463 ;
  assign n37469 = n37466 | n37468 ;
  assign n37470 = ( ~n35759 & n37467 ) | ( ~n35759 & n37469 ) | ( n37467 & n37469 ) ;
  assign n37471 = ~x8 & n37469 ;
  assign n37472 = ~x8 & n37467 ;
  assign n37473 = ( ~n35759 & n37471 ) | ( ~n35759 & n37472 ) | ( n37471 & n37472 ) ;
  assign n37474 = x8 | n37472 ;
  assign n37475 = x8 | n37471 ;
  assign n37476 = ( ~n35759 & n37474 ) | ( ~n35759 & n37475 ) | ( n37474 & n37475 ) ;
  assign n37477 = ( ~n37470 & n37473 ) | ( ~n37470 & n37476 ) | ( n37473 & n37476 ) ;
  assign n37480 = n37477 & n37479 ;
  assign n37481 = n37479 & ~n37480 ;
  assign n37482 = n37462 & n37477 ;
  assign n37483 = ~n37479 & n37482 ;
  assign n37484 = ( n37462 & n37481 ) | ( n37462 & n37483 ) | ( n37481 & n37483 ) ;
  assign n37485 = n37462 | n37477 ;
  assign n37486 = ( n37462 & ~n37479 ) | ( n37462 & n37485 ) | ( ~n37479 & n37485 ) ;
  assign n37487 = n37481 | n37486 ;
  assign n37488 = ~n37484 & n37487 ;
  assign n37489 = n36978 | n37219 ;
  assign n37490 = ( n36978 & n36980 ) | ( n36978 & n37489 ) | ( n36980 & n37489 ) ;
  assign n37491 = n37488 & n37490 ;
  assign n37492 = n37488 | n37490 ;
  assign n37493 = ~n37491 & n37492 ;
  assign n37494 = n37226 | n37229 ;
  assign n37495 = n37226 | n37227 ;
  assign n37496 = ( n36956 & n37494 ) | ( n36956 & n37495 ) | ( n37494 & n37495 ) ;
  assign n37497 = n37493 & n37496 ;
  assign n37498 = n37226 & n37493 ;
  assign n37499 = ( n37229 & n37493 ) | ( n37229 & n37498 ) | ( n37493 & n37498 ) ;
  assign n37500 = ( n36959 & n37497 ) | ( n36959 & n37499 ) | ( n37497 & n37499 ) ;
  assign n37501 = n37493 | n37496 ;
  assign n37502 = n37493 | n37494 ;
  assign n37503 = ( n36959 & n37501 ) | ( n36959 & n37502 ) | ( n37501 & n37502 ) ;
  assign n37504 = ~n37500 & n37503 ;
  assign n37505 = n37236 | n37504 ;
  assign n37506 = n37235 & n37504 ;
  assign n37507 = n36963 & n37506 ;
  assign n37508 = n37505 & ~n37507 ;
  assign n37671 = n37403 | n37405 ;
  assign n37672 = n37403 | n37404 ;
  assign n37673 = ( n37407 & n37671 ) | ( n37407 & n37672 ) | ( n37671 & n37672 ) ;
  assign n37547 = n1060 & n26017 ;
  assign n37548 = n1065 & ~n26270 ;
  assign n37549 = ~n26263 & n37548 ;
  assign n37550 = n37547 | n37549 ;
  assign n37551 = n1057 & ~n26526 ;
  assign n37552 = ~n26520 & n37551 ;
  assign n37553 = n37550 | n37552 ;
  assign n37554 = n1062 | n37552 ;
  assign n37555 = n37550 | n37554 ;
  assign n37556 = ( ~n26555 & n37553 ) | ( ~n26555 & n37555 ) | ( n37553 & n37555 ) ;
  assign n37557 = ( n26528 & n37553 ) | ( n26528 & n37555 ) | ( n37553 & n37555 ) ;
  assign n37558 = ( ~n26543 & n37556 ) | ( ~n26543 & n37557 ) | ( n37556 & n37557 ) ;
  assign n37509 = n125 | n1662 ;
  assign n37510 = n11077 | n37509 ;
  assign n37511 = n2604 | n4144 ;
  assign n37512 = n37510 | n37511 ;
  assign n37513 = n937 | n1416 ;
  assign n37514 = n37512 | n37513 ;
  assign n37515 = n1523 | n7001 ;
  assign n37516 = n7000 | n37515 ;
  assign n37517 = n37514 | n37516 ;
  assign n37518 = n1650 | n2846 ;
  assign n37519 = n12274 | n37518 ;
  assign n37520 = n1435 | n37519 ;
  assign n37521 = n249 | n602 ;
  assign n37522 = n1303 | n37521 ;
  assign n37523 = n64 | n193 ;
  assign n37524 = n37522 | n37523 ;
  assign n37525 = n37520 | n37524 ;
  assign n37526 = n37517 | n37525 ;
  assign n37527 = n914 | n3429 ;
  assign n37528 = n5100 | n37527 ;
  assign n37529 = n37526 | n37528 ;
  assign n37530 = n419 | n1675 ;
  assign n37531 = n839 | n3330 ;
  assign n37532 = n37530 | n37531 ;
  assign n37533 = n202 | n901 ;
  assign n37534 = n444 | n37533 ;
  assign n37535 = n435 | n37534 ;
  assign n37536 = n37532 | n37535 ;
  assign n37537 = n277 | n37536 ;
  assign n37538 = n5978 | n37537 ;
  assign n37539 = n37529 | n37538 ;
  assign n37540 = n332 | n37539 ;
  assign n37541 = ~n36423 & n37265 ;
  assign n37542 = n37247 & ~n37541 ;
  assign n37543 = ( n37268 & ~n37541 ) | ( n37268 & n37542 ) | ( ~n37541 & n37542 ) ;
  assign n37544 = n37540 | n37543 ;
  assign n37545 = n37540 & n37543 ;
  assign n37546 = n37544 & ~n37545 ;
  assign n37559 = n37546 & n37558 ;
  assign n37560 = n37546 & ~n37558 ;
  assign n37561 = ( n37558 & ~n37559 ) | ( n37558 & n37560 ) | ( ~n37559 & n37560 ) ;
  assign n37562 = ( n37240 & n37271 ) | ( n37240 & n37283 ) | ( n37271 & n37283 ) ;
  assign n37563 = n37561 | n37562 ;
  assign n37564 = n37561 & n37562 ;
  assign n37565 = n37563 & ~n37564 ;
  assign n37566 = n1826 & ~n27133 ;
  assign n37567 = ~n27125 & n37566 ;
  assign n37568 = n1823 & ~n27371 ;
  assign n37569 = ~n27363 & n37568 ;
  assign n37570 = n37567 | n37569 ;
  assign n37571 = n1829 & ~n27606 ;
  assign n37572 = ~n27597 & n37571 ;
  assign n37573 = n37570 | n37572 ;
  assign n37574 = n27630 | n37573 ;
  assign n37575 = ( ~n27625 & n37573 ) | ( ~n27625 & n37574 ) | ( n37573 & n37574 ) ;
  assign n37576 = n27634 & ~n37575 ;
  assign n37577 = n1821 | n37572 ;
  assign n37578 = n37570 | n37577 ;
  assign n37579 = ~n37576 & n37578 ;
  assign n37580 = x29 & n37578 ;
  assign n37581 = ~n37576 & n37580 ;
  assign n37582 = x29 & ~n37580 ;
  assign n37583 = ( x29 & n37576 ) | ( x29 & n37582 ) | ( n37576 & n37582 ) ;
  assign n37584 = ( n37579 & ~n37581 ) | ( n37579 & n37583 ) | ( ~n37581 & n37583 ) ;
  assign n37585 = n37565 & n37584 ;
  assign n37586 = n37565 | n37584 ;
  assign n37587 = ~n37585 & n37586 ;
  assign n37588 = n37290 | n37309 ;
  assign n37589 = ( n37290 & n37291 ) | ( n37290 & n37588 ) | ( n37291 & n37588 ) ;
  assign n37590 = n37587 & n37589 ;
  assign n37591 = n37587 | n37589 ;
  assign n37592 = ~n37590 & n37591 ;
  assign n37593 = n2315 & ~n28714 ;
  assign n37594 = n2308 & n28492 ;
  assign n37595 = n2312 & ~n28503 ;
  assign n37596 = n28498 & n37595 ;
  assign n37597 = n37594 | n37596 ;
  assign n37598 = n37593 | n37597 ;
  assign n37599 = n2306 & ~n28731 ;
  assign n37600 = ~n28518 & n37599 ;
  assign n37601 = n37598 | n37600 ;
  assign n37602 = n2306 | n37598 ;
  assign n37603 = ( n28720 & n37601 ) | ( n28720 & n37602 ) | ( n37601 & n37602 ) ;
  assign n37604 = x26 | n37603 ;
  assign n37605 = ~x26 & n37603 ;
  assign n37606 = ( ~n37603 & n37604 ) | ( ~n37603 & n37605 ) | ( n37604 & n37605 ) ;
  assign n37607 = n37592 & ~n37606 ;
  assign n37608 = n37592 | n37606 ;
  assign n37609 = ( ~n37592 & n37607 ) | ( ~n37592 & n37608 ) | ( n37607 & n37608 ) ;
  assign n37610 = n37331 | n37336 ;
  assign n37611 = n37609 | n37610 ;
  assign n37612 = n37609 & n37610 ;
  assign n37613 = n37611 & ~n37612 ;
  assign n37614 = n2932 & n30212 ;
  assign n37615 = n2925 & n29620 ;
  assign n37616 = n2928 & ~n30199 ;
  assign n37617 = n37615 | n37616 ;
  assign n37618 = n37614 | n37617 ;
  assign n37619 = n2936 & ~n30266 ;
  assign n37620 = ( n2936 & n30276 ) | ( n2936 & n37619 ) | ( n30276 & n37619 ) ;
  assign n37621 = n37618 | n37620 ;
  assign n37622 = x23 | n37618 ;
  assign n37623 = n37620 | n37622 ;
  assign n37624 = ~x23 & n37622 ;
  assign n37625 = ( ~x23 & n37620 ) | ( ~x23 & n37624 ) | ( n37620 & n37624 ) ;
  assign n37626 = ( ~n37621 & n37623 ) | ( ~n37621 & n37625 ) | ( n37623 & n37625 ) ;
  assign n37627 = ~n37613 & n37626 ;
  assign n37628 = n37612 | n37626 ;
  assign n37629 = n37611 & ~n37628 ;
  assign n37630 = n37627 | n37629 ;
  assign n37631 = n37353 | n37359 ;
  assign n37632 = n37630 | n37631 ;
  assign n37633 = n37630 & n37631 ;
  assign n37634 = n37632 & ~n37633 ;
  assign n37635 = n3547 & ~n31323 ;
  assign n37636 = n3544 & ~n30186 ;
  assign n37637 = n3541 & ~n31309 ;
  assign n37638 = n37636 | n37637 ;
  assign n37639 = n37635 | n37638 ;
  assign n37640 = n3537 & n31384 ;
  assign n37641 = n3537 & n31386 ;
  assign n37642 = ( ~n30232 & n37640 ) | ( ~n30232 & n37641 ) | ( n37640 & n37641 ) ;
  assign n37643 = n37639 | n37642 ;
  assign n37644 = n3537 | n37639 ;
  assign n37645 = ( ~n31376 & n37643 ) | ( ~n31376 & n37644 ) | ( n37643 & n37644 ) ;
  assign n37646 = x20 | n37645 ;
  assign n37647 = ~x20 & n37645 ;
  assign n37648 = ( ~n37645 & n37646 ) | ( ~n37645 & n37647 ) | ( n37646 & n37647 ) ;
  assign n37649 = ~n37634 & n37648 ;
  assign n37650 = n37633 | n37648 ;
  assign n37651 = n37632 & ~n37650 ;
  assign n37652 = n37649 | n37651 ;
  assign n37653 = n37378 | n37384 ;
  assign n37654 = n37652 | n37653 ;
  assign n37655 = n37652 & n37653 ;
  assign n37656 = n37654 & ~n37655 ;
  assign n37657 = n4471 & n32293 ;
  assign n37658 = n4466 & n31295 ;
  assign n37659 = n4468 & n32306 ;
  assign n37660 = n37658 | n37659 ;
  assign n37661 = n37657 | n37660 ;
  assign n37662 = n4475 & n32497 ;
  assign n37663 = ( n4475 & n32494 ) | ( n4475 & n37662 ) | ( n32494 & n37662 ) ;
  assign n37664 = n37661 | n37663 ;
  assign n37665 = x17 | n37661 ;
  assign n37666 = n37663 | n37665 ;
  assign n37667 = ~x17 & n37665 ;
  assign n37668 = ( ~x17 & n37663 ) | ( ~x17 & n37667 ) | ( n37663 & n37667 ) ;
  assign n37669 = ( ~n37664 & n37666 ) | ( ~n37664 & n37668 ) | ( n37666 & n37668 ) ;
  assign n37670 = ~n37656 & n37669 ;
  assign n37674 = n37670 & n37673 ;
  assign n37675 = n37655 | n37669 ;
  assign n37676 = n37654 & ~n37675 ;
  assign n37677 = ( n37673 & n37674 ) | ( n37673 & n37676 ) | ( n37674 & n37676 ) ;
  assign n37678 = n37670 | n37676 ;
  assign n37679 = n37673 | n37678 ;
  assign n37680 = ~n37677 & n37679 ;
  assign n37681 = n5234 & ~n33423 ;
  assign n37682 = n5237 & ~n32442 ;
  assign n37683 = n5231 & n33436 ;
  assign n37684 = n37682 | n37683 ;
  assign n37685 = n37681 | n37684 ;
  assign n37686 = n5227 & n33575 ;
  assign n37687 = n5227 & ~n33577 ;
  assign n37688 = ( ~n32456 & n37686 ) | ( ~n32456 & n37687 ) | ( n37686 & n37687 ) ;
  assign n37689 = n37685 | n37688 ;
  assign n37690 = n5227 | n37685 ;
  assign n37691 = ( n33567 & n37689 ) | ( n33567 & n37690 ) | ( n37689 & n37690 ) ;
  assign n37692 = x14 | n37691 ;
  assign n37693 = ~x14 & n37691 ;
  assign n37694 = ( ~n37691 & n37692 ) | ( ~n37691 & n37693 ) | ( n37692 & n37693 ) ;
  assign n37695 = n37679 & n37694 ;
  assign n37696 = ~n37677 & n37695 ;
  assign n37697 = n37680 & ~n37696 ;
  assign n37698 = ~n37679 & n37694 ;
  assign n37699 = ( n37677 & n37694 ) | ( n37677 & n37698 ) | ( n37694 & n37698 ) ;
  assign n37700 = n37697 | n37699 ;
  assign n37701 = n37430 & n37700 ;
  assign n37702 = ( n37435 & n37700 ) | ( n37435 & n37701 ) | ( n37700 & n37701 ) ;
  assign n37703 = n37430 | n37700 ;
  assign n37704 = n37435 | n37703 ;
  assign n37705 = ~n37702 & n37704 ;
  assign n37706 = n6122 & n35021 ;
  assign n37707 = n6125 & n33526 ;
  assign n37708 = n6119 & n34656 ;
  assign n37709 = n37707 | n37708 ;
  assign n37710 = n37706 | n37709 ;
  assign n37711 = n6115 | n37706 ;
  assign n37712 = n37709 | n37711 ;
  assign n37713 = ( n35033 & n37710 ) | ( n35033 & n37712 ) | ( n37710 & n37712 ) ;
  assign n37714 = x11 & n37712 ;
  assign n37715 = x11 & n37710 ;
  assign n37716 = ( n35033 & n37714 ) | ( n35033 & n37715 ) | ( n37714 & n37715 ) ;
  assign n37717 = x11 & ~n37715 ;
  assign n37718 = x11 & ~n37714 ;
  assign n37719 = ( ~n35033 & n37717 ) | ( ~n35033 & n37718 ) | ( n37717 & n37718 ) ;
  assign n37720 = ( n37713 & ~n37716 ) | ( n37713 & n37719 ) | ( ~n37716 & n37719 ) ;
  assign n37721 = n37705 & n37720 ;
  assign n37722 = n37705 & ~n37721 ;
  assign n37723 = n37454 | n37459 ;
  assign n37724 = ~n37705 & n37720 ;
  assign n37725 = n37454 & n37724 ;
  assign n37726 = ( n37459 & n37724 ) | ( n37459 & n37725 ) | ( n37724 & n37725 ) ;
  assign n37727 = ( n37722 & n37723 ) | ( n37722 & n37726 ) | ( n37723 & n37726 ) ;
  assign n37728 = n37454 | n37724 ;
  assign n37729 = n37459 | n37728 ;
  assign n37730 = n37722 | n37729 ;
  assign n37731 = ~n37727 & n37730 ;
  assign n37732 = n7079 & n36083 ;
  assign n37733 = n7074 & ~n35371 ;
  assign n37734 = n7068 & n35746 ;
  assign n37735 = n37733 | n37734 ;
  assign n37736 = n37732 | n37735 ;
  assign n37737 = n7078 | n37732 ;
  assign n37738 = n37735 | n37737 ;
  assign n37739 = ( n36107 & n37736 ) | ( n36107 & n37738 ) | ( n37736 & n37738 ) ;
  assign n37740 = n37736 | n37738 ;
  assign n37741 = ( n36094 & n37739 ) | ( n36094 & n37740 ) | ( n37739 & n37740 ) ;
  assign n37742 = x8 & n37741 ;
  assign n37743 = x8 & ~n37741 ;
  assign n37744 = ( n37741 & ~n37742 ) | ( n37741 & n37743 ) | ( ~n37742 & n37743 ) ;
  assign n37745 = n37731 & ~n37744 ;
  assign n37746 = n37731 | n37744 ;
  assign n37747 = ( ~n37731 & n37745 ) | ( ~n37731 & n37746 ) | ( n37745 & n37746 ) ;
  assign n37748 = n37480 | n37483 ;
  assign n37749 = n37462 | n37480 ;
  assign n37750 = ( n37481 & n37748 ) | ( n37481 & n37749 ) | ( n37748 & n37749 ) ;
  assign n37751 = ~n37747 & n37750 ;
  assign n37752 = n37747 & ~n37750 ;
  assign n37753 = n37751 | n37752 ;
  assign n37754 = n37491 | n37497 ;
  assign n37755 = n37753 | n37754 ;
  assign n37756 = n37491 | n37499 ;
  assign n37757 = n37753 | n37756 ;
  assign n37758 = ( n36959 & n37755 ) | ( n36959 & n37757 ) | ( n37755 & n37757 ) ;
  assign n37759 = n37753 & n37754 ;
  assign n37760 = n37753 & n37756 ;
  assign n37761 = ( n36959 & n37759 ) | ( n36959 & n37760 ) | ( n37759 & n37760 ) ;
  assign n37762 = n37758 & ~n37761 ;
  assign n37763 = n37507 & n37762 ;
  assign n37764 = n37507 & ~n37763 ;
  assign n37765 = ( n37762 & ~n37763 ) | ( n37762 & n37764 ) | ( ~n37763 & n37764 ) ;
  assign n37766 = n26018 & n36083 ;
  assign n37767 = n7074 & n35746 ;
  assign n37768 = n37766 | n37767 ;
  assign n37769 = n7078 | n37768 ;
  assign n37770 = ( n36103 & n37768 ) | ( n36103 & n37769 ) | ( n37768 & n37769 ) ;
  assign n37771 = ( n36105 & n37768 ) | ( n36105 & n37769 ) | ( n37768 & n37769 ) ;
  assign n37772 = ( n32456 & n37770 ) | ( n32456 & n37771 ) | ( n37770 & n37771 ) ;
  assign n37773 = x8 & n37772 ;
  assign n37774 = x8 & ~n37772 ;
  assign n37775 = ( n37772 & ~n37773 ) | ( n37772 & n37774 ) | ( ~n37773 & n37774 ) ;
  assign n37776 = n37702 | n37720 ;
  assign n37777 = ( n37702 & n37705 ) | ( n37702 & n37776 ) | ( n37705 & n37776 ) ;
  assign n37778 = n37775 & n37777 ;
  assign n37779 = n37775 | n37777 ;
  assign n37780 = ~n37778 & n37779 ;
  assign n37781 = n37677 | n37696 ;
  assign n37782 = n365 | n19243 ;
  assign n37783 = n5132 | n37782 ;
  assign n37784 = n498 | n4246 ;
  assign n37785 = n14392 | n37784 ;
  assign n37786 = n37783 | n37785 ;
  assign n37787 = n46 | n1172 ;
  assign n37788 = n272 | n309 ;
  assign n37789 = n37787 | n37788 ;
  assign n37790 = n555 | n37789 ;
  assign n37791 = n145 & ~n264 ;
  assign n37792 = ~n137 & n37791 ;
  assign n37793 = ~n37790 & n37792 ;
  assign n37794 = ~n37786 & n37793 ;
  assign n37795 = ~n4030 & n37794 ;
  assign n37796 = n28108 | n29740 ;
  assign n37797 = n13843 | n37796 ;
  assign n37798 = n13831 | n37797 ;
  assign n37799 = n37795 & ~n37798 ;
  assign n37800 = n192 | n278 ;
  assign n37801 = n159 | n469 ;
  assign n37802 = n37800 | n37801 ;
  assign n37803 = n184 | n37802 ;
  assign n37804 = n318 | n542 ;
  assign n37805 = n222 | n313 ;
  assign n37806 = n37804 | n37805 ;
  assign n37807 = n206 | n435 ;
  assign n37808 = n104 | n37807 ;
  assign n37809 = n37806 | n37808 ;
  assign n37810 = n196 | n758 ;
  assign n37811 = n37809 | n37810 ;
  assign n37812 = n18129 | n37811 ;
  assign n37813 = n18484 | n37812 ;
  assign n37814 = n483 | n591 ;
  assign n37815 = n213 | n37814 ;
  assign n37816 = n37813 | n37815 ;
  assign n37817 = n37803 | n37816 ;
  assign n37818 = n37799 & ~n37817 ;
  assign n37819 = n37540 & n37818 ;
  assign n37820 = n37540 | n37818 ;
  assign n37821 = ~n37819 & n37820 ;
  assign n37822 = n37544 & ~n37546 ;
  assign n37823 = ( n37544 & ~n37558 ) | ( n37544 & n37822 ) | ( ~n37558 & n37822 ) ;
  assign n37824 = ~n37821 & n37823 ;
  assign n37825 = ~n37540 & n37821 ;
  assign n37826 = ~n37543 & n37825 ;
  assign n37827 = ( n37546 & n37821 ) | ( n37546 & n37826 ) | ( n37821 & n37826 ) ;
  assign n37828 = n37821 & n37826 ;
  assign n37829 = ( n37558 & n37827 ) | ( n37558 & n37828 ) | ( n37827 & n37828 ) ;
  assign n37830 = n37824 | n37829 ;
  assign n37831 = n1060 & ~n26270 ;
  assign n37832 = ~n26263 & n37831 ;
  assign n37833 = n1065 & ~n26526 ;
  assign n37834 = ~n26520 & n37833 ;
  assign n37835 = n37832 | n37834 ;
  assign n37836 = n1057 & ~n27133 ;
  assign n37837 = ~n27125 & n37836 ;
  assign n37838 = n37835 | n37837 ;
  assign n37839 = n1062 & n27699 ;
  assign n37840 = ( n1062 & ~n27696 ) | ( n1062 & n37839 ) | ( ~n27696 & n37839 ) ;
  assign n37841 = n37838 | n37840 ;
  assign n37842 = ~n37829 & n37841 ;
  assign n37843 = ~n37824 & n37842 ;
  assign n37844 = n37830 | n37843 ;
  assign n37845 = n37829 & n37841 ;
  assign n37846 = ( n37824 & n37841 ) | ( n37824 & n37845 ) | ( n37841 & n37845 ) ;
  assign n37847 = n37844 & ~n37846 ;
  assign n37848 = n37564 | n37584 ;
  assign n37849 = ( n37564 & n37565 ) | ( n37564 & n37848 ) | ( n37565 & n37848 ) ;
  assign n37850 = n37847 & ~n37849 ;
  assign n37851 = ~n37847 & n37849 ;
  assign n37852 = n37850 | n37851 ;
  assign n37853 = n1826 & ~n27371 ;
  assign n37854 = ~n27363 & n37853 ;
  assign n37855 = n1823 & ~n27606 ;
  assign n37856 = ~n27597 & n37855 ;
  assign n37857 = n37854 | n37856 ;
  assign n37858 = n1829 & ~n28503 ;
  assign n37859 = n28498 & n37858 ;
  assign n37860 = n37857 | n37859 ;
  assign n37861 = n1821 & n28794 ;
  assign n37862 = ( n1821 & n28783 ) | ( n1821 & n37861 ) | ( n28783 & n37861 ) ;
  assign n37863 = n37860 | n37862 ;
  assign n37864 = x29 | n37860 ;
  assign n37865 = n37862 | n37864 ;
  assign n37866 = ~x29 & n37864 ;
  assign n37867 = ( ~x29 & n37862 ) | ( ~x29 & n37866 ) | ( n37862 & n37866 ) ;
  assign n37868 = ( ~n37863 & n37865 ) | ( ~n37863 & n37867 ) | ( n37865 & n37867 ) ;
  assign n37869 = ~n37852 & n37868 ;
  assign n37870 = n37852 | n37869 ;
  assign n37871 = n2315 & n29620 ;
  assign n37872 = n2312 & n28492 ;
  assign n37873 = n2308 & ~n28714 ;
  assign n37874 = n37872 | n37873 ;
  assign n37875 = n37871 | n37874 ;
  assign n37876 = n2306 | n37871 ;
  assign n37877 = n37874 | n37876 ;
  assign n37878 = ( ~n29642 & n37875 ) | ( ~n29642 & n37877 ) | ( n37875 & n37877 ) ;
  assign n37879 = n37875 | n37877 ;
  assign n37880 = ( n29629 & n37878 ) | ( n29629 & n37879 ) | ( n37878 & n37879 ) ;
  assign n37881 = ~x26 & n37880 ;
  assign n37882 = x26 | n37880 ;
  assign n37883 = ( ~n37880 & n37881 ) | ( ~n37880 & n37882 ) | ( n37881 & n37882 ) ;
  assign n37884 = n37852 & n37868 ;
  assign n37885 = n37883 & n37884 ;
  assign n37886 = ( ~n37870 & n37883 ) | ( ~n37870 & n37885 ) | ( n37883 & n37885 ) ;
  assign n37887 = n37883 | n37884 ;
  assign n37888 = n37870 & ~n37887 ;
  assign n37889 = n37886 | n37888 ;
  assign n37890 = n37590 | n37606 ;
  assign n37891 = ( n37590 & n37592 ) | ( n37590 & n37890 ) | ( n37592 & n37890 ) ;
  assign n37892 = n37889 & ~n37891 ;
  assign n37893 = ~n37889 & n37891 ;
  assign n37894 = n37892 | n37893 ;
  assign n37895 = n2932 & ~n30186 ;
  assign n37896 = n2925 & ~n30199 ;
  assign n37897 = n2928 & n30212 ;
  assign n37898 = n37896 | n37897 ;
  assign n37899 = n37895 | n37898 ;
  assign n37900 = n2936 | n37895 ;
  assign n37901 = n37898 | n37900 ;
  assign n37902 = ( ~n30241 & n37899 ) | ( ~n30241 & n37901 ) | ( n37899 & n37901 ) ;
  assign n37903 = ~x23 & n37901 ;
  assign n37904 = ~x23 & n37899 ;
  assign n37905 = ( ~n30241 & n37903 ) | ( ~n30241 & n37904 ) | ( n37903 & n37904 ) ;
  assign n37906 = x23 | n37904 ;
  assign n37907 = x23 | n37903 ;
  assign n37908 = ( ~n30241 & n37906 ) | ( ~n30241 & n37907 ) | ( n37906 & n37907 ) ;
  assign n37909 = ( ~n37902 & n37905 ) | ( ~n37902 & n37908 ) | ( n37905 & n37908 ) ;
  assign n37910 = n37894 & n37909 ;
  assign n37911 = n37889 & ~n37909 ;
  assign n37912 = ( n37891 & n37909 ) | ( n37891 & ~n37911 ) | ( n37909 & ~n37911 ) ;
  assign n37913 = n37892 | n37912 ;
  assign n37914 = ~n37910 & n37913 ;
  assign n37915 = ( n37612 & n37613 ) | ( n37612 & n37628 ) | ( n37613 & n37628 ) ;
  assign n37916 = n37914 & ~n37915 ;
  assign n37917 = ~n37914 & n37915 ;
  assign n37918 = n37916 | n37917 ;
  assign n37919 = n3547 & n31295 ;
  assign n37920 = n3544 & ~n31309 ;
  assign n37921 = n3541 & ~n31323 ;
  assign n37922 = n37920 | n37921 ;
  assign n37923 = n37919 | n37922 ;
  assign n37924 = n3537 | n37919 ;
  assign n37925 = n37922 | n37924 ;
  assign n37926 = ( n31355 & n37923 ) | ( n31355 & n37925 ) | ( n37923 & n37925 ) ;
  assign n37927 = x20 & n37925 ;
  assign n37928 = x20 & n37923 ;
  assign n37929 = ( n31355 & n37927 ) | ( n31355 & n37928 ) | ( n37927 & n37928 ) ;
  assign n37930 = x20 & ~n37928 ;
  assign n37931 = x20 & ~n37927 ;
  assign n37932 = ( ~n31355 & n37930 ) | ( ~n31355 & n37931 ) | ( n37930 & n37931 ) ;
  assign n37933 = ( n37926 & ~n37929 ) | ( n37926 & n37932 ) | ( ~n37929 & n37932 ) ;
  assign n37934 = n37918 & n37933 ;
  assign n37935 = n37917 | n37933 ;
  assign n37936 = n37916 | n37935 ;
  assign n37937 = ~n37934 & n37936 ;
  assign n37938 = ( n37633 & n37634 ) | ( n37633 & n37650 ) | ( n37634 & n37650 ) ;
  assign n37939 = n37937 & ~n37938 ;
  assign n37940 = ~n37937 & n37938 ;
  assign n37941 = n37939 | n37940 ;
  assign n37942 = n4471 & ~n32442 ;
  assign n37943 = n4466 & n32306 ;
  assign n37944 = n4468 & n32293 ;
  assign n37945 = n37943 | n37944 ;
  assign n37946 = n37942 | n37945 ;
  assign n37947 = n4475 | n37942 ;
  assign n37948 = n37945 | n37947 ;
  assign n37949 = ( ~n32458 & n37946 ) | ( ~n32458 & n37948 ) | ( n37946 & n37948 ) ;
  assign n37950 = ~x17 & n37948 ;
  assign n37951 = ~x17 & n37946 ;
  assign n37952 = ( ~n32458 & n37950 ) | ( ~n32458 & n37951 ) | ( n37950 & n37951 ) ;
  assign n37953 = x17 | n37951 ;
  assign n37954 = x17 | n37950 ;
  assign n37955 = ( ~n32458 & n37953 ) | ( ~n32458 & n37954 ) | ( n37953 & n37954 ) ;
  assign n37956 = ( ~n37949 & n37952 ) | ( ~n37949 & n37955 ) | ( n37952 & n37955 ) ;
  assign n37957 = n37941 & n37956 ;
  assign n37958 = n37940 | n37956 ;
  assign n37959 = n37939 | n37958 ;
  assign n37960 = ~n37957 & n37959 ;
  assign n37961 = ( n37655 & n37656 ) | ( n37655 & n37675 ) | ( n37656 & n37675 ) ;
  assign n37962 = n37960 & ~n37961 ;
  assign n37963 = ~n37960 & n37961 ;
  assign n37964 = n5234 & n33526 ;
  assign n37965 = n5237 & n33436 ;
  assign n37966 = n5231 & ~n33423 ;
  assign n37967 = n37965 | n37966 ;
  assign n37968 = n37964 | n37967 ;
  assign n37969 = n5227 & n33545 ;
  assign n37970 = n5227 & ~n33548 ;
  assign n37971 = ( ~n32456 & n37969 ) | ( ~n32456 & n37970 ) | ( n37969 & n37970 ) ;
  assign n37972 = n37968 | n37971 ;
  assign n37973 = n5227 | n37968 ;
  assign n37974 = ( n33536 & n37972 ) | ( n33536 & n37973 ) | ( n37972 & n37973 ) ;
  assign n37975 = x14 | n37974 ;
  assign n37976 = ~x14 & n37974 ;
  assign n37977 = ( ~n37974 & n37975 ) | ( ~n37974 & n37976 ) | ( n37975 & n37976 ) ;
  assign n37978 = n37963 | n37977 ;
  assign n37979 = n37962 | n37978 ;
  assign n37980 = n37962 | n37963 ;
  assign n37981 = n37977 & n37980 ;
  assign n37982 = n37677 & n37981 ;
  assign n37983 = ( n37696 & n37981 ) | ( n37696 & n37982 ) | ( n37981 & n37982 ) ;
  assign n37984 = ( n37781 & ~n37979 ) | ( n37781 & n37983 ) | ( ~n37979 & n37983 ) ;
  assign n37985 = n37677 | n37981 ;
  assign n37986 = n37696 | n37985 ;
  assign n37987 = n37979 & ~n37986 ;
  assign n37988 = n37984 | n37987 ;
  assign n37989 = n6122 & ~n35371 ;
  assign n37990 = n6125 & n34656 ;
  assign n37991 = n6119 & n35021 ;
  assign n37992 = n37990 | n37991 ;
  assign n37993 = n37989 | n37992 ;
  assign n37994 = n6115 & ~n35392 ;
  assign n37995 = n6115 & ~n35395 ;
  assign n37996 = ( ~n32456 & n37994 ) | ( ~n32456 & n37995 ) | ( n37994 & n37995 ) ;
  assign n37997 = n37993 | n37996 ;
  assign n37998 = n6115 | n37993 ;
  assign n37999 = ( n35381 & n37997 ) | ( n35381 & n37998 ) | ( n37997 & n37998 ) ;
  assign n38000 = x11 | n37999 ;
  assign n38001 = ~x11 & n37999 ;
  assign n38002 = ( ~n37999 & n38000 ) | ( ~n37999 & n38001 ) | ( n38000 & n38001 ) ;
  assign n38003 = n37988 | n38002 ;
  assign n38004 = n37988 & ~n38002 ;
  assign n38005 = ( ~n37988 & n38003 ) | ( ~n37988 & n38004 ) | ( n38003 & n38004 ) ;
  assign n38006 = n37780 & ~n38005 ;
  assign n38007 = n37780 & ~n38006 ;
  assign n38008 = n37780 | n38005 ;
  assign n38009 = ~n38007 & n38008 ;
  assign n38010 = n37727 | n37744 ;
  assign n38011 = ( n37727 & n37731 ) | ( n37727 & n38010 ) | ( n37731 & n38010 ) ;
  assign n38012 = n38009 & ~n38011 ;
  assign n38013 = ~n38009 & n38011 ;
  assign n38014 = n38012 | n38013 ;
  assign n38015 = n37747 & ~n38014 ;
  assign n38016 = n37750 & n38015 ;
  assign n38017 = ( n37753 & ~n38014 ) | ( n37753 & n38016 ) | ( ~n38014 & n38016 ) ;
  assign n38018 = ( n37754 & n38016 ) | ( n37754 & n38017 ) | ( n38016 & n38017 ) ;
  assign n38019 = ( n37756 & n38016 ) | ( n37756 & n38017 ) | ( n38016 & n38017 ) ;
  assign n38020 = ( n36959 & n38018 ) | ( n36959 & n38019 ) | ( n38018 & n38019 ) ;
  assign n38021 = ( n37747 & n37750 ) | ( n37747 & n37754 ) | ( n37750 & n37754 ) ;
  assign n38022 = n38014 & ~n38021 ;
  assign n38023 = ( n37747 & n37750 ) | ( n37747 & n37756 ) | ( n37750 & n37756 ) ;
  assign n38024 = n38014 & ~n38023 ;
  assign n38025 = ( ~n36959 & n38022 ) | ( ~n36959 & n38024 ) | ( n38022 & n38024 ) ;
  assign n38026 = n38020 | n38025 ;
  assign n38027 = ~n37763 & n38026 ;
  assign n38028 = n37762 & ~n38026 ;
  assign n38029 = n37506 & n38028 ;
  assign n38030 = n36963 & n38029 ;
  assign n38031 = n38027 | n38030 ;
  assign n38032 = ~n405 & n911 ;
  assign n38033 = n3282 | n6988 ;
  assign n38034 = n224 | n3411 ;
  assign n38035 = n38033 | n38034 ;
  assign n38036 = n3495 | n29288 ;
  assign n38037 = n38035 | n38036 ;
  assign n38038 = n2075 | n38037 ;
  assign n38039 = n2040 | n38038 ;
  assign n38040 = n38032 & ~n38039 ;
  assign n38041 = n271 | n6080 ;
  assign n38042 = n6070 | n38041 ;
  assign n38043 = n54 | n796 ;
  assign n38044 = n59 | n178 ;
  assign n38045 = n38043 | n38044 ;
  assign n38046 = n38042 | n38045 ;
  assign n38047 = n38040 & ~n38046 ;
  assign n38048 = ~n37540 & n38047 ;
  assign n38049 = n37540 & ~n38047 ;
  assign n38050 = n38048 | n38049 ;
  assign n38051 = n26303 & n36083 ;
  assign n38052 = ~x8 & n26303 ;
  assign n38053 = n36083 & n38052 ;
  assign n38054 = x8 | n38052 ;
  assign n38055 = ( x8 & n36083 ) | ( x8 & n38054 ) | ( n36083 & n38054 ) ;
  assign n38056 = ( ~n38051 & n38053 ) | ( ~n38051 & n38055 ) | ( n38053 & n38055 ) ;
  assign n38057 = n38050 | n38056 ;
  assign n38058 = n38050 & n38056 ;
  assign n38059 = n38057 & ~n38058 ;
  assign n38060 = ~n37820 & n38059 ;
  assign n38061 = ( n37829 & n38059 ) | ( n37829 & n38060 ) | ( n38059 & n38060 ) ;
  assign n38062 = n37820 & ~n38059 ;
  assign n38063 = ~n37829 & n38062 ;
  assign n38064 = n38061 | n38063 ;
  assign n38065 = n1060 & ~n26526 ;
  assign n38066 = ~n26520 & n38065 ;
  assign n38067 = n1065 & ~n27133 ;
  assign n38068 = ~n27125 & n38067 ;
  assign n38069 = n38066 | n38068 ;
  assign n38070 = n1057 & ~n27371 ;
  assign n38071 = ~n27363 & n38070 ;
  assign n38072 = n38069 | n38071 ;
  assign n38073 = n1062 | n38071 ;
  assign n38074 = n38069 | n38073 ;
  assign n38075 = ( ~n27654 & n38072 ) | ( ~n27654 & n38074 ) | ( n38072 & n38074 ) ;
  assign n38076 = n38064 & n38075 ;
  assign n38077 = n38064 | n38075 ;
  assign n38078 = ~n38076 & n38077 ;
  assign n38079 = n1829 & n28492 ;
  assign n38080 = n1826 & ~n27606 ;
  assign n38081 = ~n27597 & n38080 ;
  assign n38082 = n1823 & ~n28503 ;
  assign n38083 = n28498 & n38082 ;
  assign n38084 = n38081 | n38083 ;
  assign n38085 = n38079 | n38084 ;
  assign n38086 = n1821 | n38085 ;
  assign n38087 = ( ~n28749 & n38085 ) | ( ~n28749 & n38086 ) | ( n38085 & n38086 ) ;
  assign n38088 = ~x29 & n38086 ;
  assign n38089 = ~x29 & n38085 ;
  assign n38090 = ( ~n28749 & n38088 ) | ( ~n28749 & n38089 ) | ( n38088 & n38089 ) ;
  assign n38091 = x29 | n38088 ;
  assign n38092 = x29 | n38089 ;
  assign n38093 = ( ~n28749 & n38091 ) | ( ~n28749 & n38092 ) | ( n38091 & n38092 ) ;
  assign n38094 = ( ~n38087 & n38090 ) | ( ~n38087 & n38093 ) | ( n38090 & n38093 ) ;
  assign n38095 = ~n38078 & n38094 ;
  assign n38096 = n38078 & ~n38094 ;
  assign n38097 = n38095 | n38096 ;
  assign n38098 = n37843 | n37851 ;
  assign n38099 = n38097 & ~n38098 ;
  assign n38100 = ~n38097 & n38098 ;
  assign n38101 = n38099 | n38100 ;
  assign n38102 = n2315 & ~n30199 ;
  assign n38103 = n2312 & ~n28714 ;
  assign n38104 = n2308 & n29620 ;
  assign n38105 = n38103 | n38104 ;
  assign n38106 = n38102 | n38105 ;
  assign n38107 = n2306 | n38102 ;
  assign n38108 = n38105 | n38107 ;
  assign n38109 = ( ~n30299 & n38106 ) | ( ~n30299 & n38108 ) | ( n38106 & n38108 ) ;
  assign n38110 = ~x26 & n38108 ;
  assign n38111 = ~x26 & n38106 ;
  assign n38112 = ( ~n30299 & n38110 ) | ( ~n30299 & n38111 ) | ( n38110 & n38111 ) ;
  assign n38113 = x26 | n38111 ;
  assign n38114 = x26 | n38110 ;
  assign n38115 = ( ~n30299 & n38113 ) | ( ~n30299 & n38114 ) | ( n38113 & n38114 ) ;
  assign n38116 = ( ~n38109 & n38112 ) | ( ~n38109 & n38115 ) | ( n38112 & n38115 ) ;
  assign n38117 = ~n38101 & n38116 ;
  assign n38118 = n38101 | n38117 ;
  assign n38119 = n38101 & n38116 ;
  assign n38120 = n38118 & ~n38119 ;
  assign n38121 = n37869 | n37886 ;
  assign n38122 = n38120 & ~n38121 ;
  assign n38123 = ~n38120 & n38121 ;
  assign n38124 = n38122 | n38123 ;
  assign n38125 = n2932 & ~n31309 ;
  assign n38126 = n2925 & n30212 ;
  assign n38127 = n2928 & ~n30186 ;
  assign n38128 = n38126 | n38127 ;
  assign n38129 = n38125 | n38128 ;
  assign n38130 = n2936 | n38125 ;
  assign n38131 = n38128 | n38130 ;
  assign n38132 = ( n31404 & n38129 ) | ( n31404 & n38131 ) | ( n38129 & n38131 ) ;
  assign n38133 = x23 & n38131 ;
  assign n38134 = x23 & n38129 ;
  assign n38135 = ( n31404 & n38133 ) | ( n31404 & n38134 ) | ( n38133 & n38134 ) ;
  assign n38136 = x23 & ~n38134 ;
  assign n38137 = x23 & ~n38133 ;
  assign n38138 = ( ~n31404 & n38136 ) | ( ~n31404 & n38137 ) | ( n38136 & n38137 ) ;
  assign n38139 = ( n38132 & ~n38135 ) | ( n38132 & n38138 ) | ( ~n38135 & n38138 ) ;
  assign n38140 = ~n38124 & n38139 ;
  assign n38141 = n38124 | n38140 ;
  assign n38143 = n37893 | n37909 ;
  assign n38144 = ( n37893 & ~n37894 ) | ( n37893 & n38143 ) | ( ~n37894 & n38143 ) ;
  assign n38142 = n38124 & n38139 ;
  assign n38145 = n38142 & n38144 ;
  assign n38146 = ( ~n38141 & n38144 ) | ( ~n38141 & n38145 ) | ( n38144 & n38145 ) ;
  assign n38147 = n38142 | n38144 ;
  assign n38148 = n38141 & ~n38147 ;
  assign n38149 = n38146 | n38148 ;
  assign n38150 = n3547 & n32306 ;
  assign n38151 = n3544 & ~n31323 ;
  assign n38152 = n3541 & n31295 ;
  assign n38153 = n38151 | n38152 ;
  assign n38154 = n38150 | n38153 ;
  assign n38155 = n3537 | n38150 ;
  assign n38156 = n38153 | n38155 ;
  assign n38157 = ( ~n32525 & n38154 ) | ( ~n32525 & n38156 ) | ( n38154 & n38156 ) ;
  assign n38158 = ~x20 & n38156 ;
  assign n38159 = ~x20 & n38154 ;
  assign n38160 = ( ~n32525 & n38158 ) | ( ~n32525 & n38159 ) | ( n38158 & n38159 ) ;
  assign n38161 = x20 | n38159 ;
  assign n38162 = x20 | n38158 ;
  assign n38163 = ( ~n32525 & n38161 ) | ( ~n32525 & n38162 ) | ( n38161 & n38162 ) ;
  assign n38164 = ( ~n38157 & n38160 ) | ( ~n38157 & n38163 ) | ( n38160 & n38163 ) ;
  assign n38165 = ~n38149 & n38164 ;
  assign n38166 = n38149 | n38165 ;
  assign n38167 = n38149 & n38164 ;
  assign n38168 = ( n37917 & ~n37918 ) | ( n37917 & n37935 ) | ( ~n37918 & n37935 ) ;
  assign n38169 = n38167 | n38168 ;
  assign n38170 = n38166 & ~n38169 ;
  assign n38171 = n38167 & n38168 ;
  assign n38172 = ( ~n38166 & n38168 ) | ( ~n38166 & n38171 ) | ( n38168 & n38171 ) ;
  assign n38173 = n38170 | n38172 ;
  assign n38188 = ( n37940 & ~n37941 ) | ( n37940 & n37958 ) | ( ~n37941 & n37958 ) ;
  assign n38174 = n4471 & n33436 ;
  assign n38175 = n4466 & n32293 ;
  assign n38176 = n4468 & ~n32442 ;
  assign n38177 = n38175 | n38176 ;
  assign n38178 = n38174 | n38177 ;
  assign n38179 = n4475 & ~n33441 ;
  assign n38180 = ~n32456 & n38179 ;
  assign n38181 = ( n4475 & n34271 ) | ( n4475 & n38180 ) | ( n34271 & n38180 ) ;
  assign n38182 = n38178 | n38181 ;
  assign n38183 = x17 | n38178 ;
  assign n38184 = n38181 | n38183 ;
  assign n38185 = ~x17 & n38183 ;
  assign n38186 = ( ~x17 & n38181 ) | ( ~x17 & n38185 ) | ( n38181 & n38185 ) ;
  assign n38187 = ( ~n38182 & n38184 ) | ( ~n38182 & n38186 ) | ( n38184 & n38186 ) ;
  assign n38189 = n38187 & n38188 ;
  assign n38190 = n38188 & ~n38189 ;
  assign n38191 = ~n38173 & n38187 ;
  assign n38192 = ~n38188 & n38191 ;
  assign n38193 = ( ~n38173 & n38190 ) | ( ~n38173 & n38192 ) | ( n38190 & n38192 ) ;
  assign n38194 = n38173 & ~n38187 ;
  assign n38195 = ( n38173 & n38188 ) | ( n38173 & n38194 ) | ( n38188 & n38194 ) ;
  assign n38196 = ~n38190 & n38195 ;
  assign n38197 = n38193 | n38196 ;
  assign n38198 = n5234 & n34656 ;
  assign n38199 = n5237 & ~n33423 ;
  assign n38200 = n5231 & n33526 ;
  assign n38201 = n38199 | n38200 ;
  assign n38202 = n38198 | n38201 ;
  assign n38203 = n5227 | n38198 ;
  assign n38204 = n38201 | n38203 ;
  assign n38205 = ( n34667 & n38202 ) | ( n34667 & n38204 ) | ( n38202 & n38204 ) ;
  assign n38206 = x14 & n38204 ;
  assign n38207 = x14 & n38202 ;
  assign n38208 = ( n34667 & n38206 ) | ( n34667 & n38207 ) | ( n38206 & n38207 ) ;
  assign n38209 = x14 & ~n38207 ;
  assign n38210 = x14 & ~n38206 ;
  assign n38211 = ( ~n34667 & n38209 ) | ( ~n34667 & n38210 ) | ( n38209 & n38210 ) ;
  assign n38212 = ( n38205 & ~n38208 ) | ( n38205 & n38211 ) | ( ~n38208 & n38211 ) ;
  assign n38213 = ~n38197 & n38212 ;
  assign n38214 = n38197 | n38213 ;
  assign n38216 = ( n37963 & n37978 ) | ( n37963 & ~n37980 ) | ( n37978 & ~n37980 ) ;
  assign n38215 = n38197 & n38212 ;
  assign n38217 = n38215 & n38216 ;
  assign n38218 = ( ~n38214 & n38216 ) | ( ~n38214 & n38217 ) | ( n38216 & n38217 ) ;
  assign n38219 = n38215 | n38216 ;
  assign n38220 = n38214 & ~n38219 ;
  assign n38221 = n38218 | n38220 ;
  assign n38237 = n37984 | n38002 ;
  assign n38238 = ( n37984 & ~n37988 ) | ( n37984 & n38237 ) | ( ~n37988 & n38237 ) ;
  assign n38222 = n6122 & n35746 ;
  assign n38223 = n6125 & n35021 ;
  assign n38224 = n6119 & ~n35371 ;
  assign n38225 = n38223 | n38224 ;
  assign n38226 = n38222 | n38225 ;
  assign n38227 = n6115 | n38222 ;
  assign n38228 = n38225 | n38227 ;
  assign n38229 = ( ~n35759 & n38226 ) | ( ~n35759 & n38228 ) | ( n38226 & n38228 ) ;
  assign n38230 = ~x11 & n38228 ;
  assign n38231 = ~x11 & n38226 ;
  assign n38232 = ( ~n35759 & n38230 ) | ( ~n35759 & n38231 ) | ( n38230 & n38231 ) ;
  assign n38233 = x11 | n38231 ;
  assign n38234 = x11 | n38230 ;
  assign n38235 = ( ~n35759 & n38233 ) | ( ~n35759 & n38234 ) | ( n38233 & n38234 ) ;
  assign n38236 = ( ~n38229 & n38232 ) | ( ~n38229 & n38235 ) | ( n38232 & n38235 ) ;
  assign n38239 = n38236 & n38238 ;
  assign n38240 = n38238 & ~n38239 ;
  assign n38241 = ~n38221 & n38236 ;
  assign n38242 = ~n38238 & n38241 ;
  assign n38243 = ( ~n38221 & n38240 ) | ( ~n38221 & n38242 ) | ( n38240 & n38242 ) ;
  assign n38244 = n38221 & ~n38236 ;
  assign n38245 = ( n38221 & n38238 ) | ( n38221 & n38244 ) | ( n38238 & n38244 ) ;
  assign n38246 = ~n38240 & n38245 ;
  assign n38247 = n38243 | n38246 ;
  assign n38248 = ~n37778 & n38005 ;
  assign n38249 = ( n37778 & n37780 ) | ( n37778 & ~n38248 ) | ( n37780 & ~n38248 ) ;
  assign n38250 = ~n38247 & n38249 ;
  assign n38251 = n38247 & ~n38249 ;
  assign n38252 = n38250 | n38251 ;
  assign n38253 = n38013 | n38016 ;
  assign n38254 = ~n38013 & n38014 ;
  assign n38255 = ( n37753 & n38253 ) | ( n37753 & ~n38254 ) | ( n38253 & ~n38254 ) ;
  assign n38256 = ~n38252 & n38255 ;
  assign n38257 = n38013 & ~n38252 ;
  assign n38258 = ( n38016 & ~n38252 ) | ( n38016 & n38257 ) | ( ~n38252 & n38257 ) ;
  assign n38259 = ( n37754 & n38256 ) | ( n37754 & n38258 ) | ( n38256 & n38258 ) ;
  assign n38260 = ( n37756 & n38256 ) | ( n37756 & n38258 ) | ( n38256 & n38258 ) ;
  assign n38261 = ( n36959 & n38259 ) | ( n36959 & n38260 ) | ( n38259 & n38260 ) ;
  assign n38262 = ( n37754 & n38253 ) | ( n37754 & n38255 ) | ( n38253 & n38255 ) ;
  assign n38263 = n38252 & ~n38262 ;
  assign n38264 = ( n37756 & n38253 ) | ( n37756 & n38255 ) | ( n38253 & n38255 ) ;
  assign n38265 = n38252 & ~n38264 ;
  assign n38266 = ( ~n36959 & n38263 ) | ( ~n36959 & n38265 ) | ( n38263 & n38265 ) ;
  assign n38267 = n38261 | n38266 ;
  assign n38268 = ~n38030 & n38267 ;
  assign n38269 = n38030 & ~n38267 ;
  assign n38270 = n38268 | n38269 ;
  assign n38271 = n38213 | n38218 ;
  assign n38428 = n38189 | n38192 ;
  assign n38429 = n38173 & ~n38189 ;
  assign n38430 = ( n38190 & n38428 ) | ( n38190 & ~n38429 ) | ( n38428 & ~n38429 ) ;
  assign n38272 = n1060 & ~n27133 ;
  assign n38273 = ~n27125 & n38272 ;
  assign n38274 = n1065 & ~n27371 ;
  assign n38275 = ~n27363 & n38274 ;
  assign n38276 = n38273 | n38275 ;
  assign n38277 = n1057 & ~n27606 ;
  assign n38278 = ~n27597 & n38277 ;
  assign n38279 = n38276 | n38278 ;
  assign n38280 = n1062 & n27630 ;
  assign n38281 = ~n27625 & n38280 ;
  assign n38282 = ( n1062 & ~n27634 ) | ( n1062 & n38281 ) | ( ~n27634 & n38281 ) ;
  assign n38283 = n38279 | n38282 ;
  assign n38284 = n27386 | n27387 ;
  assign n38285 = n1114 | n3351 ;
  assign n38286 = n2743 | n38285 ;
  assign n38287 = n17712 | n38286 ;
  assign n38288 = n38284 | n38287 ;
  assign n38289 = n517 | n10379 ;
  assign n38290 = n15256 | n38289 ;
  assign n38291 = n38288 | n38290 ;
  assign n38292 = ( ~n2833 & n6938 ) | ( ~n2833 & n38291 ) | ( n6938 & n38291 ) ;
  assign n38293 = n6938 & n38291 ;
  assign n38294 = ( n2827 & n38292 ) | ( n2827 & n38293 ) | ( n38292 & n38293 ) ;
  assign n38295 = n2834 & ~n38294 ;
  assign n38296 = n112 | n283 ;
  assign n38297 = n632 | n38296 ;
  assign n38298 = n418 | n444 ;
  assign n38299 = n356 | n38298 ;
  assign n38300 = n38297 | n38299 ;
  assign n38301 = n226 | n250 ;
  assign n38302 = n758 | n38301 ;
  assign n38303 = n38300 | n38302 ;
  assign n38304 = n38295 & ~n38303 ;
  assign n38305 = ( n38049 & ~n38050 ) | ( n38049 & n38304 ) | ( ~n38050 & n38304 ) ;
  assign n38306 = n38049 & n38304 ;
  assign n38307 = ( ~n38056 & n38305 ) | ( ~n38056 & n38306 ) | ( n38305 & n38306 ) ;
  assign n38308 = ~n38049 & n38050 ;
  assign n38309 = ~n38304 & n38308 ;
  assign n38310 = n38049 | n38304 ;
  assign n38311 = ( n38056 & n38309 ) | ( n38056 & ~n38310 ) | ( n38309 & ~n38310 ) ;
  assign n38312 = n38307 | n38311 ;
  assign n38313 = n38279 | n38312 ;
  assign n38314 = n38282 | n38313 ;
  assign n38315 = ~n38312 & n38313 ;
  assign n38316 = ( n38282 & ~n38312 ) | ( n38282 & n38315 ) | ( ~n38312 & n38315 ) ;
  assign n38317 = ( ~n38283 & n38314 ) | ( ~n38283 & n38316 ) | ( n38314 & n38316 ) ;
  assign n38318 = n38061 | n38075 ;
  assign n38319 = ( n38061 & ~n38064 ) | ( n38061 & n38318 ) | ( ~n38064 & n38318 ) ;
  assign n38320 = n38317 & ~n38319 ;
  assign n38321 = ~n38317 & n38319 ;
  assign n38322 = n38320 | n38321 ;
  assign n38323 = n1823 & n28492 ;
  assign n38324 = n1826 & ~n28503 ;
  assign n38325 = n28498 & n38324 ;
  assign n38326 = n38323 | n38325 ;
  assign n38327 = n1829 & ~n28714 ;
  assign n38328 = n1821 | n38327 ;
  assign n38329 = n38326 | n38328 ;
  assign n38330 = n38326 | n38327 ;
  assign n38331 = n28731 & ~n38330 ;
  assign n38332 = ( n28518 & ~n38330 ) | ( n28518 & n38331 ) | ( ~n38330 & n38331 ) ;
  assign n38333 = n38329 & ~n38332 ;
  assign n38334 = ( n28720 & n38329 ) | ( n28720 & n38333 ) | ( n38329 & n38333 ) ;
  assign n38335 = x29 & n38334 ;
  assign n38336 = x29 & ~n38334 ;
  assign n38337 = ( n38334 & ~n38335 ) | ( n38334 & n38336 ) | ( ~n38335 & n38336 ) ;
  assign n38338 = ~n38322 & n38337 ;
  assign n38339 = n38322 & ~n38337 ;
  assign n38340 = n38338 | n38339 ;
  assign n38341 = n38095 | n38100 ;
  assign n38342 = ~n38340 & n38341 ;
  assign n38343 = n38340 & ~n38341 ;
  assign n38344 = n38342 | n38343 ;
  assign n38345 = n2315 & n30212 ;
  assign n38346 = n2312 & n29620 ;
  assign n38347 = n2308 & ~n30199 ;
  assign n38348 = n38346 | n38347 ;
  assign n38349 = n38345 | n38348 ;
  assign n38350 = n2306 & ~n30266 ;
  assign n38351 = ( n2306 & n30276 ) | ( n2306 & n38350 ) | ( n30276 & n38350 ) ;
  assign n38352 = n38349 | n38351 ;
  assign n38353 = x26 | n38349 ;
  assign n38354 = n38351 | n38353 ;
  assign n38355 = ~x26 & n38353 ;
  assign n38356 = ( ~x26 & n38351 ) | ( ~x26 & n38355 ) | ( n38351 & n38355 ) ;
  assign n38357 = ( ~n38352 & n38354 ) | ( ~n38352 & n38356 ) | ( n38354 & n38356 ) ;
  assign n38358 = n38344 | n38357 ;
  assign n38359 = n38344 & ~n38357 ;
  assign n38360 = ( ~n38344 & n38358 ) | ( ~n38344 & n38359 ) | ( n38358 & n38359 ) ;
  assign n38361 = n38117 | n38121 ;
  assign n38362 = ( n38117 & ~n38120 ) | ( n38117 & n38361 ) | ( ~n38120 & n38361 ) ;
  assign n38363 = n38360 & ~n38362 ;
  assign n38364 = ~n38360 & n38362 ;
  assign n38365 = n38363 | n38364 ;
  assign n38366 = n2932 & ~n31323 ;
  assign n38367 = n2925 & ~n30186 ;
  assign n38368 = n2928 & ~n31309 ;
  assign n38369 = n38367 | n38368 ;
  assign n38370 = n38366 | n38369 ;
  assign n38371 = n2936 & n31384 ;
  assign n38372 = n2936 & n31386 ;
  assign n38373 = ( ~n30232 & n38371 ) | ( ~n30232 & n38372 ) | ( n38371 & n38372 ) ;
  assign n38374 = n38370 | n38373 ;
  assign n38375 = n2936 | n38370 ;
  assign n38376 = ( ~n31376 & n38374 ) | ( ~n31376 & n38375 ) | ( n38374 & n38375 ) ;
  assign n38377 = x23 | n38376 ;
  assign n38378 = ~x23 & n38376 ;
  assign n38379 = ( ~n38376 & n38377 ) | ( ~n38376 & n38378 ) | ( n38377 & n38378 ) ;
  assign n38380 = n38365 & n38379 ;
  assign n38381 = n38364 | n38379 ;
  assign n38382 = n38363 | n38381 ;
  assign n38383 = ~n38380 & n38382 ;
  assign n38384 = n38140 | n38146 ;
  assign n38385 = n38383 & ~n38384 ;
  assign n38386 = ~n38383 & n38384 ;
  assign n38387 = n38385 | n38386 ;
  assign n38388 = n3547 & n32293 ;
  assign n38389 = n3544 & n31295 ;
  assign n38390 = n3541 & n32306 ;
  assign n38391 = n38389 | n38390 ;
  assign n38392 = n38388 | n38391 ;
  assign n38393 = n3537 & n32497 ;
  assign n38394 = ( n3537 & n32494 ) | ( n3537 & n38393 ) | ( n32494 & n38393 ) ;
  assign n38395 = n38392 | n38394 ;
  assign n38396 = x20 | n38392 ;
  assign n38397 = n38394 | n38396 ;
  assign n38398 = ~x20 & n38396 ;
  assign n38399 = ( ~x20 & n38394 ) | ( ~x20 & n38398 ) | ( n38394 & n38398 ) ;
  assign n38400 = ( ~n38395 & n38397 ) | ( ~n38395 & n38399 ) | ( n38397 & n38399 ) ;
  assign n38401 = n38387 & n38400 ;
  assign n38402 = n38383 & ~n38400 ;
  assign n38403 = ( n38384 & n38400 ) | ( n38384 & ~n38402 ) | ( n38400 & ~n38402 ) ;
  assign n38404 = n38385 | n38403 ;
  assign n38405 = ~n38401 & n38404 ;
  assign n38406 = n38165 | n38172 ;
  assign n38407 = n38405 & ~n38406 ;
  assign n38408 = ~n38405 & n38406 ;
  assign n38409 = n38407 | n38408 ;
  assign n38410 = n4471 & ~n33423 ;
  assign n38411 = n4466 & ~n32442 ;
  assign n38412 = n4468 & n33436 ;
  assign n38413 = n38411 | n38412 ;
  assign n38414 = n38410 | n38413 ;
  assign n38415 = n4475 & n33575 ;
  assign n38416 = n4475 & ~n33577 ;
  assign n38417 = ( ~n32456 & n38415 ) | ( ~n32456 & n38416 ) | ( n38415 & n38416 ) ;
  assign n38418 = n38414 | n38417 ;
  assign n38419 = n4475 | n38414 ;
  assign n38420 = ( n33567 & n38418 ) | ( n33567 & n38419 ) | ( n38418 & n38419 ) ;
  assign n38421 = x17 | n38420 ;
  assign n38422 = ~x17 & n38420 ;
  assign n38423 = ( ~n38420 & n38421 ) | ( ~n38420 & n38422 ) | ( n38421 & n38422 ) ;
  assign n38424 = n38409 & n38423 ;
  assign n38425 = n38408 | n38423 ;
  assign n38426 = n38407 | n38425 ;
  assign n38427 = ~n38424 & n38426 ;
  assign n38431 = ~n38427 & n38430 ;
  assign n38432 = n38430 & ~n38431 ;
  assign n38433 = n5234 & n35021 ;
  assign n38434 = n5237 & n33526 ;
  assign n38435 = n5231 & n34656 ;
  assign n38436 = n38434 | n38435 ;
  assign n38437 = n38433 | n38436 ;
  assign n38438 = n5227 | n38433 ;
  assign n38439 = n38436 | n38438 ;
  assign n38440 = ( n35033 & n38437 ) | ( n35033 & n38439 ) | ( n38437 & n38439 ) ;
  assign n38441 = x14 & n38439 ;
  assign n38442 = x14 & n38437 ;
  assign n38443 = ( n35033 & n38441 ) | ( n35033 & n38442 ) | ( n38441 & n38442 ) ;
  assign n38444 = x14 & ~n38442 ;
  assign n38445 = x14 & ~n38441 ;
  assign n38446 = ( ~n35033 & n38444 ) | ( ~n35033 & n38445 ) | ( n38444 & n38445 ) ;
  assign n38447 = ( n38440 & ~n38443 ) | ( n38440 & n38446 ) | ( ~n38443 & n38446 ) ;
  assign n38448 = n38427 | n38430 ;
  assign n38449 = n38447 & ~n38448 ;
  assign n38450 = ( n38432 & n38447 ) | ( n38432 & n38449 ) | ( n38447 & n38449 ) ;
  assign n38451 = ~n38447 & n38448 ;
  assign n38452 = ~n38432 & n38451 ;
  assign n38453 = n38450 | n38452 ;
  assign n38454 = ~n38271 & n38453 ;
  assign n38455 = n38271 & ~n38453 ;
  assign n38456 = n38454 | n38455 ;
  assign n38457 = n6122 & n36083 ;
  assign n38458 = n6125 & ~n35371 ;
  assign n38459 = n6119 & n35746 ;
  assign n38460 = n38458 | n38459 ;
  assign n38461 = n38457 | n38460 ;
  assign n38462 = n6115 | n38457 ;
  assign n38463 = n38460 | n38462 ;
  assign n38464 = ( n36107 & n38461 ) | ( n36107 & n38463 ) | ( n38461 & n38463 ) ;
  assign n38465 = n38461 | n38463 ;
  assign n38466 = ( n36094 & n38464 ) | ( n36094 & n38465 ) | ( n38464 & n38465 ) ;
  assign n38467 = x11 & n38466 ;
  assign n38468 = x11 & ~n38466 ;
  assign n38469 = ( n38466 & ~n38467 ) | ( n38466 & n38468 ) | ( ~n38467 & n38468 ) ;
  assign n38470 = n38456 & n38469 ;
  assign n38471 = n38453 & ~n38469 ;
  assign n38472 = ( n38271 & n38469 ) | ( n38271 & ~n38471 ) | ( n38469 & ~n38471 ) ;
  assign n38473 = n38454 | n38472 ;
  assign n38474 = ~n38470 & n38473 ;
  assign n38475 = n38239 | n38242 ;
  assign n38476 = n38221 & ~n38239 ;
  assign n38477 = ( n38240 & n38475 ) | ( n38240 & ~n38476 ) | ( n38475 & ~n38476 ) ;
  assign n38478 = ~n38474 & n38477 ;
  assign n38479 = n38474 | n38478 ;
  assign n38480 = n38474 & n38477 ;
  assign n38481 = n38479 & ~n38480 ;
  assign n38482 = ~n38250 & n38252 ;
  assign n38483 = n38481 | n38482 ;
  assign n38484 = n38250 & ~n38481 ;
  assign n38485 = ( n38255 & ~n38483 ) | ( n38255 & n38484 ) | ( ~n38483 & n38484 ) ;
  assign n38486 = n38250 | n38257 ;
  assign n38487 = ~n38481 & n38486 ;
  assign n38488 = ( n38016 & ~n38483 ) | ( n38016 & n38487 ) | ( ~n38483 & n38487 ) ;
  assign n38489 = ( n37754 & n38485 ) | ( n37754 & n38488 ) | ( n38485 & n38488 ) ;
  assign n38490 = ( n37756 & n38485 ) | ( n37756 & n38488 ) | ( n38485 & n38488 ) ;
  assign n38491 = ( n36959 & n38489 ) | ( n36959 & n38490 ) | ( n38489 & n38490 ) ;
  assign n38492 = ( n38250 & n38255 ) | ( n38250 & ~n38482 ) | ( n38255 & ~n38482 ) ;
  assign n38493 = ( n38016 & ~n38482 ) | ( n38016 & n38486 ) | ( ~n38482 & n38486 ) ;
  assign n38494 = ( n37754 & n38492 ) | ( n37754 & n38493 ) | ( n38492 & n38493 ) ;
  assign n38495 = n38481 & ~n38494 ;
  assign n38496 = ( n37756 & n38492 ) | ( n37756 & n38493 ) | ( n38492 & n38493 ) ;
  assign n38497 = n38481 & ~n38496 ;
  assign n38498 = ( ~n36959 & n38495 ) | ( ~n36959 & n38497 ) | ( n38495 & n38497 ) ;
  assign n38499 = n38491 | n38498 ;
  assign n38500 = n38269 & n38499 ;
  assign n38501 = n38269 | n38499 ;
  assign n38502 = ~n38500 & n38501 ;
  assign n38503 = n27136 & n36083 ;
  assign n38504 = n6125 & n35746 ;
  assign n38505 = n38503 | n38504 ;
  assign n38506 = n6115 | n38505 ;
  assign n38507 = ( n36103 & n38505 ) | ( n36103 & n38506 ) | ( n38505 & n38506 ) ;
  assign n38508 = ( n36105 & n38505 ) | ( n36105 & n38506 ) | ( n38505 & n38506 ) ;
  assign n38509 = ( n32456 & n38507 ) | ( n32456 & n38508 ) | ( n38507 & n38508 ) ;
  assign n38510 = x11 & n38509 ;
  assign n38511 = x11 & ~n38509 ;
  assign n38512 = ( n38509 & ~n38510 ) | ( n38509 & n38511 ) | ( ~n38510 & n38511 ) ;
  assign n38513 = n38431 & n38512 ;
  assign n38514 = ( n38450 & n38512 ) | ( n38450 & n38513 ) | ( n38512 & n38513 ) ;
  assign n38515 = n38431 | n38512 ;
  assign n38516 = n38450 | n38515 ;
  assign n38517 = ~n38514 & n38516 ;
  assign n38518 = ~n38307 & n38312 ;
  assign n38519 = n38279 | n38307 ;
  assign n38520 = ( n38307 & ~n38312 ) | ( n38307 & n38519 ) | ( ~n38312 & n38519 ) ;
  assign n38521 = ( n38282 & ~n38518 ) | ( n38282 & n38520 ) | ( ~n38518 & n38520 ) ;
  assign n38522 = n22920 | n22921 ;
  assign n38523 = n834 | n1499 ;
  assign n38524 = n925 | n38523 ;
  assign n38525 = n2135 | n2214 ;
  assign n38526 = n38524 | n38525 ;
  assign n38527 = n38522 | n38526 ;
  assign n38528 = ( ~n13027 & n29455 ) | ( ~n13027 & n38527 ) | ( n29455 & n38527 ) ;
  assign n38529 = n29455 & n38527 ;
  assign n38530 = ( ~n13023 & n38528 ) | ( ~n13023 & n38529 ) | ( n38528 & n38529 ) ;
  assign n38531 = n35800 | n38530 ;
  assign n38532 = n617 | n5860 ;
  assign n38533 = n414 | n38532 ;
  assign n38534 = n37516 | n37524 ;
  assign n38535 = n37514 | n38534 ;
  assign n38536 = n38533 | n38535 ;
  assign n38537 = n140 | n2053 ;
  assign n38538 = n214 | n959 ;
  assign n38539 = n666 | n38538 ;
  assign n38540 = n38537 | n38539 ;
  assign n38541 = n234 | n395 ;
  assign n38542 = n38540 | n38541 ;
  assign n38543 = n38536 | n38542 ;
  assign n38544 = n38531 | n38543 ;
  assign n38545 = n38304 | n38544 ;
  assign n38546 = n38304 & n38544 ;
  assign n38547 = n38545 & ~n38546 ;
  assign n38548 = n38520 & n38547 ;
  assign n38549 = n38307 & n38547 ;
  assign n38550 = ( ~n38312 & n38547 ) | ( ~n38312 & n38549 ) | ( n38547 & n38549 ) ;
  assign n38551 = ( n38282 & n38548 ) | ( n38282 & n38550 ) | ( n38548 & n38550 ) ;
  assign n38552 = n38521 & ~n38551 ;
  assign n38553 = n38546 | n38548 ;
  assign n38554 = n38545 & ~n38553 ;
  assign n38555 = n38546 | n38550 ;
  assign n38556 = n38545 & ~n38555 ;
  assign n38557 = ( ~n38282 & n38554 ) | ( ~n38282 & n38556 ) | ( n38554 & n38556 ) ;
  assign n38558 = n38552 | n38557 ;
  assign n38559 = n1060 & ~n27371 ;
  assign n38560 = ~n27363 & n38559 ;
  assign n38561 = n1065 & ~n27606 ;
  assign n38562 = ~n27597 & n38561 ;
  assign n38563 = n38560 | n38562 ;
  assign n38564 = n1057 & ~n28503 ;
  assign n38565 = n28498 & n38564 ;
  assign n38566 = n38563 | n38565 ;
  assign n38567 = n1062 & n28794 ;
  assign n38568 = ( n1062 & n28783 ) | ( n1062 & n38567 ) | ( n28783 & n38567 ) ;
  assign n38569 = n38566 | n38568 ;
  assign n38570 = n38558 & n38569 ;
  assign n38571 = n38558 & ~n38570 ;
  assign n38573 = n1826 & n28492 ;
  assign n38574 = n1823 & ~n28714 ;
  assign n38575 = n38573 | n38574 ;
  assign n38572 = n1829 & n29620 ;
  assign n38577 = n1821 | n38572 ;
  assign n38578 = n38575 | n38577 ;
  assign n38576 = n38572 | n38575 ;
  assign n38579 = n38576 & n38578 ;
  assign n38580 = ( ~n29642 & n38578 ) | ( ~n29642 & n38579 ) | ( n38578 & n38579 ) ;
  assign n38581 = n38578 | n38579 ;
  assign n38582 = ( n29629 & n38580 ) | ( n29629 & n38581 ) | ( n38580 & n38581 ) ;
  assign n38583 = ~x29 & n38582 ;
  assign n38584 = x29 | n38582 ;
  assign n38585 = ( ~n38582 & n38583 ) | ( ~n38582 & n38584 ) | ( n38583 & n38584 ) ;
  assign n38586 = ~n38558 & n38569 ;
  assign n38587 = n38585 & n38586 ;
  assign n38588 = ( n38571 & n38585 ) | ( n38571 & n38587 ) | ( n38585 & n38587 ) ;
  assign n38589 = n38585 | n38586 ;
  assign n38590 = n38571 | n38589 ;
  assign n38591 = ~n38588 & n38590 ;
  assign n38592 = n38321 | n38337 ;
  assign n38593 = ( n38321 & ~n38322 ) | ( n38321 & n38592 ) | ( ~n38322 & n38592 ) ;
  assign n38594 = n38591 & n38593 ;
  assign n38595 = n38591 | n38593 ;
  assign n38596 = ~n38594 & n38595 ;
  assign n38597 = n2315 & ~n30186 ;
  assign n38598 = n2312 & ~n30199 ;
  assign n38599 = n2308 & n30212 ;
  assign n38600 = n38598 | n38599 ;
  assign n38601 = n38597 | n38600 ;
  assign n38602 = n2306 | n38597 ;
  assign n38603 = n38600 | n38602 ;
  assign n38604 = ( ~n30241 & n38601 ) | ( ~n30241 & n38603 ) | ( n38601 & n38603 ) ;
  assign n38605 = ~x26 & n38603 ;
  assign n38606 = ~x26 & n38601 ;
  assign n38607 = ( ~n30241 & n38605 ) | ( ~n30241 & n38606 ) | ( n38605 & n38606 ) ;
  assign n38608 = x26 | n38606 ;
  assign n38609 = x26 | n38605 ;
  assign n38610 = ( ~n30241 & n38608 ) | ( ~n30241 & n38609 ) | ( n38608 & n38609 ) ;
  assign n38611 = ( ~n38604 & n38607 ) | ( ~n38604 & n38610 ) | ( n38607 & n38610 ) ;
  assign n38612 = n38596 & ~n38611 ;
  assign n38613 = n38596 | n38611 ;
  assign n38614 = ( ~n38596 & n38612 ) | ( ~n38596 & n38613 ) | ( n38612 & n38613 ) ;
  assign n38615 = n38342 | n38357 ;
  assign n38616 = ( n38342 & ~n38344 ) | ( n38342 & n38615 ) | ( ~n38344 & n38615 ) ;
  assign n38617 = n38614 | n38616 ;
  assign n38618 = n38614 & n38616 ;
  assign n38619 = n38617 & ~n38618 ;
  assign n38620 = n2932 & n31295 ;
  assign n38621 = n2925 & ~n31309 ;
  assign n38622 = n2928 & ~n31323 ;
  assign n38623 = n38621 | n38622 ;
  assign n38624 = n38620 | n38623 ;
  assign n38625 = n2936 | n38620 ;
  assign n38626 = n38623 | n38625 ;
  assign n38627 = ( n31355 & n38624 ) | ( n31355 & n38626 ) | ( n38624 & n38626 ) ;
  assign n38628 = x23 & n38626 ;
  assign n38629 = x23 & n38624 ;
  assign n38630 = ( n31355 & n38628 ) | ( n31355 & n38629 ) | ( n38628 & n38629 ) ;
  assign n38631 = x23 & ~n38629 ;
  assign n38632 = x23 & ~n38628 ;
  assign n38633 = ( ~n31355 & n38631 ) | ( ~n31355 & n38632 ) | ( n38631 & n38632 ) ;
  assign n38634 = ( n38627 & ~n38630 ) | ( n38627 & n38633 ) | ( ~n38630 & n38633 ) ;
  assign n38635 = ~n38619 & n38634 ;
  assign n38636 = n38614 | n38634 ;
  assign n38637 = ( n38616 & n38634 ) | ( n38616 & n38636 ) | ( n38634 & n38636 ) ;
  assign n38638 = n38617 & ~n38637 ;
  assign n38639 = n38635 | n38638 ;
  assign n38640 = ( n38364 & ~n38365 ) | ( n38364 & n38381 ) | ( ~n38365 & n38381 ) ;
  assign n38641 = n38639 | n38640 ;
  assign n38642 = n38639 & n38640 ;
  assign n38643 = n38641 & ~n38642 ;
  assign n38644 = n3547 & ~n32442 ;
  assign n38645 = n3544 & n32306 ;
  assign n38646 = n3541 & n32293 ;
  assign n38647 = n38645 | n38646 ;
  assign n38648 = n38644 | n38647 ;
  assign n38649 = n3537 | n38644 ;
  assign n38650 = n38647 | n38649 ;
  assign n38651 = ( ~n32458 & n38648 ) | ( ~n32458 & n38650 ) | ( n38648 & n38650 ) ;
  assign n38652 = ~x20 & n38650 ;
  assign n38653 = ~x20 & n38648 ;
  assign n38654 = ( ~n32458 & n38652 ) | ( ~n32458 & n38653 ) | ( n38652 & n38653 ) ;
  assign n38655 = x20 | n38653 ;
  assign n38656 = x20 | n38652 ;
  assign n38657 = ( ~n32458 & n38655 ) | ( ~n32458 & n38656 ) | ( n38655 & n38656 ) ;
  assign n38658 = ( ~n38651 & n38654 ) | ( ~n38651 & n38657 ) | ( n38654 & n38657 ) ;
  assign n38659 = ~n38643 & n38658 ;
  assign n38660 = n38642 | n38658 ;
  assign n38661 = n38641 & ~n38660 ;
  assign n38662 = n38659 | n38661 ;
  assign n38663 = n38386 | n38400 ;
  assign n38664 = ( n38386 & ~n38387 ) | ( n38386 & n38663 ) | ( ~n38387 & n38663 ) ;
  assign n38665 = n38662 | n38664 ;
  assign n38666 = n38662 & n38664 ;
  assign n38667 = n38665 & ~n38666 ;
  assign n38668 = n4471 & n33526 ;
  assign n38669 = n4466 & n33436 ;
  assign n38670 = n4468 & ~n33423 ;
  assign n38671 = n38669 | n38670 ;
  assign n38672 = n38668 | n38671 ;
  assign n38673 = n4475 & n33545 ;
  assign n38674 = n4475 & ~n33548 ;
  assign n38675 = ( ~n32456 & n38673 ) | ( ~n32456 & n38674 ) | ( n38673 & n38674 ) ;
  assign n38676 = n38672 | n38675 ;
  assign n38677 = n4475 | n38672 ;
  assign n38678 = ( n33536 & n38676 ) | ( n33536 & n38677 ) | ( n38676 & n38677 ) ;
  assign n38679 = x17 | n38678 ;
  assign n38680 = ~x17 & n38678 ;
  assign n38681 = ( ~n38678 & n38679 ) | ( ~n38678 & n38680 ) | ( n38679 & n38680 ) ;
  assign n38682 = ~n38667 & n38681 ;
  assign n38683 = n38662 | n38681 ;
  assign n38684 = ( n38664 & n38681 ) | ( n38664 & n38683 ) | ( n38681 & n38683 ) ;
  assign n38685 = n38665 & ~n38684 ;
  assign n38686 = n38682 | n38685 ;
  assign n38687 = ( n38408 & ~n38409 ) | ( n38408 & n38425 ) | ( ~n38409 & n38425 ) ;
  assign n38688 = n38686 | n38687 ;
  assign n38689 = n38686 & n38687 ;
  assign n38690 = n38688 & ~n38689 ;
  assign n38691 = n5234 & ~n35371 ;
  assign n38692 = n5237 & n34656 ;
  assign n38693 = n5231 & n35021 ;
  assign n38694 = n38692 | n38693 ;
  assign n38695 = n38691 | n38694 ;
  assign n38696 = n5227 & ~n35392 ;
  assign n38697 = n5227 & ~n35395 ;
  assign n38698 = ( ~n32456 & n38696 ) | ( ~n32456 & n38697 ) | ( n38696 & n38697 ) ;
  assign n38699 = n38695 | n38698 ;
  assign n38700 = n5227 | n38695 ;
  assign n38701 = ( n35381 & n38699 ) | ( n35381 & n38700 ) | ( n38699 & n38700 ) ;
  assign n38702 = x14 | n38701 ;
  assign n38703 = ~x14 & n38701 ;
  assign n38704 = ( ~n38701 & n38702 ) | ( ~n38701 & n38703 ) | ( n38702 & n38703 ) ;
  assign n38705 = ~n38690 & n38704 ;
  assign n38706 = n38689 | n38704 ;
  assign n38707 = n38688 & ~n38706 ;
  assign n38708 = n38705 | n38707 ;
  assign n38709 = n38517 & ~n38708 ;
  assign n38710 = n38517 | n38708 ;
  assign n38711 = ( ~n38517 & n38709 ) | ( ~n38517 & n38710 ) | ( n38709 & n38710 ) ;
  assign n38712 = ( n38455 & ~n38456 ) | ( n38455 & n38472 ) | ( ~n38456 & n38472 ) ;
  assign n38713 = n38711 | n38712 ;
  assign n38714 = n38711 & n38712 ;
  assign n38715 = n38713 & ~n38714 ;
  assign n38716 = ~n38478 & n38483 ;
  assign n38717 = n38715 & ~n38716 ;
  assign n38718 = n38478 | n38484 ;
  assign n38719 = n38715 & n38718 ;
  assign n38720 = ( n38255 & n38717 ) | ( n38255 & n38719 ) | ( n38717 & n38719 ) ;
  assign n38721 = n38478 & n38715 ;
  assign n38722 = ( n38488 & n38715 ) | ( n38488 & n38721 ) | ( n38715 & n38721 ) ;
  assign n38723 = ( n37754 & n38720 ) | ( n37754 & n38722 ) | ( n38720 & n38722 ) ;
  assign n38724 = ( n37756 & n38720 ) | ( n37756 & n38722 ) | ( n38720 & n38722 ) ;
  assign n38725 = ( n36959 & n38723 ) | ( n36959 & n38724 ) | ( n38723 & n38724 ) ;
  assign n38726 = n38478 | n38488 ;
  assign n38727 = ( n38255 & ~n38716 ) | ( n38255 & n38718 ) | ( ~n38716 & n38718 ) ;
  assign n38728 = ( n37754 & n38726 ) | ( n37754 & n38727 ) | ( n38726 & n38727 ) ;
  assign n38729 = n38715 | n38728 ;
  assign n38730 = ( n37756 & n38726 ) | ( n37756 & n38727 ) | ( n38726 & n38727 ) ;
  assign n38731 = n38715 | n38730 ;
  assign n38732 = ( n36959 & n38729 ) | ( n36959 & n38731 ) | ( n38729 & n38731 ) ;
  assign n38733 = ~n38725 & n38732 ;
  assign n38734 = n38267 | n38499 ;
  assign n38735 = n38030 & ~n38734 ;
  assign n38736 = n38733 | n38735 ;
  assign n38737 = n38733 & ~n38734 ;
  assign n38738 = n38030 & n38737 ;
  assign n38739 = n38736 & ~n38738 ;
  assign n38740 = n1057 & n28492 ;
  assign n38741 = n1060 & ~n27606 ;
  assign n38742 = ~n27597 & n38741 ;
  assign n38743 = n1065 & ~n28503 ;
  assign n38744 = n28498 & n38743 ;
  assign n38745 = n38742 | n38744 ;
  assign n38746 = n38740 | n38745 ;
  assign n38747 = n1062 | n38746 ;
  assign n38748 = ( ~n28749 & n38746 ) | ( ~n28749 & n38747 ) | ( n38746 & n38747 ) ;
  assign n38749 = n705 | n13295 ;
  assign n38750 = n1625 | n38749 ;
  assign n38751 = n931 | n38750 ;
  assign n38752 = n13327 | n38751 ;
  assign n38753 = n3407 & ~n38752 ;
  assign n38754 = n6971 | n6980 ;
  assign n38755 = n38753 & ~n38754 ;
  assign n38756 = n1352 | n1725 ;
  assign n38757 = n1348 | n38756 ;
  assign n38758 = n1785 | n2051 ;
  assign n38759 = n1398 | n38758 ;
  assign n38760 = n38757 | n38759 ;
  assign n38761 = n112 | n213 ;
  assign n38762 = n1126 | n38761 ;
  assign n38763 = n229 | n518 ;
  assign n38764 = n38762 | n38763 ;
  assign n38765 = n38760 | n38764 ;
  assign n38766 = n38755 & ~n38765 ;
  assign n38767 = n38304 & n38766 ;
  assign n38768 = n38304 | n38766 ;
  assign n38769 = ~n38767 & n38768 ;
  assign n38770 = n27400 & n36083 ;
  assign n38771 = ~x11 & n27400 ;
  assign n38772 = n36083 & n38771 ;
  assign n38773 = x11 | n38771 ;
  assign n38774 = ( x11 & n36083 ) | ( x11 & n38773 ) | ( n36083 & n38773 ) ;
  assign n38775 = ( ~n38770 & n38772 ) | ( ~n38770 & n38774 ) | ( n38772 & n38774 ) ;
  assign n38776 = n38769 & ~n38775 ;
  assign n38777 = ~n38769 & n38775 ;
  assign n38778 = n38776 | n38777 ;
  assign n38779 = n38747 & ~n38778 ;
  assign n38780 = n38746 & ~n38778 ;
  assign n38781 = ( ~n28749 & n38779 ) | ( ~n28749 & n38780 ) | ( n38779 & n38780 ) ;
  assign n38782 = n38748 & ~n38781 ;
  assign n38783 = n38747 | n38778 ;
  assign n38784 = n38746 | n38778 ;
  assign n38785 = ( ~n28749 & n38783 ) | ( ~n28749 & n38784 ) | ( n38783 & n38784 ) ;
  assign n38786 = ~n38782 & n38785 ;
  assign n38787 = ( n38282 & n38553 ) | ( n38282 & n38555 ) | ( n38553 & n38555 ) ;
  assign n38788 = ~n38785 & n38787 ;
  assign n38789 = ( n38782 & n38787 ) | ( n38782 & n38788 ) | ( n38787 & n38788 ) ;
  assign n38790 = n38786 | n38789 ;
  assign n38791 = n38787 & ~n38789 ;
  assign n38792 = n38790 & ~n38791 ;
  assign n38793 = n38570 & ~n38792 ;
  assign n38794 = ( n38588 & ~n38792 ) | ( n38588 & n38793 ) | ( ~n38792 & n38793 ) ;
  assign n38795 = ~n38570 & n38792 ;
  assign n38796 = ~n38588 & n38795 ;
  assign n38797 = n38794 | n38796 ;
  assign n38798 = n1829 & ~n30199 ;
  assign n38799 = n1826 & ~n28714 ;
  assign n38800 = n1823 & n29620 ;
  assign n38801 = n38799 | n38800 ;
  assign n38802 = n38798 | n38801 ;
  assign n38803 = n1821 | n38798 ;
  assign n38804 = n38801 | n38803 ;
  assign n38805 = ( ~n30299 & n38802 ) | ( ~n30299 & n38804 ) | ( n38802 & n38804 ) ;
  assign n38806 = ~x29 & n38804 ;
  assign n38807 = ~x29 & n38802 ;
  assign n38808 = ( ~n30299 & n38806 ) | ( ~n30299 & n38807 ) | ( n38806 & n38807 ) ;
  assign n38809 = x29 | n38807 ;
  assign n38810 = x29 | n38806 ;
  assign n38811 = ( ~n30299 & n38809 ) | ( ~n30299 & n38810 ) | ( n38809 & n38810 ) ;
  assign n38812 = ( ~n38805 & n38808 ) | ( ~n38805 & n38811 ) | ( n38808 & n38811 ) ;
  assign n38813 = ~n38797 & n38812 ;
  assign n38814 = n38797 | n38813 ;
  assign n38815 = n2315 & ~n31309 ;
  assign n38816 = n2312 & n30212 ;
  assign n38817 = n2308 & ~n30186 ;
  assign n38818 = n38816 | n38817 ;
  assign n38819 = n38815 | n38818 ;
  assign n38820 = n2306 | n38815 ;
  assign n38821 = n38818 | n38820 ;
  assign n38822 = ( n31404 & n38819 ) | ( n31404 & n38821 ) | ( n38819 & n38821 ) ;
  assign n38823 = x26 & n38821 ;
  assign n38824 = x26 & n38819 ;
  assign n38825 = ( n31404 & n38823 ) | ( n31404 & n38824 ) | ( n38823 & n38824 ) ;
  assign n38826 = x26 & ~n38824 ;
  assign n38827 = x26 & ~n38823 ;
  assign n38828 = ( ~n31404 & n38826 ) | ( ~n31404 & n38827 ) | ( n38826 & n38827 ) ;
  assign n38829 = ( n38822 & ~n38825 ) | ( n38822 & n38828 ) | ( ~n38825 & n38828 ) ;
  assign n38830 = n38797 & n38812 ;
  assign n38831 = n38829 & n38830 ;
  assign n38832 = ( ~n38814 & n38829 ) | ( ~n38814 & n38831 ) | ( n38829 & n38831 ) ;
  assign n38833 = n38829 | n38830 ;
  assign n38834 = n38814 & ~n38833 ;
  assign n38835 = n38832 | n38834 ;
  assign n38836 = n38594 | n38611 ;
  assign n38837 = ( n38594 & n38596 ) | ( n38594 & n38836 ) | ( n38596 & n38836 ) ;
  assign n38838 = n38835 & ~n38837 ;
  assign n38839 = ~n38835 & n38837 ;
  assign n38840 = n38838 | n38839 ;
  assign n38841 = n2932 & n32306 ;
  assign n38842 = n2925 & ~n31323 ;
  assign n38843 = n2928 & n31295 ;
  assign n38844 = n38842 | n38843 ;
  assign n38845 = n38841 | n38844 ;
  assign n38846 = n2936 | n38841 ;
  assign n38847 = n38844 | n38846 ;
  assign n38848 = ( ~n32525 & n38845 ) | ( ~n32525 & n38847 ) | ( n38845 & n38847 ) ;
  assign n38849 = ~x23 & n38847 ;
  assign n38850 = ~x23 & n38845 ;
  assign n38851 = ( ~n32525 & n38849 ) | ( ~n32525 & n38850 ) | ( n38849 & n38850 ) ;
  assign n38852 = x23 | n38850 ;
  assign n38853 = x23 | n38849 ;
  assign n38854 = ( ~n32525 & n38852 ) | ( ~n32525 & n38853 ) | ( n38852 & n38853 ) ;
  assign n38855 = ( ~n38848 & n38851 ) | ( ~n38848 & n38854 ) | ( n38851 & n38854 ) ;
  assign n38856 = ~n38840 & n38855 ;
  assign n38857 = n38840 | n38856 ;
  assign n38859 = n38618 | n38634 ;
  assign n38860 = ( n38618 & n38619 ) | ( n38618 & n38859 ) | ( n38619 & n38859 ) ;
  assign n38858 = n38840 & n38855 ;
  assign n38861 = n38858 & n38860 ;
  assign n38862 = ( ~n38857 & n38860 ) | ( ~n38857 & n38861 ) | ( n38860 & n38861 ) ;
  assign n38863 = n38858 | n38860 ;
  assign n38864 = n38857 & ~n38863 ;
  assign n38865 = n38862 | n38864 ;
  assign n38880 = ( n38642 & n38643 ) | ( n38642 & n38660 ) | ( n38643 & n38660 ) ;
  assign n38866 = n3547 & n33436 ;
  assign n38867 = n3544 & n32293 ;
  assign n38868 = n3541 & ~n32442 ;
  assign n38869 = n38867 | n38868 ;
  assign n38870 = n38866 | n38869 ;
  assign n38871 = n3537 & ~n33441 ;
  assign n38872 = ~n32456 & n38871 ;
  assign n38873 = ( n3537 & n34271 ) | ( n3537 & n38872 ) | ( n34271 & n38872 ) ;
  assign n38874 = n38870 | n38873 ;
  assign n38875 = x20 | n38870 ;
  assign n38876 = n38873 | n38875 ;
  assign n38877 = ~x20 & n38875 ;
  assign n38878 = ( ~x20 & n38873 ) | ( ~x20 & n38877 ) | ( n38873 & n38877 ) ;
  assign n38879 = ( ~n38874 & n38876 ) | ( ~n38874 & n38878 ) | ( n38876 & n38878 ) ;
  assign n38881 = n38879 & n38880 ;
  assign n38882 = n38880 & ~n38881 ;
  assign n38883 = ~n38865 & n38879 ;
  assign n38884 = ~n38880 & n38883 ;
  assign n38885 = ( ~n38865 & n38882 ) | ( ~n38865 & n38884 ) | ( n38882 & n38884 ) ;
  assign n38886 = n38865 & ~n38879 ;
  assign n38887 = ( n38865 & n38880 ) | ( n38865 & n38886 ) | ( n38880 & n38886 ) ;
  assign n38888 = ~n38882 & n38887 ;
  assign n38889 = n38885 | n38888 ;
  assign n38890 = n4471 & n34656 ;
  assign n38891 = n4466 & ~n33423 ;
  assign n38892 = n4468 & n33526 ;
  assign n38893 = n38891 | n38892 ;
  assign n38894 = n38890 | n38893 ;
  assign n38895 = n4475 | n38890 ;
  assign n38896 = n38893 | n38895 ;
  assign n38897 = ( n34667 & n38894 ) | ( n34667 & n38896 ) | ( n38894 & n38896 ) ;
  assign n38898 = x17 & n38896 ;
  assign n38899 = x17 & n38894 ;
  assign n38900 = ( n34667 & n38898 ) | ( n34667 & n38899 ) | ( n38898 & n38899 ) ;
  assign n38901 = x17 & ~n38899 ;
  assign n38902 = x17 & ~n38898 ;
  assign n38903 = ( ~n34667 & n38901 ) | ( ~n34667 & n38902 ) | ( n38901 & n38902 ) ;
  assign n38904 = ( n38897 & ~n38900 ) | ( n38897 & n38903 ) | ( ~n38900 & n38903 ) ;
  assign n38905 = ~n38889 & n38904 ;
  assign n38906 = n38889 | n38905 ;
  assign n38908 = n38666 | n38681 ;
  assign n38909 = ( n38666 & n38667 ) | ( n38666 & n38908 ) | ( n38667 & n38908 ) ;
  assign n38907 = n38889 & n38904 ;
  assign n38910 = n38907 & n38909 ;
  assign n38911 = ( ~n38906 & n38909 ) | ( ~n38906 & n38910 ) | ( n38909 & n38910 ) ;
  assign n38912 = n38907 | n38909 ;
  assign n38913 = n38906 & ~n38912 ;
  assign n38914 = n38911 | n38913 ;
  assign n38930 = ( n38689 & n38690 ) | ( n38689 & n38706 ) | ( n38690 & n38706 ) ;
  assign n38915 = n5234 & n35746 ;
  assign n38916 = n5237 & n35021 ;
  assign n38917 = n5231 & ~n35371 ;
  assign n38918 = n38916 | n38917 ;
  assign n38919 = n38915 | n38918 ;
  assign n38920 = n5227 | n38915 ;
  assign n38921 = n38918 | n38920 ;
  assign n38922 = ( ~n35759 & n38919 ) | ( ~n35759 & n38921 ) | ( n38919 & n38921 ) ;
  assign n38923 = ~x14 & n38921 ;
  assign n38924 = ~x14 & n38919 ;
  assign n38925 = ( ~n35759 & n38923 ) | ( ~n35759 & n38924 ) | ( n38923 & n38924 ) ;
  assign n38926 = x14 | n38924 ;
  assign n38927 = x14 | n38923 ;
  assign n38928 = ( ~n35759 & n38926 ) | ( ~n35759 & n38927 ) | ( n38926 & n38927 ) ;
  assign n38929 = ( ~n38922 & n38925 ) | ( ~n38922 & n38928 ) | ( n38925 & n38928 ) ;
  assign n38931 = n38929 & n38930 ;
  assign n38932 = n38930 & ~n38931 ;
  assign n38933 = ~n38914 & n38929 ;
  assign n38934 = ~n38930 & n38933 ;
  assign n38935 = ( ~n38914 & n38932 ) | ( ~n38914 & n38934 ) | ( n38932 & n38934 ) ;
  assign n38936 = n38914 & ~n38929 ;
  assign n38937 = ( n38914 & n38930 ) | ( n38914 & n38936 ) | ( n38930 & n38936 ) ;
  assign n38938 = ~n38932 & n38937 ;
  assign n38939 = n38935 | n38938 ;
  assign n38940 = n38514 | n38708 ;
  assign n38941 = ( n38514 & n38517 ) | ( n38514 & n38940 ) | ( n38517 & n38940 ) ;
  assign n38942 = ~n38939 & n38941 ;
  assign n38943 = n38939 & ~n38941 ;
  assign n38944 = n38942 | n38943 ;
  assign n38945 = n38714 | n38717 ;
  assign n38946 = ~n38944 & n38945 ;
  assign n38947 = n38714 | n38719 ;
  assign n38948 = ~n38944 & n38947 ;
  assign n38949 = ( n38255 & n38946 ) | ( n38255 & n38948 ) | ( n38946 & n38948 ) ;
  assign n38950 = n38714 | n38721 ;
  assign n38951 = ~n38944 & n38950 ;
  assign n38952 = n38714 | n38715 ;
  assign n38953 = ~n38944 & n38952 ;
  assign n38954 = ( n38488 & n38951 ) | ( n38488 & n38953 ) | ( n38951 & n38953 ) ;
  assign n38955 = ( n37754 & n38949 ) | ( n37754 & n38954 ) | ( n38949 & n38954 ) ;
  assign n38956 = ( n37756 & n38949 ) | ( n37756 & n38954 ) | ( n38949 & n38954 ) ;
  assign n38957 = ( n36959 & n38955 ) | ( n36959 & n38956 ) | ( n38955 & n38956 ) ;
  assign n38958 = ( n38255 & n38945 ) | ( n38255 & n38947 ) | ( n38945 & n38947 ) ;
  assign n38959 = ( n38488 & n38950 ) | ( n38488 & n38952 ) | ( n38950 & n38952 ) ;
  assign n38960 = ( n37754 & n38958 ) | ( n37754 & n38959 ) | ( n38958 & n38959 ) ;
  assign n38961 = n38944 & ~n38960 ;
  assign n38962 = ( n37756 & n38958 ) | ( n37756 & n38959 ) | ( n38958 & n38959 ) ;
  assign n38963 = n38944 & ~n38962 ;
  assign n38964 = ( ~n36959 & n38961 ) | ( ~n36959 & n38963 ) | ( n38961 & n38963 ) ;
  assign n38965 = n38957 | n38964 ;
  assign n38966 = ~n38738 & n38965 ;
  assign n38967 = n38738 & ~n38965 ;
  assign n38968 = n38966 | n38967 ;
  assign n38969 = n38905 | n38911 ;
  assign n38970 = n38781 | n38789 ;
  assign n38997 = n1057 & ~n28714 ;
  assign n38998 = n1065 & n28492 ;
  assign n38999 = n1060 & ~n28503 ;
  assign n39000 = n28498 & n38999 ;
  assign n39001 = n38998 | n39000 ;
  assign n39002 = n38997 | n39001 ;
  assign n39003 = n1062 & ~n28731 ;
  assign n39004 = ~n28518 & n39003 ;
  assign n39005 = n39002 | n39004 ;
  assign n39006 = n1062 | n39002 ;
  assign n39007 = ( n28720 & n39005 ) | ( n28720 & n39006 ) | ( n39005 & n39006 ) ;
  assign n38971 = n481 | n718 ;
  assign n38972 = n3347 | n38971 ;
  assign n38973 = n7948 | n38972 ;
  assign n38974 = n30936 | n38973 ;
  assign n38975 = n624 | n35448 ;
  assign n38976 = n38974 | n38975 ;
  assign n38977 = n30884 | n38976 ;
  assign n38978 = n513 | n22913 ;
  assign n38979 = n22923 | n38978 ;
  assign n38980 = n22911 | n38979 ;
  assign n38981 = n36138 | n38980 ;
  assign n38982 = n38977 | n38981 ;
  assign n38983 = n438 | n748 ;
  assign n38984 = n138 | n406 ;
  assign n38985 = n94 | n38984 ;
  assign n38986 = n38983 | n38985 ;
  assign n38987 = n6915 | n38986 ;
  assign n38988 = n38982 | n38987 ;
  assign n38989 = ( n38768 & ~n38769 ) | ( n38768 & n38988 ) | ( ~n38769 & n38988 ) ;
  assign n38990 = n38768 | n38988 ;
  assign n38991 = ( n38775 & n38989 ) | ( n38775 & n38990 ) | ( n38989 & n38990 ) ;
  assign n38992 = n38768 & ~n38769 ;
  assign n38993 = n38988 & n38992 ;
  assign n38994 = n38768 & n38988 ;
  assign n38995 = ( n38775 & n38993 ) | ( n38775 & n38994 ) | ( n38993 & n38994 ) ;
  assign n38996 = n38991 & ~n38995 ;
  assign n39008 = n38996 | n39007 ;
  assign n39009 = ~n38996 & n39007 ;
  assign n39010 = ( ~n39007 & n39008 ) | ( ~n39007 & n39009 ) | ( n39008 & n39009 ) ;
  assign n39011 = n38970 | n39010 ;
  assign n39012 = n38970 & n39010 ;
  assign n39013 = n39011 & ~n39012 ;
  assign n39014 = n1829 & n30212 ;
  assign n39015 = n1826 & n29620 ;
  assign n39016 = n1823 & ~n30199 ;
  assign n39017 = n39015 | n39016 ;
  assign n39018 = n39014 | n39017 ;
  assign n39019 = n30266 & ~n39018 ;
  assign n39020 = ~n30276 & n39019 ;
  assign n39021 = n1821 | n39014 ;
  assign n39022 = n39017 | n39021 ;
  assign n39023 = ~n39020 & n39022 ;
  assign n39024 = x29 & n39022 ;
  assign n39025 = ~n39020 & n39024 ;
  assign n39026 = x29 & ~n39024 ;
  assign n39027 = ( x29 & n39020 ) | ( x29 & n39026 ) | ( n39020 & n39026 ) ;
  assign n39028 = ( n39023 & ~n39025 ) | ( n39023 & n39027 ) | ( ~n39025 & n39027 ) ;
  assign n39029 = n39013 & n39028 ;
  assign n39030 = n39013 | n39028 ;
  assign n39031 = ~n39029 & n39030 ;
  assign n39032 = n38794 | n38812 ;
  assign n39033 = ( n38794 & ~n38797 ) | ( n38794 & n39032 ) | ( ~n38797 & n39032 ) ;
  assign n39034 = n39031 & n39033 ;
  assign n39035 = n39031 | n39033 ;
  assign n39036 = ~n39034 & n39035 ;
  assign n39037 = n2315 & ~n31323 ;
  assign n39038 = n2312 & ~n30186 ;
  assign n39039 = n2308 & ~n31309 ;
  assign n39040 = n39038 | n39039 ;
  assign n39041 = n39037 | n39040 ;
  assign n39042 = n2306 & n31384 ;
  assign n39043 = n2306 & n31386 ;
  assign n39044 = ( ~n30232 & n39042 ) | ( ~n30232 & n39043 ) | ( n39042 & n39043 ) ;
  assign n39045 = n39041 | n39044 ;
  assign n39046 = n2306 | n39041 ;
  assign n39047 = ( ~n31376 & n39045 ) | ( ~n31376 & n39046 ) | ( n39045 & n39046 ) ;
  assign n39048 = x26 | n39047 ;
  assign n39049 = ~x26 & n39047 ;
  assign n39050 = ( ~n39047 & n39048 ) | ( ~n39047 & n39049 ) | ( n39048 & n39049 ) ;
  assign n39051 = n39036 & ~n39050 ;
  assign n39052 = n39036 | n39050 ;
  assign n39053 = ( ~n39036 & n39051 ) | ( ~n39036 & n39052 ) | ( n39051 & n39052 ) ;
  assign n39054 = n38832 | n38837 ;
  assign n39055 = ( n38832 & ~n38835 ) | ( n38832 & n39054 ) | ( ~n38835 & n39054 ) ;
  assign n39056 = n39053 | n39055 ;
  assign n39057 = n39053 & n39055 ;
  assign n39058 = n39056 & ~n39057 ;
  assign n39059 = n2932 & n32293 ;
  assign n39060 = n2925 & n31295 ;
  assign n39061 = n2928 & n32306 ;
  assign n39062 = n39060 | n39061 ;
  assign n39063 = n39059 | n39062 ;
  assign n39064 = n2936 & n32497 ;
  assign n39065 = ( n2936 & n32494 ) | ( n2936 & n39064 ) | ( n32494 & n39064 ) ;
  assign n39066 = n39063 | n39065 ;
  assign n39067 = x23 | n39063 ;
  assign n39068 = n39065 | n39067 ;
  assign n39069 = ~x23 & n39067 ;
  assign n39070 = ( ~x23 & n39065 ) | ( ~x23 & n39069 ) | ( n39065 & n39069 ) ;
  assign n39071 = ( ~n39066 & n39068 ) | ( ~n39066 & n39070 ) | ( n39068 & n39070 ) ;
  assign n39072 = ~n39058 & n39071 ;
  assign n39073 = n39057 | n39071 ;
  assign n39074 = n39056 & ~n39073 ;
  assign n39075 = n39072 | n39074 ;
  assign n39076 = n38856 | n38862 ;
  assign n39077 = n39075 | n39076 ;
  assign n39078 = n39075 & n39076 ;
  assign n39079 = n39077 & ~n39078 ;
  assign n39080 = n3547 & ~n33423 ;
  assign n39081 = n3544 & ~n32442 ;
  assign n39082 = n3541 & n33436 ;
  assign n39083 = n39081 | n39082 ;
  assign n39084 = n39080 | n39083 ;
  assign n39085 = n3537 & n33575 ;
  assign n39086 = n3537 & ~n33577 ;
  assign n39087 = ( ~n32456 & n39085 ) | ( ~n32456 & n39086 ) | ( n39085 & n39086 ) ;
  assign n39088 = n39084 | n39087 ;
  assign n39089 = n3537 | n39084 ;
  assign n39090 = ( n33567 & n39088 ) | ( n33567 & n39089 ) | ( n39088 & n39089 ) ;
  assign n39091 = x20 | n39090 ;
  assign n39092 = ~x20 & n39090 ;
  assign n39093 = ( ~n39090 & n39091 ) | ( ~n39090 & n39092 ) | ( n39091 & n39092 ) ;
  assign n39094 = ~n39079 & n39093 ;
  assign n39095 = n39075 | n39093 ;
  assign n39096 = ( n39076 & n39093 ) | ( n39076 & n39095 ) | ( n39093 & n39095 ) ;
  assign n39097 = n39077 & ~n39096 ;
  assign n39098 = n39094 | n39097 ;
  assign n39099 = n38881 | n38884 ;
  assign n39100 = n38865 & ~n38881 ;
  assign n39101 = ( n38882 & n39099 ) | ( n38882 & ~n39100 ) | ( n39099 & ~n39100 ) ;
  assign n39102 = n39098 & n39101 ;
  assign n39103 = n39098 & ~n39102 ;
  assign n39104 = n4471 & n35021 ;
  assign n39105 = n4466 & n33526 ;
  assign n39106 = n4468 & n34656 ;
  assign n39107 = n39105 | n39106 ;
  assign n39108 = n39104 | n39107 ;
  assign n39109 = n4475 | n39104 ;
  assign n39110 = n39107 | n39109 ;
  assign n39111 = ( n35033 & n39108 ) | ( n35033 & n39110 ) | ( n39108 & n39110 ) ;
  assign n39112 = x17 & n39110 ;
  assign n39113 = x17 & n39108 ;
  assign n39114 = ( n35033 & n39112 ) | ( n35033 & n39113 ) | ( n39112 & n39113 ) ;
  assign n39115 = x17 & ~n39113 ;
  assign n39116 = x17 & ~n39112 ;
  assign n39117 = ( ~n35033 & n39115 ) | ( ~n35033 & n39116 ) | ( n39115 & n39116 ) ;
  assign n39118 = ( n39111 & ~n39114 ) | ( n39111 & n39117 ) | ( ~n39114 & n39117 ) ;
  assign n39119 = ~n39098 & n39101 ;
  assign n39120 = n39118 & n39119 ;
  assign n39121 = ( n39103 & n39118 ) | ( n39103 & n39120 ) | ( n39118 & n39120 ) ;
  assign n39122 = n39118 | n39119 ;
  assign n39123 = n39103 | n39122 ;
  assign n39124 = ~n39121 & n39123 ;
  assign n39125 = n38969 | n39124 ;
  assign n39126 = n38969 & n39124 ;
  assign n39127 = n39125 & ~n39126 ;
  assign n39128 = n5234 & n36083 ;
  assign n39129 = n5237 & ~n35371 ;
  assign n39130 = n5231 & n35746 ;
  assign n39131 = n39129 | n39130 ;
  assign n39132 = n39128 | n39131 ;
  assign n39133 = n5227 | n39128 ;
  assign n39134 = n39131 | n39133 ;
  assign n39135 = ( n36107 & n39132 ) | ( n36107 & n39134 ) | ( n39132 & n39134 ) ;
  assign n39136 = n39132 | n39134 ;
  assign n39137 = ( n36094 & n39135 ) | ( n36094 & n39136 ) | ( n39135 & n39136 ) ;
  assign n39138 = x14 & n39137 ;
  assign n39139 = x14 & ~n39137 ;
  assign n39140 = ( n39137 & ~n39138 ) | ( n39137 & n39139 ) | ( ~n39138 & n39139 ) ;
  assign n39141 = ~n39127 & n39140 ;
  assign n39142 = n39124 | n39140 ;
  assign n39143 = ( n38969 & n39140 ) | ( n38969 & n39142 ) | ( n39140 & n39142 ) ;
  assign n39144 = n39125 & ~n39143 ;
  assign n39145 = n39141 | n39144 ;
  assign n39146 = n38931 | n38934 ;
  assign n39147 = n38914 & ~n38931 ;
  assign n39148 = ( n38932 & n39146 ) | ( n38932 & ~n39147 ) | ( n39146 & ~n39147 ) ;
  assign n39149 = n39145 & n39148 ;
  assign n39150 = n39145 & ~n39149 ;
  assign n39151 = ~n39145 & n39148 ;
  assign n39152 = n39150 | n39151 ;
  assign n39153 = n38942 | n38949 ;
  assign n39154 = n38942 | n38951 ;
  assign n39155 = n38942 | n38953 ;
  assign n39156 = ( n38488 & n39154 ) | ( n38488 & n39155 ) | ( n39154 & n39155 ) ;
  assign n39157 = ( n37754 & n39153 ) | ( n37754 & n39156 ) | ( n39153 & n39156 ) ;
  assign n39158 = n39152 & n39157 ;
  assign n39159 = ( n37756 & n39153 ) | ( n37756 & n39156 ) | ( n39153 & n39156 ) ;
  assign n39160 = n39152 & n39159 ;
  assign n39161 = ( n36959 & n39158 ) | ( n36959 & n39160 ) | ( n39158 & n39160 ) ;
  assign n39162 = n39152 | n39157 ;
  assign n39163 = n39152 | n39159 ;
  assign n39164 = ( n36959 & n39162 ) | ( n36959 & n39163 ) | ( n39162 & n39163 ) ;
  assign n39165 = ~n39161 & n39164 ;
  assign n39166 = ~n38967 & n39165 ;
  assign n39167 = n38967 & ~n39165 ;
  assign n39168 = n39166 | n39167 ;
  assign n39169 = n28075 & n36083 ;
  assign n39170 = n5237 & n35746 ;
  assign n39171 = n39169 | n39170 ;
  assign n39172 = n5227 | n39171 ;
  assign n39173 = ( n36103 & n39171 ) | ( n36103 & n39172 ) | ( n39171 & n39172 ) ;
  assign n39174 = ( n36105 & n39171 ) | ( n36105 & n39172 ) | ( n39171 & n39172 ) ;
  assign n39175 = ( n32456 & n39173 ) | ( n32456 & n39174 ) | ( n39173 & n39174 ) ;
  assign n39176 = x14 & n39175 ;
  assign n39177 = x14 & ~n39175 ;
  assign n39178 = ( n39175 & ~n39176 ) | ( n39175 & n39177 ) | ( ~n39176 & n39177 ) ;
  assign n39179 = n39102 & n39178 ;
  assign n39180 = ( n39121 & n39178 ) | ( n39121 & n39179 ) | ( n39178 & n39179 ) ;
  assign n39181 = n39102 | n39178 ;
  assign n39182 = n39121 | n39181 ;
  assign n39183 = ~n39180 & n39182 ;
  assign n39184 = n1057 & n29620 ;
  assign n39185 = n1060 & n28492 ;
  assign n39186 = n1065 & ~n28714 ;
  assign n39187 = n39185 | n39186 ;
  assign n39188 = n39184 | n39187 ;
  assign n39189 = n1062 | n39184 ;
  assign n39190 = n39187 | n39189 ;
  assign n39191 = ( ~n29642 & n39188 ) | ( ~n29642 & n39190 ) | ( n39188 & n39190 ) ;
  assign n39192 = n39188 | n39190 ;
  assign n39193 = ( n29629 & n39191 ) | ( n29629 & n39192 ) | ( n39191 & n39192 ) ;
  assign n39194 = n16801 | n16806 ;
  assign n39195 = ( ~n1303 & n2874 ) | ( ~n1303 & n10344 ) | ( n2874 & n10344 ) ;
  assign n39196 = n2874 & n10344 ;
  assign n39197 = ( ~n1613 & n39195 ) | ( ~n1613 & n39196 ) | ( n39195 & n39196 ) ;
  assign n39198 = n1614 | n39197 ;
  assign n39199 = n517 | n19256 ;
  assign n39200 = n39198 | n39199 ;
  assign n39201 = n20391 | n39200 ;
  assign n39202 = n6858 | n6859 ;
  assign n39203 = n1104 & ~n39202 ;
  assign n39204 = ~n268 & n39203 ;
  assign n39205 = ~n39201 & n39204 ;
  assign n39206 = ~n39194 & n39205 ;
  assign n39207 = n94 | n608 ;
  assign n39208 = n1001 | n39207 ;
  assign n39209 = n46 | n64 ;
  assign n39210 = n444 | n39209 ;
  assign n39211 = n39208 | n39210 ;
  assign n39212 = n99 | n424 ;
  assign n39213 = n568 | n39212 ;
  assign n39214 = n39211 | n39213 ;
  assign n39215 = n39206 & ~n39214 ;
  assign n39216 = n38988 & n39215 ;
  assign n39217 = n38988 | n39215 ;
  assign n39218 = n39184 & n39217 ;
  assign n39219 = ( n39187 & n39217 ) | ( n39187 & n39218 ) | ( n39217 & n39218 ) ;
  assign n39220 = ~n39216 & n39219 ;
  assign n39221 = ~n39216 & n39217 ;
  assign n39222 = n39190 & n39221 ;
  assign n39223 = ( ~n29642 & n39220 ) | ( ~n29642 & n39222 ) | ( n39220 & n39222 ) ;
  assign n39224 = n39220 | n39222 ;
  assign n39225 = ( n29629 & n39223 ) | ( n29629 & n39224 ) | ( n39223 & n39224 ) ;
  assign n39226 = n39193 & ~n39225 ;
  assign n39227 = n38996 & n39002 ;
  assign n39228 = ( n38996 & n39004 ) | ( n38996 & n39227 ) | ( n39004 & n39227 ) ;
  assign n39229 = ( n1062 & n38996 ) | ( n1062 & n39227 ) | ( n38996 & n39227 ) ;
  assign n39230 = ( n28720 & n39228 ) | ( n28720 & n39229 ) | ( n39228 & n39229 ) ;
  assign n39231 = n38991 & ~n39230 ;
  assign n39232 = n39217 & ~n39221 ;
  assign n39233 = ( ~n39190 & n39217 ) | ( ~n39190 & n39232 ) | ( n39217 & n39232 ) ;
  assign n39234 = n39216 & n39217 ;
  assign n39235 = ( n39217 & ~n39219 ) | ( n39217 & n39234 ) | ( ~n39219 & n39234 ) ;
  assign n39236 = ( n29642 & n39233 ) | ( n29642 & n39235 ) | ( n39233 & n39235 ) ;
  assign n39237 = n39233 & n39235 ;
  assign n39238 = ( ~n29629 & n39236 ) | ( ~n29629 & n39237 ) | ( n39236 & n39237 ) ;
  assign n39239 = ~n39216 & n39238 ;
  assign n39240 = ~n39231 & n39239 ;
  assign n39241 = ( n39226 & ~n39231 ) | ( n39226 & n39240 ) | ( ~n39231 & n39240 ) ;
  assign n39242 = n39231 & ~n39239 ;
  assign n39243 = ~n39226 & n39242 ;
  assign n39244 = n39241 | n39243 ;
  assign n39245 = n39012 | n39028 ;
  assign n39246 = ( n39012 & n39013 ) | ( n39012 & n39245 ) | ( n39013 & n39245 ) ;
  assign n39247 = n39244 & ~n39246 ;
  assign n39248 = ~n39244 & n39246 ;
  assign n39249 = n39247 | n39248 ;
  assign n39250 = n1829 & ~n30186 ;
  assign n39251 = n1826 & ~n30199 ;
  assign n39252 = n1823 & n30212 ;
  assign n39253 = n39251 | n39252 ;
  assign n39254 = n39250 | n39253 ;
  assign n39255 = n1821 | n39250 ;
  assign n39256 = n39253 | n39255 ;
  assign n39257 = ( ~n30241 & n39254 ) | ( ~n30241 & n39256 ) | ( n39254 & n39256 ) ;
  assign n39258 = ~x29 & n39256 ;
  assign n39259 = ~x29 & n39254 ;
  assign n39260 = ( ~n30241 & n39258 ) | ( ~n30241 & n39259 ) | ( n39258 & n39259 ) ;
  assign n39261 = x29 | n39259 ;
  assign n39262 = x29 | n39258 ;
  assign n39263 = ( ~n30241 & n39261 ) | ( ~n30241 & n39262 ) | ( n39261 & n39262 ) ;
  assign n39264 = ( ~n39257 & n39260 ) | ( ~n39257 & n39263 ) | ( n39260 & n39263 ) ;
  assign n39265 = ~n39249 & n39264 ;
  assign n39266 = n39249 | n39265 ;
  assign n39267 = n2315 & n31295 ;
  assign n39268 = n2312 & ~n31309 ;
  assign n39269 = n2308 & ~n31323 ;
  assign n39270 = n39268 | n39269 ;
  assign n39271 = n39267 | n39270 ;
  assign n39272 = n2306 | n39267 ;
  assign n39273 = n39270 | n39272 ;
  assign n39274 = ( n31355 & n39271 ) | ( n31355 & n39273 ) | ( n39271 & n39273 ) ;
  assign n39275 = x26 & n39273 ;
  assign n39276 = x26 & n39271 ;
  assign n39277 = ( n31355 & n39275 ) | ( n31355 & n39276 ) | ( n39275 & n39276 ) ;
  assign n39278 = x26 & ~n39276 ;
  assign n39279 = x26 & ~n39275 ;
  assign n39280 = ( ~n31355 & n39278 ) | ( ~n31355 & n39279 ) | ( n39278 & n39279 ) ;
  assign n39281 = ( n39274 & ~n39277 ) | ( n39274 & n39280 ) | ( ~n39277 & n39280 ) ;
  assign n39282 = n39249 & n39264 ;
  assign n39283 = n39281 & n39282 ;
  assign n39284 = ( ~n39266 & n39281 ) | ( ~n39266 & n39283 ) | ( n39281 & n39283 ) ;
  assign n39285 = n39281 | n39282 ;
  assign n39286 = n39266 & ~n39285 ;
  assign n39287 = n39284 | n39286 ;
  assign n39288 = n39034 | n39050 ;
  assign n39289 = ( n39034 & n39036 ) | ( n39034 & n39288 ) | ( n39036 & n39288 ) ;
  assign n39290 = n39287 & ~n39289 ;
  assign n39291 = ~n39287 & n39289 ;
  assign n39292 = n39290 | n39291 ;
  assign n39293 = n2932 & ~n32442 ;
  assign n39294 = n2925 & n32306 ;
  assign n39295 = n2928 & n32293 ;
  assign n39296 = n39294 | n39295 ;
  assign n39297 = n39293 | n39296 ;
  assign n39298 = n2936 | n39293 ;
  assign n39299 = n39296 | n39298 ;
  assign n39300 = ( ~n32458 & n39297 ) | ( ~n32458 & n39299 ) | ( n39297 & n39299 ) ;
  assign n39301 = ~x23 & n39299 ;
  assign n39302 = ~x23 & n39297 ;
  assign n39303 = ( ~n32458 & n39301 ) | ( ~n32458 & n39302 ) | ( n39301 & n39302 ) ;
  assign n39304 = x23 | n39302 ;
  assign n39305 = x23 | n39301 ;
  assign n39306 = ( ~n32458 & n39304 ) | ( ~n32458 & n39305 ) | ( n39304 & n39305 ) ;
  assign n39307 = ( ~n39300 & n39303 ) | ( ~n39300 & n39306 ) | ( n39303 & n39306 ) ;
  assign n39308 = n39292 & n39307 ;
  assign n39309 = n39289 | n39307 ;
  assign n39310 = ( ~n39287 & n39307 ) | ( ~n39287 & n39309 ) | ( n39307 & n39309 ) ;
  assign n39311 = n39290 | n39310 ;
  assign n39312 = ~n39308 & n39311 ;
  assign n39313 = ( n39057 & n39058 ) | ( n39057 & n39073 ) | ( n39058 & n39073 ) ;
  assign n39314 = n39312 & ~n39313 ;
  assign n39315 = ~n39312 & n39313 ;
  assign n39316 = n39314 | n39315 ;
  assign n39317 = n3547 & n33526 ;
  assign n39318 = n3544 & n33436 ;
  assign n39319 = n3541 & ~n33423 ;
  assign n39320 = n39318 | n39319 ;
  assign n39321 = n39317 | n39320 ;
  assign n39322 = n3537 & n33545 ;
  assign n39323 = n3537 & ~n33548 ;
  assign n39324 = ( ~n32456 & n39322 ) | ( ~n32456 & n39323 ) | ( n39322 & n39323 ) ;
  assign n39325 = n39321 | n39324 ;
  assign n39326 = n3537 | n39321 ;
  assign n39327 = ( n33536 & n39325 ) | ( n33536 & n39326 ) | ( n39325 & n39326 ) ;
  assign n39328 = x20 | n39327 ;
  assign n39329 = ~x20 & n39327 ;
  assign n39330 = ( ~n39327 & n39328 ) | ( ~n39327 & n39329 ) | ( n39328 & n39329 ) ;
  assign n39331 = n39316 & n39330 ;
  assign n39332 = n39313 | n39330 ;
  assign n39333 = ( ~n39312 & n39330 ) | ( ~n39312 & n39332 ) | ( n39330 & n39332 ) ;
  assign n39334 = n39314 | n39333 ;
  assign n39335 = ~n39331 & n39334 ;
  assign n39336 = n39078 | n39093 ;
  assign n39337 = ( n39078 & n39079 ) | ( n39078 & n39336 ) | ( n39079 & n39336 ) ;
  assign n39338 = n39335 & ~n39337 ;
  assign n39339 = ~n39335 & n39337 ;
  assign n39340 = n39338 | n39339 ;
  assign n39341 = n4471 & ~n35371 ;
  assign n39342 = n4466 & n34656 ;
  assign n39343 = n4468 & n35021 ;
  assign n39344 = n39342 | n39343 ;
  assign n39345 = n39341 | n39344 ;
  assign n39346 = n4475 & ~n35392 ;
  assign n39347 = n4475 & ~n35395 ;
  assign n39348 = ( ~n32456 & n39346 ) | ( ~n32456 & n39347 ) | ( n39346 & n39347 ) ;
  assign n39349 = n39345 | n39348 ;
  assign n39350 = n4475 | n39345 ;
  assign n39351 = ( n35381 & n39349 ) | ( n35381 & n39350 ) | ( n39349 & n39350 ) ;
  assign n39352 = x17 | n39351 ;
  assign n39353 = ~x17 & n39351 ;
  assign n39354 = ( ~n39351 & n39352 ) | ( ~n39351 & n39353 ) | ( n39352 & n39353 ) ;
  assign n39355 = n39340 & n39354 ;
  assign n39356 = n39339 | n39354 ;
  assign n39357 = n39338 | n39356 ;
  assign n39358 = ~n39355 & n39357 ;
  assign n39359 = n39183 & ~n39358 ;
  assign n39360 = n39183 | n39358 ;
  assign n39361 = ( ~n39183 & n39359 ) | ( ~n39183 & n39360 ) | ( n39359 & n39360 ) ;
  assign n39362 = n39126 | n39140 ;
  assign n39363 = ( n39126 & n39127 ) | ( n39126 & n39362 ) | ( n39127 & n39362 ) ;
  assign n39364 = n39361 & ~n39363 ;
  assign n39365 = ~n39361 & n39363 ;
  assign n39366 = n39364 | n39365 ;
  assign n39367 = n39149 & ~n39366 ;
  assign n39368 = ( n39161 & ~n39366 ) | ( n39161 & n39367 ) | ( ~n39366 & n39367 ) ;
  assign n39369 = ~n39149 & n39366 ;
  assign n39370 = ~n39161 & n39369 ;
  assign n39371 = n39368 | n39370 ;
  assign n39372 = ~n38965 & n39165 ;
  assign n39373 = n38738 & n39372 ;
  assign n39374 = n39371 & ~n39373 ;
  assign n39375 = ~n39371 & n39372 ;
  assign n39376 = n38738 & n39375 ;
  assign n39377 = n39374 | n39376 ;
  assign n39378 = n4292 | n4295 ;
  assign n39379 = n28273 | n28277 ;
  assign n39380 = n810 | n18101 ;
  assign n39381 = n10721 | n39380 ;
  assign n39382 = n2614 | n28280 ;
  assign n39383 = n39381 | n39382 ;
  assign n39384 = n1402 & ~n39383 ;
  assign n39385 = ~n39379 & n39384 ;
  assign n39386 = ~n39378 & n39385 ;
  assign n39387 = n444 | n1355 ;
  assign n39388 = n1250 | n39387 ;
  assign n39389 = n183 | n434 ;
  assign n39390 = n39388 | n39389 ;
  assign n39391 = n4204 | n39390 ;
  assign n39392 = n39386 & ~n39391 ;
  assign n39393 = ~n38988 & n39392 ;
  assign n39394 = n38988 & ~n39392 ;
  assign n39395 = n39393 | n39394 ;
  assign n39396 = n28546 & n36083 ;
  assign n39397 = ~x14 & n28546 ;
  assign n39398 = n36083 & n39397 ;
  assign n39399 = x14 | n39397 ;
  assign n39400 = ( x14 & n36083 ) | ( x14 & n39399 ) | ( n36083 & n39399 ) ;
  assign n39401 = ( ~n39396 & n39398 ) | ( ~n39396 & n39400 ) | ( n39398 & n39400 ) ;
  assign n39402 = n39395 | n39401 ;
  assign n39403 = n39395 & n39401 ;
  assign n39404 = n39402 & ~n39403 ;
  assign n39405 = ~n39238 & n39404 ;
  assign n39406 = n39238 & ~n39404 ;
  assign n39407 = n39405 | n39406 ;
  assign n39408 = n1057 & ~n30199 ;
  assign n39409 = n1060 & ~n28714 ;
  assign n39410 = n1065 & n29620 ;
  assign n39411 = n39409 | n39410 ;
  assign n39412 = n39408 | n39411 ;
  assign n39413 = n1062 | n39408 ;
  assign n39414 = n39411 | n39413 ;
  assign n39415 = ( ~n30299 & n39412 ) | ( ~n30299 & n39414 ) | ( n39412 & n39414 ) ;
  assign n39416 = n39407 & n39415 ;
  assign n39417 = n39407 | n39415 ;
  assign n39418 = ~n39416 & n39417 ;
  assign n39419 = n1829 & ~n31309 ;
  assign n39420 = n1826 & n30212 ;
  assign n39421 = n1823 & ~n30186 ;
  assign n39422 = n39420 | n39421 ;
  assign n39423 = n39419 | n39422 ;
  assign n39424 = n1821 | n39419 ;
  assign n39425 = n39422 | n39424 ;
  assign n39426 = ( n31404 & n39423 ) | ( n31404 & n39425 ) | ( n39423 & n39425 ) ;
  assign n39427 = x29 & n39425 ;
  assign n39428 = x29 & n39423 ;
  assign n39429 = ( n31404 & n39427 ) | ( n31404 & n39428 ) | ( n39427 & n39428 ) ;
  assign n39430 = x29 & ~n39428 ;
  assign n39431 = x29 & ~n39427 ;
  assign n39432 = ( ~n31404 & n39430 ) | ( ~n31404 & n39431 ) | ( n39430 & n39431 ) ;
  assign n39433 = ( n39426 & ~n39429 ) | ( n39426 & n39432 ) | ( ~n39429 & n39432 ) ;
  assign n39434 = ~n39418 & n39433 ;
  assign n39435 = n39418 | n39434 ;
  assign n39436 = n39418 & n39433 ;
  assign n39437 = n39435 & ~n39436 ;
  assign n39438 = ~n39241 & n39244 ;
  assign n39439 = ( n39241 & n39246 ) | ( n39241 & ~n39438 ) | ( n39246 & ~n39438 ) ;
  assign n39440 = n39437 & ~n39439 ;
  assign n39441 = ~n39437 & n39439 ;
  assign n39442 = n39440 | n39441 ;
  assign n39443 = n2315 & n32306 ;
  assign n39444 = n2312 & ~n31323 ;
  assign n39445 = n2308 & n31295 ;
  assign n39446 = n39444 | n39445 ;
  assign n39447 = n39443 | n39446 ;
  assign n39448 = n2306 | n39443 ;
  assign n39449 = n39446 | n39448 ;
  assign n39450 = ( ~n32525 & n39447 ) | ( ~n32525 & n39449 ) | ( n39447 & n39449 ) ;
  assign n39451 = ~x26 & n39449 ;
  assign n39452 = ~x26 & n39447 ;
  assign n39453 = ( ~n32525 & n39451 ) | ( ~n32525 & n39452 ) | ( n39451 & n39452 ) ;
  assign n39454 = x26 | n39452 ;
  assign n39455 = x26 | n39451 ;
  assign n39456 = ( ~n32525 & n39454 ) | ( ~n32525 & n39455 ) | ( n39454 & n39455 ) ;
  assign n39457 = ( ~n39450 & n39453 ) | ( ~n39450 & n39456 ) | ( n39453 & n39456 ) ;
  assign n39458 = ~n39442 & n39457 ;
  assign n39459 = n39442 | n39458 ;
  assign n39460 = n39442 & n39457 ;
  assign n39461 = n39459 & ~n39460 ;
  assign n39462 = n39265 | n39284 ;
  assign n39463 = n39461 & ~n39462 ;
  assign n39464 = ~n39461 & n39462 ;
  assign n39465 = n39463 | n39464 ;
  assign n39480 = n39291 | n39307 ;
  assign n39481 = ( n39291 & ~n39292 ) | ( n39291 & n39480 ) | ( ~n39292 & n39480 ) ;
  assign n39466 = n2932 & n33436 ;
  assign n39467 = n2925 & n32293 ;
  assign n39468 = n2928 & ~n32442 ;
  assign n39469 = n39467 | n39468 ;
  assign n39470 = n39466 | n39469 ;
  assign n39471 = n2936 & ~n33441 ;
  assign n39472 = ~n32456 & n39471 ;
  assign n39473 = ( n2936 & n34271 ) | ( n2936 & n39472 ) | ( n34271 & n39472 ) ;
  assign n39474 = n39470 | n39473 ;
  assign n39475 = x23 | n39470 ;
  assign n39476 = n39473 | n39475 ;
  assign n39477 = ~x23 & n39475 ;
  assign n39478 = ( ~x23 & n39473 ) | ( ~x23 & n39477 ) | ( n39473 & n39477 ) ;
  assign n39479 = ( ~n39474 & n39476 ) | ( ~n39474 & n39478 ) | ( n39476 & n39478 ) ;
  assign n39482 = n39479 & n39481 ;
  assign n39483 = n39481 & ~n39482 ;
  assign n39484 = n39479 & ~n39481 ;
  assign n39485 = ~n39465 & n39484 ;
  assign n39486 = ( ~n39465 & n39483 ) | ( ~n39465 & n39485 ) | ( n39483 & n39485 ) ;
  assign n39487 = n39465 & ~n39484 ;
  assign n39488 = ~n39483 & n39487 ;
  assign n39489 = n39486 | n39488 ;
  assign n39490 = n3547 & n34656 ;
  assign n39491 = n3544 & ~n33423 ;
  assign n39492 = n3541 & n33526 ;
  assign n39493 = n39491 | n39492 ;
  assign n39494 = n39490 | n39493 ;
  assign n39495 = n3537 | n39490 ;
  assign n39496 = n39493 | n39495 ;
  assign n39497 = ( n34667 & n39494 ) | ( n34667 & n39496 ) | ( n39494 & n39496 ) ;
  assign n39498 = x20 & n39496 ;
  assign n39499 = x20 & n39494 ;
  assign n39500 = ( n34667 & n39498 ) | ( n34667 & n39499 ) | ( n39498 & n39499 ) ;
  assign n39501 = x20 & ~n39499 ;
  assign n39502 = x20 & ~n39498 ;
  assign n39503 = ( ~n34667 & n39501 ) | ( ~n34667 & n39502 ) | ( n39501 & n39502 ) ;
  assign n39504 = ( n39497 & ~n39500 ) | ( n39497 & n39503 ) | ( ~n39500 & n39503 ) ;
  assign n39505 = ~n39489 & n39504 ;
  assign n39506 = n39489 | n39505 ;
  assign n39508 = n39315 | n39330 ;
  assign n39509 = ( n39315 & ~n39316 ) | ( n39315 & n39508 ) | ( ~n39316 & n39508 ) ;
  assign n39507 = n39489 & n39504 ;
  assign n39510 = n39507 & n39509 ;
  assign n39511 = ( ~n39506 & n39509 ) | ( ~n39506 & n39510 ) | ( n39509 & n39510 ) ;
  assign n39512 = n39507 | n39509 ;
  assign n39513 = n39506 & ~n39512 ;
  assign n39514 = n39511 | n39513 ;
  assign n39530 = ( n39339 & ~n39340 ) | ( n39339 & n39356 ) | ( ~n39340 & n39356 ) ;
  assign n39515 = n4471 & n35746 ;
  assign n39516 = n4466 & n35021 ;
  assign n39517 = n4468 & ~n35371 ;
  assign n39518 = n39516 | n39517 ;
  assign n39519 = n39515 | n39518 ;
  assign n39520 = n4475 | n39515 ;
  assign n39521 = n39518 | n39520 ;
  assign n39522 = ( ~n35759 & n39519 ) | ( ~n35759 & n39521 ) | ( n39519 & n39521 ) ;
  assign n39523 = ~x17 & n39521 ;
  assign n39524 = ~x17 & n39519 ;
  assign n39525 = ( ~n35759 & n39523 ) | ( ~n35759 & n39524 ) | ( n39523 & n39524 ) ;
  assign n39526 = x17 | n39524 ;
  assign n39527 = x17 | n39523 ;
  assign n39528 = ( ~n35759 & n39526 ) | ( ~n35759 & n39527 ) | ( n39526 & n39527 ) ;
  assign n39529 = ( ~n39522 & n39525 ) | ( ~n39522 & n39528 ) | ( n39525 & n39528 ) ;
  assign n39531 = n39529 & n39530 ;
  assign n39532 = n39530 & ~n39531 ;
  assign n39533 = n39529 & ~n39530 ;
  assign n39534 = ~n39514 & n39533 ;
  assign n39535 = ( ~n39514 & n39532 ) | ( ~n39514 & n39534 ) | ( n39532 & n39534 ) ;
  assign n39536 = n39514 & ~n39533 ;
  assign n39537 = ~n39532 & n39536 ;
  assign n39538 = n39535 | n39537 ;
  assign n39539 = ~n39180 & n39358 ;
  assign n39540 = ( n39180 & n39183 ) | ( n39180 & ~n39539 ) | ( n39183 & ~n39539 ) ;
  assign n39541 = ~n39538 & n39540 ;
  assign n39542 = n39538 & ~n39540 ;
  assign n39543 = n39541 | n39542 ;
  assign n39544 = n39365 & ~n39543 ;
  assign n39545 = ( n39367 & ~n39543 ) | ( n39367 & n39544 ) | ( ~n39543 & n39544 ) ;
  assign n39546 = ( n39366 & n39543 ) | ( n39366 & ~n39544 ) | ( n39543 & ~n39544 ) ;
  assign n39547 = ( n39161 & n39545 ) | ( n39161 & ~n39546 ) | ( n39545 & ~n39546 ) ;
  assign n39548 = n39365 | n39367 ;
  assign n39549 = n39543 & ~n39548 ;
  assign n39550 = ~n39365 & n39366 ;
  assign n39551 = n39543 & n39550 ;
  assign n39552 = ( ~n39161 & n39549 ) | ( ~n39161 & n39551 ) | ( n39549 & n39551 ) ;
  assign n39553 = n39547 | n39552 ;
  assign n39554 = ~n39376 & n39553 ;
  assign n39555 = n39375 & ~n39553 ;
  assign n39556 = n38738 & n39555 ;
  assign n39557 = n39554 | n39556 ;
  assign n39558 = n39505 | n39511 ;
  assign n39559 = n39482 | n39486 ;
  assign n39560 = n1057 & n30212 ;
  assign n39561 = n1060 & n29620 ;
  assign n39562 = n1065 & ~n30199 ;
  assign n39563 = n39561 | n39562 ;
  assign n39564 = n39560 | n39563 ;
  assign n39565 = n1062 & ~n30266 ;
  assign n39566 = ( n1062 & n30276 ) | ( n1062 & n39565 ) | ( n30276 & n39565 ) ;
  assign n39567 = n39564 | n39566 ;
  assign n39568 = n11772 | n11773 ;
  assign n39569 = n1136 | n3422 ;
  assign n39570 = n6846 | n39569 ;
  assign n39571 = n25795 | n39570 ;
  assign n39572 = n39568 | n39571 ;
  assign n39573 = n13340 | n39572 ;
  assign n39574 = n561 | n1479 ;
  assign n39575 = n711 | n1723 ;
  assign n39576 = n39574 | n39575 ;
  assign n39577 = n39573 | n39576 ;
  assign n39578 = n405 | n5946 ;
  assign n39579 = n911 & ~n39578 ;
  assign n39580 = n233 | n1039 ;
  assign n39581 = n857 | n39580 ;
  assign n39582 = n198 | n443 ;
  assign n39583 = n39581 | n39582 ;
  assign n39584 = n39579 & ~n39583 ;
  assign n39585 = ~n39577 & n39584 ;
  assign n39586 = ( n39394 & ~n39395 ) | ( n39394 & n39585 ) | ( ~n39395 & n39585 ) ;
  assign n39587 = n39394 & n39585 ;
  assign n39588 = ( ~n39401 & n39586 ) | ( ~n39401 & n39587 ) | ( n39586 & n39587 ) ;
  assign n39589 = ~n39394 & n39395 ;
  assign n39590 = ~n39585 & n39589 ;
  assign n39591 = n39394 | n39585 ;
  assign n39592 = ( n39401 & n39590 ) | ( n39401 & ~n39591 ) | ( n39590 & ~n39591 ) ;
  assign n39593 = n39588 | n39592 ;
  assign n39594 = n39564 | n39593 ;
  assign n39595 = n39566 | n39594 ;
  assign n39596 = ~n39593 & n39594 ;
  assign n39597 = ( n39566 & ~n39593 ) | ( n39566 & n39596 ) | ( ~n39593 & n39596 ) ;
  assign n39598 = ( ~n39567 & n39595 ) | ( ~n39567 & n39597 ) | ( n39595 & n39597 ) ;
  assign n39599 = n39405 | n39415 ;
  assign n39600 = ( n39405 & ~n39407 ) | ( n39405 & n39599 ) | ( ~n39407 & n39599 ) ;
  assign n39601 = n39598 & ~n39600 ;
  assign n39602 = ~n39598 & n39600 ;
  assign n39603 = n39601 | n39602 ;
  assign n39604 = n1826 & ~n30186 ;
  assign n39605 = n1823 & ~n31309 ;
  assign n39606 = n39604 | n39605 ;
  assign n39607 = n1829 & ~n31323 ;
  assign n39608 = n1821 | n39607 ;
  assign n39609 = n39606 | n39608 ;
  assign n39610 = n39606 | n39607 ;
  assign n39611 = n31384 | n39610 ;
  assign n39612 = n31386 | n39610 ;
  assign n39613 = ( ~n30232 & n39611 ) | ( ~n30232 & n39612 ) | ( n39611 & n39612 ) ;
  assign n39614 = n39609 & n39613 ;
  assign n39615 = ( ~n31376 & n39609 ) | ( ~n31376 & n39614 ) | ( n39609 & n39614 ) ;
  assign n39616 = x29 & n39615 ;
  assign n39617 = x29 & ~n39615 ;
  assign n39618 = ( n39615 & ~n39616 ) | ( n39615 & n39617 ) | ( ~n39616 & n39617 ) ;
  assign n39619 = ~n39603 & n39618 ;
  assign n39620 = n39603 & ~n39618 ;
  assign n39621 = n39619 | n39620 ;
  assign n39622 = n39434 | n39439 ;
  assign n39623 = ( n39434 & ~n39437 ) | ( n39434 & n39622 ) | ( ~n39437 & n39622 ) ;
  assign n39624 = ~n39621 & n39623 ;
  assign n39625 = n39621 & ~n39623 ;
  assign n39626 = n39624 | n39625 ;
  assign n39627 = n2315 & n32293 ;
  assign n39628 = n2312 & n31295 ;
  assign n39629 = n2308 & n32306 ;
  assign n39630 = n39628 | n39629 ;
  assign n39631 = n39627 | n39630 ;
  assign n39632 = n2306 & n32497 ;
  assign n39633 = ( n2306 & n32494 ) | ( n2306 & n39632 ) | ( n32494 & n39632 ) ;
  assign n39634 = n39631 | n39633 ;
  assign n39635 = x26 | n39631 ;
  assign n39636 = n39633 | n39635 ;
  assign n39637 = ~x26 & n39635 ;
  assign n39638 = ( ~x26 & n39633 ) | ( ~x26 & n39637 ) | ( n39633 & n39637 ) ;
  assign n39639 = ( ~n39634 & n39636 ) | ( ~n39634 & n39638 ) | ( n39636 & n39638 ) ;
  assign n39640 = n39626 | n39639 ;
  assign n39641 = n39626 & ~n39639 ;
  assign n39642 = ( ~n39626 & n39640 ) | ( ~n39626 & n39641 ) | ( n39640 & n39641 ) ;
  assign n39643 = n39458 | n39462 ;
  assign n39644 = ( n39458 & ~n39461 ) | ( n39458 & n39643 ) | ( ~n39461 & n39643 ) ;
  assign n39645 = n39642 & ~n39644 ;
  assign n39646 = ~n39642 & n39644 ;
  assign n39647 = n39645 | n39646 ;
  assign n39648 = n2932 & ~n33423 ;
  assign n39649 = n2925 & ~n32442 ;
  assign n39650 = n2928 & n33436 ;
  assign n39651 = n39649 | n39650 ;
  assign n39652 = n39648 | n39651 ;
  assign n39653 = n2936 & n33575 ;
  assign n39654 = n2936 & ~n33577 ;
  assign n39655 = ( ~n32456 & n39653 ) | ( ~n32456 & n39654 ) | ( n39653 & n39654 ) ;
  assign n39656 = n39652 | n39655 ;
  assign n39657 = n2936 | n39652 ;
  assign n39658 = ( n33567 & n39656 ) | ( n33567 & n39657 ) | ( n39656 & n39657 ) ;
  assign n39659 = x23 | n39658 ;
  assign n39660 = ~x23 & n39658 ;
  assign n39661 = ( ~n39658 & n39659 ) | ( ~n39658 & n39660 ) | ( n39659 & n39660 ) ;
  assign n39662 = n39647 & n39661 ;
  assign n39663 = n39642 & ~n39661 ;
  assign n39664 = ( n39644 & n39661 ) | ( n39644 & ~n39663 ) | ( n39661 & ~n39663 ) ;
  assign n39665 = n39645 | n39664 ;
  assign n39666 = ~n39662 & n39665 ;
  assign n39667 = n39559 & ~n39666 ;
  assign n39668 = n39559 & ~n39667 ;
  assign n39669 = n3547 & n35021 ;
  assign n39670 = n3544 & n33526 ;
  assign n39671 = n3541 & n34656 ;
  assign n39672 = n39670 | n39671 ;
  assign n39673 = n39669 | n39672 ;
  assign n39674 = n3537 | n39669 ;
  assign n39675 = n39672 | n39674 ;
  assign n39676 = ( n35033 & n39673 ) | ( n35033 & n39675 ) | ( n39673 & n39675 ) ;
  assign n39677 = x20 & n39675 ;
  assign n39678 = x20 & n39673 ;
  assign n39679 = ( n35033 & n39677 ) | ( n35033 & n39678 ) | ( n39677 & n39678 ) ;
  assign n39680 = x20 & ~n39678 ;
  assign n39681 = x20 & ~n39677 ;
  assign n39682 = ( ~n35033 & n39680 ) | ( ~n35033 & n39681 ) | ( n39680 & n39681 ) ;
  assign n39683 = ( n39676 & ~n39679 ) | ( n39676 & n39682 ) | ( ~n39679 & n39682 ) ;
  assign n39684 = n39559 | n39666 ;
  assign n39685 = n39683 & ~n39684 ;
  assign n39686 = ( n39668 & n39683 ) | ( n39668 & n39685 ) | ( n39683 & n39685 ) ;
  assign n39687 = ~n39683 & n39684 ;
  assign n39688 = ~n39668 & n39687 ;
  assign n39689 = n39686 | n39688 ;
  assign n39690 = ~n39558 & n39689 ;
  assign n39691 = n39558 & ~n39689 ;
  assign n39692 = n39690 | n39691 ;
  assign n39693 = n4471 & n36083 ;
  assign n39694 = n4466 & ~n35371 ;
  assign n39695 = n4468 & n35746 ;
  assign n39696 = n39694 | n39695 ;
  assign n39697 = n39693 | n39696 ;
  assign n39698 = n4475 | n39693 ;
  assign n39699 = n39696 | n39698 ;
  assign n39700 = ( n36107 & n39697 ) | ( n36107 & n39699 ) | ( n39697 & n39699 ) ;
  assign n39701 = n39697 | n39699 ;
  assign n39702 = ( n36094 & n39700 ) | ( n36094 & n39701 ) | ( n39700 & n39701 ) ;
  assign n39703 = x17 & n39702 ;
  assign n39704 = x17 & ~n39702 ;
  assign n39705 = ( n39702 & ~n39703 ) | ( n39702 & n39704 ) | ( ~n39703 & n39704 ) ;
  assign n39706 = n39692 & n39705 ;
  assign n39707 = n39691 | n39705 ;
  assign n39708 = n39690 | n39707 ;
  assign n39709 = ~n39706 & n39708 ;
  assign n39710 = n39531 | n39535 ;
  assign n39711 = ~n39709 & n39710 ;
  assign n39712 = n39709 | n39711 ;
  assign n39713 = n39710 & ~n39711 ;
  assign n39714 = n39712 & ~n39713 ;
  assign n39715 = n39541 | n39544 ;
  assign n39716 = ~n39541 & n39543 ;
  assign n39717 = ( n39367 & n39715 ) | ( n39367 & ~n39716 ) | ( n39715 & ~n39716 ) ;
  assign n39718 = ~n39714 & n39717 ;
  assign n39719 = n39541 & ~n39714 ;
  assign n39720 = ( n39546 & n39714 ) | ( n39546 & ~n39719 ) | ( n39714 & ~n39719 ) ;
  assign n39721 = ( n39161 & n39718 ) | ( n39161 & ~n39720 ) | ( n39718 & ~n39720 ) ;
  assign n39722 = n39714 & ~n39717 ;
  assign n39723 = ~n39541 & n39546 ;
  assign n39724 = n39714 & n39723 ;
  assign n39725 = ( ~n39161 & n39722 ) | ( ~n39161 & n39724 ) | ( n39722 & n39724 ) ;
  assign n39726 = n39721 | n39725 ;
  assign n39727 = n39556 & ~n39726 ;
  assign n39728 = n39726 | n39727 ;
  assign n39729 = ( ~n39556 & n39727 ) | ( ~n39556 & n39728 ) | ( n39727 & n39728 ) ;
  assign n39730 = n29766 & n36083 ;
  assign n39731 = n4466 & n35746 ;
  assign n39732 = n39730 | n39731 ;
  assign n39733 = n4475 | n39732 ;
  assign n39734 = ( n36103 & n39732 ) | ( n36103 & n39733 ) | ( n39732 & n39733 ) ;
  assign n39735 = ( n36105 & n39732 ) | ( n36105 & n39733 ) | ( n39732 & n39733 ) ;
  assign n39736 = ( n32456 & n39734 ) | ( n32456 & n39735 ) | ( n39734 & n39735 ) ;
  assign n39737 = x17 & n39736 ;
  assign n39738 = x17 & ~n39736 ;
  assign n39739 = ( n39736 & ~n39737 ) | ( n39736 & n39738 ) | ( ~n39737 & n39738 ) ;
  assign n39740 = ~n39666 & n39739 ;
  assign n39741 = n39559 & n39740 ;
  assign n39742 = ( n39686 & n39739 ) | ( n39686 & n39741 ) | ( n39739 & n39741 ) ;
  assign n39743 = n39666 & ~n39739 ;
  assign n39744 = ( n39559 & n39739 ) | ( n39559 & ~n39743 ) | ( n39739 & ~n39743 ) ;
  assign n39745 = n39686 | n39744 ;
  assign n39746 = ~n39742 & n39745 ;
  assign n39747 = ~n39588 & n39593 ;
  assign n39748 = n39564 | n39588 ;
  assign n39749 = ( n39588 & ~n39593 ) | ( n39588 & n39748 ) | ( ~n39593 & n39748 ) ;
  assign n39750 = ( n39566 & ~n39747 ) | ( n39566 & n39749 ) | ( ~n39747 & n39749 ) ;
  assign n39751 = n391 | n601 ;
  assign n39752 = n112 | n288 ;
  assign n39753 = n1013 | n39752 ;
  assign n39754 = n39751 | n39753 ;
  assign n39755 = n1650 | n39754 ;
  assign n39756 = n19524 | n39755 ;
  assign n39757 = n12398 | n39756 ;
  assign n39758 = n26282 | n39757 ;
  assign n39759 = n324 | n566 ;
  assign n39760 = n254 | n39759 ;
  assign n39761 = n513 | n7842 ;
  assign n39762 = n201 | n1460 ;
  assign n39763 = n39761 | n39762 ;
  assign n39764 = n438 | n806 ;
  assign n39765 = n214 | n39764 ;
  assign n39766 = n142 | n39765 ;
  assign n39767 = n39763 | n39766 ;
  assign n39768 = n39760 | n39767 ;
  assign n39769 = n39758 | n39768 ;
  assign n39770 = n39585 & n39769 ;
  assign n39771 = n39585 | n39769 ;
  assign n39772 = n39588 & n39771 ;
  assign n39773 = ( ~n39593 & n39771 ) | ( ~n39593 & n39772 ) | ( n39771 & n39772 ) ;
  assign n39774 = ~n39770 & n39773 ;
  assign n39775 = ~n39770 & n39771 ;
  assign n39776 = n39749 & n39775 ;
  assign n39777 = ( n39566 & n39774 ) | ( n39566 & n39776 ) | ( n39774 & n39776 ) ;
  assign n39778 = n39750 & ~n39777 ;
  assign n39779 = n1057 & ~n30186 ;
  assign n39780 = n1060 & ~n30199 ;
  assign n39781 = n1065 & n30212 ;
  assign n39782 = n39780 | n39781 ;
  assign n39783 = n39779 | n39782 ;
  assign n39784 = n1062 | n39779 ;
  assign n39785 = n39782 | n39784 ;
  assign n39786 = ( ~n30241 & n39783 ) | ( ~n30241 & n39785 ) | ( n39783 & n39785 ) ;
  assign n39787 = n39770 & n39771 ;
  assign n39788 = ( n39771 & ~n39773 ) | ( n39771 & n39787 ) | ( ~n39773 & n39787 ) ;
  assign n39789 = ~n39770 & n39788 ;
  assign n39790 = n39771 & ~n39775 ;
  assign n39791 = ( ~n39749 & n39771 ) | ( ~n39749 & n39790 ) | ( n39771 & n39790 ) ;
  assign n39792 = ~n39770 & n39791 ;
  assign n39793 = ( ~n39566 & n39789 ) | ( ~n39566 & n39792 ) | ( n39789 & n39792 ) ;
  assign n39794 = n39786 & n39793 ;
  assign n39795 = ( n39778 & n39786 ) | ( n39778 & n39794 ) | ( n39786 & n39794 ) ;
  assign n39796 = n39786 | n39793 ;
  assign n39797 = n39778 | n39796 ;
  assign n39798 = ~n39795 & n39797 ;
  assign n39800 = n1826 & ~n31309 ;
  assign n39801 = n1823 & ~n31323 ;
  assign n39802 = n39800 | n39801 ;
  assign n39799 = n1829 & n31295 ;
  assign n39804 = n1821 | n39799 ;
  assign n39805 = n39802 | n39804 ;
  assign n39803 = n39799 | n39802 ;
  assign n39806 = n39803 & n39805 ;
  assign n39807 = ( n31355 & n39805 ) | ( n31355 & n39806 ) | ( n39805 & n39806 ) ;
  assign n39808 = x29 & n39806 ;
  assign n39809 = x29 & n39805 ;
  assign n39810 = ( n31355 & n39808 ) | ( n31355 & n39809 ) | ( n39808 & n39809 ) ;
  assign n39811 = x29 & ~n39808 ;
  assign n39812 = x29 & ~n39809 ;
  assign n39813 = ( ~n31355 & n39811 ) | ( ~n31355 & n39812 ) | ( n39811 & n39812 ) ;
  assign n39814 = ( n39807 & ~n39810 ) | ( n39807 & n39813 ) | ( ~n39810 & n39813 ) ;
  assign n39815 = n39798 & n39814 ;
  assign n39816 = n39798 | n39814 ;
  assign n39817 = ~n39815 & n39816 ;
  assign n39818 = n39602 | n39618 ;
  assign n39819 = ( n39602 & ~n39603 ) | ( n39602 & n39818 ) | ( ~n39603 & n39818 ) ;
  assign n39820 = n39817 & n39819 ;
  assign n39821 = n39817 | n39819 ;
  assign n39822 = ~n39820 & n39821 ;
  assign n39823 = n2315 & ~n32442 ;
  assign n39824 = n2312 & n32306 ;
  assign n39825 = n2308 & n32293 ;
  assign n39826 = n39824 | n39825 ;
  assign n39827 = n39823 | n39826 ;
  assign n39828 = n2306 | n39823 ;
  assign n39829 = n39826 | n39828 ;
  assign n39830 = ( ~n32458 & n39827 ) | ( ~n32458 & n39829 ) | ( n39827 & n39829 ) ;
  assign n39831 = ~x26 & n39829 ;
  assign n39832 = ~x26 & n39827 ;
  assign n39833 = ( ~n32458 & n39831 ) | ( ~n32458 & n39832 ) | ( n39831 & n39832 ) ;
  assign n39834 = x26 | n39832 ;
  assign n39835 = x26 | n39831 ;
  assign n39836 = ( ~n32458 & n39834 ) | ( ~n32458 & n39835 ) | ( n39834 & n39835 ) ;
  assign n39837 = ( ~n39830 & n39833 ) | ( ~n39830 & n39836 ) | ( n39833 & n39836 ) ;
  assign n39838 = n39822 & ~n39837 ;
  assign n39839 = n39822 | n39837 ;
  assign n39840 = ( ~n39822 & n39838 ) | ( ~n39822 & n39839 ) | ( n39838 & n39839 ) ;
  assign n39841 = n39624 | n39639 ;
  assign n39842 = ( n39624 & ~n39626 ) | ( n39624 & n39841 ) | ( ~n39626 & n39841 ) ;
  assign n39843 = n39840 | n39842 ;
  assign n39844 = n39840 & n39842 ;
  assign n39845 = n39843 & ~n39844 ;
  assign n39846 = n2932 & n33526 ;
  assign n39847 = n2925 & n33436 ;
  assign n39848 = n2928 & ~n33423 ;
  assign n39849 = n39847 | n39848 ;
  assign n39850 = n39846 | n39849 ;
  assign n39851 = n2936 & n33545 ;
  assign n39852 = n2936 & ~n33548 ;
  assign n39853 = ( ~n32456 & n39851 ) | ( ~n32456 & n39852 ) | ( n39851 & n39852 ) ;
  assign n39854 = n39850 | n39853 ;
  assign n39855 = n2936 | n39850 ;
  assign n39856 = ( n33536 & n39854 ) | ( n33536 & n39855 ) | ( n39854 & n39855 ) ;
  assign n39857 = x23 | n39856 ;
  assign n39858 = ~x23 & n39856 ;
  assign n39859 = ( ~n39856 & n39857 ) | ( ~n39856 & n39858 ) | ( n39857 & n39858 ) ;
  assign n39860 = ~n39845 & n39859 ;
  assign n39861 = n39840 | n39859 ;
  assign n39862 = ( n39842 & n39859 ) | ( n39842 & n39861 ) | ( n39859 & n39861 ) ;
  assign n39863 = n39843 & ~n39862 ;
  assign n39864 = n39860 | n39863 ;
  assign n39865 = n39646 | n39661 ;
  assign n39866 = ( n39646 & ~n39647 ) | ( n39646 & n39865 ) | ( ~n39647 & n39865 ) ;
  assign n39867 = n39864 | n39866 ;
  assign n39868 = n39864 & n39866 ;
  assign n39869 = n39867 & ~n39868 ;
  assign n39870 = n3547 & ~n35371 ;
  assign n39871 = n3544 & n34656 ;
  assign n39872 = n3541 & n35021 ;
  assign n39873 = n39871 | n39872 ;
  assign n39874 = n39870 | n39873 ;
  assign n39875 = n3537 & ~n35392 ;
  assign n39876 = n3537 & ~n35395 ;
  assign n39877 = ( ~n32456 & n39875 ) | ( ~n32456 & n39876 ) | ( n39875 & n39876 ) ;
  assign n39878 = n39874 | n39877 ;
  assign n39879 = n3537 | n39874 ;
  assign n39880 = ( n35381 & n39878 ) | ( n35381 & n39879 ) | ( n39878 & n39879 ) ;
  assign n39881 = x20 | n39880 ;
  assign n39882 = ~x20 & n39880 ;
  assign n39883 = ( ~n39880 & n39881 ) | ( ~n39880 & n39882 ) | ( n39881 & n39882 ) ;
  assign n39884 = ~n39869 & n39883 ;
  assign n39885 = n39864 | n39883 ;
  assign n39886 = ( n39866 & n39883 ) | ( n39866 & n39885 ) | ( n39883 & n39885 ) ;
  assign n39887 = n39867 & ~n39886 ;
  assign n39888 = n39884 | n39887 ;
  assign n39889 = n39746 & ~n39888 ;
  assign n39890 = n39746 | n39888 ;
  assign n39891 = ( ~n39746 & n39889 ) | ( ~n39746 & n39890 ) | ( n39889 & n39890 ) ;
  assign n39892 = ( n39691 & ~n39692 ) | ( n39691 & n39707 ) | ( ~n39692 & n39707 ) ;
  assign n39893 = n39891 | n39892 ;
  assign n39894 = n39891 & n39892 ;
  assign n39895 = n39893 & ~n39894 ;
  assign n39896 = ~n39711 & n39714 ;
  assign n39897 = n39711 | n39719 ;
  assign n39898 = ( n39546 & n39896 ) | ( n39546 & ~n39897 ) | ( n39896 & ~n39897 ) ;
  assign n39899 = n39895 & ~n39898 ;
  assign n39900 = n39895 & ~n39896 ;
  assign n39901 = n39711 & n39895 ;
  assign n39902 = ( n39717 & n39900 ) | ( n39717 & n39901 ) | ( n39900 & n39901 ) ;
  assign n39903 = ( n39161 & n39899 ) | ( n39161 & n39902 ) | ( n39899 & n39902 ) ;
  assign n39904 = ( n39711 & n39717 ) | ( n39711 & ~n39896 ) | ( n39717 & ~n39896 ) ;
  assign n39905 = n39895 | n39904 ;
  assign n39906 = ~n39895 & n39898 ;
  assign n39907 = ( n39161 & n39905 ) | ( n39161 & ~n39906 ) | ( n39905 & ~n39906 ) ;
  assign n39908 = ~n39903 & n39907 ;
  assign n39909 = n39727 | n39908 ;
  assign n39910 = ~n39726 & n39908 ;
  assign n39911 = n39556 & n39910 ;
  assign n39912 = n39909 & ~n39911 ;
  assign n39913 = n2315 & n33436 ;
  assign n39914 = n2312 & n32293 ;
  assign n39915 = n2308 & ~n32442 ;
  assign n39916 = n39914 | n39915 ;
  assign n39917 = n39913 | n39916 ;
  assign n39918 = n2306 & ~n33441 ;
  assign n39919 = ~n32456 & n39918 ;
  assign n39920 = ( n2306 & n34271 ) | ( n2306 & n39919 ) | ( n34271 & n39919 ) ;
  assign n39921 = n39917 | n39920 ;
  assign n39922 = x26 | n39917 ;
  assign n39923 = n39920 | n39922 ;
  assign n39924 = ~x26 & n39922 ;
  assign n39925 = ( ~x26 & n39920 ) | ( ~x26 & n39924 ) | ( n39920 & n39924 ) ;
  assign n39926 = ( ~n39921 & n39923 ) | ( ~n39921 & n39925 ) | ( n39923 & n39925 ) ;
  assign n39998 = n39820 | n39837 ;
  assign n39999 = ( n39820 & n39822 ) | ( n39820 & n39998 ) | ( n39822 & n39998 ) ;
  assign n39973 = n39795 | n39814 ;
  assign n39974 = ( n39795 & n39798 ) | ( n39795 & n39973 ) | ( n39798 & n39973 ) ;
  assign n39927 = ( ~n39566 & n39788 ) | ( ~n39566 & n39791 ) | ( n39788 & n39791 ) ;
  assign n39928 = n1057 & ~n31309 ;
  assign n39929 = n1060 & n30212 ;
  assign n39930 = n1065 & ~n30186 ;
  assign n39931 = n39929 | n39930 ;
  assign n39932 = n39928 | n39931 ;
  assign n39933 = n1062 | n39928 ;
  assign n39934 = n39931 | n39933 ;
  assign n39935 = ( n31404 & n39932 ) | ( n31404 & n39934 ) | ( n39932 & n39934 ) ;
  assign n39936 = n4307 | n23827 ;
  assign n39937 = n861 | n39936 ;
  assign n39938 = n15250 | n39937 ;
  assign n39939 = n16937 | n39938 ;
  assign n39940 = n5128 | n29912 ;
  assign n39941 = n5971 | n39940 ;
  assign n39942 = n602 | n1166 ;
  assign n39943 = n39941 | n39942 ;
  assign n39944 = n162 | n222 ;
  assign n39945 = n245 | n324 ;
  assign n39946 = n39944 | n39945 ;
  assign n39947 = n39943 | n39946 ;
  assign n39948 = n39939 | n39947 ;
  assign n39949 = n39769 | n39948 ;
  assign n39950 = n39769 & n39948 ;
  assign n39951 = n39949 & ~n39950 ;
  assign n39952 = n29768 & n36083 ;
  assign n39953 = ~x17 & n29768 ;
  assign n39954 = n36083 & n39953 ;
  assign n39955 = x17 | n39953 ;
  assign n39956 = ( x17 & n36083 ) | ( x17 & n39955 ) | ( n36083 & n39955 ) ;
  assign n39957 = ( ~n39952 & n39954 ) | ( ~n39952 & n39956 ) | ( n39954 & n39956 ) ;
  assign n39958 = n39951 & ~n39957 ;
  assign n39959 = ~n39951 & n39957 ;
  assign n39960 = n39958 | n39959 ;
  assign n39961 = n39934 & ~n39960 ;
  assign n39962 = n39932 & ~n39960 ;
  assign n39963 = ( n31404 & n39961 ) | ( n31404 & n39962 ) | ( n39961 & n39962 ) ;
  assign n39964 = n39935 & ~n39963 ;
  assign n39965 = n39934 | n39960 ;
  assign n39966 = n39932 | n39960 ;
  assign n39967 = ( n31404 & n39965 ) | ( n31404 & n39966 ) | ( n39965 & n39966 ) ;
  assign n39968 = n39927 | n39967 ;
  assign n39969 = ( n39927 & ~n39964 ) | ( n39927 & n39968 ) | ( ~n39964 & n39968 ) ;
  assign n39970 = n39927 & n39967 ;
  assign n39971 = ~n39964 & n39970 ;
  assign n39972 = n39969 & ~n39971 ;
  assign n39975 = n39972 & n39974 ;
  assign n39976 = n39974 & ~n39975 ;
  assign n39977 = n1829 & n32306 ;
  assign n39978 = n1826 & ~n31323 ;
  assign n39979 = n1823 & n31295 ;
  assign n39980 = n39978 | n39979 ;
  assign n39981 = n39977 | n39980 ;
  assign n39982 = n1821 | n39977 ;
  assign n39983 = n39980 | n39982 ;
  assign n39984 = ( ~n32525 & n39981 ) | ( ~n32525 & n39983 ) | ( n39981 & n39983 ) ;
  assign n39985 = ~x29 & n39983 ;
  assign n39986 = ~x29 & n39981 ;
  assign n39987 = ( ~n32525 & n39985 ) | ( ~n32525 & n39986 ) | ( n39985 & n39986 ) ;
  assign n39988 = x29 | n39986 ;
  assign n39989 = x29 | n39985 ;
  assign n39990 = ( ~n32525 & n39988 ) | ( ~n32525 & n39989 ) | ( n39988 & n39989 ) ;
  assign n39991 = ( ~n39984 & n39987 ) | ( ~n39984 & n39990 ) | ( n39987 & n39990 ) ;
  assign n39992 = n39972 & ~n39974 ;
  assign n39993 = n39991 & n39992 ;
  assign n39994 = ( n39976 & n39991 ) | ( n39976 & n39993 ) | ( n39991 & n39993 ) ;
  assign n39995 = n39991 | n39992 ;
  assign n39996 = n39976 | n39995 ;
  assign n39997 = ~n39994 & n39996 ;
  assign n40000 = ( n39926 & n39997 ) | ( n39926 & ~n39999 ) | ( n39997 & ~n39999 ) ;
  assign n40001 = ( ~n39926 & n39999 ) | ( ~n39926 & n40000 ) | ( n39999 & n40000 ) ;
  assign n40002 = n2932 & n34656 ;
  assign n40003 = n2925 & ~n33423 ;
  assign n40004 = n2928 & n33526 ;
  assign n40005 = n40003 | n40004 ;
  assign n40006 = n40002 | n40005 ;
  assign n40007 = n2936 | n40002 ;
  assign n40008 = n40005 | n40007 ;
  assign n40009 = ( n34667 & n40006 ) | ( n34667 & n40008 ) | ( n40006 & n40008 ) ;
  assign n40010 = x23 & n40008 ;
  assign n40011 = x23 & n40006 ;
  assign n40012 = ( n34667 & n40010 ) | ( n34667 & n40011 ) | ( n40010 & n40011 ) ;
  assign n40013 = x23 & ~n40011 ;
  assign n40014 = x23 & ~n40010 ;
  assign n40015 = ( ~n34667 & n40013 ) | ( ~n34667 & n40014 ) | ( n40013 & n40014 ) ;
  assign n40016 = ( n40009 & ~n40012 ) | ( n40009 & n40015 ) | ( ~n40012 & n40015 ) ;
  assign n40017 = n40000 & n40016 ;
  assign n40018 = ~n39997 & n40016 ;
  assign n40019 = ( n40001 & n40017 ) | ( n40001 & n40018 ) | ( n40017 & n40018 ) ;
  assign n40020 = n40000 | n40016 ;
  assign n40021 = n39997 & ~n40016 ;
  assign n40022 = ( n40001 & n40020 ) | ( n40001 & ~n40021 ) | ( n40020 & ~n40021 ) ;
  assign n40023 = ~n40019 & n40022 ;
  assign n40024 = n39844 | n39859 ;
  assign n40025 = ( n39844 & n39845 ) | ( n39844 & n40024 ) | ( n39845 & n40024 ) ;
  assign n40026 = n40023 | n40025 ;
  assign n40027 = n40023 & n40025 ;
  assign n40028 = n40026 & ~n40027 ;
  assign n40044 = n39868 | n39883 ;
  assign n40045 = ( n39868 & n39869 ) | ( n39868 & n40044 ) | ( n39869 & n40044 ) ;
  assign n40029 = n3547 & n35746 ;
  assign n40030 = n3544 & n35021 ;
  assign n40031 = n3541 & ~n35371 ;
  assign n40032 = n40030 | n40031 ;
  assign n40033 = n40029 | n40032 ;
  assign n40034 = n3537 | n40029 ;
  assign n40035 = n40032 | n40034 ;
  assign n40036 = ( ~n35759 & n40033 ) | ( ~n35759 & n40035 ) | ( n40033 & n40035 ) ;
  assign n40037 = ~x20 & n40035 ;
  assign n40038 = ~x20 & n40033 ;
  assign n40039 = ( ~n35759 & n40037 ) | ( ~n35759 & n40038 ) | ( n40037 & n40038 ) ;
  assign n40040 = x20 | n40038 ;
  assign n40041 = x20 | n40037 ;
  assign n40042 = ( ~n35759 & n40040 ) | ( ~n35759 & n40041 ) | ( n40040 & n40041 ) ;
  assign n40043 = ( ~n40036 & n40039 ) | ( ~n40036 & n40042 ) | ( n40039 & n40042 ) ;
  assign n40046 = n40043 & n40045 ;
  assign n40047 = n40045 & ~n40046 ;
  assign n40048 = n40028 & n40043 ;
  assign n40049 = ~n40045 & n40048 ;
  assign n40050 = ( n40028 & n40047 ) | ( n40028 & n40049 ) | ( n40047 & n40049 ) ;
  assign n40051 = n40028 | n40043 ;
  assign n40052 = ( n40028 & ~n40045 ) | ( n40028 & n40051 ) | ( ~n40045 & n40051 ) ;
  assign n40053 = n40047 | n40052 ;
  assign n40054 = ~n40050 & n40053 ;
  assign n40055 = n39742 | n39888 ;
  assign n40056 = ( n39742 & n39746 ) | ( n39742 & n40055 ) | ( n39746 & n40055 ) ;
  assign n40057 = n40054 & n40056 ;
  assign n40058 = n40054 | n40056 ;
  assign n40059 = ~n40057 & n40058 ;
  assign n40060 = n39894 | n39900 ;
  assign n40061 = n39894 | n39901 ;
  assign n40062 = ( n39717 & n40060 ) | ( n39717 & n40061 ) | ( n40060 & n40061 ) ;
  assign n40063 = n40059 & n40062 ;
  assign n40064 = n39894 | n39895 ;
  assign n40065 = n40059 & n40064 ;
  assign n40066 = n39894 & n40059 ;
  assign n40067 = ( ~n39898 & n40065 ) | ( ~n39898 & n40066 ) | ( n40065 & n40066 ) ;
  assign n40068 = ( n39161 & n40063 ) | ( n39161 & n40067 ) | ( n40063 & n40067 ) ;
  assign n40069 = ( n39894 & ~n39898 ) | ( n39894 & n40064 ) | ( ~n39898 & n40064 ) ;
  assign n40070 = n40059 | n40069 ;
  assign n40071 = n40059 | n40062 ;
  assign n40072 = ( n39161 & n40070 ) | ( n39161 & n40071 ) | ( n40070 & n40071 ) ;
  assign n40073 = ~n40068 & n40072 ;
  assign n40074 = n39911 | n40073 ;
  assign n40075 = n39910 & n40073 ;
  assign n40076 = n39556 & n40075 ;
  assign n40077 = n40074 & ~n40076 ;
  assign n40211 = n40046 | n40049 ;
  assign n40212 = n40028 | n40046 ;
  assign n40213 = ( n40047 & n40211 ) | ( n40047 & n40212 ) | ( n40211 & n40212 ) ;
  assign n40078 = ~n39963 & n39969 ;
  assign n40103 = n1057 & ~n31323 ;
  assign n40104 = n1060 & ~n30186 ;
  assign n40105 = n1065 & ~n31309 ;
  assign n40106 = n40104 | n40105 ;
  assign n40107 = n40103 | n40106 ;
  assign n40108 = n1062 & n31384 ;
  assign n40109 = n1062 & n31386 ;
  assign n40110 = ( ~n30232 & n40108 ) | ( ~n30232 & n40109 ) | ( n40108 & n40109 ) ;
  assign n40111 = n40107 | n40110 ;
  assign n40112 = n1062 | n40107 ;
  assign n40113 = ( ~n31376 & n40111 ) | ( ~n31376 & n40112 ) | ( n40111 & n40112 ) ;
  assign n40079 = n9161 | n9168 ;
  assign n40080 = n951 | n23174 ;
  assign n40081 = n622 | n9163 ;
  assign n40082 = n40080 | n40081 ;
  assign n40083 = n817 | n40082 ;
  assign n40084 = n6960 | n40083 ;
  assign n40085 = n40079 | n40084 ;
  assign n40086 = ~n1607 & n37794 ;
  assign n40087 = ( ~n169 & n952 ) | ( ~n169 & n15243 ) | ( n952 & n15243 ) ;
  assign n40088 = n169 | n176 ;
  assign n40089 = n40087 | n40088 ;
  assign n40090 = n257 | n820 ;
  assign n40091 = n476 | n40090 ;
  assign n40092 = n40089 | n40091 ;
  assign n40093 = n40086 & ~n40092 ;
  assign n40094 = ~n40085 & n40093 ;
  assign n40095 = ( n39950 & n39951 ) | ( n39950 & n40094 ) | ( n39951 & n40094 ) ;
  assign n40096 = n39950 & n40094 ;
  assign n40097 = ( ~n39957 & n40095 ) | ( ~n39957 & n40096 ) | ( n40095 & n40096 ) ;
  assign n40098 = n39950 | n39951 ;
  assign n40099 = n40094 | n40098 ;
  assign n40100 = n39950 | n40094 ;
  assign n40101 = ( ~n39957 & n40099 ) | ( ~n39957 & n40100 ) | ( n40099 & n40100 ) ;
  assign n40102 = ~n40097 & n40101 ;
  assign n40114 = n40102 | n40113 ;
  assign n40115 = ~n40102 & n40113 ;
  assign n40116 = ( ~n40113 & n40114 ) | ( ~n40113 & n40115 ) | ( n40114 & n40115 ) ;
  assign n40117 = n40078 & ~n40116 ;
  assign n40118 = ~n40078 & n40116 ;
  assign n40119 = n40117 | n40118 ;
  assign n40120 = n1829 & n32293 ;
  assign n40121 = n1826 & n31295 ;
  assign n40122 = n1823 & n32306 ;
  assign n40123 = n40121 | n40122 ;
  assign n40124 = n40120 | n40123 ;
  assign n40125 = n32497 | n40124 ;
  assign n40126 = n32494 | n40125 ;
  assign n40127 = n1821 | n40120 ;
  assign n40128 = n40123 | n40127 ;
  assign n40129 = n40126 & n40128 ;
  assign n40130 = ~x29 & n40128 ;
  assign n40131 = n40126 & n40130 ;
  assign n40132 = x29 | n40130 ;
  assign n40133 = ( x29 & n40126 ) | ( x29 & n40132 ) | ( n40126 & n40132 ) ;
  assign n40134 = ( ~n40129 & n40131 ) | ( ~n40129 & n40133 ) | ( n40131 & n40133 ) ;
  assign n40135 = ~n40119 & n40134 ;
  assign n40136 = n40119 & ~n40134 ;
  assign n40137 = n40135 | n40136 ;
  assign n40138 = n39975 & ~n40137 ;
  assign n40139 = ( n39994 & ~n40137 ) | ( n39994 & n40138 ) | ( ~n40137 & n40138 ) ;
  assign n40140 = ~n39975 & n40137 ;
  assign n40141 = ~n39994 & n40140 ;
  assign n40142 = n40139 | n40141 ;
  assign n40143 = n2315 & ~n33423 ;
  assign n40144 = n2312 & ~n32442 ;
  assign n40145 = n2308 & n33436 ;
  assign n40146 = n40144 | n40145 ;
  assign n40147 = n40143 | n40146 ;
  assign n40148 = n2306 & n33575 ;
  assign n40149 = n2306 & ~n33577 ;
  assign n40150 = ( ~n32456 & n40148 ) | ( ~n32456 & n40149 ) | ( n40148 & n40149 ) ;
  assign n40151 = n40147 | n40150 ;
  assign n40152 = n2306 | n40147 ;
  assign n40153 = ( n33567 & n40151 ) | ( n33567 & n40152 ) | ( n40151 & n40152 ) ;
  assign n40154 = x26 | n40153 ;
  assign n40155 = ~x26 & n40153 ;
  assign n40156 = ( ~n40153 & n40154 ) | ( ~n40153 & n40155 ) | ( n40154 & n40155 ) ;
  assign n40157 = n40142 | n40156 ;
  assign n40158 = n40142 & ~n40156 ;
  assign n40159 = ( ~n40142 & n40157 ) | ( ~n40142 & n40158 ) | ( n40157 & n40158 ) ;
  assign n40160 = n39926 & n39999 ;
  assign n40161 = n39999 & ~n40160 ;
  assign n40162 = n39926 & ~n39999 ;
  assign n40163 = n39997 & ~n40162 ;
  assign n40164 = ~n40161 & n40163 ;
  assign n40165 = ( n39997 & n40160 ) | ( n39997 & ~n40164 ) | ( n40160 & ~n40164 ) ;
  assign n40166 = ~n40159 & n40165 ;
  assign n40167 = n40159 | n40166 ;
  assign n40168 = n40165 & ~n40166 ;
  assign n40169 = n40167 & ~n40168 ;
  assign n40170 = n2932 & n35021 ;
  assign n40171 = n2925 & n33526 ;
  assign n40172 = n2928 & n34656 ;
  assign n40173 = n40171 | n40172 ;
  assign n40174 = n40170 | n40173 ;
  assign n40175 = n2936 | n40170 ;
  assign n40176 = n40173 | n40175 ;
  assign n40177 = ( n35033 & n40174 ) | ( n35033 & n40176 ) | ( n40174 & n40176 ) ;
  assign n40178 = x23 & n40176 ;
  assign n40179 = x23 & n40174 ;
  assign n40180 = ( n35033 & n40178 ) | ( n35033 & n40179 ) | ( n40178 & n40179 ) ;
  assign n40181 = x23 & ~n40179 ;
  assign n40182 = x23 & ~n40178 ;
  assign n40183 = ( ~n35033 & n40181 ) | ( ~n35033 & n40182 ) | ( n40181 & n40182 ) ;
  assign n40184 = ( n40177 & ~n40180 ) | ( n40177 & n40183 ) | ( ~n40180 & n40183 ) ;
  assign n40185 = n40169 | n40184 ;
  assign n40186 = n40019 | n40023 ;
  assign n40187 = ( n40019 & n40025 ) | ( n40019 & n40186 ) | ( n40025 & n40186 ) ;
  assign n40188 = n40184 & n40187 ;
  assign n40189 = n40169 & n40188 ;
  assign n40190 = ( ~n40185 & n40187 ) | ( ~n40185 & n40189 ) | ( n40187 & n40189 ) ;
  assign n40191 = n40184 | n40187 ;
  assign n40192 = ( n40169 & n40187 ) | ( n40169 & n40191 ) | ( n40187 & n40191 ) ;
  assign n40193 = n40185 & ~n40192 ;
  assign n40194 = n40190 | n40193 ;
  assign n40195 = n3547 & n36083 ;
  assign n40196 = n3544 & ~n35371 ;
  assign n40197 = n3541 & n35746 ;
  assign n40198 = n40196 | n40197 ;
  assign n40199 = n40195 | n40198 ;
  assign n40200 = n3537 | n40195 ;
  assign n40201 = n40198 | n40200 ;
  assign n40202 = ( n36107 & n40199 ) | ( n36107 & n40201 ) | ( n40199 & n40201 ) ;
  assign n40203 = n40199 | n40201 ;
  assign n40204 = ( n36094 & n40202 ) | ( n36094 & n40203 ) | ( n40202 & n40203 ) ;
  assign n40205 = x20 & n40204 ;
  assign n40206 = x20 & ~n40204 ;
  assign n40207 = ( n40204 & ~n40205 ) | ( n40204 & n40206 ) | ( ~n40205 & n40206 ) ;
  assign n40208 = n40194 | n40207 ;
  assign n40209 = n40194 & ~n40207 ;
  assign n40210 = ( ~n40194 & n40208 ) | ( ~n40194 & n40209 ) | ( n40208 & n40209 ) ;
  assign n40214 = ~n40210 & n40213 ;
  assign n40215 = n40213 & ~n40214 ;
  assign n40216 = n40210 | n40213 ;
  assign n40217 = ~n40215 & n40216 ;
  assign n40218 = n40057 | n40059 ;
  assign n40219 = ~n40217 & n40218 ;
  assign n40220 = n40057 & ~n40217 ;
  assign n40221 = ( n40062 & n40219 ) | ( n40062 & n40220 ) | ( n40219 & n40220 ) ;
  assign n40222 = n40057 | n40065 ;
  assign n40223 = ~n40217 & n40222 ;
  assign n40224 = n40057 | n40066 ;
  assign n40225 = ~n40217 & n40224 ;
  assign n40226 = ( ~n39898 & n40223 ) | ( ~n39898 & n40225 ) | ( n40223 & n40225 ) ;
  assign n40227 = ( n39161 & n40221 ) | ( n39161 & n40226 ) | ( n40221 & n40226 ) ;
  assign n40228 = ( n40057 & n40062 ) | ( n40057 & n40218 ) | ( n40062 & n40218 ) ;
  assign n40229 = n40217 & ~n40228 ;
  assign n40230 = ( ~n39898 & n40222 ) | ( ~n39898 & n40224 ) | ( n40222 & n40224 ) ;
  assign n40231 = n40217 & ~n40230 ;
  assign n40232 = ( ~n39161 & n40229 ) | ( ~n39161 & n40231 ) | ( n40229 & n40231 ) ;
  assign n40233 = n40227 | n40232 ;
  assign n40234 = n40076 | n40233 ;
  assign n40235 = n40076 & n40233 ;
  assign n40236 = n40234 & ~n40235 ;
  assign n40237 = n30847 & n36083 ;
  assign n40238 = n3544 & n35746 ;
  assign n40239 = n40237 | n40238 ;
  assign n40240 = n3537 | n40239 ;
  assign n40241 = ( n36103 & n40239 ) | ( n36103 & n40240 ) | ( n40239 & n40240 ) ;
  assign n40242 = ( n36105 & n40239 ) | ( n36105 & n40240 ) | ( n40239 & n40240 ) ;
  assign n40243 = ( n32456 & n40241 ) | ( n32456 & n40242 ) | ( n40241 & n40242 ) ;
  assign n40244 = x20 & n40243 ;
  assign n40245 = x20 & ~n40243 ;
  assign n40246 = ( n40243 & ~n40244 ) | ( n40243 & n40245 ) | ( ~n40244 & n40245 ) ;
  assign n40247 = n40166 | n40184 ;
  assign n40248 = n40246 & n40247 ;
  assign n40249 = n40166 & n40246 ;
  assign n40250 = ( ~n40169 & n40248 ) | ( ~n40169 & n40249 ) | ( n40248 & n40249 ) ;
  assign n40251 = n40246 | n40247 ;
  assign n40252 = n40166 | n40246 ;
  assign n40253 = ( ~n40169 & n40251 ) | ( ~n40169 & n40252 ) | ( n40251 & n40252 ) ;
  assign n40254 = ~n40250 & n40253 ;
  assign n40255 = n1057 & n31295 ;
  assign n40256 = n1060 & ~n31309 ;
  assign n40257 = n1065 & ~n31323 ;
  assign n40258 = n40256 | n40257 ;
  assign n40259 = n40255 | n40258 ;
  assign n40260 = n1062 | n40255 ;
  assign n40261 = n40258 | n40260 ;
  assign n40262 = ( n31355 & n40259 ) | ( n31355 & n40261 ) | ( n40259 & n40261 ) ;
  assign n40263 = n29918 | n39753 ;
  assign n40264 = n15505 & ~n40263 ;
  assign n40265 = ~n15501 & n40264 ;
  assign n40266 = ~n16923 & n40265 ;
  assign n40267 = ~n4043 & n40266 ;
  assign n40268 = n617 | n878 ;
  assign n40269 = n3995 | n40268 ;
  assign n40270 = n40267 & ~n40269 ;
  assign n40271 = n5978 | n36702 ;
  assign n40272 = n40270 & ~n40271 ;
  assign n40273 = n387 | n638 ;
  assign n40274 = n71 | n886 ;
  assign n40275 = n40273 | n40274 ;
  assign n40276 = n40272 & ~n40275 ;
  assign n40277 = ~n40094 & n40276 ;
  assign n40278 = n40094 & ~n40276 ;
  assign n40279 = n40255 & ~n40278 ;
  assign n40280 = ( n40258 & ~n40278 ) | ( n40258 & n40279 ) | ( ~n40278 & n40279 ) ;
  assign n40281 = ~n40277 & n40280 ;
  assign n40282 = n40277 | n40278 ;
  assign n40283 = n40261 & ~n40282 ;
  assign n40284 = ( n31355 & n40281 ) | ( n31355 & n40283 ) | ( n40281 & n40283 ) ;
  assign n40285 = n40262 & ~n40284 ;
  assign n40286 = n40102 & n40107 ;
  assign n40287 = ( n40102 & n40110 ) | ( n40102 & n40286 ) | ( n40110 & n40286 ) ;
  assign n40288 = ( n1062 & n40102 ) | ( n1062 & n40286 ) | ( n40102 & n40286 ) ;
  assign n40289 = ( ~n31376 & n40287 ) | ( ~n31376 & n40288 ) | ( n40287 & n40288 ) ;
  assign n40290 = n40097 | n40289 ;
  assign n40291 = n40277 & ~n40278 ;
  assign n40292 = ( n40278 & n40280 ) | ( n40278 & ~n40291 ) | ( n40280 & ~n40291 ) ;
  assign n40293 = n40277 | n40292 ;
  assign n40294 = ~n40278 & n40282 ;
  assign n40295 = ( n40261 & n40278 ) | ( n40261 & ~n40294 ) | ( n40278 & ~n40294 ) ;
  assign n40296 = n40277 | n40295 ;
  assign n40297 = ( n31355 & n40293 ) | ( n31355 & n40296 ) | ( n40293 & n40296 ) ;
  assign n40298 = n40290 & ~n40297 ;
  assign n40299 = ( n40285 & n40290 ) | ( n40285 & n40298 ) | ( n40290 & n40298 ) ;
  assign n40300 = ~n40290 & n40297 ;
  assign n40301 = ~n40285 & n40300 ;
  assign n40302 = n40299 | n40301 ;
  assign n40303 = n40118 | n40134 ;
  assign n40304 = ( n40118 & ~n40119 ) | ( n40118 & n40303 ) | ( ~n40119 & n40303 ) ;
  assign n40305 = n40302 & ~n40304 ;
  assign n40306 = ~n40302 & n40304 ;
  assign n40307 = n40305 | n40306 ;
  assign n40308 = n1829 & ~n32442 ;
  assign n40309 = n1826 & n32306 ;
  assign n40310 = n1823 & n32293 ;
  assign n40311 = n40309 | n40310 ;
  assign n40312 = n40308 | n40311 ;
  assign n40313 = n1821 | n40308 ;
  assign n40314 = n40311 | n40313 ;
  assign n40315 = ( ~n32458 & n40312 ) | ( ~n32458 & n40314 ) | ( n40312 & n40314 ) ;
  assign n40316 = ~x29 & n40314 ;
  assign n40317 = ~x29 & n40312 ;
  assign n40318 = ( ~n32458 & n40316 ) | ( ~n32458 & n40317 ) | ( n40316 & n40317 ) ;
  assign n40319 = x29 | n40317 ;
  assign n40320 = x29 | n40316 ;
  assign n40321 = ( ~n32458 & n40319 ) | ( ~n32458 & n40320 ) | ( n40319 & n40320 ) ;
  assign n40322 = ( ~n40315 & n40318 ) | ( ~n40315 & n40321 ) | ( n40318 & n40321 ) ;
  assign n40323 = ~n40307 & n40322 ;
  assign n40324 = n40307 | n40323 ;
  assign n40325 = n2315 & n33526 ;
  assign n40326 = n2312 & n33436 ;
  assign n40327 = n2308 & ~n33423 ;
  assign n40328 = n40326 | n40327 ;
  assign n40329 = n40325 | n40328 ;
  assign n40330 = n2306 & n33545 ;
  assign n40331 = n2306 & ~n33548 ;
  assign n40332 = ( ~n32456 & n40330 ) | ( ~n32456 & n40331 ) | ( n40330 & n40331 ) ;
  assign n40333 = n40329 | n40332 ;
  assign n40334 = n2306 | n40329 ;
  assign n40335 = ( n33536 & n40333 ) | ( n33536 & n40334 ) | ( n40333 & n40334 ) ;
  assign n40336 = x26 | n40335 ;
  assign n40337 = ~x26 & n40335 ;
  assign n40338 = ( ~n40335 & n40336 ) | ( ~n40335 & n40337 ) | ( n40336 & n40337 ) ;
  assign n40339 = n40307 & n40322 ;
  assign n40340 = n40338 & n40339 ;
  assign n40341 = ( ~n40324 & n40338 ) | ( ~n40324 & n40340 ) | ( n40338 & n40340 ) ;
  assign n40342 = n40338 | n40339 ;
  assign n40343 = n40324 & ~n40342 ;
  assign n40344 = n40341 | n40343 ;
  assign n40345 = n40139 | n40156 ;
  assign n40346 = ( n40139 & ~n40142 ) | ( n40139 & n40345 ) | ( ~n40142 & n40345 ) ;
  assign n40347 = n40344 & ~n40346 ;
  assign n40348 = ~n40344 & n40346 ;
  assign n40349 = n40347 | n40348 ;
  assign n40350 = n2932 & ~n35371 ;
  assign n40351 = n2925 & n34656 ;
  assign n40352 = n2928 & n35021 ;
  assign n40353 = n40351 | n40352 ;
  assign n40354 = n40350 | n40353 ;
  assign n40355 = n2936 & ~n35392 ;
  assign n40356 = n2936 & ~n35395 ;
  assign n40357 = ( ~n32456 & n40355 ) | ( ~n32456 & n40356 ) | ( n40355 & n40356 ) ;
  assign n40358 = n40354 | n40357 ;
  assign n40359 = n2936 | n40354 ;
  assign n40360 = ( n35381 & n40358 ) | ( n35381 & n40359 ) | ( n40358 & n40359 ) ;
  assign n40361 = x23 | n40360 ;
  assign n40362 = ~x23 & n40360 ;
  assign n40363 = ( ~n40360 & n40361 ) | ( ~n40360 & n40362 ) | ( n40361 & n40362 ) ;
  assign n40364 = n40349 & n40363 ;
  assign n40365 = n40346 | n40363 ;
  assign n40366 = ( ~n40344 & n40363 ) | ( ~n40344 & n40365 ) | ( n40363 & n40365 ) ;
  assign n40367 = n40347 | n40366 ;
  assign n40368 = ~n40364 & n40367 ;
  assign n40369 = n40254 & ~n40368 ;
  assign n40370 = n40254 & ~n40369 ;
  assign n40371 = n40254 | n40368 ;
  assign n40372 = ~n40370 & n40371 ;
  assign n40373 = n40190 | n40207 ;
  assign n40374 = ( n40190 & ~n40194 ) | ( n40190 & n40373 ) | ( ~n40194 & n40373 ) ;
  assign n40375 = n40372 & ~n40374 ;
  assign n40376 = ~n40372 & n40374 ;
  assign n40377 = n40375 | n40376 ;
  assign n40378 = n40214 | n40223 ;
  assign n40379 = n40214 | n40225 ;
  assign n40380 = ( ~n39898 & n40378 ) | ( ~n39898 & n40379 ) | ( n40378 & n40379 ) ;
  assign n40381 = ~n40377 & n40380 ;
  assign n40382 = n40214 | n40219 ;
  assign n40383 = ~n40377 & n40382 ;
  assign n40384 = n40214 | n40220 ;
  assign n40385 = ~n40377 & n40384 ;
  assign n40386 = ( n40062 & n40383 ) | ( n40062 & n40385 ) | ( n40383 & n40385 ) ;
  assign n40387 = ( n39161 & n40381 ) | ( n39161 & n40386 ) | ( n40381 & n40386 ) ;
  assign n40388 = ( n40062 & n40382 ) | ( n40062 & n40384 ) | ( n40382 & n40384 ) ;
  assign n40389 = n40377 & ~n40388 ;
  assign n40390 = n40377 & ~n40380 ;
  assign n40391 = ( ~n39161 & n40389 ) | ( ~n39161 & n40390 ) | ( n40389 & n40390 ) ;
  assign n40392 = n40387 | n40391 ;
  assign n40393 = n40073 & ~n40233 ;
  assign n40394 = n39910 & n40393 ;
  assign n40395 = n39555 & n40394 ;
  assign n40396 = n38738 & n40395 ;
  assign n40397 = ~n40392 & n40396 ;
  assign n40398 = n40392 & ~n40396 ;
  assign n40399 = n40397 | n40398 ;
  assign n40400 = n40323 | n40341 ;
  assign n40401 = n297 | n434 ;
  assign n40402 = n280 | n40401 ;
  assign n40403 = n12276 & ~n12277 ;
  assign n40404 = n988 | n6871 ;
  assign n40405 = n5923 | n40404 ;
  assign n40406 = n24261 | n40405 ;
  assign n40407 = ( n14422 & n40403 ) | ( n14422 & ~n40406 ) | ( n40403 & ~n40406 ) ;
  assign n40408 = ~n40403 & n40406 ;
  assign n40409 = ( n14413 & n40407 ) | ( n14413 & ~n40408 ) | ( n40407 & ~n40408 ) ;
  assign n40410 = ~n14423 & n40409 ;
  assign n40411 = n784 | n5154 ;
  assign n40412 = n201 | n40411 ;
  assign n40413 = n2192 | n5092 ;
  assign n40414 = n608 | n40413 ;
  assign n40415 = n209 | n40414 ;
  assign n40416 = n40412 | n40415 ;
  assign n40417 = n331 | n40416 ;
  assign n40418 = n4282 | n40417 ;
  assign n40419 = n40410 & ~n40418 ;
  assign n40420 = ~n40402 & n40419 ;
  assign n40421 = n40094 & n40420 ;
  assign n40422 = n40094 | n40420 ;
  assign n40423 = ~n40421 & n40422 ;
  assign n40424 = n30849 & n36083 ;
  assign n40425 = ~x20 & n30849 ;
  assign n40426 = n36083 & n40425 ;
  assign n40427 = x20 | n40425 ;
  assign n40428 = ( x20 & n36083 ) | ( x20 & n40427 ) | ( n36083 & n40427 ) ;
  assign n40429 = ( ~n40424 & n40426 ) | ( ~n40424 & n40428 ) | ( n40426 & n40428 ) ;
  assign n40430 = n40423 & ~n40429 ;
  assign n40431 = ~n40423 & n40429 ;
  assign n40432 = n40430 | n40431 ;
  assign n40433 = n40292 & ~n40432 ;
  assign n40434 = n40295 & ~n40432 ;
  assign n40435 = ( n31355 & n40433 ) | ( n31355 & n40434 ) | ( n40433 & n40434 ) ;
  assign n40436 = ~n40292 & n40432 ;
  assign n40437 = ~n40295 & n40432 ;
  assign n40438 = ( ~n31355 & n40436 ) | ( ~n31355 & n40437 ) | ( n40436 & n40437 ) ;
  assign n40439 = n40435 | n40438 ;
  assign n40440 = n1057 & n32306 ;
  assign n40441 = n1060 & ~n31323 ;
  assign n40442 = n1065 & n31295 ;
  assign n40443 = n40441 | n40442 ;
  assign n40444 = n40440 | n40443 ;
  assign n40445 = n1062 | n40440 ;
  assign n40446 = n40443 | n40445 ;
  assign n40447 = ( ~n32525 & n40444 ) | ( ~n32525 & n40446 ) | ( n40444 & n40446 ) ;
  assign n40448 = n40439 & n40447 ;
  assign n40449 = n40439 | n40447 ;
  assign n40450 = ~n40448 & n40449 ;
  assign n40451 = ( ~n40299 & n40302 ) | ( ~n40299 & n40450 ) | ( n40302 & n40450 ) ;
  assign n40452 = n40299 & ~n40450 ;
  assign n40453 = ( n40304 & ~n40451 ) | ( n40304 & n40452 ) | ( ~n40451 & n40452 ) ;
  assign n40454 = ~n40299 & n40302 ;
  assign n40455 = n40450 & n40454 ;
  assign n40456 = ~n40299 & n40450 ;
  assign n40457 = ( ~n40304 & n40455 ) | ( ~n40304 & n40456 ) | ( n40455 & n40456 ) ;
  assign n40458 = n40453 | n40457 ;
  assign n40459 = n1829 & n33436 ;
  assign n40460 = n1826 & n32293 ;
  assign n40461 = n1823 & ~n32442 ;
  assign n40462 = n40460 | n40461 ;
  assign n40463 = n40459 | n40462 ;
  assign n40464 = n1821 & ~n33441 ;
  assign n40465 = ~n32456 & n40464 ;
  assign n40466 = ( n1821 & n34271 ) | ( n1821 & n40465 ) | ( n34271 & n40465 ) ;
  assign n40467 = n40463 | n40466 ;
  assign n40468 = x29 | n40463 ;
  assign n40469 = n40466 | n40468 ;
  assign n40470 = ~x29 & n40468 ;
  assign n40471 = ( ~x29 & n40466 ) | ( ~x29 & n40470 ) | ( n40466 & n40470 ) ;
  assign n40472 = ( ~n40467 & n40469 ) | ( ~n40467 & n40471 ) | ( n40469 & n40471 ) ;
  assign n40473 = ~n40458 & n40472 ;
  assign n40474 = n40458 | n40473 ;
  assign n40475 = n2315 & n34656 ;
  assign n40476 = n2312 & ~n33423 ;
  assign n40477 = n2308 & n33526 ;
  assign n40478 = n40476 | n40477 ;
  assign n40479 = n40475 | n40478 ;
  assign n40480 = n2306 | n40475 ;
  assign n40481 = n40478 | n40480 ;
  assign n40482 = ( n34667 & n40479 ) | ( n34667 & n40481 ) | ( n40479 & n40481 ) ;
  assign n40483 = x26 & n40481 ;
  assign n40484 = x26 & n40479 ;
  assign n40485 = ( n34667 & n40483 ) | ( n34667 & n40484 ) | ( n40483 & n40484 ) ;
  assign n40486 = x26 & ~n40484 ;
  assign n40487 = x26 & ~n40483 ;
  assign n40488 = ( ~n34667 & n40486 ) | ( ~n34667 & n40487 ) | ( n40486 & n40487 ) ;
  assign n40489 = ( n40482 & ~n40485 ) | ( n40482 & n40488 ) | ( ~n40485 & n40488 ) ;
  assign n40490 = n40458 & n40472 ;
  assign n40491 = n40489 & n40490 ;
  assign n40492 = ( ~n40474 & n40489 ) | ( ~n40474 & n40491 ) | ( n40489 & n40491 ) ;
  assign n40493 = n40489 | n40490 ;
  assign n40494 = n40474 & ~n40493 ;
  assign n40495 = n40492 | n40494 ;
  assign n40496 = ~n40400 & n40495 ;
  assign n40497 = n40400 & ~n40495 ;
  assign n40498 = n40496 | n40497 ;
  assign n40514 = ( n40348 & ~n40349 ) | ( n40348 & n40366 ) | ( ~n40349 & n40366 ) ;
  assign n40499 = n2932 & n35746 ;
  assign n40500 = n2925 & n35021 ;
  assign n40501 = n2928 & ~n35371 ;
  assign n40502 = n40500 | n40501 ;
  assign n40503 = n40499 | n40502 ;
  assign n40504 = n2936 | n40499 ;
  assign n40505 = n40502 | n40504 ;
  assign n40506 = ( ~n35759 & n40503 ) | ( ~n35759 & n40505 ) | ( n40503 & n40505 ) ;
  assign n40507 = ~x23 & n40505 ;
  assign n40508 = ~x23 & n40503 ;
  assign n40509 = ( ~n35759 & n40507 ) | ( ~n35759 & n40508 ) | ( n40507 & n40508 ) ;
  assign n40510 = x23 | n40508 ;
  assign n40511 = x23 | n40507 ;
  assign n40512 = ( ~n35759 & n40510 ) | ( ~n35759 & n40511 ) | ( n40510 & n40511 ) ;
  assign n40513 = ( ~n40506 & n40509 ) | ( ~n40506 & n40512 ) | ( n40509 & n40512 ) ;
  assign n40515 = n40513 & n40514 ;
  assign n40516 = n40514 & ~n40515 ;
  assign n40517 = ~n40498 & n40513 ;
  assign n40518 = ~n40514 & n40517 ;
  assign n40519 = ( ~n40498 & n40516 ) | ( ~n40498 & n40518 ) | ( n40516 & n40518 ) ;
  assign n40520 = n40498 & ~n40513 ;
  assign n40521 = ( n40498 & n40514 ) | ( n40498 & n40520 ) | ( n40514 & n40520 ) ;
  assign n40522 = ~n40516 & n40521 ;
  assign n40523 = n40519 | n40522 ;
  assign n40524 = ~n40250 & n40368 ;
  assign n40525 = ( n40250 & n40254 ) | ( n40250 & ~n40524 ) | ( n40254 & ~n40524 ) ;
  assign n40526 = ~n40523 & n40525 ;
  assign n40527 = n40523 & ~n40525 ;
  assign n40528 = n40526 | n40527 ;
  assign n40529 = n40376 | n40383 ;
  assign n40530 = ~n40528 & n40529 ;
  assign n40531 = n40376 | n40385 ;
  assign n40532 = ~n40528 & n40531 ;
  assign n40533 = ( n40062 & n40530 ) | ( n40062 & n40532 ) | ( n40530 & n40532 ) ;
  assign n40534 = ~n40376 & n40377 ;
  assign n40535 = n40528 | n40534 ;
  assign n40536 = n40376 & ~n40528 ;
  assign n40537 = ( n40380 & ~n40535 ) | ( n40380 & n40536 ) | ( ~n40535 & n40536 ) ;
  assign n40538 = ( n39161 & n40533 ) | ( n39161 & n40537 ) | ( n40533 & n40537 ) ;
  assign n40539 = ( n40376 & n40380 ) | ( n40376 & ~n40534 ) | ( n40380 & ~n40534 ) ;
  assign n40540 = n40528 & ~n40539 ;
  assign n40541 = ( n40062 & n40529 ) | ( n40062 & n40531 ) | ( n40529 & n40531 ) ;
  assign n40542 = n40528 & ~n40541 ;
  assign n40543 = ( ~n39161 & n40540 ) | ( ~n39161 & n40542 ) | ( n40540 & n40542 ) ;
  assign n40544 = n40538 | n40543 ;
  assign n40545 = ~n40397 & n40544 ;
  assign n40546 = n40392 | n40544 ;
  assign n40547 = n40396 & ~n40546 ;
  assign n40548 = n40545 | n40547 ;
  assign n40655 = n40515 | n40518 ;
  assign n40656 = n40498 & ~n40515 ;
  assign n40657 = ( n40516 & n40655 ) | ( n40516 & ~n40656 ) | ( n40655 & ~n40656 ) ;
  assign n40549 = n1057 & n32293 ;
  assign n40550 = n1060 & n31295 ;
  assign n40551 = n1065 & n32306 ;
  assign n40552 = n40550 | n40551 ;
  assign n40553 = n40549 | n40552 ;
  assign n40554 = n1062 & n32497 ;
  assign n40555 = ( n1062 & n32494 ) | ( n1062 & n40554 ) | ( n32494 & n40554 ) ;
  assign n40556 = n40553 | n40555 ;
  assign n40557 = n2835 | n9150 ;
  assign n40558 = n3465 | n40557 ;
  assign n40559 = n3453 | n40558 ;
  assign n40560 = n2666 | n40559 ;
  assign n40561 = ( ~n16936 & n25788 ) | ( ~n16936 & n40560 ) | ( n25788 & n40560 ) ;
  assign n40562 = n25788 & n40560 ;
  assign n40563 = ( ~n16929 & n40561 ) | ( ~n16929 & n40562 ) | ( n40561 & n40562 ) ;
  assign n40564 = n16937 | n40563 ;
  assign n40565 = n10809 | n18116 ;
  assign n40566 = n2818 | n40565 ;
  assign n40567 = n202 | n387 ;
  assign n40568 = n1785 | n40567 ;
  assign n40569 = n131 | n223 ;
  assign n40570 = n390 | n40569 ;
  assign n40571 = n40568 | n40570 ;
  assign n40572 = n40566 | n40571 ;
  assign n40573 = n40564 | n40572 ;
  assign n40574 = ( n40422 & ~n40423 ) | ( n40422 & n40573 ) | ( ~n40423 & n40573 ) ;
  assign n40575 = n40422 | n40573 ;
  assign n40576 = ( n40429 & n40574 ) | ( n40429 & n40575 ) | ( n40574 & n40575 ) ;
  assign n40577 = n40422 & ~n40423 ;
  assign n40578 = n40573 & n40577 ;
  assign n40579 = n40422 & n40573 ;
  assign n40580 = ( n40429 & n40578 ) | ( n40429 & n40579 ) | ( n40578 & n40579 ) ;
  assign n40581 = n40576 & ~n40580 ;
  assign n40582 = n40553 | n40581 ;
  assign n40583 = n40555 | n40582 ;
  assign n40584 = ~n40581 & n40582 ;
  assign n40585 = ( n40555 & ~n40581 ) | ( n40555 & n40584 ) | ( ~n40581 & n40584 ) ;
  assign n40586 = ( ~n40556 & n40583 ) | ( ~n40556 & n40585 ) | ( n40583 & n40585 ) ;
  assign n40587 = n40435 | n40447 ;
  assign n40588 = ( n40435 & ~n40439 ) | ( n40435 & n40587 ) | ( ~n40439 & n40587 ) ;
  assign n40589 = n40586 | n40588 ;
  assign n40590 = n40586 & n40588 ;
  assign n40591 = n40589 & ~n40590 ;
  assign n40592 = n1826 & ~n32442 ;
  assign n40593 = n1823 & n33436 ;
  assign n40594 = n40592 | n40593 ;
  assign n40595 = n1829 & ~n33423 ;
  assign n40596 = n1821 | n40595 ;
  assign n40597 = n40594 | n40596 ;
  assign n40598 = n40594 | n40595 ;
  assign n40599 = n33575 | n40598 ;
  assign n40600 = n33577 & ~n40598 ;
  assign n40601 = ( n32456 & ~n40599 ) | ( n32456 & n40600 ) | ( ~n40599 & n40600 ) ;
  assign n40602 = n40597 & ~n40601 ;
  assign n40603 = ( n33567 & n40597 ) | ( n33567 & n40602 ) | ( n40597 & n40602 ) ;
  assign n40604 = x29 & n40603 ;
  assign n40605 = x29 & ~n40603 ;
  assign n40606 = ( n40603 & ~n40604 ) | ( n40603 & n40605 ) | ( ~n40604 & n40605 ) ;
  assign n40607 = n40591 & n40606 ;
  assign n40608 = n40591 | n40606 ;
  assign n40609 = ~n40607 & n40608 ;
  assign n40610 = n40453 | n40472 ;
  assign n40611 = ( n40453 & ~n40458 ) | ( n40453 & n40610 ) | ( ~n40458 & n40610 ) ;
  assign n40612 = n40609 & n40611 ;
  assign n40613 = n40609 | n40611 ;
  assign n40614 = ~n40612 & n40613 ;
  assign n40615 = n2315 & n35021 ;
  assign n40616 = n2312 & n33526 ;
  assign n40617 = n2308 & n34656 ;
  assign n40618 = n40616 | n40617 ;
  assign n40619 = n40615 | n40618 ;
  assign n40620 = n2306 | n40615 ;
  assign n40621 = n40618 | n40620 ;
  assign n40622 = ( n35033 & n40619 ) | ( n35033 & n40621 ) | ( n40619 & n40621 ) ;
  assign n40623 = x26 & n40621 ;
  assign n40624 = x26 & n40619 ;
  assign n40625 = ( n35033 & n40623 ) | ( n35033 & n40624 ) | ( n40623 & n40624 ) ;
  assign n40626 = x26 & ~n40624 ;
  assign n40627 = x26 & ~n40623 ;
  assign n40628 = ( ~n35033 & n40626 ) | ( ~n35033 & n40627 ) | ( n40626 & n40627 ) ;
  assign n40629 = ( n40622 & ~n40625 ) | ( n40622 & n40628 ) | ( ~n40625 & n40628 ) ;
  assign n40630 = n40614 & ~n40629 ;
  assign n40631 = n40614 | n40629 ;
  assign n40632 = ( ~n40614 & n40630 ) | ( ~n40614 & n40631 ) | ( n40630 & n40631 ) ;
  assign n40633 = n40492 | n40497 ;
  assign n40634 = n40632 | n40633 ;
  assign n40635 = n40632 & n40633 ;
  assign n40636 = n40634 & ~n40635 ;
  assign n40637 = n2932 & n36083 ;
  assign n40638 = n2925 & ~n35371 ;
  assign n40639 = n2928 & n35746 ;
  assign n40640 = n40638 | n40639 ;
  assign n40641 = n40637 | n40640 ;
  assign n40642 = n2936 | n40637 ;
  assign n40643 = n40640 | n40642 ;
  assign n40644 = ( n36107 & n40641 ) | ( n36107 & n40643 ) | ( n40641 & n40643 ) ;
  assign n40645 = n40641 | n40643 ;
  assign n40646 = ( n36094 & n40644 ) | ( n36094 & n40645 ) | ( n40644 & n40645 ) ;
  assign n40647 = x23 & n40646 ;
  assign n40648 = x23 & ~n40646 ;
  assign n40649 = ( n40646 & ~n40647 ) | ( n40646 & n40648 ) | ( ~n40647 & n40648 ) ;
  assign n40650 = ~n40636 & n40649 ;
  assign n40651 = n40632 | n40649 ;
  assign n40652 = ( n40633 & n40649 ) | ( n40633 & n40651 ) | ( n40649 & n40651 ) ;
  assign n40653 = n40634 & ~n40652 ;
  assign n40654 = n40650 | n40653 ;
  assign n40658 = n40654 & n40657 ;
  assign n40659 = n40657 & ~n40658 ;
  assign n40660 = n40654 & ~n40657 ;
  assign n40661 = n40659 | n40660 ;
  assign n40662 = n40526 | n40530 ;
  assign n40663 = n40526 | n40532 ;
  assign n40664 = ( n40062 & n40662 ) | ( n40062 & n40663 ) | ( n40662 & n40663 ) ;
  assign n40665 = n40661 & n40664 ;
  assign n40666 = ~n40526 & n40535 ;
  assign n40667 = n40661 & ~n40666 ;
  assign n40668 = n40526 | n40536 ;
  assign n40669 = n40661 & n40668 ;
  assign n40670 = ( n40380 & n40667 ) | ( n40380 & n40669 ) | ( n40667 & n40669 ) ;
  assign n40671 = ( n39161 & n40665 ) | ( n39161 & n40670 ) | ( n40665 & n40670 ) ;
  assign n40672 = ( n40380 & ~n40666 ) | ( n40380 & n40668 ) | ( ~n40666 & n40668 ) ;
  assign n40673 = n40661 | n40672 ;
  assign n40674 = n40661 | n40664 ;
  assign n40675 = ( n39161 & n40673 ) | ( n39161 & n40674 ) | ( n40673 & n40674 ) ;
  assign n40676 = ~n40671 & n40675 ;
  assign n40677 = n40547 & ~n40676 ;
  assign n40678 = ~n40547 & n40676 ;
  assign n40679 = n40677 | n40678 ;
  assign n40680 = n32066 & n36083 ;
  assign n40681 = n2925 & n35746 ;
  assign n40682 = n40680 | n40681 ;
  assign n40683 = n2936 | n40682 ;
  assign n40684 = ( n36103 & n40682 ) | ( n36103 & n40683 ) | ( n40682 & n40683 ) ;
  assign n40685 = ( n36105 & n40682 ) | ( n36105 & n40683 ) | ( n40682 & n40683 ) ;
  assign n40686 = ( n32456 & n40684 ) | ( n32456 & n40685 ) | ( n40684 & n40685 ) ;
  assign n40687 = x23 & n40686 ;
  assign n40688 = x23 & ~n40686 ;
  assign n40689 = ( n40686 & ~n40687 ) | ( n40686 & n40688 ) | ( ~n40687 & n40688 ) ;
  assign n40690 = n40612 | n40629 ;
  assign n40691 = ( n40612 & n40614 ) | ( n40612 & n40690 ) | ( n40614 & n40690 ) ;
  assign n40692 = n40689 & n40691 ;
  assign n40693 = n40689 | n40691 ;
  assign n40694 = ~n40692 & n40693 ;
  assign n40695 = n40576 & ~n40581 ;
  assign n40696 = ~n40553 & n40576 ;
  assign n40697 = ( n40576 & ~n40581 ) | ( n40576 & n40696 ) | ( ~n40581 & n40696 ) ;
  assign n40698 = ( ~n40555 & n40695 ) | ( ~n40555 & n40697 ) | ( n40695 & n40697 ) ;
  assign n40699 = n607 | n696 ;
  assign n40700 = n4369 | n7024 ;
  assign n40701 = n23176 | n40700 ;
  assign n40702 = n17690 | n40701 ;
  assign n40703 = ( ~n15599 & n32341 ) | ( ~n15599 & n40702 ) | ( n32341 & n40702 ) ;
  assign n40704 = n32341 & n40702 ;
  assign n40705 = ( ~n15591 & n40703 ) | ( ~n15591 & n40704 ) | ( n40703 & n40704 ) ;
  assign n40706 = n15600 | n40705 ;
  assign n40707 = n617 | n37810 ;
  assign n40708 = n4197 | n40707 ;
  assign n40709 = n37809 | n40708 ;
  assign n40710 = n274 | n1785 ;
  assign n40711 = n40709 | n40710 ;
  assign n40712 = n22490 | n22508 ;
  assign n40713 = n22486 & ~n40712 ;
  assign n40714 = n163 | n511 ;
  assign n40715 = n40713 & ~n40714 ;
  assign n40716 = ~n40711 & n40715 ;
  assign n40717 = ~n40706 & n40716 ;
  assign n40718 = ~n40699 & n40717 ;
  assign n40719 = n40573 | n40718 ;
  assign n40720 = n40573 & n40718 ;
  assign n40721 = n40576 | n40720 ;
  assign n40722 = ( ~n40581 & n40720 ) | ( ~n40581 & n40721 ) | ( n40720 & n40721 ) ;
  assign n40723 = n40719 & ~n40722 ;
  assign n40724 = n40719 & ~n40720 ;
  assign n40725 = ~n40697 & n40724 ;
  assign n40726 = ( n40555 & n40723 ) | ( n40555 & n40725 ) | ( n40723 & n40725 ) ;
  assign n40727 = n40698 | n40726 ;
  assign n40728 = n1057 & ~n32442 ;
  assign n40729 = n1060 & n32306 ;
  assign n40730 = n1065 & n32293 ;
  assign n40731 = n40729 | n40730 ;
  assign n40732 = n40728 | n40731 ;
  assign n40733 = n1062 | n40728 ;
  assign n40734 = n40731 | n40733 ;
  assign n40735 = ( ~n32458 & n40732 ) | ( ~n32458 & n40734 ) | ( n40732 & n40734 ) ;
  assign n40736 = n40719 | n40720 ;
  assign n40737 = ( n40720 & ~n40722 ) | ( n40720 & n40736 ) | ( ~n40722 & n40736 ) ;
  assign n40738 = n40719 & ~n40737 ;
  assign n40739 = n40720 | n40724 ;
  assign n40740 = ( ~n40697 & n40720 ) | ( ~n40697 & n40739 ) | ( n40720 & n40739 ) ;
  assign n40741 = n40719 & ~n40740 ;
  assign n40742 = ( ~n40555 & n40738 ) | ( ~n40555 & n40741 ) | ( n40738 & n40741 ) ;
  assign n40743 = n40735 & n40742 ;
  assign n40744 = ( ~n40727 & n40735 ) | ( ~n40727 & n40743 ) | ( n40735 & n40743 ) ;
  assign n40745 = n40735 | n40742 ;
  assign n40746 = n40727 & ~n40745 ;
  assign n40747 = n40744 | n40746 ;
  assign n40748 = n40590 | n40606 ;
  assign n40749 = ( n40590 & n40591 ) | ( n40590 & n40748 ) | ( n40591 & n40748 ) ;
  assign n40750 = n40747 & ~n40749 ;
  assign n40751 = ~n40747 & n40749 ;
  assign n40752 = n40750 | n40751 ;
  assign n40753 = n1829 & n33526 ;
  assign n40754 = n1826 & n33436 ;
  assign n40755 = n1823 & ~n33423 ;
  assign n40756 = n40754 | n40755 ;
  assign n40757 = n40753 | n40756 ;
  assign n40758 = n1821 & n33545 ;
  assign n40759 = n1821 & ~n33548 ;
  assign n40760 = ( ~n32456 & n40758 ) | ( ~n32456 & n40759 ) | ( n40758 & n40759 ) ;
  assign n40761 = n40757 | n40760 ;
  assign n40762 = n1821 | n40757 ;
  assign n40763 = ( n33536 & n40761 ) | ( n33536 & n40762 ) | ( n40761 & n40762 ) ;
  assign n40764 = x29 | n40763 ;
  assign n40765 = ~x29 & n40763 ;
  assign n40766 = ( ~n40763 & n40764 ) | ( ~n40763 & n40765 ) | ( n40764 & n40765 ) ;
  assign n40767 = ~n40752 & n40766 ;
  assign n40768 = n40752 | n40767 ;
  assign n40769 = n2315 & ~n35371 ;
  assign n40770 = n2312 & n34656 ;
  assign n40771 = n2308 & n35021 ;
  assign n40772 = n40770 | n40771 ;
  assign n40773 = n40769 | n40772 ;
  assign n40774 = n2306 & ~n35392 ;
  assign n40775 = n2306 & ~n35395 ;
  assign n40776 = ( ~n32456 & n40774 ) | ( ~n32456 & n40775 ) | ( n40774 & n40775 ) ;
  assign n40777 = n40773 | n40776 ;
  assign n40778 = n2306 | n40773 ;
  assign n40779 = ( n35381 & n40777 ) | ( n35381 & n40778 ) | ( n40777 & n40778 ) ;
  assign n40780 = x26 | n40779 ;
  assign n40781 = ~x26 & n40779 ;
  assign n40782 = ( ~n40779 & n40780 ) | ( ~n40779 & n40781 ) | ( n40780 & n40781 ) ;
  assign n40783 = n40752 & n40766 ;
  assign n40784 = n40782 & n40783 ;
  assign n40785 = ( ~n40768 & n40782 ) | ( ~n40768 & n40784 ) | ( n40782 & n40784 ) ;
  assign n40786 = n40782 | n40783 ;
  assign n40787 = n40768 & ~n40786 ;
  assign n40788 = n40785 | n40787 ;
  assign n40789 = n40694 & ~n40788 ;
  assign n40790 = n40694 & ~n40789 ;
  assign n40791 = n40694 | n40788 ;
  assign n40792 = ~n40790 & n40791 ;
  assign n40793 = ( n40635 & n40636 ) | ( n40635 & n40652 ) | ( n40636 & n40652 ) ;
  assign n40794 = n40792 & ~n40793 ;
  assign n40795 = ~n40792 & n40793 ;
  assign n40796 = n40794 | n40795 ;
  assign n40797 = n40658 | n40661 ;
  assign n40798 = ~n40796 & n40797 ;
  assign n40799 = n40658 & ~n40796 ;
  assign n40800 = ( n40664 & n40798 ) | ( n40664 & n40799 ) | ( n40798 & n40799 ) ;
  assign n40801 = n40658 | n40667 ;
  assign n40802 = ~n40796 & n40801 ;
  assign n40803 = n40658 | n40669 ;
  assign n40804 = ~n40796 & n40803 ;
  assign n40805 = ( n40380 & n40802 ) | ( n40380 & n40804 ) | ( n40802 & n40804 ) ;
  assign n40806 = ( n39161 & n40800 ) | ( n39161 & n40805 ) | ( n40800 & n40805 ) ;
  assign n40807 = ( n40658 & n40664 ) | ( n40658 & n40797 ) | ( n40664 & n40797 ) ;
  assign n40808 = n40796 & ~n40807 ;
  assign n40809 = ( n40380 & n40801 ) | ( n40380 & n40803 ) | ( n40801 & n40803 ) ;
  assign n40810 = n40796 & ~n40809 ;
  assign n40811 = ( ~n39161 & n40808 ) | ( ~n39161 & n40810 ) | ( n40808 & n40810 ) ;
  assign n40812 = n40806 | n40811 ;
  assign n40813 = ~n40546 & n40676 ;
  assign n40814 = n40396 & n40813 ;
  assign n40815 = n40812 & ~n40814 ;
  assign n40816 = n40676 & ~n40812 ;
  assign n40817 = ~n40546 & n40816 ;
  assign n40818 = n40396 & n40817 ;
  assign n40819 = n40815 | n40818 ;
  assign n40820 = n2315 & n35746 ;
  assign n40821 = n2312 & n35021 ;
  assign n40822 = n2308 & ~n35371 ;
  assign n40823 = n40821 | n40822 ;
  assign n40824 = n40820 | n40823 ;
  assign n40825 = n2306 | n40820 ;
  assign n40826 = n40823 | n40825 ;
  assign n40827 = ( ~n35759 & n40824 ) | ( ~n35759 & n40826 ) | ( n40824 & n40826 ) ;
  assign n40828 = ~x26 & n40826 ;
  assign n40829 = ~x26 & n40824 ;
  assign n40830 = ( ~n35759 & n40828 ) | ( ~n35759 & n40829 ) | ( n40828 & n40829 ) ;
  assign n40831 = x26 | n40829 ;
  assign n40832 = x26 | n40828 ;
  assign n40833 = ( ~n35759 & n40831 ) | ( ~n35759 & n40832 ) | ( n40831 & n40832 ) ;
  assign n40834 = ( ~n40827 & n40830 ) | ( ~n40827 & n40833 ) | ( n40830 & n40833 ) ;
  assign n40835 = n40767 | n40785 ;
  assign n40836 = n8988 | n8992 ;
  assign n40837 = n15188 | n20355 ;
  assign n40838 = n695 | n40837 ;
  assign n40839 = n40836 | n40838 ;
  assign n40840 = n7943 & ~n40839 ;
  assign n40841 = ~n8069 & n40840 ;
  assign n40842 = ( n357 & n3375 ) | ( n357 & ~n17678 ) | ( n3375 & ~n17678 ) ;
  assign n40843 = n574 | n17678 ;
  assign n40844 = n40842 | n40843 ;
  assign n40845 = n594 | n839 ;
  assign n40846 = n133 | n40845 ;
  assign n40847 = n123 | n40846 ;
  assign n40848 = n40844 | n40847 ;
  assign n40849 = n212 | n40848 ;
  assign n40850 = n40841 & ~n40849 ;
  assign n40851 = n40718 & n40850 ;
  assign n40852 = n40718 | n40850 ;
  assign n40853 = ~n40851 & n40852 ;
  assign n40854 = n32068 & n36083 ;
  assign n40855 = ~x23 & n32068 ;
  assign n40856 = n36083 & n40855 ;
  assign n40857 = x23 | n40855 ;
  assign n40858 = ( x23 & n36083 ) | ( x23 & n40857 ) | ( n36083 & n40857 ) ;
  assign n40859 = ( ~n40854 & n40856 ) | ( ~n40854 & n40858 ) | ( n40856 & n40858 ) ;
  assign n40860 = n40853 & ~n40859 ;
  assign n40861 = ~n40853 & n40859 ;
  assign n40862 = n40860 | n40861 ;
  assign n40863 = n40737 & ~n40862 ;
  assign n40864 = n40740 & ~n40862 ;
  assign n40865 = ( n40555 & n40863 ) | ( n40555 & n40864 ) | ( n40863 & n40864 ) ;
  assign n40866 = ~n40737 & n40862 ;
  assign n40867 = ~n40740 & n40862 ;
  assign n40868 = ( ~n40555 & n40866 ) | ( ~n40555 & n40867 ) | ( n40866 & n40867 ) ;
  assign n40869 = n40865 | n40868 ;
  assign n40870 = n1057 & n33436 ;
  assign n40871 = n1060 & n32293 ;
  assign n40872 = n1065 & ~n32442 ;
  assign n40873 = n40871 | n40872 ;
  assign n40874 = n40870 | n40873 ;
  assign n40875 = n1062 & ~n33441 ;
  assign n40876 = ~n32456 & n40875 ;
  assign n40877 = ( n1062 & n34271 ) | ( n1062 & n40876 ) | ( n34271 & n40876 ) ;
  assign n40878 = n40874 | n40877 ;
  assign n40879 = ~n40869 & n40878 ;
  assign n40880 = n40869 | n40879 ;
  assign n40881 = n40869 & n40878 ;
  assign n40882 = n40880 & ~n40881 ;
  assign n40883 = ~n40744 & n40747 ;
  assign n40884 = ( n40744 & n40749 ) | ( n40744 & ~n40883 ) | ( n40749 & ~n40883 ) ;
  assign n40885 = n40882 & ~n40884 ;
  assign n40886 = ~n40882 & n40884 ;
  assign n40887 = n40885 | n40886 ;
  assign n40888 = n1829 & n34656 ;
  assign n40889 = n1826 & ~n33423 ;
  assign n40890 = n1823 & n33526 ;
  assign n40891 = n40889 | n40890 ;
  assign n40892 = n40888 | n40891 ;
  assign n40893 = n1821 | n40888 ;
  assign n40894 = n40891 | n40893 ;
  assign n40895 = ( n34667 & n40892 ) | ( n34667 & n40894 ) | ( n40892 & n40894 ) ;
  assign n40896 = x29 & n40894 ;
  assign n40897 = x29 & n40892 ;
  assign n40898 = ( n34667 & n40896 ) | ( n34667 & n40897 ) | ( n40896 & n40897 ) ;
  assign n40899 = x29 & ~n40897 ;
  assign n40900 = x29 & ~n40896 ;
  assign n40901 = ( ~n34667 & n40899 ) | ( ~n34667 & n40900 ) | ( n40899 & n40900 ) ;
  assign n40902 = ( n40895 & ~n40898 ) | ( n40895 & n40901 ) | ( ~n40898 & n40901 ) ;
  assign n40903 = n40887 & n40902 ;
  assign n40904 = n40882 & ~n40902 ;
  assign n40905 = ( n40884 & n40902 ) | ( n40884 & ~n40904 ) | ( n40902 & ~n40904 ) ;
  assign n40906 = n40885 | n40905 ;
  assign n40907 = ~n40903 & n40906 ;
  assign n40908 = ( n40834 & ~n40835 ) | ( n40834 & n40907 ) | ( ~n40835 & n40907 ) ;
  assign n40909 = ( n40835 & ~n40907 ) | ( n40835 & n40908 ) | ( ~n40907 & n40908 ) ;
  assign n40910 = ( ~n40834 & n40908 ) | ( ~n40834 & n40909 ) | ( n40908 & n40909 ) ;
  assign n40911 = ~n40692 & n40788 ;
  assign n40912 = ( n40692 & n40694 ) | ( n40692 & ~n40911 ) | ( n40694 & ~n40911 ) ;
  assign n40913 = ~n40910 & n40912 ;
  assign n40914 = n40910 & ~n40912 ;
  assign n40915 = n40913 | n40914 ;
  assign n40916 = n40795 | n40798 ;
  assign n40917 = ~n40915 & n40916 ;
  assign n40918 = n40795 | n40799 ;
  assign n40919 = ~n40915 & n40918 ;
  assign n40920 = ( n40664 & n40917 ) | ( n40664 & n40919 ) | ( n40917 & n40919 ) ;
  assign n40921 = n40795 | n40802 ;
  assign n40922 = ~n40915 & n40921 ;
  assign n40923 = n40795 | n40804 ;
  assign n40924 = ~n40915 & n40923 ;
  assign n40925 = ( n40380 & n40922 ) | ( n40380 & n40924 ) | ( n40922 & n40924 ) ;
  assign n40926 = ( n39161 & n40920 ) | ( n39161 & n40925 ) | ( n40920 & n40925 ) ;
  assign n40927 = ( n40664 & n40916 ) | ( n40664 & n40918 ) | ( n40916 & n40918 ) ;
  assign n40928 = n40915 & ~n40927 ;
  assign n40929 = ( n40380 & n40921 ) | ( n40380 & n40923 ) | ( n40921 & n40923 ) ;
  assign n40930 = n40915 & ~n40929 ;
  assign n40931 = ( ~n39161 & n40928 ) | ( ~n39161 & n40930 ) | ( n40928 & n40930 ) ;
  assign n40932 = n40926 | n40931 ;
  assign n40933 = ~n40818 & n40932 ;
  assign n40934 = n40817 & ~n40932 ;
  assign n40935 = n40396 & n40934 ;
  assign n40936 = n40933 | n40935 ;
  assign n40937 = n40766 & n40834 ;
  assign n40938 = ~n40752 & n40937 ;
  assign n40939 = ( n40785 & n40834 ) | ( n40785 & n40938 ) | ( n40834 & n40938 ) ;
  assign n40940 = n40835 & ~n40939 ;
  assign n40941 = n40834 & ~n40937 ;
  assign n40942 = ( n40752 & n40834 ) | ( n40752 & n40941 ) | ( n40834 & n40941 ) ;
  assign n40943 = ~n40785 & n40942 ;
  assign n40944 = n40907 | n40943 ;
  assign n40945 = n40940 | n40944 ;
  assign n40946 = ( ~n40907 & n40939 ) | ( ~n40907 & n40945 ) | ( n40939 & n40945 ) ;
  assign n40974 = n1057 & ~n33423 ;
  assign n40975 = n1060 & ~n32442 ;
  assign n40976 = n1065 & n33436 ;
  assign n40977 = n40975 | n40976 ;
  assign n40978 = n40974 | n40977 ;
  assign n40979 = n1062 & n33575 ;
  assign n40980 = n1062 & ~n33577 ;
  assign n40981 = ( ~n32456 & n40979 ) | ( ~n32456 & n40980 ) | ( n40979 & n40980 ) ;
  assign n40982 = n40978 | n40981 ;
  assign n40983 = n1062 | n40978 ;
  assign n40984 = ( n33567 & n40982 ) | ( n33567 & n40983 ) | ( n40982 & n40983 ) ;
  assign n40947 = n8995 | n8999 ;
  assign n40948 = n630 | n6827 ;
  assign n40949 = n26054 | n40948 ;
  assign n40950 = n1148 | n40949 ;
  assign n40951 = n33214 | n40950 ;
  assign n40952 = n8030 | n40951 ;
  assign n40953 = n40947 | n40952 ;
  assign n40954 = n17685 | n40953 ;
  assign n40955 = n711 | n7937 ;
  assign n40956 = n7936 | n40955 ;
  assign n40957 = n1301 | n3431 ;
  assign n40958 = n2243 | n40957 ;
  assign n40959 = n1171 | n40958 ;
  assign n40960 = n40956 | n40959 ;
  assign n40961 = n209 | n278 ;
  assign n40962 = n223 | n273 ;
  assign n40963 = n40961 | n40962 ;
  assign n40964 = n40960 | n40963 ;
  assign n40965 = n40954 | n40964 ;
  assign n40966 = ( n40852 & ~n40853 ) | ( n40852 & n40965 ) | ( ~n40853 & n40965 ) ;
  assign n40967 = n40852 | n40965 ;
  assign n40968 = ( n40859 & n40966 ) | ( n40859 & n40967 ) | ( n40966 & n40967 ) ;
  assign n40969 = n40852 & ~n40853 ;
  assign n40970 = n40965 & n40969 ;
  assign n40971 = n40852 & n40965 ;
  assign n40972 = ( n40859 & n40970 ) | ( n40859 & n40971 ) | ( n40970 & n40971 ) ;
  assign n40973 = n40968 & ~n40972 ;
  assign n40985 = n40973 | n40984 ;
  assign n40986 = ~n40973 & n40984 ;
  assign n40987 = ( ~n40984 & n40985 ) | ( ~n40984 & n40986 ) | ( n40985 & n40986 ) ;
  assign n40988 = n40865 | n40878 ;
  assign n40989 = ( n40865 & ~n40869 ) | ( n40865 & n40988 ) | ( ~n40869 & n40988 ) ;
  assign n40990 = n40987 | n40989 ;
  assign n40991 = n40987 & n40989 ;
  assign n40992 = n40990 & ~n40991 ;
  assign n40993 = n1829 & n35021 ;
  assign n40994 = n1826 & n33526 ;
  assign n40995 = n1823 & n34656 ;
  assign n40996 = n40994 | n40995 ;
  assign n40997 = n40993 | n40996 ;
  assign n40998 = n1821 | n40993 ;
  assign n40999 = n40996 | n40998 ;
  assign n41000 = ( n35033 & n40997 ) | ( n35033 & n40999 ) | ( n40997 & n40999 ) ;
  assign n41001 = x29 & n40999 ;
  assign n41002 = x29 & n40997 ;
  assign n41003 = ( n35033 & n41001 ) | ( n35033 & n41002 ) | ( n41001 & n41002 ) ;
  assign n41004 = x29 & ~n41002 ;
  assign n41005 = x29 & ~n41001 ;
  assign n41006 = ( ~n35033 & n41004 ) | ( ~n35033 & n41005 ) | ( n41004 & n41005 ) ;
  assign n41007 = ( n41000 & ~n41003 ) | ( n41000 & n41006 ) | ( ~n41003 & n41006 ) ;
  assign n41008 = n40992 & n41007 ;
  assign n41009 = n40992 | n41007 ;
  assign n41010 = ~n41008 & n41009 ;
  assign n41011 = n40886 | n40902 ;
  assign n41012 = ( n40886 & ~n40887 ) | ( n40886 & n41011 ) | ( ~n40887 & n41011 ) ;
  assign n41013 = n41010 & n41012 ;
  assign n41014 = n41010 | n41012 ;
  assign n41015 = ~n41013 & n41014 ;
  assign n41016 = n2315 & n36083 ;
  assign n41017 = n2312 & ~n35371 ;
  assign n41018 = n2308 & n35746 ;
  assign n41019 = n41017 | n41018 ;
  assign n41020 = n41016 | n41019 ;
  assign n41021 = n2306 | n41016 ;
  assign n41022 = n41019 | n41021 ;
  assign n41023 = ( n36107 & n41020 ) | ( n36107 & n41022 ) | ( n41020 & n41022 ) ;
  assign n41024 = n41020 | n41022 ;
  assign n41025 = ( n36094 & n41023 ) | ( n36094 & n41024 ) | ( n41023 & n41024 ) ;
  assign n41026 = x26 & n41025 ;
  assign n41027 = x26 & ~n41025 ;
  assign n41028 = ( n41025 & ~n41026 ) | ( n41025 & n41027 ) | ( ~n41026 & n41027 ) ;
  assign n41029 = n41015 & ~n41028 ;
  assign n41030 = n41015 | n41028 ;
  assign n41031 = ( ~n41015 & n41029 ) | ( ~n41015 & n41030 ) | ( n41029 & n41030 ) ;
  assign n41032 = n40946 & n41031 ;
  assign n41033 = n40946 & ~n41032 ;
  assign n41034 = ~n40946 & n41031 ;
  assign n41035 = n41033 | n41034 ;
  assign n41036 = n40913 | n40920 ;
  assign n41037 = n41035 | n41036 ;
  assign n41038 = n40913 | n40925 ;
  assign n41039 = n41035 | n41038 ;
  assign n41040 = ( n39161 & n41037 ) | ( n39161 & n41039 ) | ( n41037 & n41039 ) ;
  assign n41041 = n41035 & n41036 ;
  assign n41042 = n41035 & n41038 ;
  assign n41043 = ( n39161 & n41041 ) | ( n39161 & n41042 ) | ( n41041 & n41042 ) ;
  assign n41044 = n41040 & ~n41043 ;
  assign n41045 = n40935 & n41044 ;
  assign n41046 = n40935 & ~n41045 ;
  assign n41047 = ( n41044 & ~n41045 ) | ( n41044 & n41046 ) | ( ~n41045 & n41046 ) ;
  assign n41048 = n40968 & ~n40973 ;
  assign n41049 = n40968 & ~n40978 ;
  assign n41050 = ( n40968 & ~n40973 ) | ( n40968 & n41049 ) | ( ~n40973 & n41049 ) ;
  assign n41051 = ( ~n40981 & n41048 ) | ( ~n40981 & n41050 ) | ( n41048 & n41050 ) ;
  assign n41052 = ( ~n1062 & n41048 ) | ( ~n1062 & n41050 ) | ( n41048 & n41050 ) ;
  assign n41053 = ( ~n33567 & n41051 ) | ( ~n33567 & n41052 ) | ( n41051 & n41052 ) ;
  assign n41054 = ~n1649 & n8982 ;
  assign n41055 = n9012 | n21523 ;
  assign n41056 = n7925 | n41055 ;
  assign n41057 = n41054 & ~n41056 ;
  assign n41058 = n133 | n8004 ;
  assign n41059 = n33455 | n41058 ;
  assign n41060 = n41057 & ~n41059 ;
  assign n41061 = n40965 & n41060 ;
  assign n41062 = n40965 | n41060 ;
  assign n41063 = ~n40968 & n41062 ;
  assign n41064 = ( n40973 & n41062 ) | ( n40973 & n41063 ) | ( n41062 & n41063 ) ;
  assign n41065 = ~n41061 & n41064 ;
  assign n41066 = ~n41061 & n41062 ;
  assign n41067 = ~n41050 & n41066 ;
  assign n41068 = ( n40981 & n41065 ) | ( n40981 & n41067 ) | ( n41065 & n41067 ) ;
  assign n41069 = ( n1062 & n41065 ) | ( n1062 & n41067 ) | ( n41065 & n41067 ) ;
  assign n41070 = ( n33567 & n41068 ) | ( n33567 & n41069 ) | ( n41068 & n41069 ) ;
  assign n41071 = n41053 | n41070 ;
  assign n41072 = n41062 & ~n41066 ;
  assign n41073 = ( n41050 & n41062 ) | ( n41050 & n41072 ) | ( n41062 & n41072 ) ;
  assign n41074 = n41061 & n41062 ;
  assign n41075 = ( n41062 & ~n41064 ) | ( n41062 & n41074 ) | ( ~n41064 & n41074 ) ;
  assign n41076 = ( ~n40981 & n41073 ) | ( ~n40981 & n41075 ) | ( n41073 & n41075 ) ;
  assign n41077 = ( ~n1062 & n41073 ) | ( ~n1062 & n41075 ) | ( n41073 & n41075 ) ;
  assign n41078 = ( ~n33567 & n41076 ) | ( ~n33567 & n41077 ) | ( n41076 & n41077 ) ;
  assign n41079 = ~n41061 & n41078 ;
  assign n41080 = n41071 & ~n41079 ;
  assign n41081 = n1057 & n33526 ;
  assign n41082 = n1060 & n33436 ;
  assign n41083 = n1065 & ~n33423 ;
  assign n41084 = n41082 | n41083 ;
  assign n41085 = n41081 | n41084 ;
  assign n41086 = n1062 & n33545 ;
  assign n41087 = n1062 & ~n33548 ;
  assign n41088 = ( ~n32456 & n41086 ) | ( ~n32456 & n41087 ) | ( n41086 & n41087 ) ;
  assign n41089 = n41085 | n41088 ;
  assign n41090 = n1062 | n41085 ;
  assign n41091 = ( n33536 & n41089 ) | ( n33536 & n41090 ) | ( n41089 & n41090 ) ;
  assign n41092 = ~n41080 & n41091 ;
  assign n41093 = n41080 & ~n41091 ;
  assign n41094 = n41092 | n41093 ;
  assign n41095 = n40991 | n41007 ;
  assign n41096 = ( n40991 & n40992 ) | ( n40991 & n41095 ) | ( n40992 & n41095 ) ;
  assign n41097 = n41094 & ~n41096 ;
  assign n41098 = ~n41094 & n41096 ;
  assign n41099 = n41097 | n41098 ;
  assign n41100 = n1829 & ~n35371 ;
  assign n41101 = n1826 & n34656 ;
  assign n41102 = n1823 & n35021 ;
  assign n41103 = n41101 | n41102 ;
  assign n41104 = n41100 | n41103 ;
  assign n41105 = n1821 & ~n35392 ;
  assign n41106 = n1821 & ~n35395 ;
  assign n41107 = ( ~n32456 & n41105 ) | ( ~n32456 & n41106 ) | ( n41105 & n41106 ) ;
  assign n41108 = n41104 | n41107 ;
  assign n41109 = n1821 | n41104 ;
  assign n41110 = ( n35381 & n41108 ) | ( n35381 & n41109 ) | ( n41108 & n41109 ) ;
  assign n41111 = ~x29 & n41110 ;
  assign n41112 = n33226 & n36083 ;
  assign n41113 = n2312 & n35746 ;
  assign n41114 = n41112 | n41113 ;
  assign n41115 = n2306 | n41114 ;
  assign n41116 = ( n36103 & n41114 ) | ( n36103 & n41115 ) | ( n41114 & n41115 ) ;
  assign n41117 = ( n36105 & n41114 ) | ( n36105 & n41115 ) | ( n41114 & n41115 ) ;
  assign n41118 = ( n32456 & n41116 ) | ( n32456 & n41117 ) | ( n41116 & n41117 ) ;
  assign n41119 = x26 & n41118 ;
  assign n41120 = x26 & ~n41118 ;
  assign n41121 = ( n41118 & ~n41119 ) | ( n41118 & n41120 ) | ( ~n41119 & n41120 ) ;
  assign n41122 = x29 & n41100 ;
  assign n41123 = ( x29 & n41103 ) | ( x29 & n41122 ) | ( n41103 & n41122 ) ;
  assign n41124 = x29 & ~n41123 ;
  assign n41125 = ~n41107 & n41124 ;
  assign n41126 = ~n1821 & n41124 ;
  assign n41127 = ( ~n35381 & n41125 ) | ( ~n35381 & n41126 ) | ( n41125 & n41126 ) ;
  assign n41128 = n41121 & n41127 ;
  assign n41129 = ( n41111 & n41121 ) | ( n41111 & n41128 ) | ( n41121 & n41128 ) ;
  assign n41130 = n41121 | n41127 ;
  assign n41131 = n41111 | n41130 ;
  assign n41132 = ~n41129 & n41131 ;
  assign n41133 = n41099 & ~n41132 ;
  assign n41134 = ~n41099 & n41132 ;
  assign n41135 = n41133 | n41134 ;
  assign n41136 = n41013 | n41028 ;
  assign n41137 = ( n41013 & n41015 ) | ( n41013 & n41136 ) | ( n41015 & n41136 ) ;
  assign n41138 = ~n41135 & n41137 ;
  assign n41139 = n41135 & ~n41137 ;
  assign n41140 = n41138 | n41139 ;
  assign n41141 = n41032 | n41034 ;
  assign n41142 = n41033 | n41141 ;
  assign n41143 = ~n41140 & n41142 ;
  assign n41144 = n41032 & ~n41140 ;
  assign n41145 = ( n41036 & n41143 ) | ( n41036 & n41144 ) | ( n41143 & n41144 ) ;
  assign n41146 = ( n41038 & n41143 ) | ( n41038 & n41144 ) | ( n41143 & n41144 ) ;
  assign n41147 = ( n39161 & n41145 ) | ( n39161 & n41146 ) | ( n41145 & n41146 ) ;
  assign n41148 = ( n40946 & n41031 ) | ( n40946 & n41036 ) | ( n41031 & n41036 ) ;
  assign n41149 = n41140 & ~n41148 ;
  assign n41150 = ( n40946 & n41031 ) | ( n40946 & n41038 ) | ( n41031 & n41038 ) ;
  assign n41151 = n41140 & ~n41150 ;
  assign n41152 = ( ~n39161 & n41149 ) | ( ~n39161 & n41151 ) | ( n41149 & n41151 ) ;
  assign n41153 = n41147 | n41152 ;
  assign n41154 = ~n41045 & n41153 ;
  assign n41155 = n41044 & ~n41153 ;
  assign n41156 = n40934 & n41155 ;
  assign n41157 = n40396 & n41156 ;
  assign n41158 = n41154 | n41157 ;
  assign n41159 = ~n41138 & n41140 ;
  assign n41160 = ( n41138 & n41142 ) | ( n41138 & ~n41159 ) | ( n41142 & ~n41159 ) ;
  assign n41161 = ( n41032 & n41138 ) | ( n41032 & ~n41159 ) | ( n41138 & ~n41159 ) ;
  assign n41162 = ( n41036 & n41160 ) | ( n41036 & n41161 ) | ( n41160 & n41161 ) ;
  assign n41163 = ( n41038 & n41160 ) | ( n41038 & n41161 ) | ( n41160 & n41161 ) ;
  assign n41164 = ( n39161 & n41162 ) | ( n39161 & n41163 ) | ( n41162 & n41163 ) ;
  assign n41165 = n1829 & n35746 ;
  assign n41166 = n1826 & n35021 ;
  assign n41167 = n1823 & ~n35371 ;
  assign n41168 = n41166 | n41167 ;
  assign n41169 = n41165 | n41168 ;
  assign n41170 = n1821 | n41165 ;
  assign n41171 = n41168 | n41170 ;
  assign n41172 = ( ~n35759 & n41169 ) | ( ~n35759 & n41171 ) | ( n41169 & n41171 ) ;
  assign n41173 = ~n41092 & n41094 ;
  assign n41174 = ( n41092 & n41096 ) | ( n41092 & ~n41173 ) | ( n41096 & ~n41173 ) ;
  assign n41175 = ( x29 & n41172 ) | ( x29 & ~n41174 ) | ( n41172 & ~n41174 ) ;
  assign n41176 = ( ~x29 & n41174 ) | ( ~x29 & n41175 ) | ( n41174 & n41175 ) ;
  assign n41177 = ( ~n41172 & n41175 ) | ( ~n41172 & n41176 ) | ( n41175 & n41176 ) ;
  assign n41178 = n1057 & n34656 ;
  assign n41179 = n1060 & ~n33423 ;
  assign n41180 = n1065 & n33526 ;
  assign n41181 = n41179 | n41180 ;
  assign n41182 = n41178 | n41181 ;
  assign n41183 = n1062 | n41178 ;
  assign n41184 = n41181 | n41183 ;
  assign n41185 = ( n34667 & n41182 ) | ( n34667 & n41184 ) | ( n41182 & n41184 ) ;
  assign n41186 = ( ~n41078 & n41175 ) | ( ~n41078 & n41185 ) | ( n41175 & n41185 ) ;
  assign n41187 = ( n41078 & n41172 ) | ( n41078 & ~n41185 ) | ( n41172 & ~n41185 ) ;
  assign n41188 = ( n41176 & n41186 ) | ( n41176 & ~n41187 ) | ( n41186 & ~n41187 ) ;
  assign n41189 = ( n41078 & ~n41177 ) | ( n41078 & n41188 ) | ( ~n41177 & n41188 ) ;
  assign n41190 = n41129 | n41132 ;
  assign n41191 = ( ~n41099 & n41129 ) | ( ~n41099 & n41190 ) | ( n41129 & n41190 ) ;
  assign n41192 = n9001 | n33457 ;
  assign n41193 = n9018 | n41192 ;
  assign n41194 = x26 & n401 ;
  assign n41195 = ( x26 & n41193 ) | ( x26 & ~n41194 ) | ( n41193 & ~n41194 ) ;
  assign n41196 = x26 | n41194 ;
  assign n41197 = n41193 & ~n41196 ;
  assign n41198 = ( ~n41193 & n41195 ) | ( ~n41193 & n41197 ) | ( n41195 & n41197 ) ;
  assign n41200 = ( n33228 & n40965 ) | ( n33228 & n41198 ) | ( n40965 & n41198 ) ;
  assign n41201 = n40965 & n41198 ;
  assign n41202 = ( n36083 & n41200 ) | ( n36083 & n41201 ) | ( n41200 & n41201 ) ;
  assign n41199 = n33228 & n36083 ;
  assign n41203 = ( n41198 & n41199 ) | ( n41198 & ~n41202 ) | ( n41199 & ~n41202 ) ;
  assign n41204 = ( n40965 & ~n41202 ) | ( n40965 & n41203 ) | ( ~n41202 & n41203 ) ;
  assign n41205 = n41190 & n41204 ;
  assign n41206 = n41129 & n41204 ;
  assign n41207 = ( ~n41099 & n41205 ) | ( ~n41099 & n41206 ) | ( n41205 & n41206 ) ;
  assign n41208 = n41204 & ~n41205 ;
  assign n41209 = n41204 & ~n41206 ;
  assign n41210 = ( n41099 & n41208 ) | ( n41099 & n41209 ) | ( n41208 & n41209 ) ;
  assign n41211 = ( n41191 & ~n41207 ) | ( n41191 & n41210 ) | ( ~n41207 & n41210 ) ;
  assign n41212 = n41188 & n41211 ;
  assign n41213 = ~n41185 & n41211 ;
  assign n41214 = ( n41189 & n41212 ) | ( n41189 & n41213 ) | ( n41212 & n41213 ) ;
  assign n41215 = n41188 | n41211 ;
  assign n41216 = n41185 & ~n41211 ;
  assign n41217 = ( n41189 & n41215 ) | ( n41189 & ~n41216 ) | ( n41215 & ~n41216 ) ;
  assign n41218 = ~n41214 & n41217 ;
  assign n41219 = n41162 & n41218 ;
  assign n41220 = n41163 & n41218 ;
  assign n41221 = ( n39161 & n41219 ) | ( n39161 & n41220 ) | ( n41219 & n41220 ) ;
  assign n41222 = n41218 & ~n41219 ;
  assign n41223 = n41218 & ~n41220 ;
  assign n41224 = ( ~n39161 & n41222 ) | ( ~n39161 & n41223 ) | ( n41222 & n41223 ) ;
  assign n41225 = ( n41164 & ~n41221 ) | ( n41164 & n41224 ) | ( ~n41221 & n41224 ) ;
  assign n41226 = n41157 & ~n41225 ;
  assign n41227 = n41157 | n41225 ;
  assign n41228 = ( ~n41157 & n41226 ) | ( ~n41157 & n41227 ) | ( n41226 & n41227 ) ;
  assign y0 = n34310 ;
  assign y1 = n34699 ;
  assign y2 = ~n35064 ;
  assign y3 = ~n35417 ;
  assign y4 = ~n35788 ;
  assign y5 = ~n36124 ;
  assign y6 = ~n36409 ;
  assign y7 = ~n36694 ;
  assign y8 = n36965 ;
  assign y9 = n37238 ;
  assign y10 = n37508 ;
  assign y11 = n37765 ;
  assign y12 = ~n38031 ;
  assign y13 = ~n38270 ;
  assign y14 = ~n38502 ;
  assign y15 = n38739 ;
  assign y16 = ~n38968 ;
  assign y17 = n39168 ;
  assign y18 = ~n39377 ;
  assign y19 = ~n39557 ;
  assign y20 = ~n39729 ;
  assign y21 = n39912 ;
  assign y22 = n40077 ;
  assign y23 = ~n40236 ;
  assign y24 = ~n40399 ;
  assign y25 = ~n40548 ;
  assign y26 = n40679 ;
  assign y27 = ~n40819 ;
  assign y28 = ~n40936 ;
  assign y29 = n41047 ;
  assign y30 = ~n41158 ;
  assign y31 = n41228 ;
endmodule
