module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 ;
  wire n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 ;
  assign n66 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n67 = ( ~x0 & x1 ) | ( ~x0 & n66 ) | ( x1 & n66 ) ;
  assign n68 = ( ~x2 & n66 ) | ( ~x2 & n67 ) | ( n66 & n67 ) ;
  assign n69 = ( x0 & x1 ) | ( x0 & x2 ) | ( x1 & x2 ) ;
  assign n70 = ( x3 & ~x4 ) | ( x3 & n69 ) | ( ~x4 & n69 ) ;
  assign n71 = ( ~x3 & x4 ) | ( ~x3 & n70 ) | ( x4 & n70 ) ;
  assign n72 = ( ~n69 & n70 ) | ( ~n69 & n71 ) | ( n70 & n71 ) ;
  assign n73 = ( x3 & x4 ) | ( x3 & n69 ) | ( x4 & n69 ) ;
  assign n74 = ( x5 & ~x6 ) | ( x5 & n73 ) | ( ~x6 & n73 ) ;
  assign n75 = ( ~x5 & x6 ) | ( ~x5 & n74 ) | ( x6 & n74 ) ;
  assign n76 = ( ~n73 & n74 ) | ( ~n73 & n75 ) | ( n74 & n75 ) ;
  assign n77 = ( x5 & x6 ) | ( x5 & n73 ) | ( x6 & n73 ) ;
  assign n78 = ( x7 & ~x8 ) | ( x7 & n77 ) | ( ~x8 & n77 ) ;
  assign n79 = ( ~x7 & x8 ) | ( ~x7 & n78 ) | ( x8 & n78 ) ;
  assign n80 = ( ~n77 & n78 ) | ( ~n77 & n79 ) | ( n78 & n79 ) ;
  assign n81 = ( x7 & x8 ) | ( x7 & n77 ) | ( x8 & n77 ) ;
  assign n82 = ( x9 & ~x10 ) | ( x9 & n81 ) | ( ~x10 & n81 ) ;
  assign n83 = ( ~x9 & x10 ) | ( ~x9 & n82 ) | ( x10 & n82 ) ;
  assign n84 = ( ~n81 & n82 ) | ( ~n81 & n83 ) | ( n82 & n83 ) ;
  assign n85 = ( x9 & x10 ) | ( x9 & n81 ) | ( x10 & n81 ) ;
  assign n86 = ( x11 & ~x12 ) | ( x11 & n85 ) | ( ~x12 & n85 ) ;
  assign n87 = ( ~x11 & x12 ) | ( ~x11 & n86 ) | ( x12 & n86 ) ;
  assign n88 = ( ~n85 & n86 ) | ( ~n85 & n87 ) | ( n86 & n87 ) ;
  assign n89 = ( x11 & x12 ) | ( x11 & n85 ) | ( x12 & n85 ) ;
  assign n90 = ( x13 & ~x14 ) | ( x13 & n89 ) | ( ~x14 & n89 ) ;
  assign n91 = ( ~x13 & x14 ) | ( ~x13 & n90 ) | ( x14 & n90 ) ;
  assign n92 = ( ~n89 & n90 ) | ( ~n89 & n91 ) | ( n90 & n91 ) ;
  assign n93 = ( x13 & x14 ) | ( x13 & n89 ) | ( x14 & n89 ) ;
  assign n94 = ( x15 & ~x16 ) | ( x15 & n93 ) | ( ~x16 & n93 ) ;
  assign n95 = ( ~x15 & x16 ) | ( ~x15 & n94 ) | ( x16 & n94 ) ;
  assign n96 = ( ~n93 & n94 ) | ( ~n93 & n95 ) | ( n94 & n95 ) ;
  assign n97 = ( x15 & x16 ) | ( x15 & n93 ) | ( x16 & n93 ) ;
  assign n98 = ( x17 & ~x18 ) | ( x17 & n97 ) | ( ~x18 & n97 ) ;
  assign n99 = ( ~x17 & x18 ) | ( ~x17 & n98 ) | ( x18 & n98 ) ;
  assign n100 = ( ~n97 & n98 ) | ( ~n97 & n99 ) | ( n98 & n99 ) ;
  assign n101 = ( x17 & x18 ) | ( x17 & n97 ) | ( x18 & n97 ) ;
  assign n102 = ( x19 & ~x20 ) | ( x19 & n101 ) | ( ~x20 & n101 ) ;
  assign n103 = ( ~x19 & x20 ) | ( ~x19 & n102 ) | ( x20 & n102 ) ;
  assign n104 = ( ~n101 & n102 ) | ( ~n101 & n103 ) | ( n102 & n103 ) ;
  assign n105 = ( x19 & x20 ) | ( x19 & n101 ) | ( x20 & n101 ) ;
  assign n106 = ( x21 & ~x22 ) | ( x21 & n105 ) | ( ~x22 & n105 ) ;
  assign n107 = ( ~x21 & x22 ) | ( ~x21 & n106 ) | ( x22 & n106 ) ;
  assign n108 = ( ~n105 & n106 ) | ( ~n105 & n107 ) | ( n106 & n107 ) ;
  assign n109 = ( x21 & x22 ) | ( x21 & n105 ) | ( x22 & n105 ) ;
  assign n110 = ( x23 & ~x24 ) | ( x23 & n109 ) | ( ~x24 & n109 ) ;
  assign n111 = ( ~x23 & x24 ) | ( ~x23 & n110 ) | ( x24 & n110 ) ;
  assign n112 = ( ~n109 & n110 ) | ( ~n109 & n111 ) | ( n110 & n111 ) ;
  assign n113 = ( x23 & x24 ) | ( x23 & n109 ) | ( x24 & n109 ) ;
  assign n114 = ( x25 & ~x26 ) | ( x25 & n113 ) | ( ~x26 & n113 ) ;
  assign n115 = ( ~x25 & x26 ) | ( ~x25 & n114 ) | ( x26 & n114 ) ;
  assign n116 = ( ~n113 & n114 ) | ( ~n113 & n115 ) | ( n114 & n115 ) ;
  assign n117 = ( x25 & x26 ) | ( x25 & n113 ) | ( x26 & n113 ) ;
  assign n118 = ( x27 & ~x28 ) | ( x27 & n117 ) | ( ~x28 & n117 ) ;
  assign n119 = ( ~x27 & x28 ) | ( ~x27 & n118 ) | ( x28 & n118 ) ;
  assign n120 = ( ~n117 & n118 ) | ( ~n117 & n119 ) | ( n118 & n119 ) ;
  assign n121 = ( x27 & x28 ) | ( x27 & n117 ) | ( x28 & n117 ) ;
  assign n122 = ( x29 & ~x30 ) | ( x29 & n121 ) | ( ~x30 & n121 ) ;
  assign n123 = ( ~x29 & x30 ) | ( ~x29 & n122 ) | ( x30 & n122 ) ;
  assign n124 = ( ~n121 & n122 ) | ( ~n121 & n123 ) | ( n122 & n123 ) ;
  assign n125 = ( x29 & x30 ) | ( x29 & n121 ) | ( x30 & n121 ) ;
  assign n126 = ( x31 & ~x32 ) | ( x31 & n125 ) | ( ~x32 & n125 ) ;
  assign n127 = ( ~x31 & x32 ) | ( ~x31 & n126 ) | ( x32 & n126 ) ;
  assign n128 = ( ~n125 & n126 ) | ( ~n125 & n127 ) | ( n126 & n127 ) ;
  assign n129 = ( x31 & x32 ) | ( x31 & n125 ) | ( x32 & n125 ) ;
  assign n130 = ( x33 & ~x34 ) | ( x33 & n129 ) | ( ~x34 & n129 ) ;
  assign n131 = ( ~x33 & x34 ) | ( ~x33 & n130 ) | ( x34 & n130 ) ;
  assign n132 = ( ~n129 & n130 ) | ( ~n129 & n131 ) | ( n130 & n131 ) ;
  assign n133 = ( x33 & x34 ) | ( x33 & n129 ) | ( x34 & n129 ) ;
  assign n134 = ( x35 & ~x36 ) | ( x35 & n133 ) | ( ~x36 & n133 ) ;
  assign n135 = ( ~x35 & x36 ) | ( ~x35 & n134 ) | ( x36 & n134 ) ;
  assign n136 = ( ~n133 & n134 ) | ( ~n133 & n135 ) | ( n134 & n135 ) ;
  assign n137 = ( x35 & x36 ) | ( x35 & n133 ) | ( x36 & n133 ) ;
  assign n138 = ( x37 & ~x38 ) | ( x37 & n137 ) | ( ~x38 & n137 ) ;
  assign n139 = ( ~x37 & x38 ) | ( ~x37 & n138 ) | ( x38 & n138 ) ;
  assign n140 = ( ~n137 & n138 ) | ( ~n137 & n139 ) | ( n138 & n139 ) ;
  assign n141 = ( x37 & x38 ) | ( x37 & n137 ) | ( x38 & n137 ) ;
  assign n142 = ( x39 & ~x40 ) | ( x39 & n141 ) | ( ~x40 & n141 ) ;
  assign n143 = ( ~x39 & x40 ) | ( ~x39 & n142 ) | ( x40 & n142 ) ;
  assign n144 = ( ~n141 & n142 ) | ( ~n141 & n143 ) | ( n142 & n143 ) ;
  assign n145 = ( x39 & x40 ) | ( x39 & n141 ) | ( x40 & n141 ) ;
  assign n146 = ( x41 & ~x42 ) | ( x41 & n145 ) | ( ~x42 & n145 ) ;
  assign n147 = ( ~x41 & x42 ) | ( ~x41 & n146 ) | ( x42 & n146 ) ;
  assign n148 = ( ~n145 & n146 ) | ( ~n145 & n147 ) | ( n146 & n147 ) ;
  assign n149 = ( x41 & x42 ) | ( x41 & n145 ) | ( x42 & n145 ) ;
  assign n150 = ( x43 & ~x44 ) | ( x43 & n149 ) | ( ~x44 & n149 ) ;
  assign n151 = ( ~x43 & x44 ) | ( ~x43 & n150 ) | ( x44 & n150 ) ;
  assign n152 = ( ~n149 & n150 ) | ( ~n149 & n151 ) | ( n150 & n151 ) ;
  assign n153 = ( x43 & x44 ) | ( x43 & n149 ) | ( x44 & n149 ) ;
  assign n154 = ( x45 & ~x46 ) | ( x45 & n153 ) | ( ~x46 & n153 ) ;
  assign n155 = ( ~x45 & x46 ) | ( ~x45 & n154 ) | ( x46 & n154 ) ;
  assign n156 = ( ~n153 & n154 ) | ( ~n153 & n155 ) | ( n154 & n155 ) ;
  assign n157 = ( x45 & x46 ) | ( x45 & n153 ) | ( x46 & n153 ) ;
  assign n158 = ( x47 & ~x48 ) | ( x47 & n157 ) | ( ~x48 & n157 ) ;
  assign n159 = ( ~x47 & x48 ) | ( ~x47 & n158 ) | ( x48 & n158 ) ;
  assign n160 = ( ~n157 & n158 ) | ( ~n157 & n159 ) | ( n158 & n159 ) ;
  assign n161 = ( x47 & x48 ) | ( x47 & n157 ) | ( x48 & n157 ) ;
  assign n162 = ( x49 & ~x50 ) | ( x49 & n161 ) | ( ~x50 & n161 ) ;
  assign n163 = ( ~x49 & x50 ) | ( ~x49 & n162 ) | ( x50 & n162 ) ;
  assign n164 = ( ~n161 & n162 ) | ( ~n161 & n163 ) | ( n162 & n163 ) ;
  assign n165 = ( x49 & x50 ) | ( x49 & n161 ) | ( x50 & n161 ) ;
  assign n166 = ( x51 & ~x52 ) | ( x51 & n165 ) | ( ~x52 & n165 ) ;
  assign n167 = ( ~x51 & x52 ) | ( ~x51 & n166 ) | ( x52 & n166 ) ;
  assign n168 = ( ~n165 & n166 ) | ( ~n165 & n167 ) | ( n166 & n167 ) ;
  assign n169 = ( x51 & x52 ) | ( x51 & n165 ) | ( x52 & n165 ) ;
  assign n170 = ( x53 & ~x54 ) | ( x53 & n169 ) | ( ~x54 & n169 ) ;
  assign n171 = ( ~x53 & x54 ) | ( ~x53 & n170 ) | ( x54 & n170 ) ;
  assign n172 = ( ~n169 & n170 ) | ( ~n169 & n171 ) | ( n170 & n171 ) ;
  assign n173 = ( x53 & x54 ) | ( x53 & n169 ) | ( x54 & n169 ) ;
  assign n174 = ( x55 & ~x56 ) | ( x55 & n173 ) | ( ~x56 & n173 ) ;
  assign n175 = ( ~x55 & x56 ) | ( ~x55 & n174 ) | ( x56 & n174 ) ;
  assign n176 = ( ~n173 & n174 ) | ( ~n173 & n175 ) | ( n174 & n175 ) ;
  assign n177 = ( x55 & x56 ) | ( x55 & n173 ) | ( x56 & n173 ) ;
  assign n178 = ( x57 & ~x58 ) | ( x57 & n177 ) | ( ~x58 & n177 ) ;
  assign n179 = ( ~x57 & x58 ) | ( ~x57 & n178 ) | ( x58 & n178 ) ;
  assign n180 = ( ~n177 & n178 ) | ( ~n177 & n179 ) | ( n178 & n179 ) ;
  assign n181 = ( x57 & x58 ) | ( x57 & n177 ) | ( x58 & n177 ) ;
  assign n182 = ( x59 & ~x60 ) | ( x59 & n181 ) | ( ~x60 & n181 ) ;
  assign n183 = ( ~x59 & x60 ) | ( ~x59 & n182 ) | ( x60 & n182 ) ;
  assign n184 = ( ~n181 & n182 ) | ( ~n181 & n183 ) | ( n182 & n183 ) ;
  assign n185 = ( x59 & x60 ) | ( x59 & n181 ) | ( x60 & n181 ) ;
  assign n186 = ( x61 & ~x62 ) | ( x61 & n185 ) | ( ~x62 & n185 ) ;
  assign n187 = ( ~x61 & x62 ) | ( ~x61 & n186 ) | ( x62 & n186 ) ;
  assign n188 = ( ~n185 & n186 ) | ( ~n185 & n187 ) | ( n186 & n187 ) ;
  assign n189 = ( x61 & x62 ) | ( x61 & n185 ) | ( x62 & n185 ) ;
  assign n190 = ( x63 & ~x64 ) | ( x63 & n189 ) | ( ~x64 & n189 ) ;
  assign n191 = ( ~x63 & x64 ) | ( ~x63 & n190 ) | ( x64 & n190 ) ;
  assign n192 = ( ~n189 & n190 ) | ( ~n189 & n191 ) | ( n190 & n191 ) ;
  assign n193 = ( x63 & x64 ) | ( x63 & n189 ) | ( x64 & n189 ) ;
  assign y0 = n68 ;
  assign y1 = n72 ;
  assign y2 = n76 ;
  assign y3 = n80 ;
  assign y4 = n84 ;
  assign y5 = n88 ;
  assign y6 = n92 ;
  assign y7 = n96 ;
  assign y8 = n100 ;
  assign y9 = n104 ;
  assign y10 = n108 ;
  assign y11 = n112 ;
  assign y12 = n116 ;
  assign y13 = n120 ;
  assign y14 = n124 ;
  assign y15 = n128 ;
  assign y16 = n132 ;
  assign y17 = n136 ;
  assign y18 = n140 ;
  assign y19 = n144 ;
  assign y20 = n148 ;
  assign y21 = n152 ;
  assign y22 = n156 ;
  assign y23 = n160 ;
  assign y24 = n164 ;
  assign y25 = n168 ;
  assign y26 = n172 ;
  assign y27 = n176 ;
  assign y28 = n180 ;
  assign y29 = n184 ;
  assign y30 = n188 ;
  assign y31 = n192 ;
  assign y32 = n193 ;
endmodule
