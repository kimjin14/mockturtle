module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 ;
  assign n11 = x3 | x5 ;
  assign n12 = ~x1 & x9 ;
  assign n13 = ~x0 & x9 ;
  assign n14 = x1 & ~n13 ;
  assign n15 = n12 | n14 ;
  assign n16 = n11 | n15 ;
  assign n17 = x0 & ~x9 ;
  assign n18 = x1 | n17 ;
  assign n19 = x1 & ~x9 ;
  assign n20 = x7 | n19 ;
  assign n21 = n18 & ~n20 ;
  assign n22 = n16 & ~n21 ;
  assign n23 = x2 | n22 ;
  assign n24 = x2 | x5 ;
  assign n25 = x1 & x2 ;
  assign n26 = ( ~x0 & n24 ) | ( ~x0 & n25 ) | ( n24 & n25 ) ;
  assign n27 = ~x9 & n26 ;
  assign n28 = x1 & ~x3 ;
  assign n29 = x0 | x9 ;
  assign n30 = x2 & ~x3 ;
  assign n31 = n12 & n30 ;
  assign n32 = ~x1 & x3 ;
  assign n33 = ( n29 & n31 ) | ( n29 & n32 ) | ( n31 & n32 ) ;
  assign n34 = n28 | n33 ;
  assign n35 = n27 | n34 ;
  assign n36 = ~x7 & n35 ;
  assign n37 = n23 & ~n36 ;
  assign n38 = x8 | n37 ;
  assign n39 = x5 | x9 ;
  assign n40 = ( ~x7 & n20 ) | ( ~x7 & n39 ) | ( n20 & n39 ) ;
  assign n41 = x7 & x8 ;
  assign n42 = ~x5 & n41 ;
  assign n43 = ( x1 & ~n20 ) | ( x1 & n42 ) | ( ~n20 & n42 ) ;
  assign n44 = n40 & ~n43 ;
  assign n45 = x0 & ~x2 ;
  assign n46 = ~n44 & n45 ;
  assign n47 = x2 & ~x9 ;
  assign n48 = x0 | x1 ;
  assign n49 = n47 & ~n48 ;
  assign n50 = n42 & n49 ;
  assign n51 = n46 | n50 ;
  assign n52 = ~x3 & n51 ;
  assign n53 = n38 & ~n52 ;
  assign n54 = x6 | n53 ;
  assign n55 = x0 | x2 ;
  assign n56 = n12 & ~n55 ;
  assign n57 = x5 | n56 ;
  assign n58 = x0 & x9 ;
  assign n59 = n29 & ~n58 ;
  assign n60 = x1 & ~n59 ;
  assign n61 = x2 & n60 ;
  assign n62 = x5 & n61 ;
  assign n63 = ( x6 & n57 ) | ( x6 & n62 ) | ( n57 & n62 ) ;
  assign n64 = x8 & n63 ;
  assign n65 = ~x1 & x2 ;
  assign n66 = n17 & n65 ;
  assign n67 = x1 & ~x8 ;
  assign n68 = ( ~x8 & n13 ) | ( ~x8 & n67 ) | ( n13 & n67 ) ;
  assign n69 = n66 | n68 ;
  assign n70 = ~x5 & n69 ;
  assign n71 = n64 | n70 ;
  assign n72 = x3 & n71 ;
  assign n73 = x2 | n17 ;
  assign n74 = x6 & n73 ;
  assign n75 = x2 | x3 ;
  assign n76 = n60 & ~n75 ;
  assign n77 = n74 | n76 ;
  assign n78 = x5 & n77 ;
  assign n79 = x2 & n13 ;
  assign n80 = ~x2 & n19 ;
  assign n81 = ~x0 & n80 ;
  assign n82 = ( ~x3 & n79 ) | ( ~x3 & n81 ) | ( n79 & n81 ) ;
  assign n83 = x6 & n82 ;
  assign n84 = n78 | n83 ;
  assign n85 = x8 & n84 ;
  assign n86 = x2 & x9 ;
  assign n87 = x1 | x9 ;
  assign n88 = x3 & ~x6 ;
  assign n89 = ( x2 & x3 ) | ( x2 & n88 ) | ( x3 & n88 ) ;
  assign n90 = n87 | n89 ;
  assign n91 = ~n86 & n90 ;
  assign n92 = x8 | n91 ;
  assign n93 = ( ~x0 & n31 ) | ( ~x0 & n67 ) | ( n31 & n67 ) ;
  assign n94 = n92 & ~n93 ;
  assign n95 = x5 | n94 ;
  assign n96 = x0 | n75 ;
  assign n97 = x8 | n87 ;
  assign n98 = n96 | n97 ;
  assign n99 = n95 & n98 ;
  assign n100 = ~n85 & n99 ;
  assign n101 = ~n72 & n100 ;
  assign n102 = x7 | n101 ;
  assign n103 = n54 & n102 ;
  assign n104 = x4 | n103 ;
  assign n105 = x4 & x8 ;
  assign n106 = ~x6 & x8 ;
  assign n107 = x8 | x9 ;
  assign n108 = x6 | n107 ;
  assign n109 = ( ~n105 & n106 ) | ( ~n105 & n108 ) | ( n106 & n108 ) ;
  assign n110 = x5 & ~n109 ;
  assign n111 = x4 & x9 ;
  assign n112 = x5 & x6 ;
  assign n113 = ~x5 & x6 ;
  assign n114 = ~x9 & n113 ;
  assign n115 = ( n111 & ~n112 ) | ( n111 & n114 ) | ( ~n112 & n114 ) ;
  assign n116 = ~x8 & n115 ;
  assign n117 = n110 | n116 ;
  assign n118 = ~x7 & n117 ;
  assign n119 = x1 | x3 ;
  assign n120 = ( n55 & n118 ) | ( n55 & ~n119 ) | ( n118 & ~n119 ) ;
  assign n121 = ~n55 & n120 ;
  assign n122 = n104 & ~n121 ;
  assign n123 = x8 | n39 ;
  assign n124 = ~x5 & x8 ;
  assign n125 = x6 & x9 ;
  assign n126 = n124 | n125 ;
  assign n127 = x6 & x8 ;
  assign n128 = n126 & ~n127 ;
  assign n129 = x0 & n128 ;
  assign n130 = ( n123 & ~n126 ) | ( n123 & n129 ) | ( ~n126 & n129 ) ;
  assign n131 = ( n17 & n123 ) | ( n17 & n130 ) | ( n123 & n130 ) ;
  assign n132 = x2 & ~n131 ;
  assign n133 = x2 | x8 ;
  assign n134 = x0 | n133 ;
  assign n135 = x8 & n58 ;
  assign n136 = ( x5 & ~n107 ) | ( x5 & n135 ) | ( ~n107 & n135 ) ;
  assign n137 = ( n86 & ~n134 ) | ( n86 & n136 ) | ( ~n134 & n136 ) ;
  assign n138 = n132 | n137 ;
  assign n139 = ~x4 & n138 ;
  assign n140 = ~x6 & x9 ;
  assign n141 = x5 & ~x8 ;
  assign n142 = ( ~x6 & n105 ) | ( ~x6 & n141 ) | ( n105 & n141 ) ;
  assign n143 = n111 | n142 ;
  assign n144 = ~n140 & n143 ;
  assign n145 = ~n55 & n144 ;
  assign n146 = n139 | n145 ;
  assign n147 = ~x1 & n146 ;
  assign n148 = ~x0 & x5 ;
  assign n149 = ~x8 & x9 ;
  assign n150 = n148 & n149 ;
  assign n151 = n129 | n150 ;
  assign n152 = ~x2 & n151 ;
  assign n153 = x6 | x8 ;
  assign n154 = ~x0 & x6 ;
  assign n155 = x2 | n154 ;
  assign n156 = n124 & n155 ;
  assign n157 = n153 & ~n156 ;
  assign n158 = x9 | n157 ;
  assign n159 = ~n152 & n158 ;
  assign n160 = x1 & ~n159 ;
  assign n161 = n47 & n106 ;
  assign n162 = n160 | n161 ;
  assign n163 = ~x4 & n162 ;
  assign n164 = n147 | n163 ;
  assign n165 = ~x3 & n164 ;
  assign n166 = x3 & n25 ;
  assign n167 = ( x5 & n75 ) | ( x5 & n166 ) | ( n75 & n166 ) ;
  assign n168 = x1 & x5 ;
  assign n169 = x1 | x8 ;
  assign n170 = ~x2 & x3 ;
  assign n171 = x0 & n170 ;
  assign n172 = ( n168 & ~n169 ) | ( n168 & n171 ) | ( ~n169 & n171 ) ;
  assign n173 = ( x0 & n168 ) | ( x0 & n172 ) | ( n168 & n172 ) ;
  assign n174 = n167 | n173 ;
  assign n175 = x6 & n174 ;
  assign n176 = n141 & n166 ;
  assign n177 = n175 | n176 ;
  assign n178 = ( x4 & x9 ) | ( x4 & ~n177 ) | ( x9 & ~n177 ) ;
  assign n179 = x5 & ~n133 ;
  assign n180 = x3 | x8 ;
  assign n181 = ~n124 & n180 ;
  assign n182 = x0 & n181 ;
  assign n183 = n179 | n182 ;
  assign n184 = ~x1 & n183 ;
  assign n185 = ~x2 & x8 ;
  assign n186 = x0 & n185 ;
  assign n187 = ( x0 & ~x5 ) | ( x0 & n186 ) | ( ~x5 & n186 ) ;
  assign n188 = ( x1 & n148 ) | ( x1 & n187 ) | ( n148 & n187 ) ;
  assign n189 = x3 & x8 ;
  assign n190 = n55 | n189 ;
  assign n191 = ( ~x0 & n188 ) | ( ~x0 & n190 ) | ( n188 & n190 ) ;
  assign n192 = n184 | n191 ;
  assign n193 = ~x6 & n192 ;
  assign n194 = ~x1 & x8 ;
  assign n195 = x6 & n194 ;
  assign n196 = ( ~x2 & n169 ) | ( ~x2 & n195 ) | ( n169 & n195 ) ;
  assign n197 = x3 & n196 ;
  assign n198 = ~x0 & x8 ;
  assign n199 = x1 | x6 ;
  assign n200 = x0 & x1 ;
  assign n201 = n199 & ~n200 ;
  assign n202 = ~n198 & n201 ;
  assign n203 = ~x2 & n202 ;
  assign n204 = n197 | n203 ;
  assign n205 = ~x5 & n204 ;
  assign n206 = n193 | n205 ;
  assign n207 = ( ~x4 & x9 ) | ( ~x4 & n206 ) | ( x9 & n206 ) ;
  assign n208 = ~n178 & n207 ;
  assign n209 = n165 | n208 ;
  assign n210 = ~x7 & n209 ;
  assign n211 = x6 | n11 ;
  assign n212 = x2 & n48 ;
  assign n213 = n73 | n200 ;
  assign n214 = ~n212 & n213 ;
  assign n215 = ~x8 & n214 ;
  assign n216 = n19 & n185 ;
  assign n217 = n215 | n216 ;
  assign n218 = x7 & n217 ;
  assign n219 = n49 | n218 ;
  assign n220 = ~x4 & n219 ;
  assign n221 = n210 | n220 ;
  assign n222 = ( n210 & ~n211 ) | ( n210 & n221 ) | ( ~n211 & n221 ) ;
  assign n223 = x3 & x5 ;
  assign n224 = ( n47 & n123 ) | ( n47 & ~n223 ) | ( n123 & ~n223 ) ;
  assign n225 = ( n24 & n97 ) | ( n24 & n224 ) | ( n97 & n224 ) ;
  assign n226 = ~x3 & x9 ;
  assign n227 = n87 & ~n226 ;
  assign n228 = ( n31 & n194 ) | ( n31 & n227 ) | ( n194 & n227 ) ;
  assign n229 = n225 & ~n228 ;
  assign n230 = x0 & ~n229 ;
  assign n231 = x1 & x9 ;
  assign n232 = x2 & ~x5 ;
  assign n233 = x5 & ~x9 ;
  assign n234 = ( n231 & n232 ) | ( n231 & n233 ) | ( n232 & n233 ) ;
  assign n235 = ( x1 & n136 ) | ( x1 & n234 ) | ( n136 & n234 ) ;
  assign n236 = x8 & x9 ;
  assign n237 = n107 & ~n236 ;
  assign n238 = ( n30 & ~n87 ) | ( n30 & n237 ) | ( ~n87 & n237 ) ;
  assign n239 = n30 & n238 ;
  assign n240 = ( ~x3 & n235 ) | ( ~x3 & n239 ) | ( n235 & n239 ) ;
  assign n241 = n230 | n240 ;
  assign n242 = ~x6 & n241 ;
  assign n243 = x0 & ~x5 ;
  assign n244 = x2 & n231 ;
  assign n245 = ( x6 & n195 ) | ( x6 & n244 ) | ( n195 & n244 ) ;
  assign n246 = x2 & x8 ;
  assign n247 = n133 & ~n246 ;
  assign n248 = ( ~n149 & n236 ) | ( ~n149 & n247 ) | ( n236 & n247 ) ;
  assign n249 = n245 | n248 ;
  assign n250 = x3 & n249 ;
  assign n251 = n87 & ~n231 ;
  assign n252 = n180 | n251 ;
  assign n253 = ( x9 & n106 ) | ( x9 & n194 ) | ( n106 & n194 ) ;
  assign n254 = ( ~x8 & n252 ) | ( ~x8 & n253 ) | ( n252 & n253 ) ;
  assign n255 = x2 | n254 ;
  assign n256 = ~n250 & n255 ;
  assign n257 = n243 & ~n256 ;
  assign n258 = n242 | n257 ;
  assign n259 = ~x4 & n258 ;
  assign n260 = ~x3 & x4 ;
  assign n261 = ~x2 & n260 ;
  assign n262 = ~x1 & n261 ;
  assign n263 = x6 & ~x8 ;
  assign n264 = ( ~x5 & n236 ) | ( ~x5 & n263 ) | ( n236 & n263 ) ;
  assign n265 = n262 & ~n264 ;
  assign n266 = ( ~x1 & n65 ) | ( ~x1 & n189 ) | ( n65 & n189 ) ;
  assign n267 = x2 & x6 ;
  assign n268 = ( x2 & n67 ) | ( x2 & n267 ) | ( n67 & n267 ) ;
  assign n269 = n266 | n268 ;
  assign n270 = x5 & n269 ;
  assign n271 = x1 & n226 ;
  assign n272 = n263 & n271 ;
  assign n273 = ( x8 & n19 ) | ( x8 & n149 ) | ( n19 & n149 ) ;
  assign n274 = ( x6 & x9 ) | ( x6 & ~n273 ) | ( x9 & ~n273 ) ;
  assign n275 = ~x2 & n274 ;
  assign n276 = ~x3 & x8 ;
  assign n277 = ( n32 & n149 ) | ( n32 & n276 ) | ( n149 & n276 ) ;
  assign n278 = ( x3 & n275 ) | ( x3 & n277 ) | ( n275 & n277 ) ;
  assign n279 = n272 | n278 ;
  assign n280 = n270 | n279 ;
  assign n281 = n28 | n149 ;
  assign n282 = x6 | n226 ;
  assign n283 = n281 & ~n282 ;
  assign n284 = ( x8 & n232 ) | ( x8 & n276 ) | ( n232 & n276 ) ;
  assign n285 = x2 & x3 ;
  assign n286 = ( x3 & ~x8 ) | ( x3 & n285 ) | ( ~x8 & n285 ) ;
  assign n287 = x5 & ~n286 ;
  assign n288 = n284 | n287 ;
  assign n289 = x1 & n288 ;
  assign n290 = ( ~x8 & n88 ) | ( ~x8 & n114 ) | ( n88 & n114 ) ;
  assign n291 = ( ~n119 & n189 ) | ( ~n119 & n290 ) | ( n189 & n290 ) ;
  assign n292 = ( ~x9 & n289 ) | ( ~x9 & n291 ) | ( n289 & n291 ) ;
  assign n293 = n283 | n292 ;
  assign n294 = n280 | n293 ;
  assign n295 = ~x4 & n294 ;
  assign n296 = ( ~x0 & n265 ) | ( ~x0 & n295 ) | ( n265 & n295 ) ;
  assign n297 = ~x7 & n296 ;
  assign n298 = ( ~x7 & n259 ) | ( ~x7 & n297 ) | ( n259 & n297 ) ;
  assign n299 = x5 | x6 ;
  assign n300 = n75 | n299 ;
  assign n301 = n17 & ~n169 ;
  assign n302 = n41 & n58 ;
  assign n303 = ( x1 & ~n29 ) | ( x1 & n302 ) | ( ~n29 & n302 ) ;
  assign n304 = ( ~x4 & n301 ) | ( ~x4 & n303 ) | ( n301 & n303 ) ;
  assign n305 = ~n300 & n304 ;
  assign n306 = n298 | n305 ;
  assign n307 = x3 & ~n140 ;
  assign n308 = n267 | n307 ;
  assign n309 = ~x4 & n308 ;
  assign n310 = x5 | n236 ;
  assign n311 = ( n112 & n128 ) | ( n112 & n310 ) | ( n128 & n310 ) ;
  assign n312 = n261 & n311 ;
  assign n313 = n309 | n312 ;
  assign n314 = ~x1 & n313 ;
  assign n315 = ~x8 & n113 ;
  assign n316 = ~n106 & n223 ;
  assign n317 = ( x3 & n315 ) | ( x3 & ~n316 ) | ( n315 & ~n316 ) ;
  assign n318 = x5 & x8 ;
  assign n319 = ( x2 & ~x9 ) | ( x2 & n318 ) | ( ~x9 & n318 ) ;
  assign n320 = ( ~n123 & n140 ) | ( ~n123 & n319 ) | ( n140 & n319 ) ;
  assign n321 = n317 | n320 ;
  assign n322 = x1 & n321 ;
  assign n323 = x2 & n113 ;
  assign n324 = n322 | n323 ;
  assign n325 = ~x4 & n324 ;
  assign n326 = n314 | n325 ;
  assign n327 = ~x0 & n326 ;
  assign n328 = x3 & ~x8 ;
  assign n329 = x6 | n328 ;
  assign n330 = x3 & ~x5 ;
  assign n331 = n329 & ~n330 ;
  assign n332 = x5 & x9 ;
  assign n333 = x8 | n332 ;
  assign n334 = ( ~n133 & n170 ) | ( ~n133 & n333 ) | ( n170 & n333 ) ;
  assign n335 = n331 | n334 ;
  assign n336 = ( x2 & x9 ) | ( x2 & n181 ) | ( x9 & n181 ) ;
  assign n337 = n319 & ~n336 ;
  assign n338 = n335 | n337 ;
  assign n339 = x1 & n338 ;
  assign n340 = ~x3 & n113 ;
  assign n341 = n179 & ~n199 ;
  assign n342 = n340 | n341 ;
  assign n343 = ~x9 & n342 ;
  assign n344 = n339 | n343 ;
  assign n345 = x0 & n344 ;
  assign n346 = x2 & n88 ;
  assign n347 = ( n75 & n113 ) | ( n75 & n346 ) | ( n113 & n346 ) ;
  assign n348 = x9 & n347 ;
  assign n349 = n290 | n348 ;
  assign n350 = ~x1 & n349 ;
  assign n351 = n39 & n153 ;
  assign n352 = x2 | n351 ;
  assign n353 = x6 | n332 ;
  assign n354 = n231 | n318 ;
  assign n355 = ~n353 & n354 ;
  assign n356 = n352 & ~n355 ;
  assign n357 = x3 & ~n356 ;
  assign n358 = n113 & n273 ;
  assign n359 = n357 | n358 ;
  assign n360 = n350 | n359 ;
  assign n361 = n345 | n360 ;
  assign n362 = ~x4 & n361 ;
  assign n363 = n327 | n362 ;
  assign n364 = ~x7 & n363 ;
  assign n365 = x3 & ~x4 ;
  assign n366 = x1 | x2 ;
  assign n367 = x0 | n366 ;
  assign n368 = ( x3 & x4 ) | ( x3 & n367 ) | ( x4 & n367 ) ;
  assign n369 = x4 | n212 ;
  assign n370 = ( n365 & ~n368 ) | ( n365 & n369 ) | ( ~n368 & n369 ) ;
  assign n371 = ~x7 & n370 ;
  assign n372 = n112 & n371 ;
  assign n373 = ~n48 & n261 ;
  assign n374 = n365 & n367 ;
  assign n375 = n373 | n374 ;
  assign n376 = ~x7 & n375 ;
  assign n377 = n112 & n376 ;
  assign n378 = ( x6 & n30 ) | ( x6 & n112 ) | ( n30 & n112 ) ;
  assign n379 = ( ~n232 & n373 ) | ( ~n232 & n378 ) | ( n373 & n378 ) ;
  assign n380 = ~x7 & n379 ;
  assign n381 = x0 | x8 ;
  assign n382 = ~n243 & n381 ;
  assign n383 = n19 & n382 ;
  assign n384 = x0 & n127 ;
  assign n385 = ( ~x2 & n67 ) | ( ~x2 & n384 ) | ( n67 & n384 ) ;
  assign n386 = ( n149 & n198 ) | ( n149 & n200 ) | ( n198 & n200 ) ;
  assign n387 = ( x9 & n385 ) | ( x9 & n386 ) | ( n385 & n386 ) ;
  assign n388 = n383 | n387 ;
  assign n389 = x0 | x6 ;
  assign n390 = n169 & ~n389 ;
  assign n391 = n251 & n390 ;
  assign n392 = ~x5 & n391 ;
  assign n393 = ( n14 & ~n80 ) | ( n14 & n301 ) | ( ~n80 & n301 ) ;
  assign n394 = ( ~x5 & n392 ) | ( ~x5 & n393 ) | ( n392 & n393 ) ;
  assign n395 = n388 | n394 ;
  assign n396 = x3 & n395 ;
  assign n397 = n13 & n246 ;
  assign n398 = x2 & ~n397 ;
  assign n399 = ~x9 & n263 ;
  assign n400 = n29 & ~n149 ;
  assign n401 = ( n263 & ~n351 ) | ( n263 & n400 ) | ( ~n351 & n400 ) ;
  assign n402 = ( n389 & n399 ) | ( n389 & n401 ) | ( n399 & n401 ) ;
  assign n403 = ( n397 & ~n398 ) | ( n397 & n402 ) | ( ~n398 & n402 ) ;
  assign n404 = ~x1 & n403 ;
  assign n405 = ~x2 & x5 ;
  assign n406 = ~n59 & n405 ;
  assign n407 = x6 | n232 ;
  assign n408 = n13 & n407 ;
  assign n409 = n406 | n408 ;
  assign n410 = ~x8 & n409 ;
  assign n411 = x0 & x8 ;
  assign n412 = n125 | n198 ;
  assign n413 = ( n267 & n411 ) | ( n267 & n412 ) | ( n411 & n412 ) ;
  assign n414 = x1 & n413 ;
  assign n415 = ( x1 & n410 ) | ( x1 & n414 ) | ( n410 & n414 ) ;
  assign n416 = n404 | n415 ;
  assign n417 = n396 | n416 ;
  assign n418 = ~x7 & n417 ;
  assign n419 = x3 | x4 ;
  assign n420 = x6 | x9 ;
  assign n421 = x1 | x5 ;
  assign n422 = ( x2 & n420 ) | ( x2 & n421 ) | ( n420 & n421 ) ;
  assign n423 = n420 | n422 ;
  assign n424 = ( n17 & n60 ) | ( n17 & n332 ) | ( n60 & n332 ) ;
  assign n425 = ( x0 & ~n423 ) | ( x0 & n424 ) | ( ~n423 & n424 ) ;
  assign n426 = ~x0 & x2 ;
  assign n427 = ( n318 & n397 ) | ( n318 & n426 ) | ( n397 & n426 ) ;
  assign n428 = ( x8 & n425 ) | ( x8 & n427 ) | ( n425 & n427 ) ;
  assign n429 = x6 & ~n237 ;
  assign n430 = ~x2 & x9 ;
  assign n431 = n47 | n430 ;
  assign n432 = n429 & ~n431 ;
  assign n433 = ( n57 & n79 ) | ( n57 & ~n97 ) | ( n79 & ~n97 ) ;
  assign n434 = n432 | n433 ;
  assign n435 = n428 | n434 ;
  assign n436 = ~x7 & n435 ;
  assign n437 = n231 & n411 ;
  assign n438 = ( x7 & ~n107 ) | ( x7 & n437 ) | ( ~n107 & n437 ) ;
  assign n439 = ~x2 & n438 ;
  assign n440 = ~x9 & n41 ;
  assign n441 = ( ~x8 & n65 ) | ( ~x8 & n440 ) | ( n65 & n440 ) ;
  assign n442 = ( ~x0 & n81 ) | ( ~x0 & n441 ) | ( n81 & n441 ) ;
  assign n443 = n439 | n442 ;
  assign n444 = ~n299 & n443 ;
  assign n445 = ( ~n419 & n436 ) | ( ~n419 & n444 ) | ( n436 & n444 ) ;
  assign n446 = ~n419 & n445 ;
  assign n447 = ( ~x4 & n418 ) | ( ~x4 & n446 ) | ( n418 & n446 ) ;
  assign n448 = n380 | n447 ;
  assign n449 = ~x6 & n180 ;
  assign n450 = ( ~n153 & n307 ) | ( ~n153 & n449 ) | ( n307 & n449 ) ;
  assign n451 = ( x0 & n449 ) | ( x0 & n450 ) | ( n449 & n450 ) ;
  assign n452 = ( n30 & n236 ) | ( n30 & n328 ) | ( n236 & n328 ) ;
  assign n453 = ( x2 & n451 ) | ( x2 & n452 ) | ( n451 & n452 ) ;
  assign n454 = x3 | n108 ;
  assign n455 = ~n453 & n454 ;
  assign n456 = ( x6 & x8 ) | ( x6 & x9 ) | ( x8 & x9 ) ;
  assign n457 = ( x9 & n282 ) | ( x9 & n451 ) | ( n282 & n451 ) ;
  assign n458 = ( n149 & n456 ) | ( n149 & ~n457 ) | ( n456 & ~n457 ) ;
  assign n459 = ( n45 & n125 ) | ( n45 & n276 ) | ( n125 & n276 ) ;
  assign n460 = n45 & n459 ;
  assign n461 = ( ~x2 & n458 ) | ( ~x2 & n460 ) | ( n458 & n460 ) ;
  assign n462 = n455 & ~n461 ;
  assign n463 = n170 & n399 ;
  assign n464 = ( x1 & ~n462 ) | ( x1 & n463 ) | ( ~n462 & n463 ) ;
  assign n465 = x2 | x6 ;
  assign n466 = n400 | n465 ;
  assign n467 = n154 & ~n237 ;
  assign n468 = n466 & ~n467 ;
  assign n469 = x3 & ~n468 ;
  assign n470 = n134 & ~n384 ;
  assign n471 = x9 | n470 ;
  assign n472 = x2 & n107 ;
  assign n473 = ~n449 & n472 ;
  assign n474 = n471 & ~n473 ;
  assign n475 = ~n469 & n474 ;
  assign n476 = ( x1 & ~n463 ) | ( x1 & n475 ) | ( ~n463 & n475 ) ;
  assign n477 = ~n464 & n476 ;
  assign n478 = x5 | n477 ;
  assign n479 = n170 & n233 ;
  assign n480 = n47 | n223 ;
  assign n481 = ~x0 & n480 ;
  assign n482 = ( x8 & n179 ) | ( x8 & n328 ) | ( n179 & n328 ) ;
  assign n483 = ( ~x8 & n481 ) | ( ~x8 & n482 ) | ( n481 & n482 ) ;
  assign n484 = n479 | n483 ;
  assign n485 = n86 & n141 ;
  assign n486 = ( x0 & x8 ) | ( x0 & n233 ) | ( x8 & n233 ) ;
  assign n487 = ( ~x0 & x8 ) | ( ~x0 & n431 ) | ( x8 & n431 ) ;
  assign n488 = n486 & n487 ;
  assign n489 = ( ~x3 & n485 ) | ( ~x3 & n488 ) | ( n485 & n488 ) ;
  assign n490 = n484 | n489 ;
  assign n491 = x1 & n490 ;
  assign n492 = x5 & n285 ;
  assign n493 = ( x2 & n171 ) | ( x2 & ~n237 ) | ( n171 & ~n237 ) ;
  assign n494 = ( x5 & n492 ) | ( x5 & n493 ) | ( n492 & n493 ) ;
  assign n495 = ( n28 & n285 ) | ( n28 & n301 ) | ( n285 & n301 ) ;
  assign n496 = ( ~x1 & n494 ) | ( ~x1 & n495 ) | ( n494 & n495 ) ;
  assign n497 = ( n179 & n236 ) | ( n179 & n492 ) | ( n236 & n492 ) ;
  assign n498 = n496 | n497 ;
  assign n499 = ~x6 & n498 ;
  assign n500 = ( ~x6 & n491 ) | ( ~x6 & n499 ) | ( n491 & n499 ) ;
  assign n501 = ~x7 & n500 ;
  assign n502 = ( x7 & n478 ) | ( x7 & ~n501 ) | ( n478 & ~n501 ) ;
  assign n503 = x4 & ~x7 ;
  assign n504 = ~n11 & n503 ;
  assign n505 = ~n367 & n504 ;
  assign n506 = ~x6 & n505 ;
  assign n507 = x4 & ~n506 ;
  assign n508 = n11 | n199 ;
  assign n509 = ( n45 & n426 ) | ( n45 & n440 ) | ( n426 & n440 ) ;
  assign n510 = ( n237 & n426 ) | ( n237 & n509 ) | ( n426 & n509 ) ;
  assign n511 = ~n508 & n510 ;
  assign n512 = ( n506 & ~n507 ) | ( n506 & n511 ) | ( ~n507 & n511 ) ;
  assign n513 = ( n502 & n507 ) | ( n502 & ~n512 ) | ( n507 & ~n512 ) ;
  assign n514 = ~n134 & n231 ;
  assign n515 = x1 & ~n514 ;
  assign n516 = x0 | n247 ;
  assign n517 = ( x9 & ~n186 ) | ( x9 & n516 ) | ( ~n186 & n516 ) ;
  assign n518 = ( n65 & n68 ) | ( n65 & n514 ) | ( n68 & n514 ) ;
  assign n519 = ( n515 & n517 ) | ( n515 & ~n518 ) | ( n517 & ~n518 ) ;
  assign n520 = n211 | n519 ;
  assign n521 = n168 | n330 ;
  assign n522 = ~x2 & n96 ;
  assign n523 = ~n521 & n522 ;
  assign n524 = ~n119 & n243 ;
  assign n525 = x8 & n524 ;
  assign n526 = ( x8 & n523 ) | ( x8 & n525 ) | ( n523 & n525 ) ;
  assign n527 = ( n289 & n426 ) | ( n289 & n524 ) | ( n426 & n524 ) ;
  assign n528 = ( n25 & n287 ) | ( n25 & n527 ) | ( n287 & n527 ) ;
  assign n529 = ~x9 & n528 ;
  assign n530 = ( ~x9 & n526 ) | ( ~x9 & n529 ) | ( n526 & n529 ) ;
  assign n531 = ( n223 & n232 ) | ( n223 & ~n286 ) | ( n232 & ~n286 ) ;
  assign n532 = x1 & n531 ;
  assign n533 = n32 & ~n148 ;
  assign n534 = n185 & n533 ;
  assign n535 = x9 & n534 ;
  assign n536 = ( x9 & n532 ) | ( x9 & n535 ) | ( n532 & n535 ) ;
  assign n537 = n530 | n536 ;
  assign n538 = n227 & ~n521 ;
  assign n539 = ~x2 & n538 ;
  assign n540 = n30 & ~n421 ;
  assign n541 = ( n30 & ~n251 ) | ( n30 & n540 ) | ( ~n251 & n540 ) ;
  assign n542 = n539 | n541 ;
  assign n543 = n233 & ~n366 ;
  assign n544 = ( n271 & ~n381 ) | ( n271 & n543 ) | ( ~n381 & n543 ) ;
  assign n545 = ~n381 & n544 ;
  assign n546 = ( ~x8 & n542 ) | ( ~x8 & n545 ) | ( n542 & n545 ) ;
  assign n547 = n537 | n546 ;
  assign n548 = x6 & ~n12 ;
  assign n549 = ( ~x8 & n273 ) | ( ~x8 & n548 ) | ( n273 & n548 ) ;
  assign n550 = n268 | n549 ;
  assign n551 = ( n200 & n301 ) | ( n200 & n465 ) | ( n301 & n465 ) ;
  assign n552 = ( x0 & n548 ) | ( x0 & n551 ) | ( n548 & n551 ) ;
  assign n553 = n550 | n552 ;
  assign n554 = n330 & n553 ;
  assign n555 = x6 & ~n554 ;
  assign n556 = ( n547 & n554 ) | ( n547 & ~n555 ) | ( n554 & ~n555 ) ;
  assign n557 = ~x7 & n520 ;
  assign n558 = n556 & n557 ;
  assign n559 = ( x4 & n520 ) | ( x4 & ~n558 ) | ( n520 & ~n558 ) ;
  assign n560 = ~n505 & n559 ;
  assign n561 = ( n125 & n353 ) | ( n125 & n412 ) | ( n353 & n412 ) ;
  assign n562 = ( x3 & n299 ) | ( x3 & n419 ) | ( n299 & n419 ) ;
  assign n563 = ~x3 & n562 ;
  assign n564 = ( ~n561 & n562 ) | ( ~n561 & n563 ) | ( n562 & n563 ) ;
  assign n565 = x2 | n564 ;
  assign n566 = ~x3 & n39 ;
  assign n567 = ( ~n65 & n333 ) | ( ~n65 & n566 ) | ( n333 & n566 ) ;
  assign n568 = n65 & n567 ;
  assign n569 = ( x1 & n565 ) | ( x1 & ~n568 ) | ( n565 & ~n568 ) ;
  assign n570 = ~n378 & n569 ;
  assign n571 = x7 & ~n30 ;
  assign n572 = ( x6 & n153 ) | ( x6 & n332 ) | ( n153 & n332 ) ;
  assign n573 = ~x3 & n572 ;
  assign n574 = ~n310 & n346 ;
  assign n575 = n573 | n574 ;
  assign n576 = ~x2 & n566 ;
  assign n577 = ( n198 & n276 ) | ( n198 & n467 ) | ( n276 & n467 ) ;
  assign n578 = ( ~x2 & n576 ) | ( ~x2 & n577 ) | ( n576 & n577 ) ;
  assign n579 = n575 | n578 ;
  assign n580 = x1 & n579 ;
  assign n581 = n571 | n580 ;
  assign n582 = n570 & ~n581 ;
  assign n583 = ~x1 & n107 ;
  assign n584 = x7 | n243 ;
  assign n585 = ( x7 & n346 ) | ( x7 & n584 ) | ( n346 & n584 ) ;
  assign n586 = ~n583 & n585 ;
  assign n587 = x2 | n119 ;
  assign n588 = ~x7 & n587 ;
  assign n589 = x0 & ~n588 ;
  assign n590 = n586 | n589 ;
  assign n591 = x4 & n587 ;
  assign n592 = n590 | n591 ;
  assign n593 = n582 & ~n592 ;
  assign n594 = ( ~x8 & n14 ) | ( ~x8 & n18 ) | ( n14 & n18 ) ;
  assign n595 = n365 & n594 ;
  assign n596 = x2 & n595 ;
  assign n597 = n373 | n596 ;
  assign n598 = ~x7 & n597 ;
  assign n599 = ~n299 & n598 ;
  assign y0 = ~n122 ;
  assign y1 = n222 ;
  assign y2 = n306 ;
  assign y3 = n364 ;
  assign y4 = n372 ;
  assign y5 = n377 ;
  assign y6 = ~n448 ;
  assign y7 = n513 ;
  assign y8 = n560 ;
  assign y9 = n593 ;
  assign y10 = n599 ;
endmodule
