module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 ;
  assign n8 = x0 & ~x1 ;
  assign n9 = x3 & x4 ;
  assign n10 = n8 & n9 ;
  assign n11 = x1 & n9 ;
  assign n12 = n10 | n11 ;
  assign n13 = ~x2 & n12 ;
  assign n14 = x3 | x4 ;
  assign n15 = ~n9 & n14 ;
  assign n16 = x1 & ~n15 ;
  assign n17 = ~x1 & n9 ;
  assign n18 = n16 | n17 ;
  assign n19 = x2 & n18 ;
  assign n20 = n13 | n19 ;
  assign n21 = ~x3 & n14 ;
  assign n22 = x1 & ~n21 ;
  assign n23 = ( x1 & ~n8 ) | ( x1 & n9 ) | ( ~n8 & n9 ) ;
  assign n24 = ~n22 & n23 ;
  assign n25 = x2 | n24 ;
  assign n26 = ~x3 & x4 ;
  assign n27 = x1 & x3 ;
  assign n28 = ( x1 & n26 ) | ( x1 & n27 ) | ( n26 & n27 ) ;
  assign n29 = x1 & ~n28 ;
  assign n30 = x2 & ~n29 ;
  assign n31 = n25 & ~n30 ;
  assign n32 = x0 | n9 ;
  assign n33 = n14 & ~n32 ;
  assign n34 = x0 & ~x3 ;
  assign n35 = ( x0 & n9 ) | ( x0 & n34 ) | ( n9 & n34 ) ;
  assign n36 = ( x0 & n33 ) | ( x0 & ~n35 ) | ( n33 & ~n35 ) ;
  assign n37 = x1 & ~n36 ;
  assign n38 = n23 & ~n37 ;
  assign n39 = ~x2 & n38 ;
  assign n40 = x0 & ~n15 ;
  assign n41 = x0 | x3 ;
  assign n42 = n26 | n41 ;
  assign n43 = ~n40 & n42 ;
  assign n44 = x1 & ~x2 ;
  assign n45 = ( x2 & n43 ) | ( x2 & ~n44 ) | ( n43 & ~n44 ) ;
  assign n46 = ( x2 & n21 ) | ( x2 & n44 ) | ( n21 & n44 ) ;
  assign n47 = ( ~x2 & n45 ) | ( ~x2 & n46 ) | ( n45 & n46 ) ;
  assign n48 = x3 & ~x5 ;
  assign n49 = ~n9 & n48 ;
  assign n50 = x3 & x5 ;
  assign n51 = x6 & n50 ;
  assign n52 = ( x6 & n49 ) | ( x6 & n51 ) | ( n49 & n51 ) ;
  assign n53 = x3 & ~x6 ;
  assign n54 = ~n9 & n53 ;
  assign n55 = x0 & n54 ;
  assign n56 = ( x0 & n52 ) | ( x0 & n55 ) | ( n52 & n55 ) ;
  assign n57 = x1 | x2 ;
  assign n58 = ~x0 & x3 ;
  assign n59 = x4 & x5 ;
  assign n60 = n58 & n59 ;
  assign n61 = ( x2 & n57 ) | ( x2 & n60 ) | ( n57 & n60 ) ;
  assign n62 = x0 & x3 ;
  assign n63 = ( x0 & ~n14 ) | ( x0 & n62 ) | ( ~n14 & n62 ) ;
  assign n64 = ~x0 & x2 ;
  assign n65 = ( x2 & n63 ) | ( x2 & n64 ) | ( n63 & n64 ) ;
  assign n66 = n61 & ~n65 ;
  assign n67 = n57 & ~n65 ;
  assign n68 = ( n56 & n66 ) | ( n56 & n67 ) | ( n66 & n67 ) ;
  assign n69 = x3 & x6 ;
  assign n70 = n54 | n69 ;
  assign n71 = ( x1 & x2 ) | ( x1 & n70 ) | ( x2 & n70 ) ;
  assign n72 = ( ~x1 & x2 ) | ( ~x1 & n22 ) | ( x2 & n22 ) ;
  assign n73 = n71 & ~n72 ;
  assign n74 = x2 & n9 ;
  assign n75 = ( x0 & n26 ) | ( x0 & n62 ) | ( n26 & n62 ) ;
  assign n76 = n33 | n75 ;
  assign n77 = x1 & n76 ;
  assign n78 = x1 | n9 ;
  assign n79 = n14 & ~n78 ;
  assign n80 = x2 | n79 ;
  assign n81 = n77 | n80 ;
  assign n82 = ( ~x2 & n74 ) | ( ~x2 & n81 ) | ( n74 & n81 ) ;
  assign n83 = x1 & ~n42 ;
  assign n84 = ( x1 & n40 ) | ( x1 & n83 ) | ( n40 & n83 ) ;
  assign n85 = n23 & ~n57 ;
  assign n86 = x2 & n10 ;
  assign n87 = n85 | n86 ;
  assign n88 = x2 | n85 ;
  assign n89 = ( n84 & n87 ) | ( n84 & n88 ) | ( n87 & n88 ) ;
  assign n90 = ( x0 & n14 ) | ( x0 & ~n58 ) | ( n14 & ~n58 ) ;
  assign n91 = ~x0 & n90 ;
  assign n92 = ( x1 & x2 ) | ( x1 & n91 ) | ( x2 & n91 ) ;
  assign n93 = ( ~x1 & x2 ) | ( ~x1 & n15 ) | ( x2 & n15 ) ;
  assign n94 = n92 & ~n93 ;
  assign n95 = x1 & ~n91 ;
  assign n96 = n78 & ~n95 ;
  assign n97 = x2 | n96 ;
  assign n98 = ~n30 & n97 ;
  assign n99 = x2 & ~n21 ;
  assign n100 = n58 | n75 ;
  assign n101 = x1 & n100 ;
  assign n102 = n80 | n101 ;
  assign n103 = ~n99 & n102 ;
  assign n104 = x3 | n26 ;
  assign n105 = ~x0 & n104 ;
  assign n106 = x0 | n105 ;
  assign n107 = x2 | n106 ;
  assign n108 = x1 | n107 ;
  assign n109 = ( x1 & x2 ) | ( x1 & x4 ) | ( x2 & x4 ) ;
  assign n110 = ( x1 & ~x2 ) | ( x1 & x3 ) | ( ~x2 & x3 ) ;
  assign n111 = ( ~n9 & n44 ) | ( ~n9 & n110 ) | ( n44 & n110 ) ;
  assign n112 = n109 & ~n111 ;
  assign n113 = ~x1 & n58 ;
  assign n114 = ( ~x1 & n75 ) | ( ~x1 & n113 ) | ( n75 & n113 ) ;
  assign n115 = ~x2 & n28 ;
  assign n116 = ( ~x2 & n114 ) | ( ~x2 & n115 ) | ( n114 & n115 ) ;
  assign n117 = n112 | n116 ;
  assign n118 = x2 & ~n75 ;
  assign n119 = x0 & n118 ;
  assign n120 = x2 & n106 ;
  assign n121 = x2 & ~n120 ;
  assign n122 = x3 & ~n9 ;
  assign n123 = ~x0 & n122 ;
  assign n124 = x2 & n123 ;
  assign n125 = ~x1 & n124 ;
  assign n126 = x0 | x1 ;
  assign n127 = x2 & n126 ;
  assign n128 = x1 & x2 ;
  assign n129 = ( ~n35 & n127 ) | ( ~n35 & n128 ) | ( n127 & n128 ) ;
  assign n130 = ~x1 & n129 ;
  assign n131 = x0 & x1 ;
  assign n132 = ( ~x2 & n35 ) | ( ~x2 & n131 ) | ( n35 & n131 ) ;
  assign n133 = n131 & ~n132 ;
  assign n134 = x1 & n124 ;
  assign n135 = x2 & ~n104 ;
  assign n136 = n49 | n50 ;
  assign n137 = n131 & n136 ;
  assign n138 = n8 & ~n35 ;
  assign n139 = x2 | n138 ;
  assign n140 = n137 | n139 ;
  assign n141 = n9 & ~n131 ;
  assign n142 = x2 & ~n141 ;
  assign n143 = n140 & ~n142 ;
  assign n144 = x0 & x5 ;
  assign n145 = ( x6 & ~n9 ) | ( x6 & n144 ) | ( ~n9 & n144 ) ;
  assign n146 = n144 & ~n145 ;
  assign n147 = x1 & ~n146 ;
  assign n148 = ( x1 & ~n35 ) | ( x1 & n126 ) | ( ~n35 & n126 ) ;
  assign n149 = ~n147 & n148 ;
  assign n150 = ~x2 & n149 ;
  assign n151 = n54 & n131 ;
  assign n152 = ( n52 & n131 ) | ( n52 & n151 ) | ( n131 & n151 ) ;
  assign n153 = x2 & ~n142 ;
  assign n154 = ( ~n142 & n152 ) | ( ~n142 & n153 ) | ( n152 & n153 ) ;
  assign n155 = ( x1 & ~n8 ) | ( x1 & n90 ) | ( ~n8 & n90 ) ;
  assign n156 = x0 & ~n63 ;
  assign n157 = x1 & ~n156 ;
  assign n158 = n155 & ~n157 ;
  assign n159 = ~x2 & n158 ;
  assign n160 = ( x2 & n8 ) | ( x2 & n63 ) | ( n8 & n63 ) ;
  assign n161 = n8 & ~n160 ;
  assign y0 = n20 ;
  assign y1 = n31 ;
  assign y2 = n39 ;
  assign y3 = n47 ;
  assign y4 = n68 ;
  assign y5 = n73 ;
  assign y6 = n82 ;
  assign y7 = n89 ;
  assign y8 = n94 ;
  assign y9 = n98 ;
  assign y10 = n103 ;
  assign y11 = ~n108 ;
  assign y12 = n117 ;
  assign y13 = n119 ;
  assign y14 = n121 ;
  assign y15 = n125 ;
  assign y16 = n130 ;
  assign y17 = n133 ;
  assign y18 = n134 ;
  assign y19 = n135 ;
  assign y20 = n143 ;
  assign y21 = n150 ;
  assign y22 = n154 ;
  assign y23 = ~1'b0 ;
  assign y24 = n159 ;
  assign y25 = n161 ;
endmodule
