module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 ;
  assign n129 = x0 & x64 ;
  assign n130 = x2 & ~n129 ;
  assign n131 = x2 | n129 ;
  assign n132 = ~n130 & n131 ;
  assign n133 = ~x0 & x1 ;
  assign n134 = x64 & n133 ;
  assign n135 = ~x1 & x2 ;
  assign n136 = x1 & ~x2 ;
  assign n137 = n135 | n136 ;
  assign n138 = x0 & x65 ;
  assign n139 = ~n137 & n138 ;
  assign n140 = n134 | n139 ;
  assign n141 = x0 & n137 ;
  assign n142 = x64 & ~x65 ;
  assign n143 = ~x64 & x65 ;
  assign n144 = n142 | n143 ;
  assign n145 = n141 & n144 ;
  assign n146 = n140 | n145 ;
  assign n147 = x2 & ~n146 ;
  assign n148 = ~x2 & n146 ;
  assign n149 = n147 | n148 ;
  assign n150 = n130 | n149 ;
  assign n151 = n130 & n149 ;
  assign n152 = n150 & ~n151 ;
  assign n153 = x65 & ~x66 ;
  assign n154 = x64 & n153 ;
  assign n155 = x65 & x66 ;
  assign n156 = x64 & x65 ;
  assign n157 = ( x66 & ~n155 ) | ( x66 & n156 ) | ( ~n155 & n156 ) ;
  assign n158 = ( x65 & ~n155 ) | ( x65 & n157 ) | ( ~n155 & n157 ) ;
  assign n159 = ~n154 & n158 ;
  assign n160 = n141 & n159 ;
  assign n161 = x65 & n133 ;
  assign n162 = x0 | x1 ;
  assign n163 = x64 & ~n162 ;
  assign n164 = ( n137 & n161 ) | ( n137 & n163 ) | ( n161 & n163 ) ;
  assign n165 = x0 & x66 ;
  assign n166 = ( ~n137 & n161 ) | ( ~n137 & n165 ) | ( n161 & n165 ) ;
  assign n167 = n164 | n166 ;
  assign n168 = x2 & ~n167 ;
  assign n169 = ~n160 & n168 ;
  assign n170 = ~x2 & n167 ;
  assign n171 = ( ~x2 & n160 ) | ( ~x2 & n170 ) | ( n160 & n170 ) ;
  assign n172 = n169 | n171 ;
  assign n173 = n151 & n172 ;
  assign n174 = n151 | n172 ;
  assign n175 = ~n173 & n174 ;
  assign n176 = x2 & ~x3 ;
  assign n177 = ~x2 & x3 ;
  assign n178 = n176 | n177 ;
  assign n179 = x64 & n178 ;
  assign n180 = n154 | n155 ;
  assign n181 = x66 | x67 ;
  assign n182 = x66 & x67 ;
  assign n183 = n181 & ~n182 ;
  assign n184 = n180 & n183 ;
  assign n185 = n180 | n183 ;
  assign n186 = ~n184 & n185 ;
  assign n187 = x66 & n133 ;
  assign n188 = x65 & ~n162 ;
  assign n189 = ( n137 & n187 ) | ( n137 & n188 ) | ( n187 & n188 ) ;
  assign n190 = x0 & x67 ;
  assign n191 = ( ~n137 & n187 ) | ( ~n137 & n190 ) | ( n187 & n190 ) ;
  assign n192 = n189 | n191 ;
  assign n193 = n141 | n192 ;
  assign n194 = ( n186 & n192 ) | ( n186 & n193 ) | ( n192 & n193 ) ;
  assign n195 = x2 | n194 ;
  assign n196 = ~x2 & n194 ;
  assign n197 = ( ~n194 & n195 ) | ( ~n194 & n196 ) | ( n195 & n196 ) ;
  assign n198 = n179 & n197 ;
  assign n199 = n179 | n197 ;
  assign n200 = ~n198 & n199 ;
  assign n201 = n173 & n200 ;
  assign n202 = n173 | n200 ;
  assign n203 = ~n201 & n202 ;
  assign n204 = ~x3 & x4 ;
  assign n205 = x3 & ~x4 ;
  assign n206 = n204 | n205 ;
  assign n207 = ~n178 & n206 ;
  assign n208 = x64 & n207 ;
  assign n209 = ~x4 & x5 ;
  assign n210 = x4 & ~x5 ;
  assign n211 = n209 | n210 ;
  assign n212 = n178 & ~n211 ;
  assign n213 = x65 & n212 ;
  assign n214 = n208 | n213 ;
  assign n215 = n178 & n211 ;
  assign n216 = x5 | n144 ;
  assign n217 = ( x5 & n215 ) | ( x5 & n216 ) | ( n215 & n216 ) ;
  assign n218 = ~x5 & n217 ;
  assign n219 = ( ~x5 & n214 ) | ( ~x5 & n218 ) | ( n214 & n218 ) ;
  assign n220 = x5 & ~x64 ;
  assign n221 = ( x5 & ~n178 ) | ( x5 & n220 ) | ( ~n178 & n220 ) ;
  assign n222 = n217 & n221 ;
  assign n223 = ( n214 & n221 ) | ( n214 & n222 ) | ( n221 & n222 ) ;
  assign n224 = n144 & n215 ;
  assign n225 = n221 & ~n224 ;
  assign n226 = ~n214 & n225 ;
  assign n227 = ( n219 & n223 ) | ( n219 & n226 ) | ( n223 & n226 ) ;
  assign n228 = n217 | n221 ;
  assign n229 = n214 | n228 ;
  assign n230 = ~n221 & n224 ;
  assign n231 = ( n214 & ~n221 ) | ( n214 & n230 ) | ( ~n221 & n230 ) ;
  assign n232 = ( n219 & n229 ) | ( n219 & ~n231 ) | ( n229 & ~n231 ) ;
  assign n233 = ~n227 & n232 ;
  assign n234 = x67 | x68 ;
  assign n235 = x67 & x68 ;
  assign n236 = n234 & ~n235 ;
  assign n237 = n182 | n183 ;
  assign n238 = ( n180 & n182 ) | ( n180 & n237 ) | ( n182 & n237 ) ;
  assign n239 = n236 & n238 ;
  assign n240 = n236 | n238 ;
  assign n241 = ~n239 & n240 ;
  assign n242 = x67 & n133 ;
  assign n243 = x66 & ~n162 ;
  assign n244 = ( n137 & n242 ) | ( n137 & n243 ) | ( n242 & n243 ) ;
  assign n245 = x0 & x68 ;
  assign n246 = ( ~n137 & n242 ) | ( ~n137 & n245 ) | ( n242 & n245 ) ;
  assign n247 = n244 | n246 ;
  assign n248 = x2 & ~n247 ;
  assign n249 = x2 & ~n141 ;
  assign n250 = ~n247 & n249 ;
  assign n251 = ( ~n241 & n248 ) | ( ~n241 & n250 ) | ( n248 & n250 ) ;
  assign n252 = ~x2 & n247 ;
  assign n253 = ~x2 & n141 ;
  assign n254 = ( ~x2 & n247 ) | ( ~x2 & n253 ) | ( n247 & n253 ) ;
  assign n255 = ( n241 & n252 ) | ( n241 & n254 ) | ( n252 & n254 ) ;
  assign n256 = n251 | n255 ;
  assign n257 = n233 & n256 ;
  assign n258 = n233 & ~n257 ;
  assign n259 = ~n233 & n256 ;
  assign n260 = n258 | n259 ;
  assign n261 = n173 | n198 ;
  assign n262 = ( n198 & n200 ) | ( n198 & n261 ) | ( n200 & n261 ) ;
  assign n263 = n260 & n262 ;
  assign n264 = n260 | n262 ;
  assign n265 = ~n263 & n264 ;
  assign n266 = x65 & n207 ;
  assign n267 = ~n178 & n211 ;
  assign n268 = x64 & ~n206 ;
  assign n269 = n267 & n268 ;
  assign n270 = n266 | n269 ;
  assign n271 = x66 & n212 ;
  assign n272 = n270 | n271 ;
  assign n273 = ( n159 & n215 ) | ( n159 & n271 ) | ( n215 & n271 ) ;
  assign n274 = n159 | n215 ;
  assign n275 = ( n270 & n273 ) | ( n270 & n274 ) | ( n273 & n274 ) ;
  assign n276 = n272 | n275 ;
  assign n277 = x5 & ~n276 ;
  assign n278 = ~x5 & n276 ;
  assign n279 = n277 | n278 ;
  assign n280 = n227 & n279 ;
  assign n281 = n227 | n279 ;
  assign n282 = ~n280 & n281 ;
  assign n283 = x68 | x69 ;
  assign n284 = x68 & x69 ;
  assign n285 = n283 & ~n284 ;
  assign n286 = n235 | n236 ;
  assign n287 = n285 & n286 ;
  assign n288 = n235 & n285 ;
  assign n289 = ( n238 & n287 ) | ( n238 & n288 ) | ( n287 & n288 ) ;
  assign n290 = n285 | n286 ;
  assign n291 = n235 | n285 ;
  assign n292 = ( n238 & n290 ) | ( n238 & n291 ) | ( n290 & n291 ) ;
  assign n293 = ~n289 & n292 ;
  assign n294 = x68 & n133 ;
  assign n295 = x67 & ~n162 ;
  assign n296 = ( n137 & n294 ) | ( n137 & n295 ) | ( n294 & n295 ) ;
  assign n297 = x0 & x69 ;
  assign n298 = ( ~n137 & n294 ) | ( ~n137 & n297 ) | ( n294 & n297 ) ;
  assign n299 = n296 | n298 ;
  assign n300 = x2 & ~n299 ;
  assign n301 = n249 & ~n299 ;
  assign n302 = ( ~n293 & n300 ) | ( ~n293 & n301 ) | ( n300 & n301 ) ;
  assign n303 = ~x2 & n299 ;
  assign n304 = ( ~x2 & n253 ) | ( ~x2 & n299 ) | ( n253 & n299 ) ;
  assign n305 = ( n293 & n303 ) | ( n293 & n304 ) | ( n303 & n304 ) ;
  assign n306 = n302 | n305 ;
  assign n307 = n282 & n306 ;
  assign n308 = n282 & ~n307 ;
  assign n309 = ~n282 & n306 ;
  assign n310 = n308 | n309 ;
  assign n311 = n257 | n262 ;
  assign n312 = ( n257 & n260 ) | ( n257 & n311 ) | ( n260 & n311 ) ;
  assign n313 = n310 & n312 ;
  assign n314 = n310 | n312 ;
  assign n315 = ~n313 & n314 ;
  assign n316 = x5 & ~x6 ;
  assign n317 = ~x5 & x6 ;
  assign n318 = n316 | n317 ;
  assign n319 = x64 & n318 ;
  assign n320 = x67 & n212 ;
  assign n321 = x66 & n207 ;
  assign n322 = x65 & ~n206 ;
  assign n323 = n267 & n322 ;
  assign n324 = n321 | n323 ;
  assign n325 = n320 | n324 ;
  assign n326 = n186 & n215 ;
  assign n327 = n325 | n326 ;
  assign n328 = x5 & ~n327 ;
  assign n329 = ~x5 & n327 ;
  assign n330 = n328 | n329 ;
  assign n331 = ( n280 & ~n319 ) | ( n280 & n330 ) | ( ~n319 & n330 ) ;
  assign n332 = ( ~n280 & n319 ) | ( ~n280 & n331 ) | ( n319 & n331 ) ;
  assign n333 = x69 | x70 ;
  assign n334 = x69 & x70 ;
  assign n335 = n333 & ~n334 ;
  assign n336 = n284 & n335 ;
  assign n337 = ( n289 & n335 ) | ( n289 & n336 ) | ( n335 & n336 ) ;
  assign n338 = n284 | n335 ;
  assign n339 = n289 | n338 ;
  assign n340 = ~n337 & n339 ;
  assign n341 = x69 & n133 ;
  assign n342 = x68 & ~n162 ;
  assign n343 = ( n137 & n341 ) | ( n137 & n342 ) | ( n341 & n342 ) ;
  assign n344 = x0 & x70 ;
  assign n345 = ( ~n137 & n341 ) | ( ~n137 & n344 ) | ( n341 & n344 ) ;
  assign n346 = n343 | n345 ;
  assign n347 = ( n141 & n340 ) | ( n141 & n346 ) | ( n340 & n346 ) ;
  assign n348 = ( x2 & n141 ) | ( x2 & ~n346 ) | ( n141 & ~n346 ) ;
  assign n349 = ( x2 & n340 ) | ( x2 & n348 ) | ( n340 & n348 ) ;
  assign n350 = ~n347 & n349 ;
  assign n351 = n346 | n348 ;
  assign n352 = x2 | n346 ;
  assign n353 = ( n340 & n351 ) | ( n340 & n352 ) | ( n351 & n352 ) ;
  assign n354 = ( ~x2 & n350 ) | ( ~x2 & n353 ) | ( n350 & n353 ) ;
  assign n355 = n331 & n354 ;
  assign n356 = ~n330 & n354 ;
  assign n357 = ( n332 & n355 ) | ( n332 & n356 ) | ( n355 & n356 ) ;
  assign n358 = n331 | n354 ;
  assign n359 = n330 & ~n354 ;
  assign n360 = ( n332 & n358 ) | ( n332 & ~n359 ) | ( n358 & ~n359 ) ;
  assign n361 = ~n357 & n360 ;
  assign n362 = n307 | n312 ;
  assign n363 = ( n307 & n310 ) | ( n307 & n362 ) | ( n310 & n362 ) ;
  assign n364 = n361 & n363 ;
  assign n365 = n361 | n363 ;
  assign n366 = ~n364 & n365 ;
  assign n367 = n215 & n241 ;
  assign n368 = x68 & n212 ;
  assign n369 = x67 & n207 ;
  assign n370 = x66 & ~n206 ;
  assign n371 = n267 & n370 ;
  assign n372 = n369 | n371 ;
  assign n373 = n368 | n372 ;
  assign n374 = n367 | n373 ;
  assign n375 = x5 | n368 ;
  assign n376 = n372 | n375 ;
  assign n377 = n367 | n376 ;
  assign n378 = ~x5 & n376 ;
  assign n379 = ( ~x5 & n367 ) | ( ~x5 & n378 ) | ( n367 & n378 ) ;
  assign n380 = ( ~n374 & n377 ) | ( ~n374 & n379 ) | ( n377 & n379 ) ;
  assign n381 = ~x6 & x7 ;
  assign n382 = x6 & ~x7 ;
  assign n383 = n381 | n382 ;
  assign n384 = ~n318 & n383 ;
  assign n385 = x64 & n384 ;
  assign n386 = ~x7 & x8 ;
  assign n387 = x7 & ~x8 ;
  assign n388 = n386 | n387 ;
  assign n389 = n318 & ~n388 ;
  assign n390 = x65 & n389 ;
  assign n391 = n385 | n390 ;
  assign n392 = n318 & n388 ;
  assign n393 = x8 | n144 ;
  assign n394 = ( x8 & n392 ) | ( x8 & n393 ) | ( n392 & n393 ) ;
  assign n395 = ~x8 & n394 ;
  assign n396 = ( ~x8 & n391 ) | ( ~x8 & n395 ) | ( n391 & n395 ) ;
  assign n397 = x8 & ~x64 ;
  assign n398 = ( x8 & ~n318 ) | ( x8 & n397 ) | ( ~n318 & n397 ) ;
  assign n399 = n394 & n398 ;
  assign n400 = ( n391 & n398 ) | ( n391 & n399 ) | ( n398 & n399 ) ;
  assign n401 = n144 & n392 ;
  assign n402 = n398 & ~n401 ;
  assign n403 = ~n391 & n402 ;
  assign n404 = ( n396 & n400 ) | ( n396 & n403 ) | ( n400 & n403 ) ;
  assign n405 = n394 | n398 ;
  assign n406 = n391 | n405 ;
  assign n407 = ~n398 & n401 ;
  assign n408 = ( n391 & ~n398 ) | ( n391 & n407 ) | ( ~n398 & n407 ) ;
  assign n409 = ( n396 & n406 ) | ( n396 & ~n408 ) | ( n406 & ~n408 ) ;
  assign n410 = ~n404 & n409 ;
  assign n411 = n380 & n410 ;
  assign n412 = n380 & ~n411 ;
  assign n413 = ~n380 & n410 ;
  assign n414 = n412 | n413 ;
  assign n415 = n227 & n319 ;
  assign n416 = n279 & n415 ;
  assign n417 = n280 & ~n416 ;
  assign n418 = ~n227 & n319 ;
  assign n419 = ( ~n279 & n319 ) | ( ~n279 & n418 ) | ( n319 & n418 ) ;
  assign n420 = n330 & ~n419 ;
  assign n421 = ~n417 & n420 ;
  assign n422 = ( n330 & n416 ) | ( n330 & ~n421 ) | ( n416 & ~n421 ) ;
  assign n423 = n414 & n422 ;
  assign n424 = n414 | n422 ;
  assign n425 = ~n423 & n424 ;
  assign n426 = x70 | x71 ;
  assign n427 = x70 & x71 ;
  assign n428 = n426 & ~n427 ;
  assign n429 = n284 | n334 ;
  assign n430 = ( n334 & n335 ) | ( n334 & n429 ) | ( n335 & n429 ) ;
  assign n431 = n428 & n430 ;
  assign n432 = n334 | n335 ;
  assign n433 = n428 & n432 ;
  assign n434 = ( n289 & n431 ) | ( n289 & n433 ) | ( n431 & n433 ) ;
  assign n435 = n428 | n430 ;
  assign n436 = n428 | n432 ;
  assign n437 = ( n289 & n435 ) | ( n289 & n436 ) | ( n435 & n436 ) ;
  assign n438 = ~n434 & n437 ;
  assign n439 = x70 & n133 ;
  assign n440 = x69 & ~n162 ;
  assign n441 = ( n137 & n439 ) | ( n137 & n440 ) | ( n439 & n440 ) ;
  assign n442 = x0 & x71 ;
  assign n443 = ( ~n137 & n439 ) | ( ~n137 & n442 ) | ( n439 & n442 ) ;
  assign n444 = n441 | n443 ;
  assign n445 = ( n141 & n438 ) | ( n141 & n444 ) | ( n438 & n444 ) ;
  assign n446 = ( x2 & n141 ) | ( x2 & ~n444 ) | ( n141 & ~n444 ) ;
  assign n447 = ( x2 & n438 ) | ( x2 & n446 ) | ( n438 & n446 ) ;
  assign n448 = ~n445 & n447 ;
  assign n449 = n444 | n446 ;
  assign n450 = x2 | n444 ;
  assign n451 = ( n438 & n449 ) | ( n438 & n450 ) | ( n449 & n450 ) ;
  assign n452 = ( ~x2 & n448 ) | ( ~x2 & n451 ) | ( n448 & n451 ) ;
  assign n453 = n425 & n452 ;
  assign n454 = n425 | n452 ;
  assign n455 = ~n453 & n454 ;
  assign n456 = n357 | n361 ;
  assign n457 = ( n357 & n363 ) | ( n357 & n456 ) | ( n363 & n456 ) ;
  assign n458 = n455 & n457 ;
  assign n459 = n455 | n457 ;
  assign n460 = ~n458 & n459 ;
  assign n461 = x66 & n389 ;
  assign n462 = x65 & n384 ;
  assign n463 = ~n318 & n388 ;
  assign n464 = x64 & ~n383 ;
  assign n465 = n463 & n464 ;
  assign n466 = n462 | n465 ;
  assign n467 = n461 | n466 ;
  assign n468 = n159 & n392 ;
  assign n469 = n467 | n468 ;
  assign n470 = x8 | n392 ;
  assign n471 = ( x8 & n159 ) | ( x8 & n470 ) | ( n159 & n470 ) ;
  assign n472 = n467 | n471 ;
  assign n473 = ~x8 & n471 ;
  assign n474 = ( ~x8 & n467 ) | ( ~x8 & n473 ) | ( n467 & n473 ) ;
  assign n475 = ( ~n469 & n472 ) | ( ~n469 & n474 ) | ( n472 & n474 ) ;
  assign n476 = n404 | n475 ;
  assign n477 = n404 & n475 ;
  assign n478 = n476 & ~n477 ;
  assign n479 = n215 & n293 ;
  assign n480 = x69 & n212 ;
  assign n481 = x68 & n207 ;
  assign n482 = x67 & ~n206 ;
  assign n483 = n267 & n482 ;
  assign n484 = n481 | n483 ;
  assign n485 = n480 | n484 ;
  assign n486 = n479 | n485 ;
  assign n487 = x5 | n480 ;
  assign n488 = n484 | n487 ;
  assign n489 = n479 | n488 ;
  assign n490 = ~x5 & n488 ;
  assign n491 = ( ~x5 & n479 ) | ( ~x5 & n490 ) | ( n479 & n490 ) ;
  assign n492 = ( ~n486 & n489 ) | ( ~n486 & n491 ) | ( n489 & n491 ) ;
  assign n493 = n478 & n492 ;
  assign n494 = n478 & ~n493 ;
  assign n495 = ~n478 & n492 ;
  assign n496 = n494 | n495 ;
  assign n497 = n411 | n414 ;
  assign n498 = ( n411 & n422 ) | ( n411 & n497 ) | ( n422 & n497 ) ;
  assign n499 = n496 | n498 ;
  assign n500 = n496 & n498 ;
  assign n501 = n499 & ~n500 ;
  assign n502 = x71 | x72 ;
  assign n503 = x71 & x72 ;
  assign n504 = n502 & ~n503 ;
  assign n505 = n427 & n504 ;
  assign n506 = ( n433 & n504 ) | ( n433 & n505 ) | ( n504 & n505 ) ;
  assign n507 = ( n431 & n504 ) | ( n431 & n505 ) | ( n504 & n505 ) ;
  assign n508 = ( n289 & n506 ) | ( n289 & n507 ) | ( n506 & n507 ) ;
  assign n509 = n427 | n504 ;
  assign n510 = n433 | n509 ;
  assign n511 = n431 | n509 ;
  assign n512 = ( n289 & n510 ) | ( n289 & n511 ) | ( n510 & n511 ) ;
  assign n513 = ~n508 & n512 ;
  assign n514 = x71 & n133 ;
  assign n515 = x70 & ~n162 ;
  assign n516 = ( n137 & n514 ) | ( n137 & n515 ) | ( n514 & n515 ) ;
  assign n517 = x0 & x72 ;
  assign n518 = ( ~n137 & n514 ) | ( ~n137 & n517 ) | ( n514 & n517 ) ;
  assign n519 = n516 | n518 ;
  assign n520 = n141 | n519 ;
  assign n521 = ( n513 & n519 ) | ( n513 & n520 ) | ( n519 & n520 ) ;
  assign n522 = x2 & n519 ;
  assign n523 = x2 & n141 ;
  assign n524 = ( x2 & n519 ) | ( x2 & n523 ) | ( n519 & n523 ) ;
  assign n525 = ( n513 & n522 ) | ( n513 & n524 ) | ( n522 & n524 ) ;
  assign n526 = x2 & ~n524 ;
  assign n527 = x2 & ~n519 ;
  assign n528 = ( ~n513 & n526 ) | ( ~n513 & n527 ) | ( n526 & n527 ) ;
  assign n529 = ( n521 & ~n525 ) | ( n521 & n528 ) | ( ~n525 & n528 ) ;
  assign n530 = n501 & n529 ;
  assign n531 = n501 & ~n530 ;
  assign n532 = ~n501 & n529 ;
  assign n533 = n531 | n532 ;
  assign n534 = n453 | n457 ;
  assign n535 = ( n453 & n455 ) | ( n453 & n534 ) | ( n455 & n534 ) ;
  assign n536 = n533 | n535 ;
  assign n537 = n532 & n535 ;
  assign n538 = ( n531 & n535 ) | ( n531 & n537 ) | ( n535 & n537 ) ;
  assign n539 = n536 & ~n538 ;
  assign n540 = x8 & ~x9 ;
  assign n541 = ~x8 & x9 ;
  assign n542 = n540 | n541 ;
  assign n543 = x64 & n542 ;
  assign n544 = ~n404 & n543 ;
  assign n545 = ( ~n475 & n543 ) | ( ~n475 & n544 ) | ( n543 & n544 ) ;
  assign n546 = n404 & ~n543 ;
  assign n547 = n475 & n546 ;
  assign n548 = n545 | n547 ;
  assign n549 = x67 & n389 ;
  assign n550 = x66 & n384 ;
  assign n551 = x65 & ~n383 ;
  assign n552 = n463 & n551 ;
  assign n553 = n550 | n552 ;
  assign n554 = n549 | n553 ;
  assign n555 = n186 & n392 ;
  assign n556 = n554 | n555 ;
  assign n557 = x8 & ~n556 ;
  assign n558 = ~x8 & n556 ;
  assign n559 = n557 | n558 ;
  assign n560 = n548 & n559 ;
  assign n561 = n548 | n559 ;
  assign n562 = ~n560 & n561 ;
  assign n563 = x69 & n207 ;
  assign n564 = x68 & ~n206 ;
  assign n565 = n267 & n564 ;
  assign n566 = n563 | n565 ;
  assign n567 = x70 & n212 ;
  assign n568 = n215 | n567 ;
  assign n569 = n566 | n568 ;
  assign n570 = x5 & ~n569 ;
  assign n571 = x5 & ~n567 ;
  assign n572 = ~n566 & n571 ;
  assign n573 = ( ~n340 & n570 ) | ( ~n340 & n572 ) | ( n570 & n572 ) ;
  assign n574 = ~x5 & n569 ;
  assign n575 = ~x5 & n567 ;
  assign n576 = ( ~x5 & n566 ) | ( ~x5 & n575 ) | ( n566 & n575 ) ;
  assign n577 = ( n340 & n574 ) | ( n340 & n576 ) | ( n574 & n576 ) ;
  assign n578 = n573 | n577 ;
  assign n579 = n562 & n578 ;
  assign n580 = n562 & ~n579 ;
  assign n581 = ~n562 & n578 ;
  assign n582 = n580 | n581 ;
  assign n583 = n493 | n495 ;
  assign n584 = n494 | n583 ;
  assign n585 = ( n493 & n498 ) | ( n493 & n584 ) | ( n498 & n584 ) ;
  assign n586 = n582 | n585 ;
  assign n587 = n582 & n585 ;
  assign n588 = n586 & ~n587 ;
  assign n589 = x72 | x73 ;
  assign n590 = x72 & x73 ;
  assign n591 = n589 & ~n590 ;
  assign n592 = n503 | n504 ;
  assign n593 = n427 | n503 ;
  assign n594 = ( n503 & n504 ) | ( n503 & n593 ) | ( n504 & n593 ) ;
  assign n595 = ( n433 & n592 ) | ( n433 & n594 ) | ( n592 & n594 ) ;
  assign n596 = ( n431 & n592 ) | ( n431 & n594 ) | ( n592 & n594 ) ;
  assign n597 = ( n289 & n595 ) | ( n289 & n596 ) | ( n595 & n596 ) ;
  assign n598 = n591 | n597 ;
  assign n599 = x72 & n133 ;
  assign n600 = x71 & ~n162 ;
  assign n601 = ( n137 & n599 ) | ( n137 & n600 ) | ( n599 & n600 ) ;
  assign n602 = x0 & x73 ;
  assign n603 = ( ~n137 & n599 ) | ( ~n137 & n602 ) | ( n599 & n602 ) ;
  assign n604 = n601 | n603 ;
  assign n605 = n141 | n604 ;
  assign n606 = n591 & n594 ;
  assign n607 = n591 & n592 ;
  assign n608 = ( n433 & n606 ) | ( n433 & n607 ) | ( n606 & n607 ) ;
  assign n609 = ( n431 & n606 ) | ( n431 & n607 ) | ( n606 & n607 ) ;
  assign n610 = ( n289 & n608 ) | ( n289 & n609 ) | ( n608 & n609 ) ;
  assign n611 = ( n604 & n605 ) | ( n604 & ~n610 ) | ( n605 & ~n610 ) ;
  assign n612 = n604 & n605 ;
  assign n613 = ( n598 & n611 ) | ( n598 & n612 ) | ( n611 & n612 ) ;
  assign n614 = x2 & n613 ;
  assign n615 = x2 & ~n613 ;
  assign n616 = ( n613 & ~n614 ) | ( n613 & n615 ) | ( ~n614 & n615 ) ;
  assign n617 = n588 & n616 ;
  assign n618 = n588 & ~n617 ;
  assign n619 = ~n588 & n616 ;
  assign n620 = n618 | n619 ;
  assign n621 = n530 | n535 ;
  assign n622 = n530 | n531 ;
  assign n623 = ( n537 & n621 ) | ( n537 & n622 ) | ( n621 & n622 ) ;
  assign n624 = n620 & n623 ;
  assign n625 = n620 | n623 ;
  assign n626 = ~n624 & n625 ;
  assign n627 = n617 | n624 ;
  assign n628 = ~x9 & x10 ;
  assign n629 = x9 & ~x10 ;
  assign n630 = n628 | n629 ;
  assign n631 = ~n542 & n630 ;
  assign n632 = x64 & n631 ;
  assign n633 = ~x10 & x11 ;
  assign n634 = x10 & ~x11 ;
  assign n635 = n633 | n634 ;
  assign n636 = n542 & ~n635 ;
  assign n637 = x65 & n636 ;
  assign n638 = n632 | n637 ;
  assign n639 = n542 & n635 ;
  assign n640 = x11 | n144 ;
  assign n641 = ( x11 & n639 ) | ( x11 & n640 ) | ( n639 & n640 ) ;
  assign n642 = ~x11 & n641 ;
  assign n643 = ( ~x11 & n638 ) | ( ~x11 & n642 ) | ( n638 & n642 ) ;
  assign n644 = x11 & ~x64 ;
  assign n645 = ( x11 & ~n542 ) | ( x11 & n644 ) | ( ~n542 & n644 ) ;
  assign n646 = n641 & n645 ;
  assign n647 = ( n638 & n645 ) | ( n638 & n646 ) | ( n645 & n646 ) ;
  assign n648 = n144 & n639 ;
  assign n649 = n645 & ~n648 ;
  assign n650 = ~n638 & n649 ;
  assign n651 = ( n643 & n647 ) | ( n643 & n650 ) | ( n647 & n650 ) ;
  assign n652 = n641 | n645 ;
  assign n653 = n638 | n652 ;
  assign n654 = ~n645 & n648 ;
  assign n655 = ( n638 & ~n645 ) | ( n638 & n654 ) | ( ~n645 & n654 ) ;
  assign n656 = ( n643 & n653 ) | ( n643 & ~n655 ) | ( n653 & ~n655 ) ;
  assign n657 = ~n651 & n656 ;
  assign n658 = n241 & n392 ;
  assign n659 = x68 & n389 ;
  assign n660 = x67 & n384 ;
  assign n661 = x66 & ~n383 ;
  assign n662 = n463 & n661 ;
  assign n663 = n660 | n662 ;
  assign n664 = n659 | n663 ;
  assign n665 = n658 | n664 ;
  assign n666 = x8 | n659 ;
  assign n667 = n663 | n666 ;
  assign n668 = n658 | n667 ;
  assign n669 = ~x8 & n667 ;
  assign n670 = ( ~x8 & n658 ) | ( ~x8 & n669 ) | ( n658 & n669 ) ;
  assign n671 = ( ~n665 & n668 ) | ( ~n665 & n670 ) | ( n668 & n670 ) ;
  assign n672 = n657 | n671 ;
  assign n673 = n657 & n671 ;
  assign n674 = n672 & ~n673 ;
  assign n675 = ( n477 & n543 ) | ( n477 & n559 ) | ( n543 & n559 ) ;
  assign n676 = n674 | n675 ;
  assign n677 = n674 & n675 ;
  assign n678 = n676 & ~n677 ;
  assign n679 = x70 & n207 ;
  assign n680 = x69 & ~n206 ;
  assign n681 = n267 & n680 ;
  assign n682 = n679 | n681 ;
  assign n683 = x71 & n212 ;
  assign n684 = n215 | n683 ;
  assign n685 = n682 | n684 ;
  assign n686 = x5 & ~n685 ;
  assign n687 = x5 & ~n683 ;
  assign n688 = ~n682 & n687 ;
  assign n689 = ( ~n438 & n686 ) | ( ~n438 & n688 ) | ( n686 & n688 ) ;
  assign n690 = ~x5 & n685 ;
  assign n691 = ~x5 & n683 ;
  assign n692 = ( ~x5 & n682 ) | ( ~x5 & n691 ) | ( n682 & n691 ) ;
  assign n693 = ( n438 & n690 ) | ( n438 & n692 ) | ( n690 & n692 ) ;
  assign n694 = n689 | n693 ;
  assign n695 = n678 & n694 ;
  assign n696 = n678 & ~n695 ;
  assign n697 = ~n678 & n694 ;
  assign n698 = n696 | n697 ;
  assign n699 = n579 | n587 ;
  assign n700 = n698 | n699 ;
  assign n701 = n698 & n699 ;
  assign n702 = n700 & ~n701 ;
  assign n703 = x73 | x74 ;
  assign n704 = x73 & x74 ;
  assign n705 = n703 & ~n704 ;
  assign n706 = n590 & n705 ;
  assign n707 = ( n610 & n705 ) | ( n610 & n706 ) | ( n705 & n706 ) ;
  assign n708 = n590 | n705 ;
  assign n709 = n610 | n708 ;
  assign n710 = ~n707 & n709 ;
  assign n711 = x73 & n133 ;
  assign n712 = x72 & ~n162 ;
  assign n713 = ( n137 & n711 ) | ( n137 & n712 ) | ( n711 & n712 ) ;
  assign n714 = x0 & x74 ;
  assign n715 = ( ~n137 & n711 ) | ( ~n137 & n714 ) | ( n711 & n714 ) ;
  assign n716 = n713 | n715 ;
  assign n717 = n141 | n716 ;
  assign n718 = ( n710 & n716 ) | ( n710 & n717 ) | ( n716 & n717 ) ;
  assign n719 = x2 & n716 ;
  assign n720 = ( x2 & n523 ) | ( x2 & n716 ) | ( n523 & n716 ) ;
  assign n721 = ( n710 & n719 ) | ( n710 & n720 ) | ( n719 & n720 ) ;
  assign n722 = x2 & ~n720 ;
  assign n723 = x2 & ~n716 ;
  assign n724 = ( ~n710 & n722 ) | ( ~n710 & n723 ) | ( n722 & n723 ) ;
  assign n725 = ( n718 & ~n721 ) | ( n718 & n724 ) | ( ~n721 & n724 ) ;
  assign n726 = n702 | n725 ;
  assign n727 = n702 & n725 ;
  assign n728 = n726 & ~n727 ;
  assign n729 = n627 | n728 ;
  assign n730 = n627 & n728 ;
  assign n731 = n729 & ~n730 ;
  assign n732 = x74 | x75 ;
  assign n733 = x74 & x75 ;
  assign n734 = n732 & ~n733 ;
  assign n735 = n704 | n705 ;
  assign n736 = n734 & n735 ;
  assign n737 = n704 & n734 ;
  assign n738 = ( n590 & n736 ) | ( n590 & n737 ) | ( n736 & n737 ) ;
  assign n739 = n736 | n737 ;
  assign n740 = ( n610 & n738 ) | ( n610 & n739 ) | ( n738 & n739 ) ;
  assign n741 = n734 | n735 ;
  assign n742 = n590 | n704 ;
  assign n743 = ( n704 & n705 ) | ( n704 & n742 ) | ( n705 & n742 ) ;
  assign n744 = n734 | n743 ;
  assign n745 = ( n610 & n741 ) | ( n610 & n744 ) | ( n741 & n744 ) ;
  assign n746 = ~n740 & n745 ;
  assign n747 = x74 & n133 ;
  assign n748 = x73 & ~n162 ;
  assign n749 = ( n137 & n747 ) | ( n137 & n748 ) | ( n747 & n748 ) ;
  assign n750 = x0 & x75 ;
  assign n751 = ( ~n137 & n747 ) | ( ~n137 & n750 ) | ( n747 & n750 ) ;
  assign n752 = n749 | n751 ;
  assign n753 = n141 | n752 ;
  assign n754 = ( n746 & n752 ) | ( n746 & n753 ) | ( n752 & n753 ) ;
  assign n755 = x2 & n752 ;
  assign n756 = ( x2 & n523 ) | ( x2 & n752 ) | ( n523 & n752 ) ;
  assign n757 = ( n746 & n755 ) | ( n746 & n756 ) | ( n755 & n756 ) ;
  assign n758 = x2 & ~n756 ;
  assign n759 = x2 & ~n752 ;
  assign n760 = ( ~n746 & n758 ) | ( ~n746 & n759 ) | ( n758 & n759 ) ;
  assign n761 = ( n754 & ~n757 ) | ( n754 & n760 ) | ( ~n757 & n760 ) ;
  assign n762 = x66 & n636 ;
  assign n763 = x65 & n631 ;
  assign n764 = ~n542 & n635 ;
  assign n765 = x64 & ~n630 ;
  assign n766 = n764 & n765 ;
  assign n767 = n763 | n766 ;
  assign n768 = n762 | n767 ;
  assign n769 = n159 & n639 ;
  assign n770 = n768 | n769 ;
  assign n771 = x11 | n639 ;
  assign n772 = ( x11 & n159 ) | ( x11 & n771 ) | ( n159 & n771 ) ;
  assign n773 = n768 | n772 ;
  assign n774 = ~x11 & n772 ;
  assign n775 = ( ~x11 & n768 ) | ( ~x11 & n774 ) | ( n768 & n774 ) ;
  assign n776 = ( ~n770 & n773 ) | ( ~n770 & n775 ) | ( n773 & n775 ) ;
  assign n777 = n651 | n776 ;
  assign n778 = n651 & n776 ;
  assign n779 = n777 & ~n778 ;
  assign n780 = n293 & n392 ;
  assign n781 = x69 & n389 ;
  assign n782 = x68 & n384 ;
  assign n783 = x67 & ~n383 ;
  assign n784 = n463 & n783 ;
  assign n785 = n782 | n784 ;
  assign n786 = n781 | n785 ;
  assign n787 = n780 | n786 ;
  assign n788 = x8 | n781 ;
  assign n789 = n785 | n788 ;
  assign n790 = n780 | n789 ;
  assign n791 = ~x8 & n789 ;
  assign n792 = ( ~x8 & n780 ) | ( ~x8 & n791 ) | ( n780 & n791 ) ;
  assign n793 = ( ~n787 & n790 ) | ( ~n787 & n792 ) | ( n790 & n792 ) ;
  assign n794 = n779 & n793 ;
  assign n795 = n779 & ~n794 ;
  assign n796 = ~n779 & n793 ;
  assign n797 = n795 | n796 ;
  assign n798 = n673 | n675 ;
  assign n799 = ( n673 & n674 ) | ( n673 & n798 ) | ( n674 & n798 ) ;
  assign n800 = n797 & n799 ;
  assign n801 = n797 | n799 ;
  assign n802 = ~n800 & n801 ;
  assign n803 = x71 & n207 ;
  assign n804 = x70 & ~n206 ;
  assign n805 = n267 & n804 ;
  assign n806 = n803 | n805 ;
  assign n807 = x72 & n212 ;
  assign n808 = n215 | n807 ;
  assign n809 = n806 | n808 ;
  assign n810 = x5 & n809 ;
  assign n811 = x5 & n807 ;
  assign n812 = ( x5 & n806 ) | ( x5 & n811 ) | ( n806 & n811 ) ;
  assign n813 = ( n513 & n810 ) | ( n513 & n812 ) | ( n810 & n812 ) ;
  assign n814 = x5 | n809 ;
  assign n815 = x5 | n807 ;
  assign n816 = n806 | n815 ;
  assign n817 = ( n513 & n814 ) | ( n513 & n816 ) | ( n814 & n816 ) ;
  assign n818 = ~n813 & n817 ;
  assign n819 = n802 & n818 ;
  assign n820 = n802 & ~n819 ;
  assign n821 = ~n802 & n818 ;
  assign n822 = n820 | n821 ;
  assign n823 = n695 | n697 ;
  assign n824 = n696 | n823 ;
  assign n825 = ( n695 & n699 ) | ( n695 & n824 ) | ( n699 & n824 ) ;
  assign n826 = ( n761 & ~n822 ) | ( n761 & n825 ) | ( ~n822 & n825 ) ;
  assign n827 = ( n822 & ~n825 ) | ( n822 & n826 ) | ( ~n825 & n826 ) ;
  assign n828 = ( ~n761 & n826 ) | ( ~n761 & n827 ) | ( n826 & n827 ) ;
  assign n829 = n727 | n728 ;
  assign n830 = ( n627 & n727 ) | ( n627 & n829 ) | ( n727 & n829 ) ;
  assign n831 = n828 & n830 ;
  assign n832 = n828 | n830 ;
  assign n833 = ~n831 & n832 ;
  assign n834 = x11 & ~x12 ;
  assign n835 = ~x11 & x12 ;
  assign n836 = n834 | n835 ;
  assign n837 = x64 & n836 ;
  assign n838 = ~n651 & n837 ;
  assign n839 = ( ~n776 & n837 ) | ( ~n776 & n838 ) | ( n837 & n838 ) ;
  assign n840 = n651 & ~n837 ;
  assign n841 = n776 & n840 ;
  assign n842 = n839 | n841 ;
  assign n843 = x67 & n636 ;
  assign n844 = x66 & n631 ;
  assign n845 = x65 & ~n630 ;
  assign n846 = n764 & n845 ;
  assign n847 = n844 | n846 ;
  assign n848 = n843 | n847 ;
  assign n849 = n186 & n639 ;
  assign n850 = n848 | n849 ;
  assign n851 = x11 & ~n850 ;
  assign n852 = ~x11 & n850 ;
  assign n853 = n851 | n852 ;
  assign n854 = n842 & n853 ;
  assign n855 = n842 | n853 ;
  assign n856 = ~n854 & n855 ;
  assign n857 = x69 & n384 ;
  assign n858 = x68 & ~n383 ;
  assign n859 = n463 & n858 ;
  assign n860 = n857 | n859 ;
  assign n861 = x70 & n389 ;
  assign n862 = n392 | n861 ;
  assign n863 = n860 | n862 ;
  assign n864 = x8 & ~n863 ;
  assign n865 = x8 & ~n861 ;
  assign n866 = ~n860 & n865 ;
  assign n867 = ( ~n340 & n864 ) | ( ~n340 & n866 ) | ( n864 & n866 ) ;
  assign n868 = ~x8 & n863 ;
  assign n869 = ~x8 & n861 ;
  assign n870 = ( ~x8 & n860 ) | ( ~x8 & n869 ) | ( n860 & n869 ) ;
  assign n871 = ( n340 & n868 ) | ( n340 & n870 ) | ( n868 & n870 ) ;
  assign n872 = n867 | n871 ;
  assign n873 = n856 & n872 ;
  assign n874 = n856 & ~n873 ;
  assign n875 = ~n856 & n872 ;
  assign n876 = n874 | n875 ;
  assign n877 = n794 | n799 ;
  assign n878 = ( n794 & n797 ) | ( n794 & n877 ) | ( n797 & n877 ) ;
  assign n879 = n876 | n878 ;
  assign n880 = n876 & n878 ;
  assign n881 = n879 & ~n880 ;
  assign n882 = x73 & n212 ;
  assign n883 = x72 & n207 ;
  assign n884 = x71 & ~n206 ;
  assign n885 = n267 & n884 ;
  assign n886 = n883 | n885 ;
  assign n887 = n882 | n886 ;
  assign n888 = ( n215 & ~n610 ) | ( n215 & n887 ) | ( ~n610 & n887 ) ;
  assign n889 = n215 & n882 ;
  assign n890 = ( n215 & n886 ) | ( n215 & n889 ) | ( n886 & n889 ) ;
  assign n891 = ( n598 & n888 ) | ( n598 & n890 ) | ( n888 & n890 ) ;
  assign n892 = ( x5 & ~n887 ) | ( x5 & n891 ) | ( ~n887 & n891 ) ;
  assign n893 = ~n891 & n892 ;
  assign n894 = x5 | n882 ;
  assign n895 = n886 | n894 ;
  assign n896 = n891 | n895 ;
  assign n897 = ( ~x5 & n893 ) | ( ~x5 & n896 ) | ( n893 & n896 ) ;
  assign n898 = n881 | n897 ;
  assign n899 = n881 & n897 ;
  assign n900 = n898 & ~n899 ;
  assign n901 = n822 & n825 ;
  assign n902 = n819 | n901 ;
  assign n903 = n900 & n902 ;
  assign n904 = n900 | n902 ;
  assign n905 = ~n903 & n904 ;
  assign n906 = x75 | x76 ;
  assign n907 = x75 & x76 ;
  assign n908 = n906 & ~n907 ;
  assign n909 = n733 | n734 ;
  assign n910 = ( n733 & n735 ) | ( n733 & n909 ) | ( n735 & n909 ) ;
  assign n911 = n908 & n910 ;
  assign n912 = n704 | n733 ;
  assign n913 = ( n733 & n734 ) | ( n733 & n912 ) | ( n734 & n912 ) ;
  assign n914 = n908 & n913 ;
  assign n915 = ( n590 & n911 ) | ( n590 & n914 ) | ( n911 & n914 ) ;
  assign n916 = n911 | n914 ;
  assign n917 = ( n610 & n915 ) | ( n610 & n916 ) | ( n915 & n916 ) ;
  assign n918 = n908 | n913 ;
  assign n919 = n910 | n918 ;
  assign n920 = n590 | n908 ;
  assign n921 = ( n910 & n918 ) | ( n910 & n920 ) | ( n918 & n920 ) ;
  assign n922 = ( n610 & n919 ) | ( n610 & n921 ) | ( n919 & n921 ) ;
  assign n923 = ~n917 & n922 ;
  assign n924 = x75 & n133 ;
  assign n925 = x74 & ~n162 ;
  assign n926 = ( n137 & n924 ) | ( n137 & n925 ) | ( n924 & n925 ) ;
  assign n927 = x0 & x76 ;
  assign n928 = ( ~n137 & n924 ) | ( ~n137 & n927 ) | ( n924 & n927 ) ;
  assign n929 = n926 | n928 ;
  assign n930 = n141 | n929 ;
  assign n931 = ( n923 & n929 ) | ( n923 & n930 ) | ( n929 & n930 ) ;
  assign n932 = x2 & n929 ;
  assign n933 = ( x2 & n523 ) | ( x2 & n929 ) | ( n523 & n929 ) ;
  assign n934 = ( n923 & n932 ) | ( n923 & n933 ) | ( n932 & n933 ) ;
  assign n935 = x2 & ~n933 ;
  assign n936 = x2 & ~n929 ;
  assign n937 = ( ~n923 & n935 ) | ( ~n923 & n936 ) | ( n935 & n936 ) ;
  assign n938 = ( n931 & ~n934 ) | ( n931 & n937 ) | ( ~n934 & n937 ) ;
  assign n939 = n905 & n938 ;
  assign n940 = n905 & ~n939 ;
  assign n941 = ~n905 & n938 ;
  assign n942 = n940 | n941 ;
  assign n943 = n825 & ~n901 ;
  assign n944 = n822 & ~n825 ;
  assign n945 = n761 & n944 ;
  assign n946 = ( n761 & n943 ) | ( n761 & n945 ) | ( n943 & n945 ) ;
  assign n947 = n828 | n946 ;
  assign n948 = ( n830 & n946 ) | ( n830 & n947 ) | ( n946 & n947 ) ;
  assign n949 = n942 & n948 ;
  assign n950 = n942 | n948 ;
  assign n951 = ~n949 & n950 ;
  assign n952 = n899 | n900 ;
  assign n953 = ( n899 & n902 ) | ( n899 & n952 ) | ( n902 & n952 ) ;
  assign n954 = ~x12 & x13 ;
  assign n955 = x12 & ~x13 ;
  assign n956 = n954 | n955 ;
  assign n957 = ~n836 & n956 ;
  assign n958 = x64 & n957 ;
  assign n959 = ~x13 & x14 ;
  assign n960 = x13 & ~x14 ;
  assign n961 = n959 | n960 ;
  assign n962 = n836 & ~n961 ;
  assign n963 = x65 & n962 ;
  assign n964 = n958 | n963 ;
  assign n965 = n836 & n961 ;
  assign n966 = x14 | n144 ;
  assign n967 = ( x14 & n965 ) | ( x14 & n966 ) | ( n965 & n966 ) ;
  assign n968 = ~x14 & n967 ;
  assign n969 = ( ~x14 & n964 ) | ( ~x14 & n968 ) | ( n964 & n968 ) ;
  assign n970 = x14 & ~x64 ;
  assign n971 = ( x14 & ~n836 ) | ( x14 & n970 ) | ( ~n836 & n970 ) ;
  assign n972 = n967 & n971 ;
  assign n973 = ( n964 & n971 ) | ( n964 & n972 ) | ( n971 & n972 ) ;
  assign n974 = n144 & n965 ;
  assign n975 = n971 & ~n974 ;
  assign n976 = ~n964 & n975 ;
  assign n977 = ( n969 & n973 ) | ( n969 & n976 ) | ( n973 & n976 ) ;
  assign n978 = n967 | n971 ;
  assign n979 = n964 | n978 ;
  assign n980 = ~n971 & n974 ;
  assign n981 = ( n964 & ~n971 ) | ( n964 & n980 ) | ( ~n971 & n980 ) ;
  assign n982 = ( n969 & n979 ) | ( n969 & ~n981 ) | ( n979 & ~n981 ) ;
  assign n983 = ~n977 & n982 ;
  assign n984 = n241 & n639 ;
  assign n985 = x68 & n636 ;
  assign n986 = x67 & n631 ;
  assign n987 = x66 & ~n630 ;
  assign n988 = n764 & n987 ;
  assign n989 = n986 | n988 ;
  assign n990 = n985 | n989 ;
  assign n991 = n984 | n990 ;
  assign n992 = x11 | n985 ;
  assign n993 = n989 | n992 ;
  assign n994 = n984 | n993 ;
  assign n995 = ~x11 & n993 ;
  assign n996 = ( ~x11 & n984 ) | ( ~x11 & n995 ) | ( n984 & n995 ) ;
  assign n997 = ( ~n991 & n994 ) | ( ~n991 & n996 ) | ( n994 & n996 ) ;
  assign n998 = n983 | n997 ;
  assign n999 = n983 & n997 ;
  assign n1000 = n998 & ~n999 ;
  assign n1001 = ( n778 & n837 ) | ( n778 & n853 ) | ( n837 & n853 ) ;
  assign n1002 = n1000 | n1001 ;
  assign n1003 = n1000 & n1001 ;
  assign n1004 = n1002 & ~n1003 ;
  assign n1005 = x70 & n384 ;
  assign n1006 = x69 & ~n383 ;
  assign n1007 = n463 & n1006 ;
  assign n1008 = n1005 | n1007 ;
  assign n1009 = x71 & n389 ;
  assign n1010 = n392 | n1009 ;
  assign n1011 = n1008 | n1010 ;
  assign n1012 = x8 & ~n1011 ;
  assign n1013 = x8 & ~n1009 ;
  assign n1014 = ~n1008 & n1013 ;
  assign n1015 = ( ~n438 & n1012 ) | ( ~n438 & n1014 ) | ( n1012 & n1014 ) ;
  assign n1016 = ~x8 & n1011 ;
  assign n1017 = ~x8 & n1009 ;
  assign n1018 = ( ~x8 & n1008 ) | ( ~x8 & n1017 ) | ( n1008 & n1017 ) ;
  assign n1019 = ( n438 & n1016 ) | ( n438 & n1018 ) | ( n1016 & n1018 ) ;
  assign n1020 = n1015 | n1019 ;
  assign n1021 = n1004 & n1020 ;
  assign n1022 = n1004 & ~n1021 ;
  assign n1023 = ~n1004 & n1020 ;
  assign n1024 = n1022 | n1023 ;
  assign n1025 = n873 | n878 ;
  assign n1026 = ( n873 & n876 ) | ( n873 & n1025 ) | ( n876 & n1025 ) ;
  assign n1027 = n1024 | n1026 ;
  assign n1028 = n1024 & n1026 ;
  assign n1029 = n1027 & ~n1028 ;
  assign n1030 = x74 & n212 ;
  assign n1031 = x73 & n207 ;
  assign n1032 = x72 & ~n206 ;
  assign n1033 = n267 & n1032 ;
  assign n1034 = n1031 | n1033 ;
  assign n1035 = n1030 | n1034 ;
  assign n1036 = n215 | n1030 ;
  assign n1037 = n1034 | n1036 ;
  assign n1038 = ( n710 & n1035 ) | ( n710 & n1037 ) | ( n1035 & n1037 ) ;
  assign n1039 = x5 & n1037 ;
  assign n1040 = x5 & n1030 ;
  assign n1041 = ( x5 & n1034 ) | ( x5 & n1040 ) | ( n1034 & n1040 ) ;
  assign n1042 = ( n710 & n1039 ) | ( n710 & n1041 ) | ( n1039 & n1041 ) ;
  assign n1043 = x5 & ~n1041 ;
  assign n1044 = x5 & ~n1037 ;
  assign n1045 = ( ~n710 & n1043 ) | ( ~n710 & n1044 ) | ( n1043 & n1044 ) ;
  assign n1046 = ( n1038 & ~n1042 ) | ( n1038 & n1045 ) | ( ~n1042 & n1045 ) ;
  assign n1047 = n1029 & n1046 ;
  assign n1048 = n1029 | n1046 ;
  assign n1049 = ~n1047 & n1048 ;
  assign n1050 = n953 & n1049 ;
  assign n1051 = n953 & ~n1050 ;
  assign n1052 = x76 | x77 ;
  assign n1053 = x76 & x77 ;
  assign n1054 = n1052 & ~n1053 ;
  assign n1055 = n907 & n1054 ;
  assign n1056 = ( n917 & n1054 ) | ( n917 & n1055 ) | ( n1054 & n1055 ) ;
  assign n1057 = n907 | n1054 ;
  assign n1058 = n917 | n1057 ;
  assign n1059 = ~n1056 & n1058 ;
  assign n1060 = x76 & n133 ;
  assign n1061 = x75 & ~n162 ;
  assign n1062 = ( n137 & n1060 ) | ( n137 & n1061 ) | ( n1060 & n1061 ) ;
  assign n1063 = x0 & x77 ;
  assign n1064 = ( ~n137 & n1060 ) | ( ~n137 & n1063 ) | ( n1060 & n1063 ) ;
  assign n1065 = n1062 | n1064 ;
  assign n1066 = n141 | n1065 ;
  assign n1067 = ( n1059 & n1065 ) | ( n1059 & n1066 ) | ( n1065 & n1066 ) ;
  assign n1068 = x2 & n1065 ;
  assign n1069 = ( x2 & n523 ) | ( x2 & n1065 ) | ( n523 & n1065 ) ;
  assign n1070 = ( n1059 & n1068 ) | ( n1059 & n1069 ) | ( n1068 & n1069 ) ;
  assign n1071 = x2 & ~n1069 ;
  assign n1072 = x2 & ~n1065 ;
  assign n1073 = ( ~n1059 & n1071 ) | ( ~n1059 & n1072 ) | ( n1071 & n1072 ) ;
  assign n1074 = ( n1067 & ~n1070 ) | ( n1067 & n1073 ) | ( ~n1070 & n1073 ) ;
  assign n1075 = ~n1048 & n1049 ;
  assign n1076 = ( ~n953 & n1049 ) | ( ~n953 & n1075 ) | ( n1049 & n1075 ) ;
  assign n1077 = ~n1074 & n1076 ;
  assign n1078 = ( n1051 & ~n1074 ) | ( n1051 & n1077 ) | ( ~n1074 & n1077 ) ;
  assign n1079 = n1074 & ~n1076 ;
  assign n1080 = ~n1051 & n1079 ;
  assign n1081 = n1078 | n1080 ;
  assign n1082 = n939 | n948 ;
  assign n1083 = ( n939 & n942 ) | ( n939 & n1082 ) | ( n942 & n1082 ) ;
  assign n1084 = n1081 & n1083 ;
  assign n1085 = n1081 | n1083 ;
  assign n1086 = ~n1084 & n1085 ;
  assign n1087 = x71 & n384 ;
  assign n1088 = x70 & ~n383 ;
  assign n1089 = n463 & n1088 ;
  assign n1090 = n1087 | n1089 ;
  assign n1091 = x72 & n389 ;
  assign n1092 = n392 | n1091 ;
  assign n1093 = n1090 | n1092 ;
  assign n1094 = x8 & n1093 ;
  assign n1095 = x8 & n1091 ;
  assign n1096 = ( x8 & n1090 ) | ( x8 & n1095 ) | ( n1090 & n1095 ) ;
  assign n1097 = ( n513 & n1094 ) | ( n513 & n1096 ) | ( n1094 & n1096 ) ;
  assign n1098 = x8 | n1093 ;
  assign n1099 = x8 | n1091 ;
  assign n1100 = n1090 | n1099 ;
  assign n1101 = ( n513 & n1098 ) | ( n513 & n1100 ) | ( n1098 & n1100 ) ;
  assign n1102 = ~n1097 & n1101 ;
  assign n1103 = x66 & n962 ;
  assign n1104 = x65 & n957 ;
  assign n1105 = ~n836 & n961 ;
  assign n1106 = x64 & ~n956 ;
  assign n1107 = n1105 & n1106 ;
  assign n1108 = n1104 | n1107 ;
  assign n1109 = n1103 | n1108 ;
  assign n1110 = n159 & n965 ;
  assign n1111 = n1109 | n1110 ;
  assign n1112 = x14 | n965 ;
  assign n1113 = ( x14 & n159 ) | ( x14 & n1112 ) | ( n159 & n1112 ) ;
  assign n1114 = n1109 | n1113 ;
  assign n1115 = ~x14 & n1113 ;
  assign n1116 = ( ~x14 & n1109 ) | ( ~x14 & n1115 ) | ( n1109 & n1115 ) ;
  assign n1117 = ( ~n1111 & n1114 ) | ( ~n1111 & n1116 ) | ( n1114 & n1116 ) ;
  assign n1118 = n977 | n1117 ;
  assign n1119 = n977 & n1117 ;
  assign n1120 = n1118 & ~n1119 ;
  assign n1121 = n293 & n639 ;
  assign n1122 = x69 & n636 ;
  assign n1123 = x68 & n631 ;
  assign n1124 = x67 & ~n630 ;
  assign n1125 = n764 & n1124 ;
  assign n1126 = n1123 | n1125 ;
  assign n1127 = n1122 | n1126 ;
  assign n1128 = n1121 | n1127 ;
  assign n1129 = x11 | n1122 ;
  assign n1130 = n1126 | n1129 ;
  assign n1131 = n1121 | n1130 ;
  assign n1132 = ~x11 & n1130 ;
  assign n1133 = ( ~x11 & n1121 ) | ( ~x11 & n1132 ) | ( n1121 & n1132 ) ;
  assign n1134 = ( ~n1128 & n1131 ) | ( ~n1128 & n1133 ) | ( n1131 & n1133 ) ;
  assign n1135 = n1120 | n1134 ;
  assign n1136 = n1120 & n1134 ;
  assign n1137 = n1135 & ~n1136 ;
  assign n1138 = n999 | n1001 ;
  assign n1139 = ( n999 & n1000 ) | ( n999 & n1138 ) | ( n1000 & n1138 ) ;
  assign n1140 = n1137 & n1139 ;
  assign n1141 = n1137 & ~n1140 ;
  assign n1142 = ~n1137 & n1139 ;
  assign n1143 = n1102 & n1142 ;
  assign n1144 = ( n1102 & n1141 ) | ( n1102 & n1143 ) | ( n1141 & n1143 ) ;
  assign n1145 = n1102 | n1142 ;
  assign n1146 = n1141 | n1145 ;
  assign n1147 = ~n1144 & n1146 ;
  assign n1148 = n1021 & n1147 ;
  assign n1149 = ( n1028 & n1147 ) | ( n1028 & n1148 ) | ( n1147 & n1148 ) ;
  assign n1150 = n1021 | n1147 ;
  assign n1151 = n1028 | n1150 ;
  assign n1152 = ~n1149 & n1151 ;
  assign n1153 = x75 & n212 ;
  assign n1154 = x74 & n207 ;
  assign n1155 = x73 & ~n206 ;
  assign n1156 = n267 & n1155 ;
  assign n1157 = n1154 | n1156 ;
  assign n1158 = n1153 | n1157 ;
  assign n1159 = n215 | n1153 ;
  assign n1160 = n1157 | n1159 ;
  assign n1161 = ( n746 & n1158 ) | ( n746 & n1160 ) | ( n1158 & n1160 ) ;
  assign n1162 = x5 & n1160 ;
  assign n1163 = x5 & n1153 ;
  assign n1164 = ( x5 & n1157 ) | ( x5 & n1163 ) | ( n1157 & n1163 ) ;
  assign n1165 = ( n746 & n1162 ) | ( n746 & n1164 ) | ( n1162 & n1164 ) ;
  assign n1166 = x5 & ~n1164 ;
  assign n1167 = x5 & ~n1160 ;
  assign n1168 = ( ~n746 & n1166 ) | ( ~n746 & n1167 ) | ( n1166 & n1167 ) ;
  assign n1169 = ( n1161 & ~n1165 ) | ( n1161 & n1168 ) | ( ~n1165 & n1168 ) ;
  assign n1170 = n1152 | n1169 ;
  assign n1171 = n1152 & n1169 ;
  assign n1172 = n1170 & ~n1171 ;
  assign n1173 = n1047 | n1048 ;
  assign n1174 = ( n953 & n1047 ) | ( n953 & n1173 ) | ( n1047 & n1173 ) ;
  assign n1175 = n1172 & n1174 ;
  assign n1176 = n1172 | n1174 ;
  assign n1177 = ~n1175 & n1176 ;
  assign n1178 = x77 | x78 ;
  assign n1179 = x77 & x78 ;
  assign n1180 = n1178 & ~n1179 ;
  assign n1181 = n1053 | n1054 ;
  assign n1182 = n1180 & n1181 ;
  assign n1183 = n1053 & n1180 ;
  assign n1184 = ( n907 & n1182 ) | ( n907 & n1183 ) | ( n1182 & n1183 ) ;
  assign n1185 = n1182 | n1183 ;
  assign n1186 = ( n917 & n1184 ) | ( n917 & n1185 ) | ( n1184 & n1185 ) ;
  assign n1187 = n1180 | n1181 ;
  assign n1188 = n907 | n1053 ;
  assign n1189 = ( n1053 & n1054 ) | ( n1053 & n1188 ) | ( n1054 & n1188 ) ;
  assign n1190 = n1180 | n1189 ;
  assign n1191 = ( n917 & n1187 ) | ( n917 & n1190 ) | ( n1187 & n1190 ) ;
  assign n1192 = ~n1186 & n1191 ;
  assign n1193 = x77 & n133 ;
  assign n1194 = x76 & ~n162 ;
  assign n1195 = ( n137 & n1193 ) | ( n137 & n1194 ) | ( n1193 & n1194 ) ;
  assign n1196 = x0 & x78 ;
  assign n1197 = ( ~n137 & n1193 ) | ( ~n137 & n1196 ) | ( n1193 & n1196 ) ;
  assign n1198 = n1195 | n1197 ;
  assign n1199 = n141 | n1198 ;
  assign n1200 = ( n1192 & n1198 ) | ( n1192 & n1199 ) | ( n1198 & n1199 ) ;
  assign n1201 = x2 & n1198 ;
  assign n1202 = ( x2 & n523 ) | ( x2 & n1198 ) | ( n523 & n1198 ) ;
  assign n1203 = ( n1192 & n1201 ) | ( n1192 & n1202 ) | ( n1201 & n1202 ) ;
  assign n1204 = x2 & ~n1202 ;
  assign n1205 = x2 & ~n1198 ;
  assign n1206 = ( ~n1192 & n1204 ) | ( ~n1192 & n1205 ) | ( n1204 & n1205 ) ;
  assign n1207 = ( n1200 & ~n1203 ) | ( n1200 & n1206 ) | ( ~n1203 & n1206 ) ;
  assign n1208 = n1177 & ~n1207 ;
  assign n1209 = ~n1177 & n1207 ;
  assign n1210 = n1208 | n1209 ;
  assign n1211 = n1051 | n1076 ;
  assign n1212 = ( n1074 & n1083 ) | ( n1074 & n1211 ) | ( n1083 & n1211 ) ;
  assign n1213 = n1210 & n1212 ;
  assign n1214 = n1210 | n1212 ;
  assign n1215 = ~n1213 & n1214 ;
  assign n1216 = n1136 | n1140 ;
  assign n1217 = x14 & ~x15 ;
  assign n1218 = ~x14 & x15 ;
  assign n1219 = n1217 | n1218 ;
  assign n1220 = x64 & n1219 ;
  assign n1221 = ~n977 & n1220 ;
  assign n1222 = ( ~n1117 & n1220 ) | ( ~n1117 & n1221 ) | ( n1220 & n1221 ) ;
  assign n1223 = n977 & ~n1220 ;
  assign n1224 = n1117 & n1223 ;
  assign n1225 = n1222 | n1224 ;
  assign n1226 = x67 & n962 ;
  assign n1227 = x66 & n957 ;
  assign n1228 = x65 & ~n956 ;
  assign n1229 = n1105 & n1228 ;
  assign n1230 = n1227 | n1229 ;
  assign n1231 = n1226 | n1230 ;
  assign n1232 = n186 & n965 ;
  assign n1233 = n1231 | n1232 ;
  assign n1234 = x14 & ~n1233 ;
  assign n1235 = ~x14 & n1233 ;
  assign n1236 = n1234 | n1235 ;
  assign n1237 = n1225 & n1236 ;
  assign n1238 = n1225 | n1236 ;
  assign n1239 = ~n1237 & n1238 ;
  assign n1240 = x69 & n631 ;
  assign n1241 = x68 & ~n630 ;
  assign n1242 = n764 & n1241 ;
  assign n1243 = n1240 | n1242 ;
  assign n1244 = x70 & n636 ;
  assign n1245 = n639 | n1244 ;
  assign n1246 = n1243 | n1245 ;
  assign n1247 = x11 & ~n1246 ;
  assign n1248 = x11 & ~n1244 ;
  assign n1249 = ~n1243 & n1248 ;
  assign n1250 = ( ~n340 & n1247 ) | ( ~n340 & n1249 ) | ( n1247 & n1249 ) ;
  assign n1251 = ~x11 & n1246 ;
  assign n1252 = ~x11 & n1244 ;
  assign n1253 = ( ~x11 & n1243 ) | ( ~x11 & n1252 ) | ( n1243 & n1252 ) ;
  assign n1254 = ( n340 & n1251 ) | ( n340 & n1253 ) | ( n1251 & n1253 ) ;
  assign n1255 = n1250 | n1254 ;
  assign n1256 = n1239 & n1255 ;
  assign n1257 = n1239 & ~n1256 ;
  assign n1258 = ~n1239 & n1255 ;
  assign n1259 = n1216 & n1258 ;
  assign n1260 = ( n1216 & n1257 ) | ( n1216 & n1259 ) | ( n1257 & n1259 ) ;
  assign n1261 = n1216 | n1258 ;
  assign n1262 = n1257 | n1261 ;
  assign n1263 = ~n1260 & n1262 ;
  assign n1264 = x73 & n389 ;
  assign n1265 = x72 & n384 ;
  assign n1266 = x71 & ~n383 ;
  assign n1267 = n463 & n1266 ;
  assign n1268 = n1265 | n1267 ;
  assign n1269 = n1264 | n1268 ;
  assign n1270 = ( n392 & ~n610 ) | ( n392 & n1269 ) | ( ~n610 & n1269 ) ;
  assign n1271 = n392 & n1264 ;
  assign n1272 = ( n392 & n1268 ) | ( n392 & n1271 ) | ( n1268 & n1271 ) ;
  assign n1273 = ( n598 & n1270 ) | ( n598 & n1272 ) | ( n1270 & n1272 ) ;
  assign n1274 = ( x8 & ~n1269 ) | ( x8 & n1273 ) | ( ~n1269 & n1273 ) ;
  assign n1275 = ~n1273 & n1274 ;
  assign n1276 = x8 | n1264 ;
  assign n1277 = n1268 | n1276 ;
  assign n1278 = n1273 | n1277 ;
  assign n1279 = ( ~x8 & n1275 ) | ( ~x8 & n1278 ) | ( n1275 & n1278 ) ;
  assign n1280 = n1263 & n1279 ;
  assign n1281 = n1263 & ~n1280 ;
  assign n1282 = ~n1263 & n1279 ;
  assign n1283 = n1281 | n1282 ;
  assign n1284 = n1144 | n1149 ;
  assign n1285 = n1283 & n1284 ;
  assign n1286 = n1283 | n1284 ;
  assign n1287 = ~n1285 & n1286 ;
  assign n1288 = x76 & n212 ;
  assign n1289 = x75 & n207 ;
  assign n1290 = x74 & ~n206 ;
  assign n1291 = n267 & n1290 ;
  assign n1292 = n1289 | n1291 ;
  assign n1293 = n1288 | n1292 ;
  assign n1294 = n215 | n1288 ;
  assign n1295 = n1292 | n1294 ;
  assign n1296 = ( n923 & n1293 ) | ( n923 & n1295 ) | ( n1293 & n1295 ) ;
  assign n1297 = x5 & n1295 ;
  assign n1298 = x5 & n1288 ;
  assign n1299 = ( x5 & n1292 ) | ( x5 & n1298 ) | ( n1292 & n1298 ) ;
  assign n1300 = ( n923 & n1297 ) | ( n923 & n1299 ) | ( n1297 & n1299 ) ;
  assign n1301 = x5 & ~n1299 ;
  assign n1302 = x5 & ~n1295 ;
  assign n1303 = ( ~n923 & n1301 ) | ( ~n923 & n1302 ) | ( n1301 & n1302 ) ;
  assign n1304 = ( n1296 & ~n1300 ) | ( n1296 & n1303 ) | ( ~n1300 & n1303 ) ;
  assign n1305 = n1287 & n1304 ;
  assign n1306 = n1287 & ~n1305 ;
  assign n1307 = n1171 | n1172 ;
  assign n1308 = ( n1171 & n1174 ) | ( n1171 & n1307 ) | ( n1174 & n1307 ) ;
  assign n1309 = ~n1287 & n1304 ;
  assign n1310 = n1308 & n1309 ;
  assign n1311 = ( n1306 & n1308 ) | ( n1306 & n1310 ) | ( n1308 & n1310 ) ;
  assign n1312 = n1308 | n1309 ;
  assign n1313 = n1306 | n1312 ;
  assign n1314 = ~n1311 & n1313 ;
  assign n1315 = x78 | x79 ;
  assign n1316 = x78 & x79 ;
  assign n1317 = n1315 & ~n1316 ;
  assign n1318 = n1179 | n1180 ;
  assign n1319 = ( n1179 & n1181 ) | ( n1179 & n1318 ) | ( n1181 & n1318 ) ;
  assign n1320 = n1317 & n1319 ;
  assign n1321 = n1053 | n1179 ;
  assign n1322 = ( n1179 & n1180 ) | ( n1179 & n1321 ) | ( n1180 & n1321 ) ;
  assign n1323 = n1317 & n1322 ;
  assign n1324 = ( n907 & n1320 ) | ( n907 & n1323 ) | ( n1320 & n1323 ) ;
  assign n1325 = n1320 | n1323 ;
  assign n1326 = ( n917 & n1324 ) | ( n917 & n1325 ) | ( n1324 & n1325 ) ;
  assign n1327 = n1317 | n1322 ;
  assign n1328 = n1319 | n1327 ;
  assign n1329 = n907 | n1317 ;
  assign n1330 = ( n1319 & n1327 ) | ( n1319 & n1329 ) | ( n1327 & n1329 ) ;
  assign n1331 = ( n917 & n1328 ) | ( n917 & n1330 ) | ( n1328 & n1330 ) ;
  assign n1332 = ~n1326 & n1331 ;
  assign n1333 = x78 & n133 ;
  assign n1334 = x77 & ~n162 ;
  assign n1335 = ( n137 & n1333 ) | ( n137 & n1334 ) | ( n1333 & n1334 ) ;
  assign n1336 = x0 & x79 ;
  assign n1337 = ( ~n137 & n1333 ) | ( ~n137 & n1336 ) | ( n1333 & n1336 ) ;
  assign n1338 = n1335 | n1337 ;
  assign n1339 = n141 | n1338 ;
  assign n1340 = ( n1332 & n1338 ) | ( n1332 & n1339 ) | ( n1338 & n1339 ) ;
  assign n1341 = x2 & n1338 ;
  assign n1342 = ( x2 & n523 ) | ( x2 & n1338 ) | ( n523 & n1338 ) ;
  assign n1343 = ( n1332 & n1341 ) | ( n1332 & n1342 ) | ( n1341 & n1342 ) ;
  assign n1344 = x2 & ~n1342 ;
  assign n1345 = x2 & ~n1338 ;
  assign n1346 = ( ~n1332 & n1344 ) | ( ~n1332 & n1345 ) | ( n1344 & n1345 ) ;
  assign n1347 = ( n1340 & ~n1343 ) | ( n1340 & n1346 ) | ( ~n1343 & n1346 ) ;
  assign n1348 = n1314 & n1347 ;
  assign n1349 = n1314 & ~n1348 ;
  assign n1350 = ~n1314 & n1347 ;
  assign n1351 = n1349 | n1350 ;
  assign n1352 = ( n1177 & n1207 ) | ( n1177 & n1211 ) | ( n1207 & n1211 ) ;
  assign n1353 = ( n1074 & n1177 ) | ( n1074 & n1207 ) | ( n1177 & n1207 ) ;
  assign n1354 = ( n1083 & n1352 ) | ( n1083 & n1353 ) | ( n1352 & n1353 ) ;
  assign n1355 = n1351 | n1354 ;
  assign n1356 = ~n1354 & n1355 ;
  assign n1357 = ( ~n1351 & n1355 ) | ( ~n1351 & n1356 ) | ( n1355 & n1356 ) ;
  assign n1358 = n1305 | n1311 ;
  assign n1359 = x70 & n631 ;
  assign n1360 = x69 & ~n630 ;
  assign n1361 = n764 & n1360 ;
  assign n1362 = n1359 | n1361 ;
  assign n1363 = x71 & n636 ;
  assign n1364 = n639 | n1363 ;
  assign n1365 = n1362 | n1364 ;
  assign n1366 = x11 & ~n1365 ;
  assign n1367 = x11 & ~n1363 ;
  assign n1368 = ~n1362 & n1367 ;
  assign n1369 = ( ~n438 & n1366 ) | ( ~n438 & n1368 ) | ( n1366 & n1368 ) ;
  assign n1370 = ~x11 & n1365 ;
  assign n1371 = ~x11 & n1363 ;
  assign n1372 = ( ~x11 & n1362 ) | ( ~x11 & n1371 ) | ( n1362 & n1371 ) ;
  assign n1373 = ( n438 & n1370 ) | ( n438 & n1372 ) | ( n1370 & n1372 ) ;
  assign n1374 = n1369 | n1373 ;
  assign n1375 = ~x15 & x16 ;
  assign n1376 = x15 & ~x16 ;
  assign n1377 = n1375 | n1376 ;
  assign n1378 = ~n1219 & n1377 ;
  assign n1379 = x64 & n1378 ;
  assign n1380 = ~x16 & x17 ;
  assign n1381 = x16 & ~x17 ;
  assign n1382 = n1380 | n1381 ;
  assign n1383 = n1219 & ~n1382 ;
  assign n1384 = x65 & n1383 ;
  assign n1385 = n1379 | n1384 ;
  assign n1386 = n1219 & n1382 ;
  assign n1387 = x17 | n144 ;
  assign n1388 = ( x17 & n1386 ) | ( x17 & n1387 ) | ( n1386 & n1387 ) ;
  assign n1389 = ~x17 & n1388 ;
  assign n1390 = ( ~x17 & n1385 ) | ( ~x17 & n1389 ) | ( n1385 & n1389 ) ;
  assign n1391 = x17 & ~x64 ;
  assign n1392 = ( x17 & ~n1219 ) | ( x17 & n1391 ) | ( ~n1219 & n1391 ) ;
  assign n1393 = n1388 & n1392 ;
  assign n1394 = ( n1385 & n1392 ) | ( n1385 & n1393 ) | ( n1392 & n1393 ) ;
  assign n1395 = n144 & n1386 ;
  assign n1396 = n1392 & ~n1395 ;
  assign n1397 = ~n1385 & n1396 ;
  assign n1398 = ( n1390 & n1394 ) | ( n1390 & n1397 ) | ( n1394 & n1397 ) ;
  assign n1399 = n1388 | n1392 ;
  assign n1400 = n1385 | n1399 ;
  assign n1401 = ~n1392 & n1395 ;
  assign n1402 = ( n1385 & ~n1392 ) | ( n1385 & n1401 ) | ( ~n1392 & n1401 ) ;
  assign n1403 = ( n1390 & n1400 ) | ( n1390 & ~n1402 ) | ( n1400 & ~n1402 ) ;
  assign n1404 = ~n1398 & n1403 ;
  assign n1405 = n241 & n965 ;
  assign n1406 = x68 & n962 ;
  assign n1407 = x67 & n957 ;
  assign n1408 = x66 & ~n956 ;
  assign n1409 = n1105 & n1408 ;
  assign n1410 = n1407 | n1409 ;
  assign n1411 = n1406 | n1410 ;
  assign n1412 = n1405 | n1411 ;
  assign n1413 = x14 | n1406 ;
  assign n1414 = n1410 | n1413 ;
  assign n1415 = n1405 | n1414 ;
  assign n1416 = ~x14 & n1414 ;
  assign n1417 = ( ~x14 & n1405 ) | ( ~x14 & n1416 ) | ( n1405 & n1416 ) ;
  assign n1418 = ( ~n1412 & n1415 ) | ( ~n1412 & n1417 ) | ( n1415 & n1417 ) ;
  assign n1419 = n1404 | n1418 ;
  assign n1420 = n1404 & n1418 ;
  assign n1421 = n1419 & ~n1420 ;
  assign n1422 = ( n1119 & n1220 ) | ( n1119 & n1236 ) | ( n1220 & n1236 ) ;
  assign n1423 = n1421 | n1422 ;
  assign n1424 = n1421 & n1422 ;
  assign n1425 = n1423 & ~n1424 ;
  assign n1426 = n1374 | n1425 ;
  assign n1427 = n1374 & n1425 ;
  assign n1428 = n1426 & ~n1427 ;
  assign n1429 = n1256 | n1257 ;
  assign n1430 = n1216 | n1256 ;
  assign n1431 = ( n1259 & n1429 ) | ( n1259 & n1430 ) | ( n1429 & n1430 ) ;
  assign n1432 = n1428 & n1431 ;
  assign n1433 = n1428 | n1431 ;
  assign n1434 = ~n1432 & n1433 ;
  assign n1435 = x74 & n389 ;
  assign n1436 = x73 & n384 ;
  assign n1437 = x72 & ~n383 ;
  assign n1438 = n463 & n1437 ;
  assign n1439 = n1436 | n1438 ;
  assign n1440 = n1435 | n1439 ;
  assign n1441 = n392 | n1435 ;
  assign n1442 = n1439 | n1441 ;
  assign n1443 = ( n710 & n1440 ) | ( n710 & n1442 ) | ( n1440 & n1442 ) ;
  assign n1444 = x8 & n1442 ;
  assign n1445 = x8 & n1435 ;
  assign n1446 = ( x8 & n1439 ) | ( x8 & n1445 ) | ( n1439 & n1445 ) ;
  assign n1447 = ( n710 & n1444 ) | ( n710 & n1446 ) | ( n1444 & n1446 ) ;
  assign n1448 = x8 & ~n1446 ;
  assign n1449 = x8 & ~n1442 ;
  assign n1450 = ( ~n710 & n1448 ) | ( ~n710 & n1449 ) | ( n1448 & n1449 ) ;
  assign n1451 = ( n1443 & ~n1447 ) | ( n1443 & n1450 ) | ( ~n1447 & n1450 ) ;
  assign n1452 = n1434 | n1451 ;
  assign n1453 = n1434 & n1451 ;
  assign n1454 = n1452 & ~n1453 ;
  assign n1455 = n1280 | n1284 ;
  assign n1456 = ( n1280 & n1283 ) | ( n1280 & n1455 ) | ( n1283 & n1455 ) ;
  assign n1457 = n1454 & n1456 ;
  assign n1458 = n1454 | n1456 ;
  assign n1459 = ~n1457 & n1458 ;
  assign n1460 = x77 & n212 ;
  assign n1461 = x76 & n207 ;
  assign n1462 = x75 & ~n206 ;
  assign n1463 = n267 & n1462 ;
  assign n1464 = n1461 | n1463 ;
  assign n1465 = n1460 | n1464 ;
  assign n1466 = n215 | n1460 ;
  assign n1467 = n1464 | n1466 ;
  assign n1468 = ( n1059 & n1465 ) | ( n1059 & n1467 ) | ( n1465 & n1467 ) ;
  assign n1469 = x5 & n1467 ;
  assign n1470 = x5 & n1460 ;
  assign n1471 = ( x5 & n1464 ) | ( x5 & n1470 ) | ( n1464 & n1470 ) ;
  assign n1472 = ( n1059 & n1469 ) | ( n1059 & n1471 ) | ( n1469 & n1471 ) ;
  assign n1473 = x5 & ~n1471 ;
  assign n1474 = x5 & ~n1467 ;
  assign n1475 = ( ~n1059 & n1473 ) | ( ~n1059 & n1474 ) | ( n1473 & n1474 ) ;
  assign n1476 = ( n1468 & ~n1472 ) | ( n1468 & n1475 ) | ( ~n1472 & n1475 ) ;
  assign n1477 = n1459 | n1476 ;
  assign n1478 = n1459 & n1476 ;
  assign n1479 = n1477 & ~n1478 ;
  assign n1480 = n1358 & n1479 ;
  assign n1481 = n1358 | n1479 ;
  assign n1482 = ~n1480 & n1481 ;
  assign n1483 = x79 | x80 ;
  assign n1484 = x79 & x80 ;
  assign n1485 = n1483 & ~n1484 ;
  assign n1486 = n1316 | n1317 ;
  assign n1487 = ( n1316 & n1319 ) | ( n1316 & n1486 ) | ( n1319 & n1486 ) ;
  assign n1488 = ( n1316 & n1322 ) | ( n1316 & n1486 ) | ( n1322 & n1486 ) ;
  assign n1489 = n1485 & n1488 ;
  assign n1490 = ( n1485 & n1487 ) | ( n1485 & n1489 ) | ( n1487 & n1489 ) ;
  assign n1491 = n907 & n1485 ;
  assign n1492 = ( n1487 & n1489 ) | ( n1487 & n1491 ) | ( n1489 & n1491 ) ;
  assign n1493 = ( n917 & n1490 ) | ( n917 & n1492 ) | ( n1490 & n1492 ) ;
  assign n1494 = n1485 | n1488 ;
  assign n1495 = n1487 | n1494 ;
  assign n1496 = n907 | n1485 ;
  assign n1497 = ( n1487 & n1494 ) | ( n1487 & n1496 ) | ( n1494 & n1496 ) ;
  assign n1498 = ( n917 & n1495 ) | ( n917 & n1497 ) | ( n1495 & n1497 ) ;
  assign n1499 = ~n1493 & n1498 ;
  assign n1500 = x79 & n133 ;
  assign n1501 = x78 & ~n162 ;
  assign n1502 = ( n137 & n1500 ) | ( n137 & n1501 ) | ( n1500 & n1501 ) ;
  assign n1503 = x0 & x80 ;
  assign n1504 = ( ~n137 & n1500 ) | ( ~n137 & n1503 ) | ( n1500 & n1503 ) ;
  assign n1505 = n1502 | n1504 ;
  assign n1506 = n141 | n1505 ;
  assign n1507 = ( n1499 & n1505 ) | ( n1499 & n1506 ) | ( n1505 & n1506 ) ;
  assign n1508 = x2 & n1505 ;
  assign n1509 = ( x2 & n523 ) | ( x2 & n1505 ) | ( n523 & n1505 ) ;
  assign n1510 = ( n1499 & n1508 ) | ( n1499 & n1509 ) | ( n1508 & n1509 ) ;
  assign n1511 = x2 & ~n1509 ;
  assign n1512 = x2 & ~n1505 ;
  assign n1513 = ( ~n1499 & n1511 ) | ( ~n1499 & n1512 ) | ( n1511 & n1512 ) ;
  assign n1514 = ( n1507 & ~n1510 ) | ( n1507 & n1513 ) | ( ~n1510 & n1513 ) ;
  assign n1515 = n1482 & n1514 ;
  assign n1516 = ~n1482 & n1514 ;
  assign n1517 = ( n1482 & ~n1515 ) | ( n1482 & n1516 ) | ( ~n1515 & n1516 ) ;
  assign n1518 = n1350 & n1354 ;
  assign n1519 = ( n1349 & n1354 ) | ( n1349 & n1518 ) | ( n1354 & n1518 ) ;
  assign n1520 = n1348 | n1519 ;
  assign n1521 = n1517 & n1520 ;
  assign n1522 = n1517 | n1520 ;
  assign n1523 = ~n1521 & n1522 ;
  assign n1524 = x72 & n636 ;
  assign n1525 = x71 & n631 ;
  assign n1526 = x70 & ~n630 ;
  assign n1527 = n764 & n1526 ;
  assign n1528 = n1525 | n1527 ;
  assign n1529 = n1524 | n1528 ;
  assign n1530 = ( n513 & n639 ) | ( n513 & n1529 ) | ( n639 & n1529 ) ;
  assign n1531 = ( x11 & n639 ) | ( x11 & ~n1524 ) | ( n639 & ~n1524 ) ;
  assign n1532 = x11 & n639 ;
  assign n1533 = ( ~n1528 & n1531 ) | ( ~n1528 & n1532 ) | ( n1531 & n1532 ) ;
  assign n1534 = ( x11 & n513 ) | ( x11 & n1533 ) | ( n513 & n1533 ) ;
  assign n1535 = ~n1530 & n1534 ;
  assign n1536 = n1529 | n1533 ;
  assign n1537 = x11 | n1529 ;
  assign n1538 = ( n513 & n1536 ) | ( n513 & n1537 ) | ( n1536 & n1537 ) ;
  assign n1539 = ( ~x11 & n1535 ) | ( ~x11 & n1538 ) | ( n1535 & n1538 ) ;
  assign n1540 = x66 & n1383 ;
  assign n1541 = x65 & n1378 ;
  assign n1542 = ~n1219 & n1382 ;
  assign n1543 = x64 & ~n1377 ;
  assign n1544 = n1542 & n1543 ;
  assign n1545 = n1541 | n1544 ;
  assign n1546 = n1540 | n1545 ;
  assign n1547 = n159 & n1386 ;
  assign n1548 = n1546 | n1547 ;
  assign n1549 = x17 | n1386 ;
  assign n1550 = ( x17 & n159 ) | ( x17 & n1549 ) | ( n159 & n1549 ) ;
  assign n1551 = n1546 | n1550 ;
  assign n1552 = ~x17 & n1550 ;
  assign n1553 = ( ~x17 & n1546 ) | ( ~x17 & n1552 ) | ( n1546 & n1552 ) ;
  assign n1554 = ( ~n1548 & n1551 ) | ( ~n1548 & n1553 ) | ( n1551 & n1553 ) ;
  assign n1555 = n1398 | n1554 ;
  assign n1556 = n1398 & n1554 ;
  assign n1557 = n1555 & ~n1556 ;
  assign n1558 = n293 & n965 ;
  assign n1559 = x69 & n962 ;
  assign n1560 = x68 & n957 ;
  assign n1561 = x67 & ~n956 ;
  assign n1562 = n1105 & n1561 ;
  assign n1563 = n1560 | n1562 ;
  assign n1564 = n1559 | n1563 ;
  assign n1565 = n1558 | n1564 ;
  assign n1566 = x14 | n1559 ;
  assign n1567 = n1563 | n1566 ;
  assign n1568 = n1558 | n1567 ;
  assign n1569 = ~x14 & n1567 ;
  assign n1570 = ( ~x14 & n1558 ) | ( ~x14 & n1569 ) | ( n1558 & n1569 ) ;
  assign n1571 = ( ~n1565 & n1568 ) | ( ~n1565 & n1570 ) | ( n1568 & n1570 ) ;
  assign n1572 = n1557 | n1571 ;
  assign n1573 = n1557 & n1571 ;
  assign n1574 = n1572 & ~n1573 ;
  assign n1575 = n1420 | n1422 ;
  assign n1576 = ( n1420 & n1421 ) | ( n1420 & n1575 ) | ( n1421 & n1575 ) ;
  assign n1577 = n1574 & n1576 ;
  assign n1578 = n1574 & ~n1577 ;
  assign n1579 = ~n1574 & n1576 ;
  assign n1580 = n1539 & n1579 ;
  assign n1581 = ( n1539 & n1578 ) | ( n1539 & n1580 ) | ( n1578 & n1580 ) ;
  assign n1582 = n1539 | n1579 ;
  assign n1583 = n1578 | n1582 ;
  assign n1584 = ~n1581 & n1583 ;
  assign n1585 = n1427 | n1428 ;
  assign n1586 = ( n1427 & n1431 ) | ( n1427 & n1585 ) | ( n1431 & n1585 ) ;
  assign n1587 = n1584 & n1586 ;
  assign n1588 = n1584 | n1586 ;
  assign n1589 = ~n1587 & n1588 ;
  assign n1590 = x75 & n389 ;
  assign n1591 = x74 & n384 ;
  assign n1592 = x73 & ~n383 ;
  assign n1593 = n463 & n1592 ;
  assign n1594 = n1591 | n1593 ;
  assign n1595 = n1590 | n1594 ;
  assign n1596 = n392 | n1590 ;
  assign n1597 = n1594 | n1596 ;
  assign n1598 = ( n746 & n1595 ) | ( n746 & n1597 ) | ( n1595 & n1597 ) ;
  assign n1599 = x8 & n1597 ;
  assign n1600 = x8 & n1590 ;
  assign n1601 = ( x8 & n1594 ) | ( x8 & n1600 ) | ( n1594 & n1600 ) ;
  assign n1602 = ( n746 & n1599 ) | ( n746 & n1601 ) | ( n1599 & n1601 ) ;
  assign n1603 = x8 & ~n1601 ;
  assign n1604 = x8 & ~n1597 ;
  assign n1605 = ( ~n746 & n1603 ) | ( ~n746 & n1604 ) | ( n1603 & n1604 ) ;
  assign n1606 = ( n1598 & ~n1602 ) | ( n1598 & n1605 ) | ( ~n1602 & n1605 ) ;
  assign n1607 = n1589 | n1606 ;
  assign n1608 = n1589 & n1606 ;
  assign n1609 = n1607 & ~n1608 ;
  assign n1610 = n1453 | n1454 ;
  assign n1611 = ( n1453 & n1456 ) | ( n1453 & n1610 ) | ( n1456 & n1610 ) ;
  assign n1612 = n1609 & n1611 ;
  assign n1613 = n1609 | n1611 ;
  assign n1614 = ~n1612 & n1613 ;
  assign n1615 = x78 & n212 ;
  assign n1616 = x77 & n207 ;
  assign n1617 = x76 & ~n206 ;
  assign n1618 = n267 & n1617 ;
  assign n1619 = n1616 | n1618 ;
  assign n1620 = n1615 | n1619 ;
  assign n1621 = n215 | n1615 ;
  assign n1622 = n1619 | n1621 ;
  assign n1623 = ( n1192 & n1620 ) | ( n1192 & n1622 ) | ( n1620 & n1622 ) ;
  assign n1624 = x5 & n1622 ;
  assign n1625 = x5 & n1615 ;
  assign n1626 = ( x5 & n1619 ) | ( x5 & n1625 ) | ( n1619 & n1625 ) ;
  assign n1627 = ( n1192 & n1624 ) | ( n1192 & n1626 ) | ( n1624 & n1626 ) ;
  assign n1628 = x5 & ~n1626 ;
  assign n1629 = x5 & ~n1622 ;
  assign n1630 = ( ~n1192 & n1628 ) | ( ~n1192 & n1629 ) | ( n1628 & n1629 ) ;
  assign n1631 = ( n1623 & ~n1627 ) | ( n1623 & n1630 ) | ( ~n1627 & n1630 ) ;
  assign n1632 = n1614 | n1631 ;
  assign n1633 = n1614 & n1631 ;
  assign n1634 = n1632 & ~n1633 ;
  assign n1635 = n1478 | n1479 ;
  assign n1636 = ( n1358 & n1478 ) | ( n1358 & n1635 ) | ( n1478 & n1635 ) ;
  assign n1637 = n1634 & n1636 ;
  assign n1638 = n1634 | n1636 ;
  assign n1639 = ~n1637 & n1638 ;
  assign n1640 = x80 | x81 ;
  assign n1641 = x80 & x81 ;
  assign n1642 = n1640 & ~n1641 ;
  assign n1643 = n1484 & n1642 ;
  assign n1644 = ( n1492 & n1642 ) | ( n1492 & n1643 ) | ( n1642 & n1643 ) ;
  assign n1645 = ( n1490 & n1642 ) | ( n1490 & n1643 ) | ( n1642 & n1643 ) ;
  assign n1646 = ( n917 & n1644 ) | ( n917 & n1645 ) | ( n1644 & n1645 ) ;
  assign n1647 = n1484 | n1642 ;
  assign n1648 = n1492 | n1647 ;
  assign n1649 = n1490 | n1647 ;
  assign n1650 = ( n917 & n1648 ) | ( n917 & n1649 ) | ( n1648 & n1649 ) ;
  assign n1651 = ~n1646 & n1650 ;
  assign n1652 = x80 & n133 ;
  assign n1653 = x79 & ~n162 ;
  assign n1654 = ( n137 & n1652 ) | ( n137 & n1653 ) | ( n1652 & n1653 ) ;
  assign n1655 = x0 & x81 ;
  assign n1656 = ( ~n137 & n1652 ) | ( ~n137 & n1655 ) | ( n1652 & n1655 ) ;
  assign n1657 = n1654 | n1656 ;
  assign n1658 = n141 | n1657 ;
  assign n1659 = ( n1651 & n1657 ) | ( n1651 & n1658 ) | ( n1657 & n1658 ) ;
  assign n1660 = x2 & n1657 ;
  assign n1661 = ( x2 & n523 ) | ( x2 & n1657 ) | ( n523 & n1657 ) ;
  assign n1662 = ( n1651 & n1660 ) | ( n1651 & n1661 ) | ( n1660 & n1661 ) ;
  assign n1663 = x2 & ~n1661 ;
  assign n1664 = x2 & ~n1657 ;
  assign n1665 = ( ~n1651 & n1663 ) | ( ~n1651 & n1664 ) | ( n1663 & n1664 ) ;
  assign n1666 = ( n1659 & ~n1662 ) | ( n1659 & n1665 ) | ( ~n1662 & n1665 ) ;
  assign n1667 = n1639 & n1666 ;
  assign n1668 = n1639 & ~n1667 ;
  assign n1669 = ~n1639 & n1666 ;
  assign n1670 = n1668 | n1669 ;
  assign n1671 = n1515 | n1521 ;
  assign n1672 = n1670 & n1671 ;
  assign n1673 = n1670 | n1671 ;
  assign n1674 = ~n1672 & n1673 ;
  assign n1675 = n1573 | n1577 ;
  assign n1676 = x17 & ~x18 ;
  assign n1677 = ~x17 & x18 ;
  assign n1678 = n1676 | n1677 ;
  assign n1679 = x64 & n1678 ;
  assign n1680 = ~n1398 & n1679 ;
  assign n1681 = ( ~n1554 & n1679 ) | ( ~n1554 & n1680 ) | ( n1679 & n1680 ) ;
  assign n1682 = n1398 & ~n1679 ;
  assign n1683 = n1554 & n1682 ;
  assign n1684 = n1681 | n1683 ;
  assign n1685 = x67 & n1383 ;
  assign n1686 = x66 & n1378 ;
  assign n1687 = x65 & ~n1377 ;
  assign n1688 = n1542 & n1687 ;
  assign n1689 = n1686 | n1688 ;
  assign n1690 = n1685 | n1689 ;
  assign n1691 = n186 & n1386 ;
  assign n1692 = n1690 | n1691 ;
  assign n1693 = x17 & ~n1692 ;
  assign n1694 = ~x17 & n1692 ;
  assign n1695 = n1693 | n1694 ;
  assign n1696 = n1684 & n1695 ;
  assign n1697 = n1684 | n1695 ;
  assign n1698 = ~n1696 & n1697 ;
  assign n1699 = x69 & n957 ;
  assign n1700 = x68 & ~n956 ;
  assign n1701 = n1105 & n1700 ;
  assign n1702 = n1699 | n1701 ;
  assign n1703 = x70 & n962 ;
  assign n1704 = n965 | n1703 ;
  assign n1705 = n1702 | n1704 ;
  assign n1706 = x14 & ~n1705 ;
  assign n1707 = x14 & ~n1703 ;
  assign n1708 = ~n1702 & n1707 ;
  assign n1709 = ( ~n340 & n1706 ) | ( ~n340 & n1708 ) | ( n1706 & n1708 ) ;
  assign n1710 = ~x14 & n1705 ;
  assign n1711 = ~x14 & n1703 ;
  assign n1712 = ( ~x14 & n1702 ) | ( ~x14 & n1711 ) | ( n1702 & n1711 ) ;
  assign n1713 = ( n340 & n1710 ) | ( n340 & n1712 ) | ( n1710 & n1712 ) ;
  assign n1714 = n1709 | n1713 ;
  assign n1715 = ( n1573 & ~n1698 ) | ( n1573 & n1714 ) | ( ~n1698 & n1714 ) ;
  assign n1716 = n1698 & ~n1714 ;
  assign n1717 = ( n1577 & n1715 ) | ( n1577 & ~n1716 ) | ( n1715 & ~n1716 ) ;
  assign n1718 = ( ~n1675 & n1698 ) | ( ~n1675 & n1717 ) | ( n1698 & n1717 ) ;
  assign n1719 = x73 & n636 ;
  assign n1720 = x72 & n631 ;
  assign n1721 = x71 & ~n630 ;
  assign n1722 = n764 & n1721 ;
  assign n1723 = n1720 | n1722 ;
  assign n1724 = n1719 | n1723 ;
  assign n1725 = n639 | n1719 ;
  assign n1726 = n1723 | n1725 ;
  assign n1727 = ( ~n610 & n1724 ) | ( ~n610 & n1726 ) | ( n1724 & n1726 ) ;
  assign n1728 = n1724 & n1726 ;
  assign n1729 = ( n598 & n1727 ) | ( n598 & n1728 ) | ( n1727 & n1728 ) ;
  assign n1730 = x11 & n1729 ;
  assign n1731 = x11 | n1729 ;
  assign n1732 = ~n1730 & n1731 ;
  assign n1733 = n1717 & n1732 ;
  assign n1734 = ~n1714 & n1732 ;
  assign n1735 = ( n1718 & n1733 ) | ( n1718 & n1734 ) | ( n1733 & n1734 ) ;
  assign n1736 = n1717 | n1732 ;
  assign n1737 = n1714 & ~n1732 ;
  assign n1738 = ( n1718 & n1736 ) | ( n1718 & ~n1737 ) | ( n1736 & ~n1737 ) ;
  assign n1739 = ~n1735 & n1738 ;
  assign n1740 = n1581 | n1584 ;
  assign n1741 = ( n1581 & n1586 ) | ( n1581 & n1740 ) | ( n1586 & n1740 ) ;
  assign n1742 = n1739 & n1741 ;
  assign n1743 = n1739 | n1741 ;
  assign n1744 = ~n1742 & n1743 ;
  assign n1745 = x76 & n389 ;
  assign n1746 = x75 & n384 ;
  assign n1747 = x74 & ~n383 ;
  assign n1748 = n463 & n1747 ;
  assign n1749 = n1746 | n1748 ;
  assign n1750 = n1745 | n1749 ;
  assign n1751 = n392 | n1745 ;
  assign n1752 = n1749 | n1751 ;
  assign n1753 = ( n923 & n1750 ) | ( n923 & n1752 ) | ( n1750 & n1752 ) ;
  assign n1754 = x8 & n1752 ;
  assign n1755 = x8 & n1745 ;
  assign n1756 = ( x8 & n1749 ) | ( x8 & n1755 ) | ( n1749 & n1755 ) ;
  assign n1757 = ( n923 & n1754 ) | ( n923 & n1756 ) | ( n1754 & n1756 ) ;
  assign n1758 = x8 & ~n1756 ;
  assign n1759 = x8 & ~n1752 ;
  assign n1760 = ( ~n923 & n1758 ) | ( ~n923 & n1759 ) | ( n1758 & n1759 ) ;
  assign n1761 = ( n1753 & ~n1757 ) | ( n1753 & n1760 ) | ( ~n1757 & n1760 ) ;
  assign n1762 = n1744 | n1761 ;
  assign n1763 = n1744 & n1761 ;
  assign n1764 = n1762 & ~n1763 ;
  assign n1765 = n1608 | n1609 ;
  assign n1766 = ( n1608 & n1611 ) | ( n1608 & n1765 ) | ( n1611 & n1765 ) ;
  assign n1767 = n1764 & n1766 ;
  assign n1768 = n1764 | n1766 ;
  assign n1769 = ~n1767 & n1768 ;
  assign n1770 = x79 & n212 ;
  assign n1771 = x78 & n207 ;
  assign n1772 = x77 & ~n206 ;
  assign n1773 = n267 & n1772 ;
  assign n1774 = n1771 | n1773 ;
  assign n1775 = n1770 | n1774 ;
  assign n1776 = n215 | n1770 ;
  assign n1777 = n1774 | n1776 ;
  assign n1778 = ( n1332 & n1775 ) | ( n1332 & n1777 ) | ( n1775 & n1777 ) ;
  assign n1779 = x5 & n1777 ;
  assign n1780 = x5 & n1770 ;
  assign n1781 = ( x5 & n1774 ) | ( x5 & n1780 ) | ( n1774 & n1780 ) ;
  assign n1782 = ( n1332 & n1779 ) | ( n1332 & n1781 ) | ( n1779 & n1781 ) ;
  assign n1783 = x5 & ~n1781 ;
  assign n1784 = x5 & ~n1777 ;
  assign n1785 = ( ~n1332 & n1783 ) | ( ~n1332 & n1784 ) | ( n1783 & n1784 ) ;
  assign n1786 = ( n1778 & ~n1782 ) | ( n1778 & n1785 ) | ( ~n1782 & n1785 ) ;
  assign n1787 = n1769 & n1786 ;
  assign n1788 = n1769 | n1786 ;
  assign n1789 = ~n1787 & n1788 ;
  assign n1790 = n1633 | n1634 ;
  assign n1791 = ( n1633 & n1636 ) | ( n1633 & n1790 ) | ( n1636 & n1790 ) ;
  assign n1792 = n1789 & n1791 ;
  assign n1793 = n1789 | n1791 ;
  assign n1794 = ~n1792 & n1793 ;
  assign n1795 = x81 | x82 ;
  assign n1796 = x81 & x82 ;
  assign n1797 = n1795 & ~n1796 ;
  assign n1798 = n1484 | n1641 ;
  assign n1799 = ( n1641 & n1642 ) | ( n1641 & n1798 ) | ( n1642 & n1798 ) ;
  assign n1800 = n1797 & n1799 ;
  assign n1801 = n1641 | n1642 ;
  assign n1802 = n1797 & n1801 ;
  assign n1803 = ( n1492 & n1800 ) | ( n1492 & n1802 ) | ( n1800 & n1802 ) ;
  assign n1804 = ( n1490 & n1800 ) | ( n1490 & n1802 ) | ( n1800 & n1802 ) ;
  assign n1805 = ( n917 & n1803 ) | ( n917 & n1804 ) | ( n1803 & n1804 ) ;
  assign n1806 = n1797 | n1799 ;
  assign n1807 = n1797 | n1801 ;
  assign n1808 = ( n1492 & n1806 ) | ( n1492 & n1807 ) | ( n1806 & n1807 ) ;
  assign n1809 = ( n1490 & n1806 ) | ( n1490 & n1807 ) | ( n1806 & n1807 ) ;
  assign n1810 = ( n917 & n1808 ) | ( n917 & n1809 ) | ( n1808 & n1809 ) ;
  assign n1811 = ~n1805 & n1810 ;
  assign n1812 = x81 & n133 ;
  assign n1813 = x80 & ~n162 ;
  assign n1814 = ( n137 & n1812 ) | ( n137 & n1813 ) | ( n1812 & n1813 ) ;
  assign n1815 = x0 & x82 ;
  assign n1816 = ( ~n137 & n1812 ) | ( ~n137 & n1815 ) | ( n1812 & n1815 ) ;
  assign n1817 = n1814 | n1816 ;
  assign n1818 = n141 | n1817 ;
  assign n1819 = ( n1811 & n1817 ) | ( n1811 & n1818 ) | ( n1817 & n1818 ) ;
  assign n1820 = x2 & n1817 ;
  assign n1821 = ( x2 & n523 ) | ( x2 & n1817 ) | ( n523 & n1817 ) ;
  assign n1822 = ( n1811 & n1820 ) | ( n1811 & n1821 ) | ( n1820 & n1821 ) ;
  assign n1823 = x2 & ~n1821 ;
  assign n1824 = x2 & ~n1817 ;
  assign n1825 = ( ~n1811 & n1823 ) | ( ~n1811 & n1824 ) | ( n1823 & n1824 ) ;
  assign n1826 = ( n1819 & ~n1822 ) | ( n1819 & n1825 ) | ( ~n1822 & n1825 ) ;
  assign n1827 = n1794 & n1826 ;
  assign n1828 = n1794 & ~n1827 ;
  assign n1829 = ~n1794 & n1826 ;
  assign n1830 = n1828 | n1829 ;
  assign n1831 = n1667 | n1672 ;
  assign n1832 = n1830 & n1831 ;
  assign n1833 = n1830 | n1831 ;
  assign n1834 = ~n1832 & n1833 ;
  assign n1835 = x70 & n957 ;
  assign n1836 = x69 & ~n956 ;
  assign n1837 = n1105 & n1836 ;
  assign n1838 = n1835 | n1837 ;
  assign n1839 = x71 & n962 ;
  assign n1840 = n965 | n1839 ;
  assign n1841 = n1838 | n1840 ;
  assign n1842 = x14 & ~n1841 ;
  assign n1843 = x14 & ~n1839 ;
  assign n1844 = ~n1838 & n1843 ;
  assign n1845 = ( ~n438 & n1842 ) | ( ~n438 & n1844 ) | ( n1842 & n1844 ) ;
  assign n1846 = ~x14 & n1841 ;
  assign n1847 = ~x14 & n1839 ;
  assign n1848 = ( ~x14 & n1838 ) | ( ~x14 & n1847 ) | ( n1838 & n1847 ) ;
  assign n1849 = ( n438 & n1846 ) | ( n438 & n1848 ) | ( n1846 & n1848 ) ;
  assign n1850 = n1845 | n1849 ;
  assign n1851 = ~x18 & x19 ;
  assign n1852 = x18 & ~x19 ;
  assign n1853 = n1851 | n1852 ;
  assign n1854 = ~n1678 & n1853 ;
  assign n1855 = x64 & n1854 ;
  assign n1856 = ~x19 & x20 ;
  assign n1857 = x19 & ~x20 ;
  assign n1858 = n1856 | n1857 ;
  assign n1859 = n1678 & ~n1858 ;
  assign n1860 = x65 & n1859 ;
  assign n1861 = n1855 | n1860 ;
  assign n1862 = n1678 & n1858 ;
  assign n1863 = x20 | n144 ;
  assign n1864 = ( x20 & n1862 ) | ( x20 & n1863 ) | ( n1862 & n1863 ) ;
  assign n1865 = ~x20 & n1864 ;
  assign n1866 = ( ~x20 & n1861 ) | ( ~x20 & n1865 ) | ( n1861 & n1865 ) ;
  assign n1867 = x20 & ~x64 ;
  assign n1868 = ( x20 & ~n1678 ) | ( x20 & n1867 ) | ( ~n1678 & n1867 ) ;
  assign n1869 = n1864 & n1868 ;
  assign n1870 = ( n1861 & n1868 ) | ( n1861 & n1869 ) | ( n1868 & n1869 ) ;
  assign n1871 = n144 & n1862 ;
  assign n1872 = n1868 & ~n1871 ;
  assign n1873 = ~n1861 & n1872 ;
  assign n1874 = ( n1866 & n1870 ) | ( n1866 & n1873 ) | ( n1870 & n1873 ) ;
  assign n1875 = n1864 | n1868 ;
  assign n1876 = n1861 | n1875 ;
  assign n1877 = ~n1868 & n1871 ;
  assign n1878 = ( n1861 & ~n1868 ) | ( n1861 & n1877 ) | ( ~n1868 & n1877 ) ;
  assign n1879 = ( n1866 & n1876 ) | ( n1866 & ~n1878 ) | ( n1876 & ~n1878 ) ;
  assign n1880 = ~n1874 & n1879 ;
  assign n1881 = n241 & n1386 ;
  assign n1882 = x68 & n1383 ;
  assign n1883 = x67 & n1378 ;
  assign n1884 = x66 & ~n1377 ;
  assign n1885 = n1542 & n1884 ;
  assign n1886 = n1883 | n1885 ;
  assign n1887 = n1882 | n1886 ;
  assign n1888 = n1881 | n1887 ;
  assign n1889 = x17 | n1882 ;
  assign n1890 = n1886 | n1889 ;
  assign n1891 = n1881 | n1890 ;
  assign n1892 = ~x17 & n1890 ;
  assign n1893 = ( ~x17 & n1881 ) | ( ~x17 & n1892 ) | ( n1881 & n1892 ) ;
  assign n1894 = ( ~n1888 & n1891 ) | ( ~n1888 & n1893 ) | ( n1891 & n1893 ) ;
  assign n1895 = n1880 & ~n1894 ;
  assign n1896 = ~n1880 & n1894 ;
  assign n1897 = n1895 | n1896 ;
  assign n1898 = ( n1556 & n1679 ) | ( n1556 & n1695 ) | ( n1679 & n1695 ) ;
  assign n1899 = n1897 | n1898 ;
  assign n1900 = n1897 & n1898 ;
  assign n1901 = n1899 & ~n1900 ;
  assign n1902 = n1850 & n1901 ;
  assign n1903 = n1850 | n1901 ;
  assign n1904 = ~n1902 & n1903 ;
  assign n1905 = ~n1698 & n1714 ;
  assign n1906 = n1675 & ~n1905 ;
  assign n1907 = n1698 & n1714 ;
  assign n1908 = n1698 & ~n1907 ;
  assign n1909 = ( n1675 & n1907 ) | ( n1675 & n1908 ) | ( n1907 & n1908 ) ;
  assign n1910 = n1675 | n1907 ;
  assign n1911 = ( ~n1906 & n1909 ) | ( ~n1906 & n1910 ) | ( n1909 & n1910 ) ;
  assign n1912 = n1904 & n1911 ;
  assign n1913 = n1904 | n1911 ;
  assign n1914 = ~n1912 & n1913 ;
  assign n1915 = x74 & n636 ;
  assign n1916 = x73 & n631 ;
  assign n1917 = x72 & ~n630 ;
  assign n1918 = n764 & n1917 ;
  assign n1919 = n1916 | n1918 ;
  assign n1920 = n1915 | n1919 ;
  assign n1921 = n639 | n1915 ;
  assign n1922 = n1919 | n1921 ;
  assign n1923 = ( n710 & n1920 ) | ( n710 & n1922 ) | ( n1920 & n1922 ) ;
  assign n1924 = x11 & n1922 ;
  assign n1925 = x11 & n1915 ;
  assign n1926 = ( x11 & n1919 ) | ( x11 & n1925 ) | ( n1919 & n1925 ) ;
  assign n1927 = ( n710 & n1924 ) | ( n710 & n1926 ) | ( n1924 & n1926 ) ;
  assign n1928 = x11 & ~n1926 ;
  assign n1929 = x11 & ~n1922 ;
  assign n1930 = ( ~n710 & n1928 ) | ( ~n710 & n1929 ) | ( n1928 & n1929 ) ;
  assign n1931 = ( n1923 & ~n1927 ) | ( n1923 & n1930 ) | ( ~n1927 & n1930 ) ;
  assign n1932 = n1914 & n1931 ;
  assign n1933 = n1914 & ~n1932 ;
  assign n1934 = n1735 | n1739 ;
  assign n1935 = ( n1735 & n1741 ) | ( n1735 & n1934 ) | ( n1741 & n1934 ) ;
  assign n1936 = ~n1914 & n1931 ;
  assign n1937 = n1935 & n1936 ;
  assign n1938 = ( n1933 & n1935 ) | ( n1933 & n1937 ) | ( n1935 & n1937 ) ;
  assign n1939 = n1935 | n1936 ;
  assign n1940 = n1933 | n1939 ;
  assign n1941 = ~n1938 & n1940 ;
  assign n1942 = x77 & n389 ;
  assign n1943 = x76 & n384 ;
  assign n1944 = x75 & ~n383 ;
  assign n1945 = n463 & n1944 ;
  assign n1946 = n1943 | n1945 ;
  assign n1947 = n1942 | n1946 ;
  assign n1948 = n392 | n1942 ;
  assign n1949 = n1946 | n1948 ;
  assign n1950 = ( n1059 & n1947 ) | ( n1059 & n1949 ) | ( n1947 & n1949 ) ;
  assign n1951 = x8 & n1949 ;
  assign n1952 = x8 & n1942 ;
  assign n1953 = ( x8 & n1946 ) | ( x8 & n1952 ) | ( n1946 & n1952 ) ;
  assign n1954 = ( n1059 & n1951 ) | ( n1059 & n1953 ) | ( n1951 & n1953 ) ;
  assign n1955 = x8 & ~n1953 ;
  assign n1956 = x8 & ~n1949 ;
  assign n1957 = ( ~n1059 & n1955 ) | ( ~n1059 & n1956 ) | ( n1955 & n1956 ) ;
  assign n1958 = ( n1950 & ~n1954 ) | ( n1950 & n1957 ) | ( ~n1954 & n1957 ) ;
  assign n1959 = n1941 | n1958 ;
  assign n1960 = n1941 & n1958 ;
  assign n1961 = n1959 & ~n1960 ;
  assign n1962 = n1763 | n1764 ;
  assign n1963 = ( n1763 & n1766 ) | ( n1763 & n1962 ) | ( n1766 & n1962 ) ;
  assign n1964 = n1961 & n1963 ;
  assign n1965 = n1961 | n1963 ;
  assign n1966 = ~n1964 & n1965 ;
  assign n1967 = x80 & n212 ;
  assign n1968 = x79 & n207 ;
  assign n1969 = x78 & ~n206 ;
  assign n1970 = n267 & n1969 ;
  assign n1971 = n1968 | n1970 ;
  assign n1972 = n1967 | n1971 ;
  assign n1973 = n215 | n1967 ;
  assign n1974 = n1971 | n1973 ;
  assign n1975 = ( n1499 & n1972 ) | ( n1499 & n1974 ) | ( n1972 & n1974 ) ;
  assign n1976 = x5 & n1974 ;
  assign n1977 = x5 & n1967 ;
  assign n1978 = ( x5 & n1971 ) | ( x5 & n1977 ) | ( n1971 & n1977 ) ;
  assign n1979 = ( n1499 & n1976 ) | ( n1499 & n1978 ) | ( n1976 & n1978 ) ;
  assign n1980 = x5 & ~n1978 ;
  assign n1981 = x5 & ~n1974 ;
  assign n1982 = ( ~n1499 & n1980 ) | ( ~n1499 & n1981 ) | ( n1980 & n1981 ) ;
  assign n1983 = ( n1975 & ~n1979 ) | ( n1975 & n1982 ) | ( ~n1979 & n1982 ) ;
  assign n1984 = n1966 & n1983 ;
  assign n1985 = n1966 & ~n1984 ;
  assign n1986 = ~n1966 & n1983 ;
  assign n1987 = n1985 | n1986 ;
  assign n1988 = n1787 | n1789 ;
  assign n1989 = ( n1787 & n1791 ) | ( n1787 & n1988 ) | ( n1791 & n1988 ) ;
  assign n1990 = n1987 | n1989 ;
  assign n1991 = n1987 & n1989 ;
  assign n1992 = n1990 & ~n1991 ;
  assign n1993 = x82 | x83 ;
  assign n1994 = x82 & x83 ;
  assign n1995 = n1993 & ~n1994 ;
  assign n1996 = n1796 | n1797 ;
  assign n1997 = ( n1796 & n1799 ) | ( n1796 & n1996 ) | ( n1799 & n1996 ) ;
  assign n1998 = n1995 & n1997 ;
  assign n1999 = ( n1796 & n1801 ) | ( n1796 & n1996 ) | ( n1801 & n1996 ) ;
  assign n2000 = n1995 & n1999 ;
  assign n2001 = ( n1492 & n1998 ) | ( n1492 & n2000 ) | ( n1998 & n2000 ) ;
  assign n2002 = ( n1490 & n1998 ) | ( n1490 & n2000 ) | ( n1998 & n2000 ) ;
  assign n2003 = ( n917 & n2001 ) | ( n917 & n2002 ) | ( n2001 & n2002 ) ;
  assign n2004 = n1995 | n1999 ;
  assign n2005 = n1995 | n1997 ;
  assign n2006 = ( n1492 & n2004 ) | ( n1492 & n2005 ) | ( n2004 & n2005 ) ;
  assign n2007 = ( n1490 & n2004 ) | ( n1490 & n2005 ) | ( n2004 & n2005 ) ;
  assign n2008 = ( n917 & n2006 ) | ( n917 & n2007 ) | ( n2006 & n2007 ) ;
  assign n2009 = ~n2003 & n2008 ;
  assign n2010 = x82 & n133 ;
  assign n2011 = x81 & ~n162 ;
  assign n2012 = ( n137 & n2010 ) | ( n137 & n2011 ) | ( n2010 & n2011 ) ;
  assign n2013 = x0 & x83 ;
  assign n2014 = ( ~n137 & n2010 ) | ( ~n137 & n2013 ) | ( n2010 & n2013 ) ;
  assign n2015 = n2012 | n2014 ;
  assign n2016 = n141 | n2015 ;
  assign n2017 = ( n2009 & n2015 ) | ( n2009 & n2016 ) | ( n2015 & n2016 ) ;
  assign n2018 = x2 & n2015 ;
  assign n2019 = ( x2 & n523 ) | ( x2 & n2015 ) | ( n523 & n2015 ) ;
  assign n2020 = ( n2009 & n2018 ) | ( n2009 & n2019 ) | ( n2018 & n2019 ) ;
  assign n2021 = x2 & ~n2019 ;
  assign n2022 = x2 & ~n2015 ;
  assign n2023 = ( ~n2009 & n2021 ) | ( ~n2009 & n2022 ) | ( n2021 & n2022 ) ;
  assign n2024 = ( n2017 & ~n2020 ) | ( n2017 & n2023 ) | ( ~n2020 & n2023 ) ;
  assign n2025 = n1992 & n2024 ;
  assign n2026 = n1992 & ~n2025 ;
  assign n2027 = ~n1992 & n2024 ;
  assign n2028 = n2026 | n2027 ;
  assign n2029 = n1827 | n1829 ;
  assign n2030 = n1828 | n2029 ;
  assign n2031 = ( n1827 & n1831 ) | ( n1827 & n2030 ) | ( n1831 & n2030 ) ;
  assign n2032 = n2028 & n2031 ;
  assign n2033 = n2028 | n2031 ;
  assign n2034 = ~n2032 & n2033 ;
  assign n2035 = x66 & n1859 ;
  assign n2036 = x65 & n1854 ;
  assign n2037 = ~n1678 & n1858 ;
  assign n2038 = x64 & ~n1853 ;
  assign n2039 = n2037 & n2038 ;
  assign n2040 = n2036 | n2039 ;
  assign n2041 = n2035 | n2040 ;
  assign n2042 = n159 & n1862 ;
  assign n2043 = n2041 | n2042 ;
  assign n2044 = x20 | n1862 ;
  assign n2045 = ( x20 & n159 ) | ( x20 & n2044 ) | ( n159 & n2044 ) ;
  assign n2046 = n2041 | n2045 ;
  assign n2047 = ~x20 & n2045 ;
  assign n2048 = ( ~x20 & n2041 ) | ( ~x20 & n2047 ) | ( n2041 & n2047 ) ;
  assign n2049 = ( ~n2043 & n2046 ) | ( ~n2043 & n2048 ) | ( n2046 & n2048 ) ;
  assign n2050 = n1874 | n2049 ;
  assign n2051 = n1874 & n2049 ;
  assign n2052 = n2050 & ~n2051 ;
  assign n2053 = n293 & n1386 ;
  assign n2054 = x69 & n1383 ;
  assign n2055 = x68 & n1378 ;
  assign n2056 = x67 & ~n1377 ;
  assign n2057 = n1542 & n2056 ;
  assign n2058 = n2055 | n2057 ;
  assign n2059 = n2054 | n2058 ;
  assign n2060 = n2053 | n2059 ;
  assign n2061 = x17 | n2054 ;
  assign n2062 = n2058 | n2061 ;
  assign n2063 = n2053 | n2062 ;
  assign n2064 = ~x17 & n2062 ;
  assign n2065 = ( ~x17 & n2053 ) | ( ~x17 & n2064 ) | ( n2053 & n2064 ) ;
  assign n2066 = ( ~n2060 & n2063 ) | ( ~n2060 & n2065 ) | ( n2063 & n2065 ) ;
  assign n2067 = n2052 | n2066 ;
  assign n2068 = n2052 & n2066 ;
  assign n2069 = n2067 & ~n2068 ;
  assign n2070 = ( n1880 & n1894 ) | ( n1880 & n1898 ) | ( n1894 & n1898 ) ;
  assign n2071 = n2068 | n2070 ;
  assign n2072 = ( n2068 & n2069 ) | ( n2068 & n2071 ) | ( n2069 & n2071 ) ;
  assign n2073 = n2067 & ~n2072 ;
  assign n2074 = x72 & n962 ;
  assign n2075 = x71 & n957 ;
  assign n2076 = x70 & ~n956 ;
  assign n2077 = n1105 & n2076 ;
  assign n2078 = n2075 | n2077 ;
  assign n2079 = n2074 | n2078 ;
  assign n2080 = ( n513 & n965 ) | ( n513 & n2079 ) | ( n965 & n2079 ) ;
  assign n2081 = ( x14 & n965 ) | ( x14 & ~n2074 ) | ( n965 & ~n2074 ) ;
  assign n2082 = x14 & n965 ;
  assign n2083 = ( ~n2078 & n2081 ) | ( ~n2078 & n2082 ) | ( n2081 & n2082 ) ;
  assign n2084 = ( x14 & n513 ) | ( x14 & n2083 ) | ( n513 & n2083 ) ;
  assign n2085 = ~n2080 & n2084 ;
  assign n2086 = n2079 | n2083 ;
  assign n2087 = x14 | n2079 ;
  assign n2088 = ( n513 & n2086 ) | ( n513 & n2087 ) | ( n2086 & n2087 ) ;
  assign n2089 = ( ~x14 & n2085 ) | ( ~x14 & n2088 ) | ( n2085 & n2088 ) ;
  assign n2090 = n2070 & n2089 ;
  assign n2091 = ~n2069 & n2090 ;
  assign n2092 = ( n2073 & n2089 ) | ( n2073 & n2091 ) | ( n2089 & n2091 ) ;
  assign n2093 = n2070 | n2089 ;
  assign n2094 = ( ~n2069 & n2089 ) | ( ~n2069 & n2093 ) | ( n2089 & n2093 ) ;
  assign n2095 = n2073 | n2094 ;
  assign n2096 = ~n2092 & n2095 ;
  assign n2097 = n1902 | n1904 ;
  assign n2098 = ( n1902 & n1911 ) | ( n1902 & n2097 ) | ( n1911 & n2097 ) ;
  assign n2099 = n2096 & n2098 ;
  assign n2100 = n2096 | n2098 ;
  assign n2101 = ~n2099 & n2100 ;
  assign n2102 = x75 & n636 ;
  assign n2103 = x74 & n631 ;
  assign n2104 = x73 & ~n630 ;
  assign n2105 = n764 & n2104 ;
  assign n2106 = n2103 | n2105 ;
  assign n2107 = n2102 | n2106 ;
  assign n2108 = n639 | n2102 ;
  assign n2109 = n2106 | n2108 ;
  assign n2110 = ( n746 & n2107 ) | ( n746 & n2109 ) | ( n2107 & n2109 ) ;
  assign n2111 = x11 & n2109 ;
  assign n2112 = x11 & n2102 ;
  assign n2113 = ( x11 & n2106 ) | ( x11 & n2112 ) | ( n2106 & n2112 ) ;
  assign n2114 = ( n746 & n2111 ) | ( n746 & n2113 ) | ( n2111 & n2113 ) ;
  assign n2115 = x11 & ~n2113 ;
  assign n2116 = x11 & ~n2109 ;
  assign n2117 = ( ~n746 & n2115 ) | ( ~n746 & n2116 ) | ( n2115 & n2116 ) ;
  assign n2118 = ( n2110 & ~n2114 ) | ( n2110 & n2117 ) | ( ~n2114 & n2117 ) ;
  assign n2119 = n2101 | n2118 ;
  assign n2120 = n2101 & n2118 ;
  assign n2121 = n2119 & ~n2120 ;
  assign n2122 = n1932 | n1938 ;
  assign n2123 = n2121 & n2122 ;
  assign n2124 = n2121 | n2122 ;
  assign n2125 = ~n2123 & n2124 ;
  assign n2126 = x78 & n389 ;
  assign n2127 = x77 & n384 ;
  assign n2128 = x76 & ~n383 ;
  assign n2129 = n463 & n2128 ;
  assign n2130 = n2127 | n2129 ;
  assign n2131 = n2126 | n2130 ;
  assign n2132 = n392 | n2126 ;
  assign n2133 = n2130 | n2132 ;
  assign n2134 = ( n1192 & n2131 ) | ( n1192 & n2133 ) | ( n2131 & n2133 ) ;
  assign n2135 = x8 & n2133 ;
  assign n2136 = x8 & n2126 ;
  assign n2137 = ( x8 & n2130 ) | ( x8 & n2136 ) | ( n2130 & n2136 ) ;
  assign n2138 = ( n1192 & n2135 ) | ( n1192 & n2137 ) | ( n2135 & n2137 ) ;
  assign n2139 = x8 & ~n2137 ;
  assign n2140 = x8 & ~n2133 ;
  assign n2141 = ( ~n1192 & n2139 ) | ( ~n1192 & n2140 ) | ( n2139 & n2140 ) ;
  assign n2142 = ( n2134 & ~n2138 ) | ( n2134 & n2141 ) | ( ~n2138 & n2141 ) ;
  assign n2143 = n2125 & n2142 ;
  assign n2144 = n2125 & ~n2143 ;
  assign n2145 = ~n2125 & n2142 ;
  assign n2146 = n2144 | n2145 ;
  assign n2147 = n1960 | n1964 ;
  assign n2148 = n2146 & n2147 ;
  assign n2149 = n2146 | n2147 ;
  assign n2150 = ~n2148 & n2149 ;
  assign n2151 = x81 & n212 ;
  assign n2152 = x80 & n207 ;
  assign n2153 = x79 & ~n206 ;
  assign n2154 = n267 & n2153 ;
  assign n2155 = n2152 | n2154 ;
  assign n2156 = n2151 | n2155 ;
  assign n2157 = n215 | n2151 ;
  assign n2158 = n2155 | n2157 ;
  assign n2159 = ( n1651 & n2156 ) | ( n1651 & n2158 ) | ( n2156 & n2158 ) ;
  assign n2160 = x5 & n2158 ;
  assign n2161 = x5 & n2151 ;
  assign n2162 = ( x5 & n2155 ) | ( x5 & n2161 ) | ( n2155 & n2161 ) ;
  assign n2163 = ( n1651 & n2160 ) | ( n1651 & n2162 ) | ( n2160 & n2162 ) ;
  assign n2164 = x5 & ~n2162 ;
  assign n2165 = x5 & ~n2158 ;
  assign n2166 = ( ~n1651 & n2164 ) | ( ~n1651 & n2165 ) | ( n2164 & n2165 ) ;
  assign n2167 = ( n2159 & ~n2163 ) | ( n2159 & n2166 ) | ( ~n2163 & n2166 ) ;
  assign n2168 = n2150 & n2167 ;
  assign n2169 = n2150 & ~n2168 ;
  assign n2170 = ~n2150 & n2167 ;
  assign n2171 = n2169 | n2170 ;
  assign n2172 = n1984 | n1991 ;
  assign n2173 = ~n2171 & n2172 ;
  assign n2174 = n2171 & ~n2172 ;
  assign n2175 = n2173 | n2174 ;
  assign n2176 = x83 | x84 ;
  assign n2177 = x83 & x84 ;
  assign n2178 = n2176 & ~n2177 ;
  assign n2179 = n1994 | n1995 ;
  assign n2180 = n2178 & n2179 ;
  assign n2181 = n1994 & n2178 ;
  assign n2182 = ( n1999 & n2180 ) | ( n1999 & n2181 ) | ( n2180 & n2181 ) ;
  assign n2183 = ( n1997 & n2180 ) | ( n1997 & n2181 ) | ( n2180 & n2181 ) ;
  assign n2184 = ( n1492 & n2182 ) | ( n1492 & n2183 ) | ( n2182 & n2183 ) ;
  assign n2185 = ( n1490 & n2182 ) | ( n1490 & n2183 ) | ( n2182 & n2183 ) ;
  assign n2186 = ( n917 & n2184 ) | ( n917 & n2185 ) | ( n2184 & n2185 ) ;
  assign n2187 = n2178 | n2179 ;
  assign n2188 = n1994 | n2178 ;
  assign n2189 = ( n1999 & n2187 ) | ( n1999 & n2188 ) | ( n2187 & n2188 ) ;
  assign n2190 = ( n1997 & n2187 ) | ( n1997 & n2188 ) | ( n2187 & n2188 ) ;
  assign n2191 = ( n1492 & n2189 ) | ( n1492 & n2190 ) | ( n2189 & n2190 ) ;
  assign n2192 = ( n1490 & n2189 ) | ( n1490 & n2190 ) | ( n2189 & n2190 ) ;
  assign n2193 = ( n917 & n2191 ) | ( n917 & n2192 ) | ( n2191 & n2192 ) ;
  assign n2194 = ~n2186 & n2193 ;
  assign n2195 = x83 & n133 ;
  assign n2196 = x82 & ~n162 ;
  assign n2197 = ( n137 & n2195 ) | ( n137 & n2196 ) | ( n2195 & n2196 ) ;
  assign n2198 = x0 & x84 ;
  assign n2199 = ( ~n137 & n2195 ) | ( ~n137 & n2198 ) | ( n2195 & n2198 ) ;
  assign n2200 = n2197 | n2199 ;
  assign n2201 = n141 | n2200 ;
  assign n2202 = ( n2194 & n2200 ) | ( n2194 & n2201 ) | ( n2200 & n2201 ) ;
  assign n2203 = x2 & n2200 ;
  assign n2204 = ( x2 & n523 ) | ( x2 & n2200 ) | ( n523 & n2200 ) ;
  assign n2205 = ( n2194 & n2203 ) | ( n2194 & n2204 ) | ( n2203 & n2204 ) ;
  assign n2206 = x2 & ~n2204 ;
  assign n2207 = x2 & ~n2200 ;
  assign n2208 = ( ~n2194 & n2206 ) | ( ~n2194 & n2207 ) | ( n2206 & n2207 ) ;
  assign n2209 = ( n2202 & ~n2205 ) | ( n2202 & n2208 ) | ( ~n2205 & n2208 ) ;
  assign n2210 = n2175 & n2209 ;
  assign n2211 = n2175 | n2209 ;
  assign n2212 = ~n2210 & n2211 ;
  assign n2213 = n2025 | n2027 ;
  assign n2214 = n2026 | n2213 ;
  assign n2215 = ( n2025 & n2031 ) | ( n2025 & n2214 ) | ( n2031 & n2214 ) ;
  assign n2216 = n2212 & n2215 ;
  assign n2217 = n2212 | n2215 ;
  assign n2218 = ~n2216 & n2217 ;
  assign n2219 = x20 & ~x21 ;
  assign n2220 = ~x20 & x21 ;
  assign n2221 = n2219 | n2220 ;
  assign n2222 = x64 & n2221 ;
  assign n2223 = ~n1874 & n2222 ;
  assign n2224 = ( ~n2049 & n2222 ) | ( ~n2049 & n2223 ) | ( n2222 & n2223 ) ;
  assign n2225 = n1874 & ~n2222 ;
  assign n2226 = n2049 & n2225 ;
  assign n2227 = n2224 | n2226 ;
  assign n2228 = x67 & n1859 ;
  assign n2229 = x66 & n1854 ;
  assign n2230 = x65 & ~n1853 ;
  assign n2231 = n2037 & n2230 ;
  assign n2232 = n2229 | n2231 ;
  assign n2233 = n2228 | n2232 ;
  assign n2234 = n186 & n1862 ;
  assign n2235 = n2233 | n2234 ;
  assign n2236 = x20 & ~n2235 ;
  assign n2237 = ~x20 & n2235 ;
  assign n2238 = n2236 | n2237 ;
  assign n2239 = n2227 & n2238 ;
  assign n2240 = n2227 | n2238 ;
  assign n2241 = ~n2239 & n2240 ;
  assign n2242 = x69 & n1378 ;
  assign n2243 = x68 & ~n1377 ;
  assign n2244 = n1542 & n2243 ;
  assign n2245 = n2242 | n2244 ;
  assign n2246 = x70 & n1383 ;
  assign n2247 = n1386 | n2246 ;
  assign n2248 = n2245 | n2247 ;
  assign n2249 = x17 & ~n2248 ;
  assign n2250 = x17 & ~n2246 ;
  assign n2251 = ~n2245 & n2250 ;
  assign n2252 = ( ~n340 & n2249 ) | ( ~n340 & n2251 ) | ( n2249 & n2251 ) ;
  assign n2253 = ~x17 & n2248 ;
  assign n2254 = ~x17 & n2246 ;
  assign n2255 = ( ~x17 & n2245 ) | ( ~x17 & n2254 ) | ( n2245 & n2254 ) ;
  assign n2256 = ( n340 & n2253 ) | ( n340 & n2255 ) | ( n2253 & n2255 ) ;
  assign n2257 = n2252 | n2256 ;
  assign n2258 = ( n2072 & ~n2241 ) | ( n2072 & n2257 ) | ( ~n2241 & n2257 ) ;
  assign n2259 = ( ~n2072 & n2241 ) | ( ~n2072 & n2258 ) | ( n2241 & n2258 ) ;
  assign n2260 = x73 & n962 ;
  assign n2261 = x72 & n957 ;
  assign n2262 = x71 & ~n956 ;
  assign n2263 = n1105 & n2262 ;
  assign n2264 = n2261 | n2263 ;
  assign n2265 = n2260 | n2264 ;
  assign n2266 = n965 | n2260 ;
  assign n2267 = n2264 | n2266 ;
  assign n2268 = ( ~n610 & n2265 ) | ( ~n610 & n2267 ) | ( n2265 & n2267 ) ;
  assign n2269 = n2265 & n2267 ;
  assign n2270 = ( n598 & n2268 ) | ( n598 & n2269 ) | ( n2268 & n2269 ) ;
  assign n2271 = x14 & n2270 ;
  assign n2272 = x14 | n2270 ;
  assign n2273 = ~n2271 & n2272 ;
  assign n2274 = ~n2257 & n2273 ;
  assign n2275 = ~n2241 & n2273 ;
  assign n2276 = n2257 & n2273 ;
  assign n2277 = ( n2072 & n2275 ) | ( n2072 & n2276 ) | ( n2275 & n2276 ) ;
  assign n2278 = ( n2259 & n2274 ) | ( n2259 & n2277 ) | ( n2274 & n2277 ) ;
  assign n2279 = n2257 & ~n2273 ;
  assign n2280 = n2241 & ~n2273 ;
  assign n2281 = n2257 | n2273 ;
  assign n2282 = ( n2072 & ~n2280 ) | ( n2072 & n2281 ) | ( ~n2280 & n2281 ) ;
  assign n2283 = ( n2259 & ~n2279 ) | ( n2259 & n2282 ) | ( ~n2279 & n2282 ) ;
  assign n2284 = ~n2278 & n2283 ;
  assign n2285 = n2092 | n2096 ;
  assign n2286 = ( n2092 & n2098 ) | ( n2092 & n2285 ) | ( n2098 & n2285 ) ;
  assign n2287 = n2284 & n2286 ;
  assign n2288 = n2284 | n2286 ;
  assign n2289 = ~n2287 & n2288 ;
  assign n2290 = x76 & n636 ;
  assign n2291 = x75 & n631 ;
  assign n2292 = x74 & ~n630 ;
  assign n2293 = n764 & n2292 ;
  assign n2294 = n2291 | n2293 ;
  assign n2295 = n2290 | n2294 ;
  assign n2296 = n639 | n2290 ;
  assign n2297 = n2294 | n2296 ;
  assign n2298 = ( n923 & n2295 ) | ( n923 & n2297 ) | ( n2295 & n2297 ) ;
  assign n2299 = x11 & n2297 ;
  assign n2300 = x11 & n2290 ;
  assign n2301 = ( x11 & n2294 ) | ( x11 & n2300 ) | ( n2294 & n2300 ) ;
  assign n2302 = ( n923 & n2299 ) | ( n923 & n2301 ) | ( n2299 & n2301 ) ;
  assign n2303 = x11 & ~n2301 ;
  assign n2304 = x11 & ~n2297 ;
  assign n2305 = ( ~n923 & n2303 ) | ( ~n923 & n2304 ) | ( n2303 & n2304 ) ;
  assign n2306 = ( n2298 & ~n2302 ) | ( n2298 & n2305 ) | ( ~n2302 & n2305 ) ;
  assign n2307 = n2289 | n2306 ;
  assign n2308 = n2289 & n2306 ;
  assign n2309 = n2307 & ~n2308 ;
  assign n2310 = n2120 | n2121 ;
  assign n2311 = ( n2120 & n2122 ) | ( n2120 & n2310 ) | ( n2122 & n2310 ) ;
  assign n2312 = n2309 & n2311 ;
  assign n2313 = n2309 | n2311 ;
  assign n2314 = ~n2312 & n2313 ;
  assign n2315 = x79 & n389 ;
  assign n2316 = x78 & n384 ;
  assign n2317 = x77 & ~n383 ;
  assign n2318 = n463 & n2317 ;
  assign n2319 = n2316 | n2318 ;
  assign n2320 = n2315 | n2319 ;
  assign n2321 = n392 | n2315 ;
  assign n2322 = n2319 | n2321 ;
  assign n2323 = ( n1332 & n2320 ) | ( n1332 & n2322 ) | ( n2320 & n2322 ) ;
  assign n2324 = x8 & n2322 ;
  assign n2325 = x8 & n2315 ;
  assign n2326 = ( x8 & n2319 ) | ( x8 & n2325 ) | ( n2319 & n2325 ) ;
  assign n2327 = ( n1332 & n2324 ) | ( n1332 & n2326 ) | ( n2324 & n2326 ) ;
  assign n2328 = x8 & ~n2326 ;
  assign n2329 = x8 & ~n2322 ;
  assign n2330 = ( ~n1332 & n2328 ) | ( ~n1332 & n2329 ) | ( n2328 & n2329 ) ;
  assign n2331 = ( n2323 & ~n2327 ) | ( n2323 & n2330 ) | ( ~n2327 & n2330 ) ;
  assign n2332 = n2314 & n2331 ;
  assign n2333 = n2314 | n2331 ;
  assign n2334 = ~n2332 & n2333 ;
  assign n2335 = n2143 & n2334 ;
  assign n2336 = ( n2148 & n2334 ) | ( n2148 & n2335 ) | ( n2334 & n2335 ) ;
  assign n2337 = n2143 | n2334 ;
  assign n2338 = n2148 | n2337 ;
  assign n2339 = ~n2336 & n2338 ;
  assign n2340 = x82 & n212 ;
  assign n2341 = x81 & n207 ;
  assign n2342 = x80 & ~n206 ;
  assign n2343 = n267 & n2342 ;
  assign n2344 = n2341 | n2343 ;
  assign n2345 = n2340 | n2344 ;
  assign n2346 = n215 | n2340 ;
  assign n2347 = n2344 | n2346 ;
  assign n2348 = ( n1811 & n2345 ) | ( n1811 & n2347 ) | ( n2345 & n2347 ) ;
  assign n2349 = x5 & n2347 ;
  assign n2350 = x5 & n2340 ;
  assign n2351 = ( x5 & n2344 ) | ( x5 & n2350 ) | ( n2344 & n2350 ) ;
  assign n2352 = ( n1811 & n2349 ) | ( n1811 & n2351 ) | ( n2349 & n2351 ) ;
  assign n2353 = x5 & ~n2351 ;
  assign n2354 = x5 & ~n2347 ;
  assign n2355 = ( ~n1811 & n2353 ) | ( ~n1811 & n2354 ) | ( n2353 & n2354 ) ;
  assign n2356 = ( n2348 & ~n2352 ) | ( n2348 & n2355 ) | ( ~n2352 & n2355 ) ;
  assign n2357 = n2339 & n2356 ;
  assign n2358 = n2339 & ~n2357 ;
  assign n2359 = ~n2339 & n2356 ;
  assign n2360 = n2358 | n2359 ;
  assign n2361 = n2168 | n2172 ;
  assign n2362 = ( n2168 & n2171 ) | ( n2168 & n2361 ) | ( n2171 & n2361 ) ;
  assign n2363 = n2360 | n2362 ;
  assign n2364 = n2360 & n2362 ;
  assign n2365 = n2363 & ~n2364 ;
  assign n2366 = x84 | x85 ;
  assign n2367 = x84 & x85 ;
  assign n2368 = n2366 & ~n2367 ;
  assign n2369 = n2177 & n2368 ;
  assign n2370 = ( n2183 & n2368 ) | ( n2183 & n2369 ) | ( n2368 & n2369 ) ;
  assign n2371 = ( n2182 & n2368 ) | ( n2182 & n2369 ) | ( n2368 & n2369 ) ;
  assign n2372 = ( n1492 & n2370 ) | ( n1492 & n2371 ) | ( n2370 & n2371 ) ;
  assign n2373 = ( n1490 & n2370 ) | ( n1490 & n2371 ) | ( n2370 & n2371 ) ;
  assign n2374 = ( n917 & n2372 ) | ( n917 & n2373 ) | ( n2372 & n2373 ) ;
  assign n2375 = n2177 | n2368 ;
  assign n2376 = n2183 | n2375 ;
  assign n2377 = n2182 | n2375 ;
  assign n2378 = ( n1492 & n2376 ) | ( n1492 & n2377 ) | ( n2376 & n2377 ) ;
  assign n2379 = ( n1490 & n2376 ) | ( n1490 & n2377 ) | ( n2376 & n2377 ) ;
  assign n2380 = ( n917 & n2378 ) | ( n917 & n2379 ) | ( n2378 & n2379 ) ;
  assign n2381 = ~n2374 & n2380 ;
  assign n2382 = x84 & n133 ;
  assign n2383 = x83 & ~n162 ;
  assign n2384 = ( n137 & n2382 ) | ( n137 & n2383 ) | ( n2382 & n2383 ) ;
  assign n2385 = x0 & x85 ;
  assign n2386 = ( ~n137 & n2382 ) | ( ~n137 & n2385 ) | ( n2382 & n2385 ) ;
  assign n2387 = n2384 | n2386 ;
  assign n2388 = n141 | n2387 ;
  assign n2389 = ( n2381 & n2387 ) | ( n2381 & n2388 ) | ( n2387 & n2388 ) ;
  assign n2390 = x2 & n2387 ;
  assign n2391 = ( x2 & n523 ) | ( x2 & n2387 ) | ( n523 & n2387 ) ;
  assign n2392 = ( n2381 & n2390 ) | ( n2381 & n2391 ) | ( n2390 & n2391 ) ;
  assign n2393 = x2 & ~n2391 ;
  assign n2394 = x2 & ~n2387 ;
  assign n2395 = ( ~n2381 & n2393 ) | ( ~n2381 & n2394 ) | ( n2393 & n2394 ) ;
  assign n2396 = ( n2389 & ~n2392 ) | ( n2389 & n2395 ) | ( ~n2392 & n2395 ) ;
  assign n2397 = n2365 & n2396 ;
  assign n2398 = n2365 & ~n2397 ;
  assign n2399 = ~n2365 & n2396 ;
  assign n2400 = n2398 | n2399 ;
  assign n2401 = n2210 | n2216 ;
  assign n2402 = n2400 & n2401 ;
  assign n2403 = n2400 | n2401 ;
  assign n2404 = ~n2402 & n2403 ;
  assign n2405 = x70 & n1378 ;
  assign n2406 = x69 & ~n1377 ;
  assign n2407 = n1542 & n2406 ;
  assign n2408 = n2405 | n2407 ;
  assign n2409 = x71 & n1383 ;
  assign n2410 = n1386 | n2409 ;
  assign n2411 = n2408 | n2410 ;
  assign n2412 = x17 & ~n2411 ;
  assign n2413 = x17 & ~n2409 ;
  assign n2414 = ~n2408 & n2413 ;
  assign n2415 = ( ~n438 & n2412 ) | ( ~n438 & n2414 ) | ( n2412 & n2414 ) ;
  assign n2416 = ~x17 & n2411 ;
  assign n2417 = ~x17 & n2409 ;
  assign n2418 = ( ~x17 & n2408 ) | ( ~x17 & n2417 ) | ( n2408 & n2417 ) ;
  assign n2419 = ( n438 & n2416 ) | ( n438 & n2418 ) | ( n2416 & n2418 ) ;
  assign n2420 = n2415 | n2419 ;
  assign n2421 = ~x21 & x22 ;
  assign n2422 = x21 & ~x22 ;
  assign n2423 = n2421 | n2422 ;
  assign n2424 = ~n2221 & n2423 ;
  assign n2425 = x64 & n2424 ;
  assign n2426 = ~x22 & x23 ;
  assign n2427 = x22 & ~x23 ;
  assign n2428 = n2426 | n2427 ;
  assign n2429 = n2221 & ~n2428 ;
  assign n2430 = x65 & n2429 ;
  assign n2431 = n2425 | n2430 ;
  assign n2432 = n2221 & n2428 ;
  assign n2433 = x23 | n144 ;
  assign n2434 = ( x23 & n2432 ) | ( x23 & n2433 ) | ( n2432 & n2433 ) ;
  assign n2435 = ~x23 & n2434 ;
  assign n2436 = ( ~x23 & n2431 ) | ( ~x23 & n2435 ) | ( n2431 & n2435 ) ;
  assign n2437 = x23 & ~x64 ;
  assign n2438 = ( x23 & ~n2221 ) | ( x23 & n2437 ) | ( ~n2221 & n2437 ) ;
  assign n2439 = n2434 & n2438 ;
  assign n2440 = ( n2431 & n2438 ) | ( n2431 & n2439 ) | ( n2438 & n2439 ) ;
  assign n2441 = n144 & n2432 ;
  assign n2442 = n2438 & ~n2441 ;
  assign n2443 = ~n2431 & n2442 ;
  assign n2444 = ( n2436 & n2440 ) | ( n2436 & n2443 ) | ( n2440 & n2443 ) ;
  assign n2445 = n2434 | n2438 ;
  assign n2446 = n2431 | n2445 ;
  assign n2447 = ~n2438 & n2441 ;
  assign n2448 = ( n2431 & ~n2438 ) | ( n2431 & n2447 ) | ( ~n2438 & n2447 ) ;
  assign n2449 = ( n2436 & n2446 ) | ( n2436 & ~n2448 ) | ( n2446 & ~n2448 ) ;
  assign n2450 = ~n2444 & n2449 ;
  assign n2451 = n241 & n1862 ;
  assign n2452 = x68 & n1859 ;
  assign n2453 = x67 & n1854 ;
  assign n2454 = x66 & ~n1853 ;
  assign n2455 = n2037 & n2454 ;
  assign n2456 = n2453 | n2455 ;
  assign n2457 = n2452 | n2456 ;
  assign n2458 = n2451 | n2457 ;
  assign n2459 = x20 | n2452 ;
  assign n2460 = n2456 | n2459 ;
  assign n2461 = n2451 | n2460 ;
  assign n2462 = ~x20 & n2460 ;
  assign n2463 = ( ~x20 & n2451 ) | ( ~x20 & n2462 ) | ( n2451 & n2462 ) ;
  assign n2464 = ( ~n2458 & n2461 ) | ( ~n2458 & n2463 ) | ( n2461 & n2463 ) ;
  assign n2465 = n2450 & ~n2464 ;
  assign n2466 = ~n2450 & n2464 ;
  assign n2467 = n2465 | n2466 ;
  assign n2468 = ( n2051 & n2222 ) | ( n2051 & n2238 ) | ( n2222 & n2238 ) ;
  assign n2469 = n2467 | n2468 ;
  assign n2470 = n2467 & n2468 ;
  assign n2471 = n2469 & ~n2470 ;
  assign n2472 = n2420 & n2471 ;
  assign n2473 = n2420 | n2471 ;
  assign n2474 = ~n2472 & n2473 ;
  assign n2475 = n2241 & n2257 ;
  assign n2476 = n2241 & ~n2475 ;
  assign n2477 = ~n2241 & n2257 ;
  assign n2478 = n2072 & ~n2477 ;
  assign n2479 = ~n2476 & n2478 ;
  assign n2480 = ( n2072 & n2475 ) | ( n2072 & ~n2479 ) | ( n2475 & ~n2479 ) ;
  assign n2481 = n2474 & n2480 ;
  assign n2482 = n2474 | n2480 ;
  assign n2483 = ~n2481 & n2482 ;
  assign n2484 = x74 & n962 ;
  assign n2485 = x73 & n957 ;
  assign n2486 = x72 & ~n956 ;
  assign n2487 = n1105 & n2486 ;
  assign n2488 = n2485 | n2487 ;
  assign n2489 = n2484 | n2488 ;
  assign n2490 = n965 | n2484 ;
  assign n2491 = n2488 | n2490 ;
  assign n2492 = ( n710 & n2489 ) | ( n710 & n2491 ) | ( n2489 & n2491 ) ;
  assign n2493 = x14 & n2491 ;
  assign n2494 = x14 & n2484 ;
  assign n2495 = ( x14 & n2488 ) | ( x14 & n2494 ) | ( n2488 & n2494 ) ;
  assign n2496 = ( n710 & n2493 ) | ( n710 & n2495 ) | ( n2493 & n2495 ) ;
  assign n2497 = x14 & ~n2495 ;
  assign n2498 = x14 & ~n2491 ;
  assign n2499 = ( ~n710 & n2497 ) | ( ~n710 & n2498 ) | ( n2497 & n2498 ) ;
  assign n2500 = ( n2492 & ~n2496 ) | ( n2492 & n2499 ) | ( ~n2496 & n2499 ) ;
  assign n2501 = n2483 & n2500 ;
  assign n2502 = n2483 & ~n2501 ;
  assign n2503 = n2278 | n2284 ;
  assign n2504 = ( n2278 & n2286 ) | ( n2278 & n2503 ) | ( n2286 & n2503 ) ;
  assign n2505 = ~n2483 & n2500 ;
  assign n2506 = n2504 & n2505 ;
  assign n2507 = ( n2502 & n2504 ) | ( n2502 & n2506 ) | ( n2504 & n2506 ) ;
  assign n2508 = n2504 | n2505 ;
  assign n2509 = n2502 | n2508 ;
  assign n2510 = ~n2507 & n2509 ;
  assign n2511 = x77 & n636 ;
  assign n2512 = x76 & n631 ;
  assign n2513 = x75 & ~n630 ;
  assign n2514 = n764 & n2513 ;
  assign n2515 = n2512 | n2514 ;
  assign n2516 = n2511 | n2515 ;
  assign n2517 = n639 | n2511 ;
  assign n2518 = n2515 | n2517 ;
  assign n2519 = ( n1059 & n2516 ) | ( n1059 & n2518 ) | ( n2516 & n2518 ) ;
  assign n2520 = x11 & n2518 ;
  assign n2521 = x11 & n2511 ;
  assign n2522 = ( x11 & n2515 ) | ( x11 & n2521 ) | ( n2515 & n2521 ) ;
  assign n2523 = ( n1059 & n2520 ) | ( n1059 & n2522 ) | ( n2520 & n2522 ) ;
  assign n2524 = x11 & ~n2522 ;
  assign n2525 = x11 & ~n2518 ;
  assign n2526 = ( ~n1059 & n2524 ) | ( ~n1059 & n2525 ) | ( n2524 & n2525 ) ;
  assign n2527 = ( n2519 & ~n2523 ) | ( n2519 & n2526 ) | ( ~n2523 & n2526 ) ;
  assign n2528 = n2510 | n2527 ;
  assign n2529 = n2510 & n2527 ;
  assign n2530 = n2528 & ~n2529 ;
  assign n2531 = n2308 | n2309 ;
  assign n2532 = ( n2308 & n2311 ) | ( n2308 & n2531 ) | ( n2311 & n2531 ) ;
  assign n2533 = n2530 & n2532 ;
  assign n2534 = n2530 | n2532 ;
  assign n2535 = ~n2533 & n2534 ;
  assign n2536 = x80 & n389 ;
  assign n2537 = x79 & n384 ;
  assign n2538 = x78 & ~n383 ;
  assign n2539 = n463 & n2538 ;
  assign n2540 = n2537 | n2539 ;
  assign n2541 = n2536 | n2540 ;
  assign n2542 = n392 | n2536 ;
  assign n2543 = n2540 | n2542 ;
  assign n2544 = ( n1499 & n2541 ) | ( n1499 & n2543 ) | ( n2541 & n2543 ) ;
  assign n2545 = x8 & n2543 ;
  assign n2546 = x8 & n2536 ;
  assign n2547 = ( x8 & n2540 ) | ( x8 & n2546 ) | ( n2540 & n2546 ) ;
  assign n2548 = ( n1499 & n2545 ) | ( n1499 & n2547 ) | ( n2545 & n2547 ) ;
  assign n2549 = x8 & ~n2547 ;
  assign n2550 = x8 & ~n2543 ;
  assign n2551 = ( ~n1499 & n2549 ) | ( ~n1499 & n2550 ) | ( n2549 & n2550 ) ;
  assign n2552 = ( n2544 & ~n2548 ) | ( n2544 & n2551 ) | ( ~n2548 & n2551 ) ;
  assign n2553 = n2535 & n2552 ;
  assign n2554 = n2535 | n2552 ;
  assign n2555 = ~n2553 & n2554 ;
  assign n2556 = n2332 & n2555 ;
  assign n2557 = ( n2336 & n2555 ) | ( n2336 & n2556 ) | ( n2555 & n2556 ) ;
  assign n2558 = n2332 | n2555 ;
  assign n2559 = n2336 | n2558 ;
  assign n2560 = ~n2557 & n2559 ;
  assign n2561 = x83 & n212 ;
  assign n2562 = x82 & n207 ;
  assign n2563 = x81 & ~n206 ;
  assign n2564 = n267 & n2563 ;
  assign n2565 = n2562 | n2564 ;
  assign n2566 = n2561 | n2565 ;
  assign n2567 = n215 | n2561 ;
  assign n2568 = n2565 | n2567 ;
  assign n2569 = ( n2009 & n2566 ) | ( n2009 & n2568 ) | ( n2566 & n2568 ) ;
  assign n2570 = x5 & n2568 ;
  assign n2571 = x5 & n2561 ;
  assign n2572 = ( x5 & n2565 ) | ( x5 & n2571 ) | ( n2565 & n2571 ) ;
  assign n2573 = ( n2009 & n2570 ) | ( n2009 & n2572 ) | ( n2570 & n2572 ) ;
  assign n2574 = x5 & ~n2572 ;
  assign n2575 = x5 & ~n2568 ;
  assign n2576 = ( ~n2009 & n2574 ) | ( ~n2009 & n2575 ) | ( n2574 & n2575 ) ;
  assign n2577 = ( n2569 & ~n2573 ) | ( n2569 & n2576 ) | ( ~n2573 & n2576 ) ;
  assign n2578 = n2560 & n2577 ;
  assign n2579 = n2560 & ~n2578 ;
  assign n2580 = ~n2560 & n2577 ;
  assign n2581 = n2579 | n2580 ;
  assign n2582 = n2357 | n2364 ;
  assign n2583 = n2581 | n2582 ;
  assign n2584 = n2581 & n2582 ;
  assign n2585 = n2583 & ~n2584 ;
  assign n2586 = x85 | x86 ;
  assign n2587 = x85 & x86 ;
  assign n2588 = n2586 & ~n2587 ;
  assign n2589 = n2177 | n2367 ;
  assign n2590 = ( n2367 & n2368 ) | ( n2367 & n2589 ) | ( n2368 & n2589 ) ;
  assign n2591 = n2588 & n2590 ;
  assign n2592 = n2367 | n2368 ;
  assign n2593 = n2588 & n2592 ;
  assign n2594 = ( n2183 & n2591 ) | ( n2183 & n2593 ) | ( n2591 & n2593 ) ;
  assign n2595 = ( n2182 & n2591 ) | ( n2182 & n2593 ) | ( n2591 & n2593 ) ;
  assign n2596 = ( n1492 & n2594 ) | ( n1492 & n2595 ) | ( n2594 & n2595 ) ;
  assign n2597 = ( n1490 & n2594 ) | ( n1490 & n2595 ) | ( n2594 & n2595 ) ;
  assign n2598 = ( n917 & n2596 ) | ( n917 & n2597 ) | ( n2596 & n2597 ) ;
  assign n2599 = n2588 | n2590 ;
  assign n2600 = n2588 | n2592 ;
  assign n2601 = ( n2182 & n2599 ) | ( n2182 & n2600 ) | ( n2599 & n2600 ) ;
  assign n2602 = ( n2183 & n2599 ) | ( n2183 & n2600 ) | ( n2599 & n2600 ) ;
  assign n2603 = ( n1492 & n2601 ) | ( n1492 & n2602 ) | ( n2601 & n2602 ) ;
  assign n2604 = ( n1490 & n2601 ) | ( n1490 & n2602 ) | ( n2601 & n2602 ) ;
  assign n2605 = ( n917 & n2603 ) | ( n917 & n2604 ) | ( n2603 & n2604 ) ;
  assign n2606 = ~n2598 & n2605 ;
  assign n2607 = x85 & n133 ;
  assign n2608 = x84 & ~n162 ;
  assign n2609 = ( n137 & n2607 ) | ( n137 & n2608 ) | ( n2607 & n2608 ) ;
  assign n2610 = x0 & x86 ;
  assign n2611 = ( ~n137 & n2607 ) | ( ~n137 & n2610 ) | ( n2607 & n2610 ) ;
  assign n2612 = n2609 | n2611 ;
  assign n2613 = n141 | n2612 ;
  assign n2614 = ( n2606 & n2612 ) | ( n2606 & n2613 ) | ( n2612 & n2613 ) ;
  assign n2615 = x2 & n2612 ;
  assign n2616 = ( x2 & n523 ) | ( x2 & n2612 ) | ( n523 & n2612 ) ;
  assign n2617 = ( n2606 & n2615 ) | ( n2606 & n2616 ) | ( n2615 & n2616 ) ;
  assign n2618 = x2 & ~n2616 ;
  assign n2619 = x2 & ~n2612 ;
  assign n2620 = ( ~n2606 & n2618 ) | ( ~n2606 & n2619 ) | ( n2618 & n2619 ) ;
  assign n2621 = ( n2614 & ~n2617 ) | ( n2614 & n2620 ) | ( ~n2617 & n2620 ) ;
  assign n2622 = n2585 | n2621 ;
  assign n2623 = n2585 & n2621 ;
  assign n2624 = n2622 & ~n2623 ;
  assign n2625 = n2397 | n2402 ;
  assign n2626 = n2624 & n2625 ;
  assign n2627 = n2624 | n2625 ;
  assign n2628 = ~n2626 & n2627 ;
  assign n2629 = x66 & n2429 ;
  assign n2630 = x65 & n2424 ;
  assign n2631 = ~n2221 & n2428 ;
  assign n2632 = x64 & ~n2423 ;
  assign n2633 = n2631 & n2632 ;
  assign n2634 = n2630 | n2633 ;
  assign n2635 = n2629 | n2634 ;
  assign n2636 = n159 & n2432 ;
  assign n2637 = n2635 | n2636 ;
  assign n2638 = x23 | n2432 ;
  assign n2639 = ( x23 & n159 ) | ( x23 & n2638 ) | ( n159 & n2638 ) ;
  assign n2640 = n2635 | n2639 ;
  assign n2641 = ~x23 & n2639 ;
  assign n2642 = ( ~x23 & n2635 ) | ( ~x23 & n2641 ) | ( n2635 & n2641 ) ;
  assign n2643 = ( ~n2637 & n2640 ) | ( ~n2637 & n2642 ) | ( n2640 & n2642 ) ;
  assign n2644 = n2444 | n2643 ;
  assign n2645 = n2444 & n2643 ;
  assign n2646 = n2644 & ~n2645 ;
  assign n2647 = n293 & n1862 ;
  assign n2648 = x69 & n1859 ;
  assign n2649 = x68 & n1854 ;
  assign n2650 = x67 & ~n1853 ;
  assign n2651 = n2037 & n2650 ;
  assign n2652 = n2649 | n2651 ;
  assign n2653 = n2648 | n2652 ;
  assign n2654 = n2647 | n2653 ;
  assign n2655 = x20 | n2648 ;
  assign n2656 = n2652 | n2655 ;
  assign n2657 = n2647 | n2656 ;
  assign n2658 = ~x20 & n2656 ;
  assign n2659 = ( ~x20 & n2647 ) | ( ~x20 & n2658 ) | ( n2647 & n2658 ) ;
  assign n2660 = ( ~n2654 & n2657 ) | ( ~n2654 & n2659 ) | ( n2657 & n2659 ) ;
  assign n2661 = n2646 | n2660 ;
  assign n2662 = n2646 & n2660 ;
  assign n2663 = n2661 & ~n2662 ;
  assign n2664 = ( n2450 & n2464 ) | ( n2450 & n2468 ) | ( n2464 & n2468 ) ;
  assign n2665 = n2662 | n2664 ;
  assign n2666 = ( n2662 & n2663 ) | ( n2662 & n2665 ) | ( n2663 & n2665 ) ;
  assign n2667 = n2661 & ~n2666 ;
  assign n2668 = x72 & n1383 ;
  assign n2669 = x71 & n1378 ;
  assign n2670 = x70 & ~n1377 ;
  assign n2671 = n1542 & n2670 ;
  assign n2672 = n2669 | n2671 ;
  assign n2673 = n2668 | n2672 ;
  assign n2674 = ( n513 & n1386 ) | ( n513 & n2673 ) | ( n1386 & n2673 ) ;
  assign n2675 = ( x17 & n1386 ) | ( x17 & ~n2668 ) | ( n1386 & ~n2668 ) ;
  assign n2676 = x17 & n1386 ;
  assign n2677 = ( ~n2672 & n2675 ) | ( ~n2672 & n2676 ) | ( n2675 & n2676 ) ;
  assign n2678 = ( x17 & n513 ) | ( x17 & n2677 ) | ( n513 & n2677 ) ;
  assign n2679 = ~n2674 & n2678 ;
  assign n2680 = n2673 | n2677 ;
  assign n2681 = x17 | n2673 ;
  assign n2682 = ( n513 & n2680 ) | ( n513 & n2681 ) | ( n2680 & n2681 ) ;
  assign n2683 = ( ~x17 & n2679 ) | ( ~x17 & n2682 ) | ( n2679 & n2682 ) ;
  assign n2684 = n2664 & n2683 ;
  assign n2685 = ~n2663 & n2684 ;
  assign n2686 = ( n2667 & n2683 ) | ( n2667 & n2685 ) | ( n2683 & n2685 ) ;
  assign n2687 = n2664 | n2683 ;
  assign n2688 = ( ~n2663 & n2683 ) | ( ~n2663 & n2687 ) | ( n2683 & n2687 ) ;
  assign n2689 = n2667 | n2688 ;
  assign n2690 = ~n2686 & n2689 ;
  assign n2691 = n2472 | n2474 ;
  assign n2692 = ( n2472 & n2480 ) | ( n2472 & n2691 ) | ( n2480 & n2691 ) ;
  assign n2693 = n2690 & n2692 ;
  assign n2694 = n2690 | n2692 ;
  assign n2695 = ~n2693 & n2694 ;
  assign n2696 = x75 & n962 ;
  assign n2697 = x74 & n957 ;
  assign n2698 = x73 & ~n956 ;
  assign n2699 = n1105 & n2698 ;
  assign n2700 = n2697 | n2699 ;
  assign n2701 = n2696 | n2700 ;
  assign n2702 = n965 | n2696 ;
  assign n2703 = n2700 | n2702 ;
  assign n2704 = ( n746 & n2701 ) | ( n746 & n2703 ) | ( n2701 & n2703 ) ;
  assign n2705 = x14 & n2703 ;
  assign n2706 = x14 & n2696 ;
  assign n2707 = ( x14 & n2700 ) | ( x14 & n2706 ) | ( n2700 & n2706 ) ;
  assign n2708 = ( n746 & n2705 ) | ( n746 & n2707 ) | ( n2705 & n2707 ) ;
  assign n2709 = x14 & ~n2707 ;
  assign n2710 = x14 & ~n2703 ;
  assign n2711 = ( ~n746 & n2709 ) | ( ~n746 & n2710 ) | ( n2709 & n2710 ) ;
  assign n2712 = ( n2704 & ~n2708 ) | ( n2704 & n2711 ) | ( ~n2708 & n2711 ) ;
  assign n2713 = n2695 | n2712 ;
  assign n2714 = n2695 & n2712 ;
  assign n2715 = n2713 & ~n2714 ;
  assign n2716 = n2501 | n2507 ;
  assign n2717 = n2715 & n2716 ;
  assign n2718 = n2715 | n2716 ;
  assign n2719 = ~n2717 & n2718 ;
  assign n2720 = x78 & n636 ;
  assign n2721 = x77 & n631 ;
  assign n2722 = x76 & ~n630 ;
  assign n2723 = n764 & n2722 ;
  assign n2724 = n2721 | n2723 ;
  assign n2725 = n2720 | n2724 ;
  assign n2726 = n639 | n2720 ;
  assign n2727 = n2724 | n2726 ;
  assign n2728 = ( n1192 & n2725 ) | ( n1192 & n2727 ) | ( n2725 & n2727 ) ;
  assign n2729 = x11 & n2727 ;
  assign n2730 = x11 & n2720 ;
  assign n2731 = ( x11 & n2724 ) | ( x11 & n2730 ) | ( n2724 & n2730 ) ;
  assign n2732 = ( n1192 & n2729 ) | ( n1192 & n2731 ) | ( n2729 & n2731 ) ;
  assign n2733 = x11 & ~n2731 ;
  assign n2734 = x11 & ~n2727 ;
  assign n2735 = ( ~n1192 & n2733 ) | ( ~n1192 & n2734 ) | ( n2733 & n2734 ) ;
  assign n2736 = ( n2728 & ~n2732 ) | ( n2728 & n2735 ) | ( ~n2732 & n2735 ) ;
  assign n2737 = n2719 & n2736 ;
  assign n2738 = n2719 & ~n2737 ;
  assign n2739 = ~n2719 & n2736 ;
  assign n2740 = n2738 | n2739 ;
  assign n2741 = n2529 | n2533 ;
  assign n2742 = n2740 & n2741 ;
  assign n2743 = n2740 | n2741 ;
  assign n2744 = ~n2742 & n2743 ;
  assign n2745 = x81 & n389 ;
  assign n2746 = x80 & n384 ;
  assign n2747 = x79 & ~n383 ;
  assign n2748 = n463 & n2747 ;
  assign n2749 = n2746 | n2748 ;
  assign n2750 = n2745 | n2749 ;
  assign n2751 = n392 | n2745 ;
  assign n2752 = n2749 | n2751 ;
  assign n2753 = ( n1651 & n2750 ) | ( n1651 & n2752 ) | ( n2750 & n2752 ) ;
  assign n2754 = x8 & n2752 ;
  assign n2755 = x8 & n2745 ;
  assign n2756 = ( x8 & n2749 ) | ( x8 & n2755 ) | ( n2749 & n2755 ) ;
  assign n2757 = ( n1651 & n2754 ) | ( n1651 & n2756 ) | ( n2754 & n2756 ) ;
  assign n2758 = x8 & ~n2756 ;
  assign n2759 = x8 & ~n2752 ;
  assign n2760 = ( ~n1651 & n2758 ) | ( ~n1651 & n2759 ) | ( n2758 & n2759 ) ;
  assign n2761 = ( n2753 & ~n2757 ) | ( n2753 & n2760 ) | ( ~n2757 & n2760 ) ;
  assign n2762 = n2744 & n2761 ;
  assign n2763 = n2744 & ~n2762 ;
  assign n2764 = ~n2744 & n2761 ;
  assign n2765 = n2763 | n2764 ;
  assign n2766 = n2553 | n2557 ;
  assign n2767 = ~n2765 & n2766 ;
  assign n2768 = n2765 & ~n2766 ;
  assign n2769 = n2767 | n2768 ;
  assign n2770 = x84 & n212 ;
  assign n2771 = x83 & n207 ;
  assign n2772 = x82 & ~n206 ;
  assign n2773 = n267 & n2772 ;
  assign n2774 = n2771 | n2773 ;
  assign n2775 = n2770 | n2774 ;
  assign n2776 = n215 | n2770 ;
  assign n2777 = n2774 | n2776 ;
  assign n2778 = ( n2194 & n2775 ) | ( n2194 & n2777 ) | ( n2775 & n2777 ) ;
  assign n2779 = x5 & n2777 ;
  assign n2780 = x5 & n2770 ;
  assign n2781 = ( x5 & n2774 ) | ( x5 & n2780 ) | ( n2774 & n2780 ) ;
  assign n2782 = ( n2194 & n2779 ) | ( n2194 & n2781 ) | ( n2779 & n2781 ) ;
  assign n2783 = x5 & ~n2781 ;
  assign n2784 = x5 & ~n2777 ;
  assign n2785 = ( ~n2194 & n2783 ) | ( ~n2194 & n2784 ) | ( n2783 & n2784 ) ;
  assign n2786 = ( n2778 & ~n2782 ) | ( n2778 & n2785 ) | ( ~n2782 & n2785 ) ;
  assign n2787 = n2769 & n2786 ;
  assign n2788 = n2769 | n2786 ;
  assign n2789 = ~n2787 & n2788 ;
  assign n2790 = n2578 | n2580 ;
  assign n2791 = n2579 | n2790 ;
  assign n2792 = ( n2578 & n2582 ) | ( n2578 & n2791 ) | ( n2582 & n2791 ) ;
  assign n2793 = n2789 | n2792 ;
  assign n2794 = n2789 & n2792 ;
  assign n2795 = n2793 & ~n2794 ;
  assign n2796 = x86 | x87 ;
  assign n2797 = x86 & x87 ;
  assign n2798 = n2796 & ~n2797 ;
  assign n2799 = n2587 | n2588 ;
  assign n2800 = ( n2587 & n2590 ) | ( n2587 & n2799 ) | ( n2590 & n2799 ) ;
  assign n2801 = n2798 & n2800 ;
  assign n2802 = ( n2587 & n2592 ) | ( n2587 & n2799 ) | ( n2592 & n2799 ) ;
  assign n2803 = n2798 & n2802 ;
  assign n2804 = ( n2183 & n2801 ) | ( n2183 & n2803 ) | ( n2801 & n2803 ) ;
  assign n2805 = ( n2182 & n2801 ) | ( n2182 & n2803 ) | ( n2801 & n2803 ) ;
  assign n2806 = ( n1492 & n2804 ) | ( n1492 & n2805 ) | ( n2804 & n2805 ) ;
  assign n2807 = ( n1490 & n2804 ) | ( n1490 & n2805 ) | ( n2804 & n2805 ) ;
  assign n2808 = ( n917 & n2806 ) | ( n917 & n2807 ) | ( n2806 & n2807 ) ;
  assign n2809 = n2798 | n2802 ;
  assign n2810 = n2798 | n2800 ;
  assign n2811 = ( n2182 & n2809 ) | ( n2182 & n2810 ) | ( n2809 & n2810 ) ;
  assign n2812 = ( n2183 & n2809 ) | ( n2183 & n2810 ) | ( n2809 & n2810 ) ;
  assign n2813 = ( n1492 & n2811 ) | ( n1492 & n2812 ) | ( n2811 & n2812 ) ;
  assign n2814 = ( n1490 & n2811 ) | ( n1490 & n2812 ) | ( n2811 & n2812 ) ;
  assign n2815 = ( n917 & n2813 ) | ( n917 & n2814 ) | ( n2813 & n2814 ) ;
  assign n2816 = ~n2808 & n2815 ;
  assign n2817 = x86 & n133 ;
  assign n2818 = x85 & ~n162 ;
  assign n2819 = ( n137 & n2817 ) | ( n137 & n2818 ) | ( n2817 & n2818 ) ;
  assign n2820 = x0 & x87 ;
  assign n2821 = ( ~n137 & n2817 ) | ( ~n137 & n2820 ) | ( n2817 & n2820 ) ;
  assign n2822 = n2819 | n2821 ;
  assign n2823 = n141 | n2822 ;
  assign n2824 = ( n2816 & n2822 ) | ( n2816 & n2823 ) | ( n2822 & n2823 ) ;
  assign n2825 = x2 & n2822 ;
  assign n2826 = ( x2 & n523 ) | ( x2 & n2822 ) | ( n523 & n2822 ) ;
  assign n2827 = ( n2816 & n2825 ) | ( n2816 & n2826 ) | ( n2825 & n2826 ) ;
  assign n2828 = x2 & ~n2826 ;
  assign n2829 = x2 & ~n2822 ;
  assign n2830 = ( ~n2816 & n2828 ) | ( ~n2816 & n2829 ) | ( n2828 & n2829 ) ;
  assign n2831 = ( n2824 & ~n2827 ) | ( n2824 & n2830 ) | ( ~n2827 & n2830 ) ;
  assign n2832 = n2795 & n2831 ;
  assign n2833 = n2795 & ~n2832 ;
  assign n2834 = ~n2795 & n2831 ;
  assign n2835 = n2833 | n2834 ;
  assign n2836 = n2623 | n2624 ;
  assign n2837 = ( n2623 & n2625 ) | ( n2623 & n2836 ) | ( n2625 & n2836 ) ;
  assign n2838 = n2835 & n2837 ;
  assign n2839 = n2835 | n2837 ;
  assign n2840 = ~n2838 & n2839 ;
  assign n2841 = n2787 | n2794 ;
  assign n2842 = x23 & ~x24 ;
  assign n2843 = ~x23 & x24 ;
  assign n2844 = n2842 | n2843 ;
  assign n2845 = x64 & n2844 ;
  assign n2846 = ~n2444 & n2845 ;
  assign n2847 = ( ~n2643 & n2845 ) | ( ~n2643 & n2846 ) | ( n2845 & n2846 ) ;
  assign n2848 = n2444 & ~n2845 ;
  assign n2849 = n2643 & n2848 ;
  assign n2850 = n2847 | n2849 ;
  assign n2851 = x67 & n2429 ;
  assign n2852 = x66 & n2424 ;
  assign n2853 = x65 & ~n2423 ;
  assign n2854 = n2631 & n2853 ;
  assign n2855 = n2852 | n2854 ;
  assign n2856 = n2851 | n2855 ;
  assign n2857 = n186 & n2432 ;
  assign n2858 = n2856 | n2857 ;
  assign n2859 = x23 & ~n2858 ;
  assign n2860 = ~x23 & n2858 ;
  assign n2861 = n2859 | n2860 ;
  assign n2862 = n2850 & n2861 ;
  assign n2863 = n2850 | n2861 ;
  assign n2864 = ~n2862 & n2863 ;
  assign n2865 = x69 & n1854 ;
  assign n2866 = x68 & ~n1853 ;
  assign n2867 = n2037 & n2866 ;
  assign n2868 = n2865 | n2867 ;
  assign n2869 = x70 & n1859 ;
  assign n2870 = n1862 | n2869 ;
  assign n2871 = n2868 | n2870 ;
  assign n2872 = x20 & ~n2871 ;
  assign n2873 = x20 & ~n2869 ;
  assign n2874 = ~n2868 & n2873 ;
  assign n2875 = ( ~n340 & n2872 ) | ( ~n340 & n2874 ) | ( n2872 & n2874 ) ;
  assign n2876 = ~x20 & n2871 ;
  assign n2877 = ~x20 & n2869 ;
  assign n2878 = ( ~x20 & n2868 ) | ( ~x20 & n2877 ) | ( n2868 & n2877 ) ;
  assign n2879 = ( n340 & n2876 ) | ( n340 & n2878 ) | ( n2876 & n2878 ) ;
  assign n2880 = n2875 | n2879 ;
  assign n2881 = ( n2666 & ~n2864 ) | ( n2666 & n2880 ) | ( ~n2864 & n2880 ) ;
  assign n2882 = ( ~n2666 & n2864 ) | ( ~n2666 & n2881 ) | ( n2864 & n2881 ) ;
  assign n2883 = x73 & n1383 ;
  assign n2884 = x72 & n1378 ;
  assign n2885 = x71 & ~n1377 ;
  assign n2886 = n1542 & n2885 ;
  assign n2887 = n2884 | n2886 ;
  assign n2888 = n2883 | n2887 ;
  assign n2889 = n1386 | n2883 ;
  assign n2890 = n2887 | n2889 ;
  assign n2891 = ( ~n610 & n2888 ) | ( ~n610 & n2890 ) | ( n2888 & n2890 ) ;
  assign n2892 = n2888 & n2890 ;
  assign n2893 = ( n598 & n2891 ) | ( n598 & n2892 ) | ( n2891 & n2892 ) ;
  assign n2894 = x17 & n2893 ;
  assign n2895 = x17 | n2893 ;
  assign n2896 = ~n2894 & n2895 ;
  assign n2897 = ~n2880 & n2896 ;
  assign n2898 = ~n2864 & n2896 ;
  assign n2899 = n2880 & n2896 ;
  assign n2900 = ( n2666 & n2898 ) | ( n2666 & n2899 ) | ( n2898 & n2899 ) ;
  assign n2901 = ( n2882 & n2897 ) | ( n2882 & n2900 ) | ( n2897 & n2900 ) ;
  assign n2902 = n2880 & ~n2896 ;
  assign n2903 = n2864 & ~n2896 ;
  assign n2904 = n2880 | n2896 ;
  assign n2905 = ( n2666 & ~n2903 ) | ( n2666 & n2904 ) | ( ~n2903 & n2904 ) ;
  assign n2906 = ( n2882 & ~n2902 ) | ( n2882 & n2905 ) | ( ~n2902 & n2905 ) ;
  assign n2907 = ~n2901 & n2906 ;
  assign n2908 = n2686 | n2690 ;
  assign n2909 = ( n2686 & n2692 ) | ( n2686 & n2908 ) | ( n2692 & n2908 ) ;
  assign n2910 = n2907 & n2909 ;
  assign n2911 = n2907 | n2909 ;
  assign n2912 = ~n2910 & n2911 ;
  assign n2913 = x76 & n962 ;
  assign n2914 = x75 & n957 ;
  assign n2915 = x74 & ~n956 ;
  assign n2916 = n1105 & n2915 ;
  assign n2917 = n2914 | n2916 ;
  assign n2918 = n2913 | n2917 ;
  assign n2919 = n965 | n2913 ;
  assign n2920 = n2917 | n2919 ;
  assign n2921 = ( n923 & n2918 ) | ( n923 & n2920 ) | ( n2918 & n2920 ) ;
  assign n2922 = x14 & n2920 ;
  assign n2923 = x14 & n2913 ;
  assign n2924 = ( x14 & n2917 ) | ( x14 & n2923 ) | ( n2917 & n2923 ) ;
  assign n2925 = ( n923 & n2922 ) | ( n923 & n2924 ) | ( n2922 & n2924 ) ;
  assign n2926 = x14 & ~n2924 ;
  assign n2927 = x14 & ~n2920 ;
  assign n2928 = ( ~n923 & n2926 ) | ( ~n923 & n2927 ) | ( n2926 & n2927 ) ;
  assign n2929 = ( n2921 & ~n2925 ) | ( n2921 & n2928 ) | ( ~n2925 & n2928 ) ;
  assign n2930 = n2912 | n2929 ;
  assign n2931 = n2912 & n2929 ;
  assign n2932 = n2930 & ~n2931 ;
  assign n2933 = n2714 | n2715 ;
  assign n2934 = ( n2714 & n2716 ) | ( n2714 & n2933 ) | ( n2716 & n2933 ) ;
  assign n2935 = n2932 & n2934 ;
  assign n2936 = n2932 | n2934 ;
  assign n2937 = ~n2935 & n2936 ;
  assign n2938 = x79 & n636 ;
  assign n2939 = x78 & n631 ;
  assign n2940 = x77 & ~n630 ;
  assign n2941 = n764 & n2940 ;
  assign n2942 = n2939 | n2941 ;
  assign n2943 = n2938 | n2942 ;
  assign n2944 = n639 | n2938 ;
  assign n2945 = n2942 | n2944 ;
  assign n2946 = ( n1332 & n2943 ) | ( n1332 & n2945 ) | ( n2943 & n2945 ) ;
  assign n2947 = x11 & n2945 ;
  assign n2948 = x11 & n2938 ;
  assign n2949 = ( x11 & n2942 ) | ( x11 & n2948 ) | ( n2942 & n2948 ) ;
  assign n2950 = ( n1332 & n2947 ) | ( n1332 & n2949 ) | ( n2947 & n2949 ) ;
  assign n2951 = x11 & ~n2949 ;
  assign n2952 = x11 & ~n2945 ;
  assign n2953 = ( ~n1332 & n2951 ) | ( ~n1332 & n2952 ) | ( n2951 & n2952 ) ;
  assign n2954 = ( n2946 & ~n2950 ) | ( n2946 & n2953 ) | ( ~n2950 & n2953 ) ;
  assign n2955 = n2937 & n2954 ;
  assign n2956 = n2937 & ~n2955 ;
  assign n2957 = ~n2937 & n2954 ;
  assign n2958 = n2956 | n2957 ;
  assign n2959 = n2737 | n2741 ;
  assign n2960 = ( n2737 & n2740 ) | ( n2737 & n2959 ) | ( n2740 & n2959 ) ;
  assign n2961 = n2958 | n2960 ;
  assign n2962 = n2958 & n2960 ;
  assign n2963 = n2961 & ~n2962 ;
  assign n2964 = x82 & n389 ;
  assign n2965 = x81 & n384 ;
  assign n2966 = x80 & ~n383 ;
  assign n2967 = n463 & n2966 ;
  assign n2968 = n2965 | n2967 ;
  assign n2969 = n2964 | n2968 ;
  assign n2970 = n392 | n2964 ;
  assign n2971 = n2968 | n2970 ;
  assign n2972 = ( n1811 & n2969 ) | ( n1811 & n2971 ) | ( n2969 & n2971 ) ;
  assign n2973 = x8 & n2971 ;
  assign n2974 = x8 & n2964 ;
  assign n2975 = ( x8 & n2968 ) | ( x8 & n2974 ) | ( n2968 & n2974 ) ;
  assign n2976 = ( n1811 & n2973 ) | ( n1811 & n2975 ) | ( n2973 & n2975 ) ;
  assign n2977 = x8 & ~n2975 ;
  assign n2978 = x8 & ~n2971 ;
  assign n2979 = ( ~n1811 & n2977 ) | ( ~n1811 & n2978 ) | ( n2977 & n2978 ) ;
  assign n2980 = ( n2972 & ~n2976 ) | ( n2972 & n2979 ) | ( ~n2976 & n2979 ) ;
  assign n2981 = n2963 | n2980 ;
  assign n2982 = n2963 & n2980 ;
  assign n2983 = n2981 & ~n2982 ;
  assign n2984 = n2762 | n2766 ;
  assign n2985 = ( n2762 & n2765 ) | ( n2762 & n2984 ) | ( n2765 & n2984 ) ;
  assign n2986 = n2983 & n2985 ;
  assign n2987 = n2983 | n2985 ;
  assign n2988 = ~n2986 & n2987 ;
  assign n2989 = x85 & n212 ;
  assign n2990 = x84 & n207 ;
  assign n2991 = x83 & ~n206 ;
  assign n2992 = n267 & n2991 ;
  assign n2993 = n2990 | n2992 ;
  assign n2994 = n2989 | n2993 ;
  assign n2995 = n215 | n2989 ;
  assign n2996 = n2993 | n2995 ;
  assign n2997 = ( n2381 & n2994 ) | ( n2381 & n2996 ) | ( n2994 & n2996 ) ;
  assign n2998 = x5 & n2996 ;
  assign n2999 = x5 & n2989 ;
  assign n3000 = ( x5 & n2993 ) | ( x5 & n2999 ) | ( n2993 & n2999 ) ;
  assign n3001 = ( n2381 & n2998 ) | ( n2381 & n3000 ) | ( n2998 & n3000 ) ;
  assign n3002 = x5 & ~n3000 ;
  assign n3003 = x5 & ~n2996 ;
  assign n3004 = ( ~n2381 & n3002 ) | ( ~n2381 & n3003 ) | ( n3002 & n3003 ) ;
  assign n3005 = ( n2997 & ~n3001 ) | ( n2997 & n3004 ) | ( ~n3001 & n3004 ) ;
  assign n3006 = n2988 & n3005 ;
  assign n3007 = n2988 & ~n3006 ;
  assign n3008 = ~n2988 & n3005 ;
  assign n3009 = n3007 | n3008 ;
  assign n3010 = ~n2841 & n3009 ;
  assign n3011 = n2841 & ~n3009 ;
  assign n3012 = n3010 | n3011 ;
  assign n3013 = x87 | x88 ;
  assign n3014 = x87 & x88 ;
  assign n3015 = n3013 & ~n3014 ;
  assign n3016 = n2797 | n2798 ;
  assign n3017 = ( n2797 & n2800 ) | ( n2797 & n3016 ) | ( n2800 & n3016 ) ;
  assign n3018 = ( n2797 & n2802 ) | ( n2797 & n3016 ) | ( n2802 & n3016 ) ;
  assign n3019 = ( n2182 & n3017 ) | ( n2182 & n3018 ) | ( n3017 & n3018 ) ;
  assign n3020 = n3015 | n3019 ;
  assign n3021 = ( n2183 & n3017 ) | ( n2183 & n3018 ) | ( n3017 & n3018 ) ;
  assign n3022 = n3015 | n3021 ;
  assign n3023 = ( n1493 & n3020 ) | ( n1493 & n3022 ) | ( n3020 & n3022 ) ;
  assign n3024 = x87 & n133 ;
  assign n3025 = x86 & ~n162 ;
  assign n3026 = ( n137 & n3024 ) | ( n137 & n3025 ) | ( n3024 & n3025 ) ;
  assign n3027 = x0 & x88 ;
  assign n3028 = ( ~n137 & n3024 ) | ( ~n137 & n3027 ) | ( n3024 & n3027 ) ;
  assign n3029 = n3026 | n3028 ;
  assign n3030 = n141 | n3029 ;
  assign n3031 = n3015 & n3016 ;
  assign n3032 = n2797 & n3015 ;
  assign n3033 = ( n2800 & n3031 ) | ( n2800 & n3032 ) | ( n3031 & n3032 ) ;
  assign n3034 = ( n2802 & n3031 ) | ( n2802 & n3032 ) | ( n3031 & n3032 ) ;
  assign n3035 = ( n2183 & n3033 ) | ( n2183 & n3034 ) | ( n3033 & n3034 ) ;
  assign n3036 = ( n2182 & n3033 ) | ( n2182 & n3034 ) | ( n3033 & n3034 ) ;
  assign n3037 = ( n1492 & n3035 ) | ( n1492 & n3036 ) | ( n3035 & n3036 ) ;
  assign n3038 = ( n1490 & n3035 ) | ( n1490 & n3036 ) | ( n3035 & n3036 ) ;
  assign n3039 = ( n917 & n3037 ) | ( n917 & n3038 ) | ( n3037 & n3038 ) ;
  assign n3040 = ( n3029 & n3030 ) | ( n3029 & ~n3039 ) | ( n3030 & ~n3039 ) ;
  assign n3041 = n3029 & n3030 ;
  assign n3042 = ( n3023 & n3040 ) | ( n3023 & n3041 ) | ( n3040 & n3041 ) ;
  assign n3043 = x2 & n3029 ;
  assign n3044 = ( x2 & n523 ) | ( x2 & n3029 ) | ( n523 & n3029 ) ;
  assign n3045 = ( ~n3039 & n3043 ) | ( ~n3039 & n3044 ) | ( n3043 & n3044 ) ;
  assign n3046 = n3043 & n3044 ;
  assign n3047 = ( n3023 & n3045 ) | ( n3023 & n3046 ) | ( n3045 & n3046 ) ;
  assign n3048 = x2 & ~n3044 ;
  assign n3049 = x2 & ~n3029 ;
  assign n3050 = ( n3039 & n3048 ) | ( n3039 & n3049 ) | ( n3048 & n3049 ) ;
  assign n3051 = n3048 | n3049 ;
  assign n3052 = ( ~n3023 & n3050 ) | ( ~n3023 & n3051 ) | ( n3050 & n3051 ) ;
  assign n3053 = ( n3042 & ~n3047 ) | ( n3042 & n3052 ) | ( ~n3047 & n3052 ) ;
  assign n3054 = n3012 & n3053 ;
  assign n3055 = n3012 | n3053 ;
  assign n3056 = ~n3054 & n3055 ;
  assign n3057 = n2832 | n2838 ;
  assign n3058 = n3056 & n3057 ;
  assign n3059 = n3056 | n3057 ;
  assign n3060 = ~n3058 & n3059 ;
  assign n3061 = x70 & n1854 ;
  assign n3062 = x69 & ~n1853 ;
  assign n3063 = n2037 & n3062 ;
  assign n3064 = n3061 | n3063 ;
  assign n3065 = x71 & n1859 ;
  assign n3066 = n1862 | n3065 ;
  assign n3067 = n3064 | n3066 ;
  assign n3068 = x20 & ~n3067 ;
  assign n3069 = x20 & ~n3065 ;
  assign n3070 = ~n3064 & n3069 ;
  assign n3071 = ( ~n438 & n3068 ) | ( ~n438 & n3070 ) | ( n3068 & n3070 ) ;
  assign n3072 = ~x20 & n3067 ;
  assign n3073 = ~x20 & n3065 ;
  assign n3074 = ( ~x20 & n3064 ) | ( ~x20 & n3073 ) | ( n3064 & n3073 ) ;
  assign n3075 = ( n438 & n3072 ) | ( n438 & n3074 ) | ( n3072 & n3074 ) ;
  assign n3076 = n3071 | n3075 ;
  assign n3077 = ~x24 & x25 ;
  assign n3078 = x24 & ~x25 ;
  assign n3079 = n3077 | n3078 ;
  assign n3080 = ~n2844 & n3079 ;
  assign n3081 = x64 & n3080 ;
  assign n3082 = ~x25 & x26 ;
  assign n3083 = x25 & ~x26 ;
  assign n3084 = n3082 | n3083 ;
  assign n3085 = n2844 & ~n3084 ;
  assign n3086 = x65 & n3085 ;
  assign n3087 = n3081 | n3086 ;
  assign n3088 = n2844 & n3084 ;
  assign n3089 = x26 | n144 ;
  assign n3090 = ( x26 & n3088 ) | ( x26 & n3089 ) | ( n3088 & n3089 ) ;
  assign n3091 = ~x26 & n3090 ;
  assign n3092 = ( ~x26 & n3087 ) | ( ~x26 & n3091 ) | ( n3087 & n3091 ) ;
  assign n3093 = x26 & ~x64 ;
  assign n3094 = ( x26 & ~n2844 ) | ( x26 & n3093 ) | ( ~n2844 & n3093 ) ;
  assign n3095 = n3090 & n3094 ;
  assign n3096 = ( n3087 & n3094 ) | ( n3087 & n3095 ) | ( n3094 & n3095 ) ;
  assign n3097 = n144 & n3088 ;
  assign n3098 = n3094 & ~n3097 ;
  assign n3099 = ~n3087 & n3098 ;
  assign n3100 = ( n3092 & n3096 ) | ( n3092 & n3099 ) | ( n3096 & n3099 ) ;
  assign n3101 = n3090 | n3094 ;
  assign n3102 = n3087 | n3101 ;
  assign n3103 = ~n3094 & n3097 ;
  assign n3104 = ( n3087 & ~n3094 ) | ( n3087 & n3103 ) | ( ~n3094 & n3103 ) ;
  assign n3105 = ( n3092 & n3102 ) | ( n3092 & ~n3104 ) | ( n3102 & ~n3104 ) ;
  assign n3106 = ~n3100 & n3105 ;
  assign n3107 = n241 & n2432 ;
  assign n3108 = x68 & n2429 ;
  assign n3109 = x67 & n2424 ;
  assign n3110 = x66 & ~n2423 ;
  assign n3111 = n2631 & n3110 ;
  assign n3112 = n3109 | n3111 ;
  assign n3113 = n3108 | n3112 ;
  assign n3114 = n3107 | n3113 ;
  assign n3115 = x23 | n3108 ;
  assign n3116 = n3112 | n3115 ;
  assign n3117 = n3107 | n3116 ;
  assign n3118 = ~x23 & n3116 ;
  assign n3119 = ( ~x23 & n3107 ) | ( ~x23 & n3118 ) | ( n3107 & n3118 ) ;
  assign n3120 = ( ~n3114 & n3117 ) | ( ~n3114 & n3119 ) | ( n3117 & n3119 ) ;
  assign n3121 = n3106 & ~n3120 ;
  assign n3122 = ~n3106 & n3120 ;
  assign n3123 = n3121 | n3122 ;
  assign n3124 = ( n2645 & n2845 ) | ( n2645 & n2861 ) | ( n2845 & n2861 ) ;
  assign n3125 = n3123 | n3124 ;
  assign n3126 = n3123 & n3124 ;
  assign n3127 = n3125 & ~n3126 ;
  assign n3128 = n3076 & n3127 ;
  assign n3129 = n3076 | n3127 ;
  assign n3130 = ~n3128 & n3129 ;
  assign n3131 = n2864 & n2880 ;
  assign n3132 = n2864 & ~n3131 ;
  assign n3133 = ~n2864 & n2880 ;
  assign n3134 = n2666 & ~n3133 ;
  assign n3135 = ~n3132 & n3134 ;
  assign n3136 = ( n2666 & n3131 ) | ( n2666 & ~n3135 ) | ( n3131 & ~n3135 ) ;
  assign n3137 = n3130 & n3136 ;
  assign n3138 = n3130 | n3136 ;
  assign n3139 = ~n3137 & n3138 ;
  assign n3140 = x74 & n1383 ;
  assign n3141 = x73 & n1378 ;
  assign n3142 = x72 & ~n1377 ;
  assign n3143 = n1542 & n3142 ;
  assign n3144 = n3141 | n3143 ;
  assign n3145 = n3140 | n3144 ;
  assign n3146 = n1386 | n3140 ;
  assign n3147 = n3144 | n3146 ;
  assign n3148 = ( n710 & n3145 ) | ( n710 & n3147 ) | ( n3145 & n3147 ) ;
  assign n3149 = x17 & n3147 ;
  assign n3150 = x17 & n3140 ;
  assign n3151 = ( x17 & n3144 ) | ( x17 & n3150 ) | ( n3144 & n3150 ) ;
  assign n3152 = ( n710 & n3149 ) | ( n710 & n3151 ) | ( n3149 & n3151 ) ;
  assign n3153 = x17 & ~n3151 ;
  assign n3154 = x17 & ~n3147 ;
  assign n3155 = ( ~n710 & n3153 ) | ( ~n710 & n3154 ) | ( n3153 & n3154 ) ;
  assign n3156 = ( n3148 & ~n3152 ) | ( n3148 & n3155 ) | ( ~n3152 & n3155 ) ;
  assign n3157 = n3139 & n3156 ;
  assign n3158 = n3139 & ~n3157 ;
  assign n3159 = n2901 | n2907 ;
  assign n3160 = ( n2901 & n2909 ) | ( n2901 & n3159 ) | ( n2909 & n3159 ) ;
  assign n3161 = ~n3139 & n3156 ;
  assign n3162 = n3160 & n3161 ;
  assign n3163 = ( n3158 & n3160 ) | ( n3158 & n3162 ) | ( n3160 & n3162 ) ;
  assign n3164 = n3160 | n3161 ;
  assign n3165 = n3158 | n3164 ;
  assign n3166 = ~n3163 & n3165 ;
  assign n3167 = x77 & n962 ;
  assign n3168 = x76 & n957 ;
  assign n3169 = x75 & ~n956 ;
  assign n3170 = n1105 & n3169 ;
  assign n3171 = n3168 | n3170 ;
  assign n3172 = n3167 | n3171 ;
  assign n3173 = n965 | n3167 ;
  assign n3174 = n3171 | n3173 ;
  assign n3175 = ( n1059 & n3172 ) | ( n1059 & n3174 ) | ( n3172 & n3174 ) ;
  assign n3176 = x14 & n3174 ;
  assign n3177 = x14 & n3167 ;
  assign n3178 = ( x14 & n3171 ) | ( x14 & n3177 ) | ( n3171 & n3177 ) ;
  assign n3179 = ( n1059 & n3176 ) | ( n1059 & n3178 ) | ( n3176 & n3178 ) ;
  assign n3180 = x14 & ~n3178 ;
  assign n3181 = x14 & ~n3174 ;
  assign n3182 = ( ~n1059 & n3180 ) | ( ~n1059 & n3181 ) | ( n3180 & n3181 ) ;
  assign n3183 = ( n3175 & ~n3179 ) | ( n3175 & n3182 ) | ( ~n3179 & n3182 ) ;
  assign n3184 = n3166 | n3183 ;
  assign n3185 = n3166 & n3183 ;
  assign n3186 = n3184 & ~n3185 ;
  assign n3187 = n2931 | n2932 ;
  assign n3188 = ( n2931 & n2934 ) | ( n2931 & n3187 ) | ( n2934 & n3187 ) ;
  assign n3189 = n3186 & n3188 ;
  assign n3190 = n3186 | n3188 ;
  assign n3191 = ~n3189 & n3190 ;
  assign n3192 = x80 & n636 ;
  assign n3193 = x79 & n631 ;
  assign n3194 = x78 & ~n630 ;
  assign n3195 = n764 & n3194 ;
  assign n3196 = n3193 | n3195 ;
  assign n3197 = n3192 | n3196 ;
  assign n3198 = n639 | n3192 ;
  assign n3199 = n3196 | n3198 ;
  assign n3200 = ( n1499 & n3197 ) | ( n1499 & n3199 ) | ( n3197 & n3199 ) ;
  assign n3201 = x11 & n3199 ;
  assign n3202 = x11 & n3192 ;
  assign n3203 = ( x11 & n3196 ) | ( x11 & n3202 ) | ( n3196 & n3202 ) ;
  assign n3204 = ( n1499 & n3201 ) | ( n1499 & n3203 ) | ( n3201 & n3203 ) ;
  assign n3205 = x11 & ~n3203 ;
  assign n3206 = x11 & ~n3199 ;
  assign n3207 = ( ~n1499 & n3205 ) | ( ~n1499 & n3206 ) | ( n3205 & n3206 ) ;
  assign n3208 = ( n3200 & ~n3204 ) | ( n3200 & n3207 ) | ( ~n3204 & n3207 ) ;
  assign n3209 = n3191 & n3208 ;
  assign n3210 = n3191 & ~n3209 ;
  assign n3211 = ~n3191 & n3208 ;
  assign n3212 = n3210 | n3211 ;
  assign n3213 = n2955 | n2962 ;
  assign n3214 = n3212 | n3213 ;
  assign n3215 = n3212 & n3213 ;
  assign n3216 = n3214 & ~n3215 ;
  assign n3217 = x83 & n389 ;
  assign n3218 = x82 & n384 ;
  assign n3219 = x81 & ~n383 ;
  assign n3220 = n463 & n3219 ;
  assign n3221 = n3218 | n3220 ;
  assign n3222 = n3217 | n3221 ;
  assign n3223 = n392 | n3217 ;
  assign n3224 = n3221 | n3223 ;
  assign n3225 = ( n2009 & n3222 ) | ( n2009 & n3224 ) | ( n3222 & n3224 ) ;
  assign n3226 = x8 & n3224 ;
  assign n3227 = x8 & n3217 ;
  assign n3228 = ( x8 & n3221 ) | ( x8 & n3227 ) | ( n3221 & n3227 ) ;
  assign n3229 = ( n2009 & n3226 ) | ( n2009 & n3228 ) | ( n3226 & n3228 ) ;
  assign n3230 = x8 & ~n3228 ;
  assign n3231 = x8 & ~n3224 ;
  assign n3232 = ( ~n2009 & n3230 ) | ( ~n2009 & n3231 ) | ( n3230 & n3231 ) ;
  assign n3233 = ( n3225 & ~n3229 ) | ( n3225 & n3232 ) | ( ~n3229 & n3232 ) ;
  assign n3234 = n3216 & n3233 ;
  assign n3235 = n3216 & ~n3234 ;
  assign n3236 = ~n3216 & n3233 ;
  assign n3237 = n3235 | n3236 ;
  assign n3238 = n2982 | n2983 ;
  assign n3239 = ( n2982 & n2985 ) | ( n2982 & n3238 ) | ( n2985 & n3238 ) ;
  assign n3240 = n3237 & n3239 ;
  assign n3241 = n3237 & ~n3240 ;
  assign n3242 = x86 & n212 ;
  assign n3243 = x85 & n207 ;
  assign n3244 = x84 & ~n206 ;
  assign n3245 = n267 & n3244 ;
  assign n3246 = n3243 | n3245 ;
  assign n3247 = n3242 | n3246 ;
  assign n3248 = n215 | n3242 ;
  assign n3249 = n3246 | n3248 ;
  assign n3250 = ( n2606 & n3247 ) | ( n2606 & n3249 ) | ( n3247 & n3249 ) ;
  assign n3251 = x5 & n3249 ;
  assign n3252 = x5 & n3242 ;
  assign n3253 = ( x5 & n3246 ) | ( x5 & n3252 ) | ( n3246 & n3252 ) ;
  assign n3254 = ( n2606 & n3251 ) | ( n2606 & n3253 ) | ( n3251 & n3253 ) ;
  assign n3255 = x5 & ~n3253 ;
  assign n3256 = x5 & ~n3249 ;
  assign n3257 = ( ~n2606 & n3255 ) | ( ~n2606 & n3256 ) | ( n3255 & n3256 ) ;
  assign n3258 = ( n3250 & ~n3254 ) | ( n3250 & n3257 ) | ( ~n3254 & n3257 ) ;
  assign n3259 = n3239 & ~n3258 ;
  assign n3260 = ~n3237 & n3259 ;
  assign n3261 = ( n3241 & ~n3258 ) | ( n3241 & n3260 ) | ( ~n3258 & n3260 ) ;
  assign n3262 = ~n3239 & n3258 ;
  assign n3263 = ( n3237 & n3258 ) | ( n3237 & n3262 ) | ( n3258 & n3262 ) ;
  assign n3264 = ~n3241 & n3263 ;
  assign n3265 = n3261 | n3264 ;
  assign n3266 = n2841 & n3009 ;
  assign n3267 = n3006 | n3266 ;
  assign n3268 = n3265 & n3267 ;
  assign n3269 = n3265 | n3267 ;
  assign n3270 = ~n3268 & n3269 ;
  assign n3271 = x88 | x89 ;
  assign n3272 = x88 & x89 ;
  assign n3273 = n3271 & ~n3272 ;
  assign n3274 = n3014 | n3035 ;
  assign n3275 = n3273 & n3274 ;
  assign n3276 = n3014 | n3036 ;
  assign n3277 = n3273 & n3276 ;
  assign n3278 = ( n1493 & n3275 ) | ( n1493 & n3277 ) | ( n3275 & n3277 ) ;
  assign n3279 = n3273 | n3274 ;
  assign n3280 = n3273 | n3276 ;
  assign n3281 = ( n1493 & n3279 ) | ( n1493 & n3280 ) | ( n3279 & n3280 ) ;
  assign n3282 = ~n3278 & n3281 ;
  assign n3283 = x88 & n133 ;
  assign n3284 = x87 & ~n162 ;
  assign n3285 = ( n137 & n3283 ) | ( n137 & n3284 ) | ( n3283 & n3284 ) ;
  assign n3286 = x0 & x89 ;
  assign n3287 = ( ~n137 & n3283 ) | ( ~n137 & n3286 ) | ( n3283 & n3286 ) ;
  assign n3288 = n3285 | n3287 ;
  assign n3289 = n141 | n3288 ;
  assign n3290 = ( n3282 & n3288 ) | ( n3282 & n3289 ) | ( n3288 & n3289 ) ;
  assign n3291 = x2 & n3288 ;
  assign n3292 = ( x2 & n523 ) | ( x2 & n3288 ) | ( n523 & n3288 ) ;
  assign n3293 = ( n3282 & n3291 ) | ( n3282 & n3292 ) | ( n3291 & n3292 ) ;
  assign n3294 = x2 & ~n3292 ;
  assign n3295 = x2 & ~n3288 ;
  assign n3296 = ( ~n3282 & n3294 ) | ( ~n3282 & n3295 ) | ( n3294 & n3295 ) ;
  assign n3297 = ( n3290 & ~n3293 ) | ( n3290 & n3296 ) | ( ~n3293 & n3296 ) ;
  assign n3298 = n3270 & n3297 ;
  assign n3299 = n3270 | n3297 ;
  assign n3300 = ~n3298 & n3299 ;
  assign n3301 = n3054 | n3056 ;
  assign n3302 = ( n3054 & n3057 ) | ( n3054 & n3301 ) | ( n3057 & n3301 ) ;
  assign n3303 = n3300 & n3302 ;
  assign n3304 = n3300 | n3302 ;
  assign n3305 = ~n3303 & n3304 ;
  assign n3306 = n3185 | n3189 ;
  assign n3307 = x66 & n3085 ;
  assign n3308 = x65 & n3080 ;
  assign n3309 = ~n2844 & n3084 ;
  assign n3310 = x64 & ~n3079 ;
  assign n3311 = n3309 & n3310 ;
  assign n3312 = n3308 | n3311 ;
  assign n3313 = n3307 | n3312 ;
  assign n3314 = n159 & n3088 ;
  assign n3315 = n3313 | n3314 ;
  assign n3316 = x26 | n3088 ;
  assign n3317 = ( x26 & n159 ) | ( x26 & n3316 ) | ( n159 & n3316 ) ;
  assign n3318 = n3313 | n3317 ;
  assign n3319 = ~x26 & n3317 ;
  assign n3320 = ( ~x26 & n3313 ) | ( ~x26 & n3319 ) | ( n3313 & n3319 ) ;
  assign n3321 = ( ~n3315 & n3318 ) | ( ~n3315 & n3320 ) | ( n3318 & n3320 ) ;
  assign n3322 = n3100 | n3321 ;
  assign n3323 = n3100 & n3321 ;
  assign n3324 = n3322 & ~n3323 ;
  assign n3325 = n293 & n2432 ;
  assign n3326 = x69 & n2429 ;
  assign n3327 = x68 & n2424 ;
  assign n3328 = x67 & ~n2423 ;
  assign n3329 = n2631 & n3328 ;
  assign n3330 = n3327 | n3329 ;
  assign n3331 = n3326 | n3330 ;
  assign n3332 = n3325 | n3331 ;
  assign n3333 = x23 | n3326 ;
  assign n3334 = n3330 | n3333 ;
  assign n3335 = n3325 | n3334 ;
  assign n3336 = ~x23 & n3334 ;
  assign n3337 = ( ~x23 & n3325 ) | ( ~x23 & n3336 ) | ( n3325 & n3336 ) ;
  assign n3338 = ( ~n3332 & n3335 ) | ( ~n3332 & n3337 ) | ( n3335 & n3337 ) ;
  assign n3339 = n3324 | n3338 ;
  assign n3340 = n3324 & n3338 ;
  assign n3341 = n3339 & ~n3340 ;
  assign n3342 = ( n3106 & n3120 ) | ( n3106 & n3124 ) | ( n3120 & n3124 ) ;
  assign n3343 = n3340 | n3342 ;
  assign n3344 = ( n3340 & n3341 ) | ( n3340 & n3343 ) | ( n3341 & n3343 ) ;
  assign n3345 = n3339 & ~n3344 ;
  assign n3346 = x72 & n1859 ;
  assign n3347 = x71 & n1854 ;
  assign n3348 = x70 & ~n1853 ;
  assign n3349 = n2037 & n3348 ;
  assign n3350 = n3347 | n3349 ;
  assign n3351 = n3346 | n3350 ;
  assign n3352 = ( n513 & n1862 ) | ( n513 & n3351 ) | ( n1862 & n3351 ) ;
  assign n3353 = ( x20 & n1862 ) | ( x20 & ~n3346 ) | ( n1862 & ~n3346 ) ;
  assign n3354 = x20 & n1862 ;
  assign n3355 = ( ~n3350 & n3353 ) | ( ~n3350 & n3354 ) | ( n3353 & n3354 ) ;
  assign n3356 = ( x20 & n513 ) | ( x20 & n3355 ) | ( n513 & n3355 ) ;
  assign n3357 = ~n3352 & n3356 ;
  assign n3358 = n3351 | n3355 ;
  assign n3359 = x20 | n3351 ;
  assign n3360 = ( n513 & n3358 ) | ( n513 & n3359 ) | ( n3358 & n3359 ) ;
  assign n3361 = ( ~x20 & n3357 ) | ( ~x20 & n3360 ) | ( n3357 & n3360 ) ;
  assign n3362 = n3342 & n3361 ;
  assign n3363 = ~n3341 & n3362 ;
  assign n3364 = ( n3345 & n3361 ) | ( n3345 & n3363 ) | ( n3361 & n3363 ) ;
  assign n3365 = n3342 | n3361 ;
  assign n3366 = ( ~n3341 & n3361 ) | ( ~n3341 & n3365 ) | ( n3361 & n3365 ) ;
  assign n3367 = n3345 | n3366 ;
  assign n3368 = ~n3364 & n3367 ;
  assign n3369 = n3128 | n3130 ;
  assign n3370 = ( n3128 & n3136 ) | ( n3128 & n3369 ) | ( n3136 & n3369 ) ;
  assign n3371 = n3368 & n3370 ;
  assign n3372 = n3368 | n3370 ;
  assign n3373 = ~n3371 & n3372 ;
  assign n3374 = x75 & n1383 ;
  assign n3375 = x74 & n1378 ;
  assign n3376 = x73 & ~n1377 ;
  assign n3377 = n1542 & n3376 ;
  assign n3378 = n3375 | n3377 ;
  assign n3379 = n3374 | n3378 ;
  assign n3380 = n1386 | n3374 ;
  assign n3381 = n3378 | n3380 ;
  assign n3382 = ( n746 & n3379 ) | ( n746 & n3381 ) | ( n3379 & n3381 ) ;
  assign n3383 = x17 & n3381 ;
  assign n3384 = x17 & n3374 ;
  assign n3385 = ( x17 & n3378 ) | ( x17 & n3384 ) | ( n3378 & n3384 ) ;
  assign n3386 = ( n746 & n3383 ) | ( n746 & n3385 ) | ( n3383 & n3385 ) ;
  assign n3387 = x17 & ~n3385 ;
  assign n3388 = x17 & ~n3381 ;
  assign n3389 = ( ~n746 & n3387 ) | ( ~n746 & n3388 ) | ( n3387 & n3388 ) ;
  assign n3390 = ( n3382 & ~n3386 ) | ( n3382 & n3389 ) | ( ~n3386 & n3389 ) ;
  assign n3391 = n3373 | n3390 ;
  assign n3392 = n3373 & n3390 ;
  assign n3393 = n3391 & ~n3392 ;
  assign n3394 = n3157 | n3163 ;
  assign n3395 = n3393 & n3394 ;
  assign n3396 = n3393 | n3394 ;
  assign n3397 = ~n3395 & n3396 ;
  assign n3398 = x78 & n962 ;
  assign n3399 = x77 & n957 ;
  assign n3400 = x76 & ~n956 ;
  assign n3401 = n1105 & n3400 ;
  assign n3402 = n3399 | n3401 ;
  assign n3403 = n3398 | n3402 ;
  assign n3404 = n965 | n3398 ;
  assign n3405 = n3402 | n3404 ;
  assign n3406 = ( n1192 & n3403 ) | ( n1192 & n3405 ) | ( n3403 & n3405 ) ;
  assign n3407 = x14 & n3405 ;
  assign n3408 = x14 & n3398 ;
  assign n3409 = ( x14 & n3402 ) | ( x14 & n3408 ) | ( n3402 & n3408 ) ;
  assign n3410 = ( n1192 & n3407 ) | ( n1192 & n3409 ) | ( n3407 & n3409 ) ;
  assign n3411 = x14 & ~n3409 ;
  assign n3412 = x14 & ~n3405 ;
  assign n3413 = ( ~n1192 & n3411 ) | ( ~n1192 & n3412 ) | ( n3411 & n3412 ) ;
  assign n3414 = ( n3406 & ~n3410 ) | ( n3406 & n3413 ) | ( ~n3410 & n3413 ) ;
  assign n3415 = n3397 & n3414 ;
  assign n3416 = n3397 & ~n3415 ;
  assign n3417 = ~n3397 & n3414 ;
  assign n3418 = n3416 | n3417 ;
  assign n3419 = n3306 & ~n3418 ;
  assign n3420 = ~n3306 & n3418 ;
  assign n3421 = n3419 | n3420 ;
  assign n3422 = x81 & n636 ;
  assign n3423 = x80 & n631 ;
  assign n3424 = x79 & ~n630 ;
  assign n3425 = n764 & n3424 ;
  assign n3426 = n3423 | n3425 ;
  assign n3427 = n3422 | n3426 ;
  assign n3428 = n639 | n3422 ;
  assign n3429 = n3426 | n3428 ;
  assign n3430 = ( n1651 & n3427 ) | ( n1651 & n3429 ) | ( n3427 & n3429 ) ;
  assign n3431 = x11 & n3429 ;
  assign n3432 = x11 & n3422 ;
  assign n3433 = ( x11 & n3426 ) | ( x11 & n3432 ) | ( n3426 & n3432 ) ;
  assign n3434 = ( n1651 & n3431 ) | ( n1651 & n3433 ) | ( n3431 & n3433 ) ;
  assign n3435 = x11 & ~n3433 ;
  assign n3436 = x11 & ~n3429 ;
  assign n3437 = ( ~n1651 & n3435 ) | ( ~n1651 & n3436 ) | ( n3435 & n3436 ) ;
  assign n3438 = ( n3430 & ~n3434 ) | ( n3430 & n3437 ) | ( ~n3434 & n3437 ) ;
  assign n3439 = n3421 & n3438 ;
  assign n3440 = n3421 | n3438 ;
  assign n3441 = ~n3439 & n3440 ;
  assign n3442 = n3209 | n3211 ;
  assign n3443 = n3210 | n3442 ;
  assign n3444 = ( n3209 & n3213 ) | ( n3209 & n3443 ) | ( n3213 & n3443 ) ;
  assign n3445 = n3441 | n3444 ;
  assign n3446 = n3441 & n3444 ;
  assign n3447 = n3445 & ~n3446 ;
  assign n3448 = x84 & n389 ;
  assign n3449 = x83 & n384 ;
  assign n3450 = x82 & ~n383 ;
  assign n3451 = n463 & n3450 ;
  assign n3452 = n3449 | n3451 ;
  assign n3453 = n3448 | n3452 ;
  assign n3454 = n392 | n3448 ;
  assign n3455 = n3452 | n3454 ;
  assign n3456 = ( n2194 & n3453 ) | ( n2194 & n3455 ) | ( n3453 & n3455 ) ;
  assign n3457 = x8 & n3455 ;
  assign n3458 = x8 & n3448 ;
  assign n3459 = ( x8 & n3452 ) | ( x8 & n3458 ) | ( n3452 & n3458 ) ;
  assign n3460 = ( n2194 & n3457 ) | ( n2194 & n3459 ) | ( n3457 & n3459 ) ;
  assign n3461 = x8 & ~n3459 ;
  assign n3462 = x8 & ~n3455 ;
  assign n3463 = ( ~n2194 & n3461 ) | ( ~n2194 & n3462 ) | ( n3461 & n3462 ) ;
  assign n3464 = ( n3456 & ~n3460 ) | ( n3456 & n3463 ) | ( ~n3460 & n3463 ) ;
  assign n3465 = n3447 & n3464 ;
  assign n3466 = n3447 & ~n3465 ;
  assign n3467 = ~n3447 & n3464 ;
  assign n3468 = n3466 | n3467 ;
  assign n3469 = n3234 | n3239 ;
  assign n3470 = ( n3234 & n3237 ) | ( n3234 & n3469 ) | ( n3237 & n3469 ) ;
  assign n3471 = n3468 | n3470 ;
  assign n3472 = n3468 & n3470 ;
  assign n3473 = n3471 & ~n3472 ;
  assign n3474 = x87 & n212 ;
  assign n3475 = x86 & n207 ;
  assign n3476 = x85 & ~n206 ;
  assign n3477 = n267 & n3476 ;
  assign n3478 = n3475 | n3477 ;
  assign n3479 = n3474 | n3478 ;
  assign n3480 = n215 | n3474 ;
  assign n3481 = n3478 | n3480 ;
  assign n3482 = ( n2816 & n3479 ) | ( n2816 & n3481 ) | ( n3479 & n3481 ) ;
  assign n3483 = x5 & n3481 ;
  assign n3484 = x5 & n3474 ;
  assign n3485 = ( x5 & n3478 ) | ( x5 & n3484 ) | ( n3478 & n3484 ) ;
  assign n3486 = ( n2816 & n3483 ) | ( n2816 & n3485 ) | ( n3483 & n3485 ) ;
  assign n3487 = x5 & ~n3485 ;
  assign n3488 = x5 & ~n3481 ;
  assign n3489 = ( ~n2816 & n3487 ) | ( ~n2816 & n3488 ) | ( n3487 & n3488 ) ;
  assign n3490 = ( n3482 & ~n3486 ) | ( n3482 & n3489 ) | ( ~n3486 & n3489 ) ;
  assign n3491 = n3473 & n3490 ;
  assign n3492 = n3473 & ~n3491 ;
  assign n3493 = ~n3473 & n3490 ;
  assign n3494 = n3492 | n3493 ;
  assign n3495 = ~n3237 & n3239 ;
  assign n3496 = ( n3006 & n3258 ) | ( n3006 & n3495 ) | ( n3258 & n3495 ) ;
  assign n3497 = n3006 | n3258 ;
  assign n3498 = ( n3241 & n3496 ) | ( n3241 & n3497 ) | ( n3496 & n3497 ) ;
  assign n3499 = n3258 | n3495 ;
  assign n3500 = n3241 | n3499 ;
  assign n3501 = ( n3266 & n3498 ) | ( n3266 & n3500 ) | ( n3498 & n3500 ) ;
  assign n3502 = ~n3494 & n3501 ;
  assign n3503 = n3494 & ~n3501 ;
  assign n3504 = n3502 | n3503 ;
  assign n3505 = x89 | x90 ;
  assign n3506 = x89 & x90 ;
  assign n3507 = n3505 & ~n3506 ;
  assign n3508 = n3272 | n3273 ;
  assign n3509 = n3507 & n3508 ;
  assign n3510 = n3272 & n3507 ;
  assign n3511 = ( n3274 & n3509 ) | ( n3274 & n3510 ) | ( n3509 & n3510 ) ;
  assign n3512 = ( n3276 & n3509 ) | ( n3276 & n3510 ) | ( n3509 & n3510 ) ;
  assign n3513 = ( n1493 & n3511 ) | ( n1493 & n3512 ) | ( n3511 & n3512 ) ;
  assign n3514 = n3507 | n3508 ;
  assign n3515 = n3272 | n3507 ;
  assign n3516 = ( n3274 & n3514 ) | ( n3274 & n3515 ) | ( n3514 & n3515 ) ;
  assign n3517 = ( n3276 & n3514 ) | ( n3276 & n3515 ) | ( n3514 & n3515 ) ;
  assign n3518 = ( n1493 & n3516 ) | ( n1493 & n3517 ) | ( n3516 & n3517 ) ;
  assign n3519 = ~n3513 & n3518 ;
  assign n3520 = x89 & n133 ;
  assign n3521 = x88 & ~n162 ;
  assign n3522 = ( n137 & n3520 ) | ( n137 & n3521 ) | ( n3520 & n3521 ) ;
  assign n3523 = x0 & x90 ;
  assign n3524 = ( ~n137 & n3520 ) | ( ~n137 & n3523 ) | ( n3520 & n3523 ) ;
  assign n3525 = n3522 | n3524 ;
  assign n3526 = n141 | n3525 ;
  assign n3527 = ( n3519 & n3525 ) | ( n3519 & n3526 ) | ( n3525 & n3526 ) ;
  assign n3528 = x2 & n3525 ;
  assign n3529 = ( x2 & n523 ) | ( x2 & n3525 ) | ( n523 & n3525 ) ;
  assign n3530 = ( n3519 & n3528 ) | ( n3519 & n3529 ) | ( n3528 & n3529 ) ;
  assign n3531 = x2 & ~n3529 ;
  assign n3532 = x2 & ~n3525 ;
  assign n3533 = ( ~n3519 & n3531 ) | ( ~n3519 & n3532 ) | ( n3531 & n3532 ) ;
  assign n3534 = ( n3527 & ~n3530 ) | ( n3527 & n3533 ) | ( ~n3530 & n3533 ) ;
  assign n3535 = n3504 & n3534 ;
  assign n3536 = n3504 | n3534 ;
  assign n3537 = ~n3535 & n3536 ;
  assign n3538 = n3298 | n3303 ;
  assign n3539 = n3537 & n3538 ;
  assign n3540 = n3537 | n3538 ;
  assign n3541 = ~n3539 & n3540 ;
  assign n3542 = x26 & ~x27 ;
  assign n3543 = ~x26 & x27 ;
  assign n3544 = n3542 | n3543 ;
  assign n3545 = x64 & n3544 ;
  assign n3546 = ~n3100 & n3545 ;
  assign n3547 = ( ~n3321 & n3545 ) | ( ~n3321 & n3546 ) | ( n3545 & n3546 ) ;
  assign n3548 = n3100 & ~n3545 ;
  assign n3549 = n3321 & n3548 ;
  assign n3550 = n3547 | n3549 ;
  assign n3551 = x67 & n3085 ;
  assign n3552 = x66 & n3080 ;
  assign n3553 = x65 & ~n3079 ;
  assign n3554 = n3309 & n3553 ;
  assign n3555 = n3552 | n3554 ;
  assign n3556 = n3551 | n3555 ;
  assign n3557 = n186 & n3088 ;
  assign n3558 = n3556 | n3557 ;
  assign n3559 = x26 & ~n3558 ;
  assign n3560 = ~x26 & n3558 ;
  assign n3561 = n3559 | n3560 ;
  assign n3562 = n3550 & n3561 ;
  assign n3563 = n3550 | n3561 ;
  assign n3564 = ~n3562 & n3563 ;
  assign n3565 = x69 & n2424 ;
  assign n3566 = x68 & ~n2423 ;
  assign n3567 = n2631 & n3566 ;
  assign n3568 = n3565 | n3567 ;
  assign n3569 = x70 & n2429 ;
  assign n3570 = n2432 | n3569 ;
  assign n3571 = n3568 | n3570 ;
  assign n3572 = x23 & ~n3571 ;
  assign n3573 = x23 & ~n3569 ;
  assign n3574 = ~n3568 & n3573 ;
  assign n3575 = ( ~n340 & n3572 ) | ( ~n340 & n3574 ) | ( n3572 & n3574 ) ;
  assign n3576 = ~x23 & n3571 ;
  assign n3577 = ~x23 & n3569 ;
  assign n3578 = ( ~x23 & n3568 ) | ( ~x23 & n3577 ) | ( n3568 & n3577 ) ;
  assign n3579 = ( n340 & n3576 ) | ( n340 & n3578 ) | ( n3576 & n3578 ) ;
  assign n3580 = n3575 | n3579 ;
  assign n3581 = n3564 & n3580 ;
  assign n3582 = n3564 & ~n3581 ;
  assign n3583 = ~n3564 & n3580 ;
  assign n3584 = n3344 | n3583 ;
  assign n3585 = n3582 | n3584 ;
  assign n3586 = ~n3344 & n3585 ;
  assign n3587 = x73 & n1859 ;
  assign n3588 = x72 & n1854 ;
  assign n3589 = x71 & ~n1853 ;
  assign n3590 = n2037 & n3589 ;
  assign n3591 = n3588 | n3590 ;
  assign n3592 = n3587 | n3591 ;
  assign n3593 = n1862 | n3587 ;
  assign n3594 = n3591 | n3593 ;
  assign n3595 = ( ~n610 & n3592 ) | ( ~n610 & n3594 ) | ( n3592 & n3594 ) ;
  assign n3596 = n3592 & n3594 ;
  assign n3597 = ( n598 & n3595 ) | ( n598 & n3596 ) | ( n3595 & n3596 ) ;
  assign n3598 = x20 & n3597 ;
  assign n3599 = x20 | n3597 ;
  assign n3600 = ~n3598 & n3599 ;
  assign n3601 = n3585 & n3600 ;
  assign n3602 = ~n3583 & n3600 ;
  assign n3603 = ~n3582 & n3602 ;
  assign n3604 = ( n3586 & n3601 ) | ( n3586 & n3603 ) | ( n3601 & n3603 ) ;
  assign n3605 = n3585 | n3600 ;
  assign n3606 = n3583 & ~n3600 ;
  assign n3607 = ( n3582 & ~n3600 ) | ( n3582 & n3606 ) | ( ~n3600 & n3606 ) ;
  assign n3608 = ( n3586 & n3605 ) | ( n3586 & ~n3607 ) | ( n3605 & ~n3607 ) ;
  assign n3609 = ~n3604 & n3608 ;
  assign n3610 = n3364 | n3368 ;
  assign n3611 = ( n3364 & n3370 ) | ( n3364 & n3610 ) | ( n3370 & n3610 ) ;
  assign n3612 = n3609 & n3611 ;
  assign n3613 = n3609 | n3611 ;
  assign n3614 = ~n3612 & n3613 ;
  assign n3615 = x76 & n1383 ;
  assign n3616 = x75 & n1378 ;
  assign n3617 = x74 & ~n1377 ;
  assign n3618 = n1542 & n3617 ;
  assign n3619 = n3616 | n3618 ;
  assign n3620 = n3615 | n3619 ;
  assign n3621 = n1386 | n3615 ;
  assign n3622 = n3619 | n3621 ;
  assign n3623 = ( n923 & n3620 ) | ( n923 & n3622 ) | ( n3620 & n3622 ) ;
  assign n3624 = x17 & n3622 ;
  assign n3625 = x17 & n3615 ;
  assign n3626 = ( x17 & n3619 ) | ( x17 & n3625 ) | ( n3619 & n3625 ) ;
  assign n3627 = ( n923 & n3624 ) | ( n923 & n3626 ) | ( n3624 & n3626 ) ;
  assign n3628 = x17 & ~n3626 ;
  assign n3629 = x17 & ~n3622 ;
  assign n3630 = ( ~n923 & n3628 ) | ( ~n923 & n3629 ) | ( n3628 & n3629 ) ;
  assign n3631 = ( n3623 & ~n3627 ) | ( n3623 & n3630 ) | ( ~n3627 & n3630 ) ;
  assign n3632 = n3614 | n3631 ;
  assign n3633 = n3614 & n3631 ;
  assign n3634 = n3632 & ~n3633 ;
  assign n3635 = n3392 | n3393 ;
  assign n3636 = ( n3392 & n3394 ) | ( n3392 & n3635 ) | ( n3394 & n3635 ) ;
  assign n3637 = n3634 & n3636 ;
  assign n3638 = n3634 | n3636 ;
  assign n3639 = ~n3637 & n3638 ;
  assign n3640 = x79 & n962 ;
  assign n3641 = x78 & n957 ;
  assign n3642 = x77 & ~n956 ;
  assign n3643 = n1105 & n3642 ;
  assign n3644 = n3641 | n3643 ;
  assign n3645 = n3640 | n3644 ;
  assign n3646 = n965 | n3640 ;
  assign n3647 = n3644 | n3646 ;
  assign n3648 = ( n1332 & n3645 ) | ( n1332 & n3647 ) | ( n3645 & n3647 ) ;
  assign n3649 = x14 & n3647 ;
  assign n3650 = x14 & n3640 ;
  assign n3651 = ( x14 & n3644 ) | ( x14 & n3650 ) | ( n3644 & n3650 ) ;
  assign n3652 = ( n1332 & n3649 ) | ( n1332 & n3651 ) | ( n3649 & n3651 ) ;
  assign n3653 = x14 & ~n3651 ;
  assign n3654 = x14 & ~n3647 ;
  assign n3655 = ( ~n1332 & n3653 ) | ( ~n1332 & n3654 ) | ( n3653 & n3654 ) ;
  assign n3656 = ( n3648 & ~n3652 ) | ( n3648 & n3655 ) | ( ~n3652 & n3655 ) ;
  assign n3657 = n3639 & n3656 ;
  assign n3658 = n3639 & ~n3657 ;
  assign n3659 = ( n3185 & n3397 ) | ( n3185 & n3414 ) | ( n3397 & n3414 ) ;
  assign n3660 = n3397 | n3414 ;
  assign n3661 = ( n3189 & n3659 ) | ( n3189 & n3660 ) | ( n3659 & n3660 ) ;
  assign n3662 = ~n3639 & n3656 ;
  assign n3663 = n3661 & n3662 ;
  assign n3664 = ( n3658 & n3661 ) | ( n3658 & n3663 ) | ( n3661 & n3663 ) ;
  assign n3665 = n3661 | n3662 ;
  assign n3666 = n3658 | n3665 ;
  assign n3667 = ~n3664 & n3666 ;
  assign n3668 = x82 & n636 ;
  assign n3669 = x81 & n631 ;
  assign n3670 = x80 & ~n630 ;
  assign n3671 = n764 & n3670 ;
  assign n3672 = n3669 | n3671 ;
  assign n3673 = n3668 | n3672 ;
  assign n3674 = n639 | n3668 ;
  assign n3675 = n3672 | n3674 ;
  assign n3676 = ( n1811 & n3673 ) | ( n1811 & n3675 ) | ( n3673 & n3675 ) ;
  assign n3677 = x11 & n3675 ;
  assign n3678 = x11 & n3668 ;
  assign n3679 = ( x11 & n3672 ) | ( x11 & n3678 ) | ( n3672 & n3678 ) ;
  assign n3680 = ( n1811 & n3677 ) | ( n1811 & n3679 ) | ( n3677 & n3679 ) ;
  assign n3681 = x11 & ~n3679 ;
  assign n3682 = x11 & ~n3675 ;
  assign n3683 = ( ~n1811 & n3681 ) | ( ~n1811 & n3682 ) | ( n3681 & n3682 ) ;
  assign n3684 = ( n3676 & ~n3680 ) | ( n3676 & n3683 ) | ( ~n3680 & n3683 ) ;
  assign n3685 = n3667 & n3684 ;
  assign n3686 = n3667 & ~n3685 ;
  assign n3687 = ~n3667 & n3684 ;
  assign n3688 = n3686 | n3687 ;
  assign n3689 = n3439 | n3446 ;
  assign n3690 = n3688 | n3689 ;
  assign n3691 = n3688 & n3689 ;
  assign n3692 = n3690 & ~n3691 ;
  assign n3693 = x85 & n389 ;
  assign n3694 = x84 & n384 ;
  assign n3695 = x83 & ~n383 ;
  assign n3696 = n463 & n3695 ;
  assign n3697 = n3694 | n3696 ;
  assign n3698 = n3693 | n3697 ;
  assign n3699 = n392 | n3693 ;
  assign n3700 = n3697 | n3699 ;
  assign n3701 = ( n2381 & n3698 ) | ( n2381 & n3700 ) | ( n3698 & n3700 ) ;
  assign n3702 = x8 & n3700 ;
  assign n3703 = x8 & n3693 ;
  assign n3704 = ( x8 & n3697 ) | ( x8 & n3703 ) | ( n3697 & n3703 ) ;
  assign n3705 = ( n2381 & n3702 ) | ( n2381 & n3704 ) | ( n3702 & n3704 ) ;
  assign n3706 = x8 & ~n3704 ;
  assign n3707 = x8 & ~n3700 ;
  assign n3708 = ( ~n2381 & n3706 ) | ( ~n2381 & n3707 ) | ( n3706 & n3707 ) ;
  assign n3709 = ( n3701 & ~n3705 ) | ( n3701 & n3708 ) | ( ~n3705 & n3708 ) ;
  assign n3710 = n3692 | n3709 ;
  assign n3711 = n3692 & n3709 ;
  assign n3712 = n3710 & ~n3711 ;
  assign n3713 = n3465 | n3472 ;
  assign n3714 = n3712 & n3713 ;
  assign n3715 = n3712 | n3713 ;
  assign n3716 = ~n3714 & n3715 ;
  assign n3717 = x88 & n212 ;
  assign n3718 = x87 & n207 ;
  assign n3719 = x86 & ~n206 ;
  assign n3720 = n267 & n3719 ;
  assign n3721 = n3718 | n3720 ;
  assign n3722 = n3717 | n3721 ;
  assign n3723 = n215 | n3717 ;
  assign n3724 = n3721 | n3723 ;
  assign n3725 = ( ~n3039 & n3722 ) | ( ~n3039 & n3724 ) | ( n3722 & n3724 ) ;
  assign n3726 = n3722 & n3724 ;
  assign n3727 = ( n3023 & n3725 ) | ( n3023 & n3726 ) | ( n3725 & n3726 ) ;
  assign n3728 = x5 & n3724 ;
  assign n3729 = x5 & n3717 ;
  assign n3730 = ( x5 & n3721 ) | ( x5 & n3729 ) | ( n3721 & n3729 ) ;
  assign n3731 = ( ~n3039 & n3728 ) | ( ~n3039 & n3730 ) | ( n3728 & n3730 ) ;
  assign n3732 = n3728 & n3730 ;
  assign n3733 = ( n3023 & n3731 ) | ( n3023 & n3732 ) | ( n3731 & n3732 ) ;
  assign n3734 = x5 & ~n3730 ;
  assign n3735 = x5 & ~n3724 ;
  assign n3736 = ( n3039 & n3734 ) | ( n3039 & n3735 ) | ( n3734 & n3735 ) ;
  assign n3737 = n3734 | n3735 ;
  assign n3738 = ( ~n3023 & n3736 ) | ( ~n3023 & n3737 ) | ( n3736 & n3737 ) ;
  assign n3739 = ( n3727 & ~n3733 ) | ( n3727 & n3738 ) | ( ~n3733 & n3738 ) ;
  assign n3740 = n3716 & n3739 ;
  assign n3741 = n3716 & ~n3740 ;
  assign n3743 = ( n3473 & n3490 ) | ( n3473 & n3500 ) | ( n3490 & n3500 ) ;
  assign n3744 = ( n3473 & n3490 ) | ( n3473 & n3498 ) | ( n3490 & n3498 ) ;
  assign n3745 = ( n3266 & n3743 ) | ( n3266 & n3744 ) | ( n3743 & n3744 ) ;
  assign n3742 = ~n3716 & n3739 ;
  assign n3746 = n3742 & n3745 ;
  assign n3747 = ( n3741 & n3745 ) | ( n3741 & n3746 ) | ( n3745 & n3746 ) ;
  assign n3748 = n3742 | n3745 ;
  assign n3749 = n3741 | n3748 ;
  assign n3750 = ~n3747 & n3749 ;
  assign n3751 = x90 | x91 ;
  assign n3752 = x90 & x91 ;
  assign n3753 = n3751 & ~n3752 ;
  assign n3754 = n3506 | n3507 ;
  assign n3755 = ( n3506 & n3508 ) | ( n3506 & n3754 ) | ( n3508 & n3754 ) ;
  assign n3756 = n3753 & n3755 ;
  assign n3757 = n3272 | n3506 ;
  assign n3758 = ( n3506 & n3507 ) | ( n3506 & n3757 ) | ( n3507 & n3757 ) ;
  assign n3759 = n3753 & n3758 ;
  assign n3760 = ( n3274 & n3756 ) | ( n3274 & n3759 ) | ( n3756 & n3759 ) ;
  assign n3761 = ( n3276 & n3756 ) | ( n3276 & n3759 ) | ( n3756 & n3759 ) ;
  assign n3762 = ( n1493 & n3760 ) | ( n1493 & n3761 ) | ( n3760 & n3761 ) ;
  assign n3763 = n3753 | n3755 ;
  assign n3764 = n3753 | n3758 ;
  assign n3765 = ( n3274 & n3763 ) | ( n3274 & n3764 ) | ( n3763 & n3764 ) ;
  assign n3766 = ( n3276 & n3763 ) | ( n3276 & n3764 ) | ( n3763 & n3764 ) ;
  assign n3767 = ( n1493 & n3765 ) | ( n1493 & n3766 ) | ( n3765 & n3766 ) ;
  assign n3768 = ~n3762 & n3767 ;
  assign n3769 = x90 & n133 ;
  assign n3770 = x89 & ~n162 ;
  assign n3771 = ( n137 & n3769 ) | ( n137 & n3770 ) | ( n3769 & n3770 ) ;
  assign n3772 = x0 & x91 ;
  assign n3773 = ( ~n137 & n3769 ) | ( ~n137 & n3772 ) | ( n3769 & n3772 ) ;
  assign n3774 = n3771 | n3773 ;
  assign n3775 = n141 | n3774 ;
  assign n3776 = ( n3768 & n3774 ) | ( n3768 & n3775 ) | ( n3774 & n3775 ) ;
  assign n3777 = x2 & n3774 ;
  assign n3778 = ( x2 & n523 ) | ( x2 & n3774 ) | ( n523 & n3774 ) ;
  assign n3779 = ( n3768 & n3777 ) | ( n3768 & n3778 ) | ( n3777 & n3778 ) ;
  assign n3780 = x2 & ~n3778 ;
  assign n3781 = x2 & ~n3774 ;
  assign n3782 = ( ~n3768 & n3780 ) | ( ~n3768 & n3781 ) | ( n3780 & n3781 ) ;
  assign n3783 = ( n3776 & ~n3779 ) | ( n3776 & n3782 ) | ( ~n3779 & n3782 ) ;
  assign n3784 = n3750 | n3783 ;
  assign n3785 = n3750 & n3783 ;
  assign n3786 = n3784 & ~n3785 ;
  assign n3787 = n3535 | n3537 ;
  assign n3788 = ( n3535 & n3538 ) | ( n3535 & n3787 ) | ( n3538 & n3787 ) ;
  assign n3789 = n3786 & n3788 ;
  assign n3790 = n3786 | n3788 ;
  assign n3791 = ~n3789 & n3790 ;
  assign n3792 = x70 & n2424 ;
  assign n3793 = x69 & ~n2423 ;
  assign n3794 = n2631 & n3793 ;
  assign n3795 = n3792 | n3794 ;
  assign n3796 = x71 & n2429 ;
  assign n3797 = n2432 | n3796 ;
  assign n3798 = n3795 | n3797 ;
  assign n3799 = x23 & ~n3798 ;
  assign n3800 = x23 & ~n3796 ;
  assign n3801 = ~n3795 & n3800 ;
  assign n3802 = ( ~n438 & n3799 ) | ( ~n438 & n3801 ) | ( n3799 & n3801 ) ;
  assign n3803 = ~x23 & n3798 ;
  assign n3804 = ~x23 & n3796 ;
  assign n3805 = ( ~x23 & n3795 ) | ( ~x23 & n3804 ) | ( n3795 & n3804 ) ;
  assign n3806 = ( n438 & n3803 ) | ( n438 & n3805 ) | ( n3803 & n3805 ) ;
  assign n3807 = n3802 | n3806 ;
  assign n3808 = ~x27 & x28 ;
  assign n3809 = x27 & ~x28 ;
  assign n3810 = n3808 | n3809 ;
  assign n3811 = ~n3544 & n3810 ;
  assign n3812 = x64 & n3811 ;
  assign n3813 = ~x28 & x29 ;
  assign n3814 = x28 & ~x29 ;
  assign n3815 = n3813 | n3814 ;
  assign n3816 = n3544 & ~n3815 ;
  assign n3817 = x65 & n3816 ;
  assign n3818 = n3812 | n3817 ;
  assign n3819 = n3544 & n3815 ;
  assign n3820 = x29 | n144 ;
  assign n3821 = ( x29 & n3819 ) | ( x29 & n3820 ) | ( n3819 & n3820 ) ;
  assign n3822 = ~x29 & n3821 ;
  assign n3823 = ( ~x29 & n3818 ) | ( ~x29 & n3822 ) | ( n3818 & n3822 ) ;
  assign n3824 = x29 & ~x64 ;
  assign n3825 = ( x29 & ~n3544 ) | ( x29 & n3824 ) | ( ~n3544 & n3824 ) ;
  assign n3826 = n3821 & n3825 ;
  assign n3827 = ( n3818 & n3825 ) | ( n3818 & n3826 ) | ( n3825 & n3826 ) ;
  assign n3828 = n144 & n3819 ;
  assign n3829 = n3825 & ~n3828 ;
  assign n3830 = ~n3818 & n3829 ;
  assign n3831 = ( n3823 & n3827 ) | ( n3823 & n3830 ) | ( n3827 & n3830 ) ;
  assign n3832 = n3821 | n3825 ;
  assign n3833 = n3818 | n3832 ;
  assign n3834 = ~n3825 & n3828 ;
  assign n3835 = ( n3818 & ~n3825 ) | ( n3818 & n3834 ) | ( ~n3825 & n3834 ) ;
  assign n3836 = ( n3823 & n3833 ) | ( n3823 & ~n3835 ) | ( n3833 & ~n3835 ) ;
  assign n3837 = ~n3831 & n3836 ;
  assign n3838 = n241 & n3088 ;
  assign n3839 = x68 & n3085 ;
  assign n3840 = x67 & n3080 ;
  assign n3841 = x66 & ~n3079 ;
  assign n3842 = n3309 & n3841 ;
  assign n3843 = n3840 | n3842 ;
  assign n3844 = n3839 | n3843 ;
  assign n3845 = n3838 | n3844 ;
  assign n3846 = x26 | n3839 ;
  assign n3847 = n3843 | n3846 ;
  assign n3848 = n3838 | n3847 ;
  assign n3849 = ~x26 & n3847 ;
  assign n3850 = ( ~x26 & n3838 ) | ( ~x26 & n3849 ) | ( n3838 & n3849 ) ;
  assign n3851 = ( ~n3845 & n3848 ) | ( ~n3845 & n3850 ) | ( n3848 & n3850 ) ;
  assign n3852 = n3837 & ~n3851 ;
  assign n3853 = ~n3837 & n3851 ;
  assign n3854 = n3852 | n3853 ;
  assign n3855 = ( n3323 & n3545 ) | ( n3323 & n3561 ) | ( n3545 & n3561 ) ;
  assign n3856 = n3854 | n3855 ;
  assign n3857 = n3854 & n3855 ;
  assign n3858 = n3856 & ~n3857 ;
  assign n3859 = n3807 & n3858 ;
  assign n3860 = n3807 | n3858 ;
  assign n3861 = ~n3859 & n3860 ;
  assign n3862 = n3344 & ~n3583 ;
  assign n3863 = ~n3582 & n3862 ;
  assign n3864 = ( n3344 & n3581 ) | ( n3344 & ~n3863 ) | ( n3581 & ~n3863 ) ;
  assign n3865 = n3861 & n3864 ;
  assign n3866 = n3861 | n3864 ;
  assign n3867 = ~n3865 & n3866 ;
  assign n3868 = x74 & n1859 ;
  assign n3869 = x73 & n1854 ;
  assign n3870 = x72 & ~n1853 ;
  assign n3871 = n2037 & n3870 ;
  assign n3872 = n3869 | n3871 ;
  assign n3873 = n3868 | n3872 ;
  assign n3874 = n1862 | n3868 ;
  assign n3875 = n3872 | n3874 ;
  assign n3876 = ( n710 & n3873 ) | ( n710 & n3875 ) | ( n3873 & n3875 ) ;
  assign n3877 = x20 & n3875 ;
  assign n3878 = x20 & n3868 ;
  assign n3879 = ( x20 & n3872 ) | ( x20 & n3878 ) | ( n3872 & n3878 ) ;
  assign n3880 = ( n710 & n3877 ) | ( n710 & n3879 ) | ( n3877 & n3879 ) ;
  assign n3881 = x20 & ~n3879 ;
  assign n3882 = x20 & ~n3875 ;
  assign n3883 = ( ~n710 & n3881 ) | ( ~n710 & n3882 ) | ( n3881 & n3882 ) ;
  assign n3884 = ( n3876 & ~n3880 ) | ( n3876 & n3883 ) | ( ~n3880 & n3883 ) ;
  assign n3885 = n3867 & n3884 ;
  assign n3886 = n3867 & ~n3885 ;
  assign n3887 = ~n3867 & n3884 ;
  assign n3888 = n3886 | n3887 ;
  assign n3889 = n3604 | n3612 ;
  assign n3890 = n3888 | n3889 ;
  assign n3891 = n3888 & n3889 ;
  assign n3892 = n3890 & ~n3891 ;
  assign n3893 = x77 & n1383 ;
  assign n3894 = x76 & n1378 ;
  assign n3895 = x75 & ~n1377 ;
  assign n3896 = n1542 & n3895 ;
  assign n3897 = n3894 | n3896 ;
  assign n3898 = n3893 | n3897 ;
  assign n3899 = n1386 | n3893 ;
  assign n3900 = n3897 | n3899 ;
  assign n3901 = ( n1059 & n3898 ) | ( n1059 & n3900 ) | ( n3898 & n3900 ) ;
  assign n3902 = x17 & n3900 ;
  assign n3903 = x17 & n3893 ;
  assign n3904 = ( x17 & n3897 ) | ( x17 & n3903 ) | ( n3897 & n3903 ) ;
  assign n3905 = ( n1059 & n3902 ) | ( n1059 & n3904 ) | ( n3902 & n3904 ) ;
  assign n3906 = x17 & ~n3904 ;
  assign n3907 = x17 & ~n3900 ;
  assign n3908 = ( ~n1059 & n3906 ) | ( ~n1059 & n3907 ) | ( n3906 & n3907 ) ;
  assign n3909 = ( n3901 & ~n3905 ) | ( n3901 & n3908 ) | ( ~n3905 & n3908 ) ;
  assign n3910 = n3892 & n3909 ;
  assign n3911 = n3892 & ~n3910 ;
  assign n3912 = ~n3892 & n3909 ;
  assign n3913 = n3633 | n3634 ;
  assign n3914 = ( n3633 & n3636 ) | ( n3633 & n3913 ) | ( n3636 & n3913 ) ;
  assign n3915 = ~n3912 & n3914 ;
  assign n3916 = ~n3911 & n3915 ;
  assign n3917 = n3912 & ~n3914 ;
  assign n3918 = ( n3911 & ~n3914 ) | ( n3911 & n3917 ) | ( ~n3914 & n3917 ) ;
  assign n3919 = n3916 | n3918 ;
  assign n3920 = x80 & n962 ;
  assign n3921 = x79 & n957 ;
  assign n3922 = x78 & ~n956 ;
  assign n3923 = n1105 & n3922 ;
  assign n3924 = n3921 | n3923 ;
  assign n3925 = n3920 | n3924 ;
  assign n3926 = n965 | n3920 ;
  assign n3927 = n3924 | n3926 ;
  assign n3928 = ( n1499 & n3925 ) | ( n1499 & n3927 ) | ( n3925 & n3927 ) ;
  assign n3929 = x14 & n3927 ;
  assign n3930 = x14 & n3920 ;
  assign n3931 = ( x14 & n3924 ) | ( x14 & n3930 ) | ( n3924 & n3930 ) ;
  assign n3932 = ( n1499 & n3929 ) | ( n1499 & n3931 ) | ( n3929 & n3931 ) ;
  assign n3933 = x14 & ~n3931 ;
  assign n3934 = x14 & ~n3927 ;
  assign n3935 = ( ~n1499 & n3933 ) | ( ~n1499 & n3934 ) | ( n3933 & n3934 ) ;
  assign n3936 = ( n3928 & ~n3932 ) | ( n3928 & n3935 ) | ( ~n3932 & n3935 ) ;
  assign n3937 = n3919 & n3936 ;
  assign n3938 = n3919 | n3936 ;
  assign n3939 = ~n3937 & n3938 ;
  assign n3940 = n3657 | n3664 ;
  assign n3941 = n3939 | n3940 ;
  assign n3942 = n3939 & n3940 ;
  assign n3943 = n3941 & ~n3942 ;
  assign n3944 = x83 & n636 ;
  assign n3945 = x82 & n631 ;
  assign n3946 = x81 & ~n630 ;
  assign n3947 = n764 & n3946 ;
  assign n3948 = n3945 | n3947 ;
  assign n3949 = n3944 | n3948 ;
  assign n3950 = n639 | n3944 ;
  assign n3951 = n3948 | n3950 ;
  assign n3952 = ( n2009 & n3949 ) | ( n2009 & n3951 ) | ( n3949 & n3951 ) ;
  assign n3953 = x11 & n3951 ;
  assign n3954 = x11 & n3944 ;
  assign n3955 = ( x11 & n3948 ) | ( x11 & n3954 ) | ( n3948 & n3954 ) ;
  assign n3956 = ( n2009 & n3953 ) | ( n2009 & n3955 ) | ( n3953 & n3955 ) ;
  assign n3957 = x11 & ~n3955 ;
  assign n3958 = x11 & ~n3951 ;
  assign n3959 = ( ~n2009 & n3957 ) | ( ~n2009 & n3958 ) | ( n3957 & n3958 ) ;
  assign n3960 = ( n3952 & ~n3956 ) | ( n3952 & n3959 ) | ( ~n3956 & n3959 ) ;
  assign n3961 = n3943 & n3960 ;
  assign n3962 = n3943 & ~n3961 ;
  assign n3963 = ~n3943 & n3960 ;
  assign n3964 = n3962 | n3963 ;
  assign n3965 = n3685 | n3687 ;
  assign n3966 = n3686 | n3965 ;
  assign n3967 = ( n3685 & n3689 ) | ( n3685 & n3966 ) | ( n3689 & n3966 ) ;
  assign n3968 = n3964 | n3967 ;
  assign n3969 = n3964 & n3967 ;
  assign n3970 = n3968 & ~n3969 ;
  assign n3971 = x86 & n389 ;
  assign n3972 = x85 & n384 ;
  assign n3973 = x84 & ~n383 ;
  assign n3974 = n463 & n3973 ;
  assign n3975 = n3972 | n3974 ;
  assign n3976 = n3971 | n3975 ;
  assign n3977 = n392 | n3971 ;
  assign n3978 = n3975 | n3977 ;
  assign n3979 = ( n2606 & n3976 ) | ( n2606 & n3978 ) | ( n3976 & n3978 ) ;
  assign n3980 = x8 & n3978 ;
  assign n3981 = x8 & n3971 ;
  assign n3982 = ( x8 & n3975 ) | ( x8 & n3981 ) | ( n3975 & n3981 ) ;
  assign n3983 = ( n2606 & n3980 ) | ( n2606 & n3982 ) | ( n3980 & n3982 ) ;
  assign n3984 = x8 & ~n3982 ;
  assign n3985 = x8 & ~n3978 ;
  assign n3986 = ( ~n2606 & n3984 ) | ( ~n2606 & n3985 ) | ( n3984 & n3985 ) ;
  assign n3987 = ( n3979 & ~n3983 ) | ( n3979 & n3986 ) | ( ~n3983 & n3986 ) ;
  assign n3988 = n3970 | n3987 ;
  assign n3989 = n3970 & n3987 ;
  assign n3990 = n3988 & ~n3989 ;
  assign n3991 = n3711 | n3712 ;
  assign n3992 = ( n3711 & n3713 ) | ( n3711 & n3991 ) | ( n3713 & n3991 ) ;
  assign n3993 = n3990 & n3992 ;
  assign n3994 = n3990 | n3992 ;
  assign n3995 = ~n3993 & n3994 ;
  assign n3996 = x89 & n212 ;
  assign n3997 = x88 & n207 ;
  assign n3998 = x87 & ~n206 ;
  assign n3999 = n267 & n3998 ;
  assign n4000 = n3997 | n3999 ;
  assign n4001 = n3996 | n4000 ;
  assign n4002 = n215 | n3996 ;
  assign n4003 = n4000 | n4002 ;
  assign n4004 = ( n3282 & n4001 ) | ( n3282 & n4003 ) | ( n4001 & n4003 ) ;
  assign n4005 = x5 & n4003 ;
  assign n4006 = x5 & n3996 ;
  assign n4007 = ( x5 & n4000 ) | ( x5 & n4006 ) | ( n4000 & n4006 ) ;
  assign n4008 = ( n3282 & n4005 ) | ( n3282 & n4007 ) | ( n4005 & n4007 ) ;
  assign n4009 = x5 & ~n4007 ;
  assign n4010 = x5 & ~n4003 ;
  assign n4011 = ( ~n3282 & n4009 ) | ( ~n3282 & n4010 ) | ( n4009 & n4010 ) ;
  assign n4012 = ( n4004 & ~n4008 ) | ( n4004 & n4011 ) | ( ~n4008 & n4011 ) ;
  assign n4013 = n3995 & n4012 ;
  assign n4014 = n3995 & ~n4013 ;
  assign n4015 = ~n3995 & n4012 ;
  assign n4016 = n4014 | n4015 ;
  assign n4017 = n3740 | n3747 ;
  assign n4018 = n4016 | n4017 ;
  assign n4019 = n4016 & n4017 ;
  assign n4020 = n4018 & ~n4019 ;
  assign n4021 = x91 | x92 ;
  assign n4022 = x91 & x92 ;
  assign n4023 = n4021 & ~n4022 ;
  assign n4024 = n3752 | n3753 ;
  assign n4025 = ( n3752 & n3758 ) | ( n3752 & n4024 ) | ( n3758 & n4024 ) ;
  assign n4026 = n4023 & n4025 ;
  assign n4027 = n4023 & n4024 ;
  assign n4028 = n3752 & n4023 ;
  assign n4029 = ( n3755 & n4027 ) | ( n3755 & n4028 ) | ( n4027 & n4028 ) ;
  assign n4030 = ( n3274 & n4026 ) | ( n3274 & n4029 ) | ( n4026 & n4029 ) ;
  assign n4031 = ( n3276 & n4026 ) | ( n3276 & n4029 ) | ( n4026 & n4029 ) ;
  assign n4032 = ( n1493 & n4030 ) | ( n1493 & n4031 ) | ( n4030 & n4031 ) ;
  assign n4033 = n4023 | n4025 ;
  assign n4034 = n4023 | n4024 ;
  assign n4035 = n3752 | n4023 ;
  assign n4036 = ( n3755 & n4034 ) | ( n3755 & n4035 ) | ( n4034 & n4035 ) ;
  assign n4037 = ( n3274 & n4033 ) | ( n3274 & n4036 ) | ( n4033 & n4036 ) ;
  assign n4038 = ( n3276 & n4033 ) | ( n3276 & n4036 ) | ( n4033 & n4036 ) ;
  assign n4039 = ( n1493 & n4037 ) | ( n1493 & n4038 ) | ( n4037 & n4038 ) ;
  assign n4040 = ~n4032 & n4039 ;
  assign n4041 = x91 & n133 ;
  assign n4042 = x90 & ~n162 ;
  assign n4043 = ( n137 & n4041 ) | ( n137 & n4042 ) | ( n4041 & n4042 ) ;
  assign n4044 = x0 & x92 ;
  assign n4045 = ( ~n137 & n4041 ) | ( ~n137 & n4044 ) | ( n4041 & n4044 ) ;
  assign n4046 = n4043 | n4045 ;
  assign n4047 = n141 | n4046 ;
  assign n4048 = ( n4040 & n4046 ) | ( n4040 & n4047 ) | ( n4046 & n4047 ) ;
  assign n4049 = x2 & n4046 ;
  assign n4050 = ( x2 & n523 ) | ( x2 & n4046 ) | ( n523 & n4046 ) ;
  assign n4051 = ( n4040 & n4049 ) | ( n4040 & n4050 ) | ( n4049 & n4050 ) ;
  assign n4052 = x2 & ~n4050 ;
  assign n4053 = x2 & ~n4046 ;
  assign n4054 = ( ~n4040 & n4052 ) | ( ~n4040 & n4053 ) | ( n4052 & n4053 ) ;
  assign n4055 = ( n4048 & ~n4051 ) | ( n4048 & n4054 ) | ( ~n4051 & n4054 ) ;
  assign n4056 = n4020 | n4055 ;
  assign n4057 = n4020 & n4055 ;
  assign n4058 = n4056 & ~n4057 ;
  assign n4059 = n3785 | n3786 ;
  assign n4060 = ( n3785 & n3788 ) | ( n3785 & n4059 ) | ( n3788 & n4059 ) ;
  assign n4061 = n4058 & n4060 ;
  assign n4062 = n4058 | n4060 ;
  assign n4063 = ~n4061 & n4062 ;
  assign n4064 = n4057 | n4061 ;
  assign n4065 = x66 & n3816 ;
  assign n4066 = x65 & n3811 ;
  assign n4067 = ~n3544 & n3815 ;
  assign n4068 = x64 & ~n3810 ;
  assign n4069 = n4067 & n4068 ;
  assign n4070 = n4066 | n4069 ;
  assign n4071 = n4065 | n4070 ;
  assign n4072 = n159 & n3819 ;
  assign n4073 = n4071 | n4072 ;
  assign n4074 = x29 | n3819 ;
  assign n4075 = ( x29 & n159 ) | ( x29 & n4074 ) | ( n159 & n4074 ) ;
  assign n4076 = n4071 | n4075 ;
  assign n4077 = ~x29 & n4075 ;
  assign n4078 = ( ~x29 & n4071 ) | ( ~x29 & n4077 ) | ( n4071 & n4077 ) ;
  assign n4079 = ( ~n4073 & n4076 ) | ( ~n4073 & n4078 ) | ( n4076 & n4078 ) ;
  assign n4080 = n3831 | n4079 ;
  assign n4081 = n3831 & n4079 ;
  assign n4082 = n4080 & ~n4081 ;
  assign n4083 = n293 & n3088 ;
  assign n4084 = x69 & n3085 ;
  assign n4085 = x68 & n3080 ;
  assign n4086 = x67 & ~n3079 ;
  assign n4087 = n3309 & n4086 ;
  assign n4088 = n4085 | n4087 ;
  assign n4089 = n4084 | n4088 ;
  assign n4090 = n4083 | n4089 ;
  assign n4091 = x26 | n4084 ;
  assign n4092 = n4088 | n4091 ;
  assign n4093 = n4083 | n4092 ;
  assign n4094 = ~x26 & n4092 ;
  assign n4095 = ( ~x26 & n4083 ) | ( ~x26 & n4094 ) | ( n4083 & n4094 ) ;
  assign n4096 = ( ~n4090 & n4093 ) | ( ~n4090 & n4095 ) | ( n4093 & n4095 ) ;
  assign n4097 = n4082 | n4096 ;
  assign n4098 = n4082 & n4096 ;
  assign n4099 = n4097 & ~n4098 ;
  assign n4100 = ( n3837 & n3851 ) | ( n3837 & n3855 ) | ( n3851 & n3855 ) ;
  assign n4101 = n4098 | n4100 ;
  assign n4102 = ( n4098 & n4099 ) | ( n4098 & n4101 ) | ( n4099 & n4101 ) ;
  assign n4103 = n4097 & ~n4102 ;
  assign n4104 = x72 & n2429 ;
  assign n4105 = x71 & n2424 ;
  assign n4106 = x70 & ~n2423 ;
  assign n4107 = n2631 & n4106 ;
  assign n4108 = n4105 | n4107 ;
  assign n4109 = n4104 | n4108 ;
  assign n4110 = ( n513 & n2432 ) | ( n513 & n4109 ) | ( n2432 & n4109 ) ;
  assign n4111 = ( x23 & n2432 ) | ( x23 & ~n4104 ) | ( n2432 & ~n4104 ) ;
  assign n4112 = x23 & n2432 ;
  assign n4113 = ( ~n4108 & n4111 ) | ( ~n4108 & n4112 ) | ( n4111 & n4112 ) ;
  assign n4114 = ( x23 & n513 ) | ( x23 & n4113 ) | ( n513 & n4113 ) ;
  assign n4115 = ~n4110 & n4114 ;
  assign n4116 = n4109 | n4113 ;
  assign n4117 = x23 | n4109 ;
  assign n4118 = ( n513 & n4116 ) | ( n513 & n4117 ) | ( n4116 & n4117 ) ;
  assign n4119 = ( ~x23 & n4115 ) | ( ~x23 & n4118 ) | ( n4115 & n4118 ) ;
  assign n4120 = n4100 & n4119 ;
  assign n4121 = ~n4099 & n4120 ;
  assign n4122 = ( n4103 & n4119 ) | ( n4103 & n4121 ) | ( n4119 & n4121 ) ;
  assign n4123 = n4100 | n4119 ;
  assign n4124 = ( ~n4099 & n4119 ) | ( ~n4099 & n4123 ) | ( n4119 & n4123 ) ;
  assign n4125 = n4103 | n4124 ;
  assign n4126 = ~n4122 & n4125 ;
  assign n4127 = n3859 | n3861 ;
  assign n4128 = ( n3859 & n3864 ) | ( n3859 & n4127 ) | ( n3864 & n4127 ) ;
  assign n4129 = n4126 & n4128 ;
  assign n4130 = n4126 | n4128 ;
  assign n4131 = ~n4129 & n4130 ;
  assign n4132 = x75 & n1859 ;
  assign n4133 = x74 & n1854 ;
  assign n4134 = x73 & ~n1853 ;
  assign n4135 = n2037 & n4134 ;
  assign n4136 = n4133 | n4135 ;
  assign n4137 = n4132 | n4136 ;
  assign n4138 = n1862 | n4132 ;
  assign n4139 = n4136 | n4138 ;
  assign n4140 = ( n746 & n4137 ) | ( n746 & n4139 ) | ( n4137 & n4139 ) ;
  assign n4141 = x20 & n4139 ;
  assign n4142 = x20 & n4132 ;
  assign n4143 = ( x20 & n4136 ) | ( x20 & n4142 ) | ( n4136 & n4142 ) ;
  assign n4144 = ( n746 & n4141 ) | ( n746 & n4143 ) | ( n4141 & n4143 ) ;
  assign n4145 = x20 & ~n4143 ;
  assign n4146 = x20 & ~n4139 ;
  assign n4147 = ( ~n746 & n4145 ) | ( ~n746 & n4146 ) | ( n4145 & n4146 ) ;
  assign n4148 = ( n4140 & ~n4144 ) | ( n4140 & n4147 ) | ( ~n4144 & n4147 ) ;
  assign n4149 = n4131 | n4148 ;
  assign n4150 = n4131 & n4148 ;
  assign n4151 = n4149 & ~n4150 ;
  assign n4152 = n3885 | n3889 ;
  assign n4153 = ( n3885 & n3888 ) | ( n3885 & n4152 ) | ( n3888 & n4152 ) ;
  assign n4154 = n4151 & n4153 ;
  assign n4155 = n4151 | n4153 ;
  assign n4156 = ~n4154 & n4155 ;
  assign n4157 = x78 & n1383 ;
  assign n4158 = x77 & n1378 ;
  assign n4159 = x76 & ~n1377 ;
  assign n4160 = n1542 & n4159 ;
  assign n4161 = n4158 | n4160 ;
  assign n4162 = n4157 | n4161 ;
  assign n4163 = n1386 | n4157 ;
  assign n4164 = n4161 | n4163 ;
  assign n4165 = ( n1192 & n4162 ) | ( n1192 & n4164 ) | ( n4162 & n4164 ) ;
  assign n4166 = x17 & n4164 ;
  assign n4167 = x17 & n4157 ;
  assign n4168 = ( x17 & n4161 ) | ( x17 & n4167 ) | ( n4161 & n4167 ) ;
  assign n4169 = ( n1192 & n4166 ) | ( n1192 & n4168 ) | ( n4166 & n4168 ) ;
  assign n4170 = x17 & ~n4168 ;
  assign n4171 = x17 & ~n4164 ;
  assign n4172 = ( ~n1192 & n4170 ) | ( ~n1192 & n4171 ) | ( n4170 & n4171 ) ;
  assign n4173 = ( n4165 & ~n4169 ) | ( n4165 & n4172 ) | ( ~n4169 & n4172 ) ;
  assign n4174 = n4156 & n4173 ;
  assign n4175 = n4156 & ~n4174 ;
  assign n4176 = ~n4156 & n4173 ;
  assign n4177 = n4175 | n4176 ;
  assign n4178 = n3912 & n3914 ;
  assign n4179 = ( n3911 & n3914 ) | ( n3911 & n4178 ) | ( n3914 & n4178 ) ;
  assign n4180 = n3910 | n4179 ;
  assign n4181 = n4177 | n4180 ;
  assign n4182 = n4177 & n4180 ;
  assign n4183 = n4181 & ~n4182 ;
  assign n4184 = x81 & n962 ;
  assign n4185 = x80 & n957 ;
  assign n4186 = x79 & ~n956 ;
  assign n4187 = n1105 & n4186 ;
  assign n4188 = n4185 | n4187 ;
  assign n4189 = n4184 | n4188 ;
  assign n4190 = n965 | n4184 ;
  assign n4191 = n4188 | n4190 ;
  assign n4192 = ( n1651 & n4189 ) | ( n1651 & n4191 ) | ( n4189 & n4191 ) ;
  assign n4193 = x14 & n4191 ;
  assign n4194 = x14 & n4184 ;
  assign n4195 = ( x14 & n4188 ) | ( x14 & n4194 ) | ( n4188 & n4194 ) ;
  assign n4196 = ( n1651 & n4193 ) | ( n1651 & n4195 ) | ( n4193 & n4195 ) ;
  assign n4197 = x14 & ~n4195 ;
  assign n4198 = x14 & ~n4191 ;
  assign n4199 = ( ~n1651 & n4197 ) | ( ~n1651 & n4198 ) | ( n4197 & n4198 ) ;
  assign n4200 = ( n4192 & ~n4196 ) | ( n4192 & n4199 ) | ( ~n4196 & n4199 ) ;
  assign n4201 = n4183 & n4200 ;
  assign n4202 = n4183 & ~n4201 ;
  assign n4203 = ~n4183 & n4200 ;
  assign n4204 = n4202 | n4203 ;
  assign n4205 = n3937 | n3942 ;
  assign n4206 = n4204 | n4205 ;
  assign n4207 = n4204 & n4205 ;
  assign n4208 = n4206 & ~n4207 ;
  assign n4209 = x84 & n636 ;
  assign n4210 = x83 & n631 ;
  assign n4211 = x82 & ~n630 ;
  assign n4212 = n764 & n4211 ;
  assign n4213 = n4210 | n4212 ;
  assign n4214 = n4209 | n4213 ;
  assign n4215 = n639 | n4209 ;
  assign n4216 = n4213 | n4215 ;
  assign n4217 = ( n2194 & n4214 ) | ( n2194 & n4216 ) | ( n4214 & n4216 ) ;
  assign n4218 = x11 & n4216 ;
  assign n4219 = x11 & n4209 ;
  assign n4220 = ( x11 & n4213 ) | ( x11 & n4219 ) | ( n4213 & n4219 ) ;
  assign n4221 = ( n2194 & n4218 ) | ( n2194 & n4220 ) | ( n4218 & n4220 ) ;
  assign n4222 = x11 & ~n4220 ;
  assign n4223 = x11 & ~n4216 ;
  assign n4224 = ( ~n2194 & n4222 ) | ( ~n2194 & n4223 ) | ( n4222 & n4223 ) ;
  assign n4225 = ( n4217 & ~n4221 ) | ( n4217 & n4224 ) | ( ~n4221 & n4224 ) ;
  assign n4226 = n4208 | n4225 ;
  assign n4227 = n4208 & n4225 ;
  assign n4228 = n4226 & ~n4227 ;
  assign n4229 = n3961 | n3969 ;
  assign n4230 = ~n4228 & n4229 ;
  assign n4231 = n4228 & n4229 ;
  assign n4232 = n4228 & ~n4231 ;
  assign n4233 = n4230 | n4232 ;
  assign n4234 = x87 & n389 ;
  assign n4235 = x86 & n384 ;
  assign n4236 = x85 & ~n383 ;
  assign n4237 = n463 & n4236 ;
  assign n4238 = n4235 | n4237 ;
  assign n4239 = n4234 | n4238 ;
  assign n4240 = n392 | n4234 ;
  assign n4241 = n4238 | n4240 ;
  assign n4242 = ( n2816 & n4239 ) | ( n2816 & n4241 ) | ( n4239 & n4241 ) ;
  assign n4243 = x8 & n4241 ;
  assign n4244 = x8 & n4234 ;
  assign n4245 = ( x8 & n4238 ) | ( x8 & n4244 ) | ( n4238 & n4244 ) ;
  assign n4246 = ( n2816 & n4243 ) | ( n2816 & n4245 ) | ( n4243 & n4245 ) ;
  assign n4247 = x8 & ~n4245 ;
  assign n4248 = x8 & ~n4241 ;
  assign n4249 = ( ~n2816 & n4247 ) | ( ~n2816 & n4248 ) | ( n4247 & n4248 ) ;
  assign n4250 = ( n4242 & ~n4246 ) | ( n4242 & n4249 ) | ( ~n4246 & n4249 ) ;
  assign n4251 = n4230 & n4250 ;
  assign n4252 = ( n4232 & n4250 ) | ( n4232 & n4251 ) | ( n4250 & n4251 ) ;
  assign n4253 = n4233 & ~n4252 ;
  assign n4254 = ~n4230 & n4250 ;
  assign n4255 = ~n4232 & n4254 ;
  assign n4256 = n4253 | n4255 ;
  assign n4257 = n3989 | n3990 ;
  assign n4258 = ( n3989 & n3992 ) | ( n3989 & n4257 ) | ( n3992 & n4257 ) ;
  assign n4259 = n4256 & n4258 ;
  assign n4260 = n4256 | n4258 ;
  assign n4261 = ~n4259 & n4260 ;
  assign n4262 = x90 & n212 ;
  assign n4263 = x89 & n207 ;
  assign n4264 = x88 & ~n206 ;
  assign n4265 = n267 & n4264 ;
  assign n4266 = n4263 | n4265 ;
  assign n4267 = n4262 | n4266 ;
  assign n4268 = n215 | n4262 ;
  assign n4269 = n4266 | n4268 ;
  assign n4270 = ( n3519 & n4267 ) | ( n3519 & n4269 ) | ( n4267 & n4269 ) ;
  assign n4271 = x5 & n4269 ;
  assign n4272 = x5 & n4262 ;
  assign n4273 = ( x5 & n4266 ) | ( x5 & n4272 ) | ( n4266 & n4272 ) ;
  assign n4274 = ( n3519 & n4271 ) | ( n3519 & n4273 ) | ( n4271 & n4273 ) ;
  assign n4275 = x5 & ~n4273 ;
  assign n4276 = x5 & ~n4269 ;
  assign n4277 = ( ~n3519 & n4275 ) | ( ~n3519 & n4276 ) | ( n4275 & n4276 ) ;
  assign n4278 = ( n4270 & ~n4274 ) | ( n4270 & n4277 ) | ( ~n4274 & n4277 ) ;
  assign n4279 = n4261 & n4278 ;
  assign n4280 = n4261 & ~n4279 ;
  assign n4281 = ~n4261 & n4278 ;
  assign n4282 = n4280 | n4281 ;
  assign n4283 = n4013 | n4019 ;
  assign n4284 = ~n4282 & n4283 ;
  assign n4285 = n4282 & ~n4283 ;
  assign n4286 = n4284 | n4285 ;
  assign n4287 = x92 | x93 ;
  assign n4288 = x92 & x93 ;
  assign n4289 = n4287 & ~n4288 ;
  assign n4290 = n4022 & n4289 ;
  assign n4291 = ( n4029 & n4289 ) | ( n4029 & n4290 ) | ( n4289 & n4290 ) ;
  assign n4292 = n4022 | n4023 ;
  assign n4293 = n4289 & n4292 ;
  assign n4294 = ( n4025 & n4290 ) | ( n4025 & n4293 ) | ( n4290 & n4293 ) ;
  assign n4295 = ( n3274 & n4291 ) | ( n3274 & n4294 ) | ( n4291 & n4294 ) ;
  assign n4296 = ( n3276 & n4291 ) | ( n3276 & n4294 ) | ( n4291 & n4294 ) ;
  assign n4297 = ( n1493 & n4295 ) | ( n1493 & n4296 ) | ( n4295 & n4296 ) ;
  assign n4298 = n4022 | n4289 ;
  assign n4299 = n4029 | n4298 ;
  assign n4300 = n4289 | n4292 ;
  assign n4301 = ( n4025 & n4298 ) | ( n4025 & n4300 ) | ( n4298 & n4300 ) ;
  assign n4302 = ( n3274 & n4299 ) | ( n3274 & n4301 ) | ( n4299 & n4301 ) ;
  assign n4303 = ( n3276 & n4299 ) | ( n3276 & n4301 ) | ( n4299 & n4301 ) ;
  assign n4304 = ( n1493 & n4302 ) | ( n1493 & n4303 ) | ( n4302 & n4303 ) ;
  assign n4305 = ~n4297 & n4304 ;
  assign n4306 = x92 & n133 ;
  assign n4307 = x91 & ~n162 ;
  assign n4308 = ( n137 & n4306 ) | ( n137 & n4307 ) | ( n4306 & n4307 ) ;
  assign n4309 = x0 & x93 ;
  assign n4310 = ( ~n137 & n4306 ) | ( ~n137 & n4309 ) | ( n4306 & n4309 ) ;
  assign n4311 = n4308 | n4310 ;
  assign n4312 = n141 | n4311 ;
  assign n4313 = ( n4305 & n4311 ) | ( n4305 & n4312 ) | ( n4311 & n4312 ) ;
  assign n4314 = x2 & n4311 ;
  assign n4315 = ( x2 & n523 ) | ( x2 & n4311 ) | ( n523 & n4311 ) ;
  assign n4316 = ( n4305 & n4314 ) | ( n4305 & n4315 ) | ( n4314 & n4315 ) ;
  assign n4317 = x2 & ~n4315 ;
  assign n4318 = x2 & ~n4311 ;
  assign n4319 = ( ~n4305 & n4317 ) | ( ~n4305 & n4318 ) | ( n4317 & n4318 ) ;
  assign n4320 = ( n4313 & ~n4316 ) | ( n4313 & n4319 ) | ( ~n4316 & n4319 ) ;
  assign n4321 = n4286 & n4320 ;
  assign n4322 = n4286 | n4320 ;
  assign n4323 = ~n4321 & n4322 ;
  assign n4324 = n4064 & n4323 ;
  assign n4325 = n4064 | n4323 ;
  assign n4326 = ~n4324 & n4325 ;
  assign n4327 = n4227 | n4231 ;
  assign n4328 = x29 & ~x30 ;
  assign n4329 = ~x29 & x30 ;
  assign n4330 = n4328 | n4329 ;
  assign n4331 = x64 & n4330 ;
  assign n4332 = ~n3831 & n4331 ;
  assign n4333 = ( ~n4079 & n4331 ) | ( ~n4079 & n4332 ) | ( n4331 & n4332 ) ;
  assign n4334 = n3831 & ~n4331 ;
  assign n4335 = n4079 & n4334 ;
  assign n4336 = n4333 | n4335 ;
  assign n4337 = x67 & n3816 ;
  assign n4338 = x66 & n3811 ;
  assign n4339 = x65 & ~n3810 ;
  assign n4340 = n4067 & n4339 ;
  assign n4341 = n4338 | n4340 ;
  assign n4342 = n4337 | n4341 ;
  assign n4343 = n186 & n3819 ;
  assign n4344 = n4342 | n4343 ;
  assign n4345 = x29 & ~n4344 ;
  assign n4346 = ~x29 & n4344 ;
  assign n4347 = n4345 | n4346 ;
  assign n4348 = n4336 & n4347 ;
  assign n4349 = n4336 | n4347 ;
  assign n4350 = ~n4348 & n4349 ;
  assign n4351 = x69 & n3080 ;
  assign n4352 = x68 & ~n3079 ;
  assign n4353 = n3309 & n4352 ;
  assign n4354 = n4351 | n4353 ;
  assign n4355 = x70 & n3085 ;
  assign n4356 = n3088 | n4355 ;
  assign n4357 = n4354 | n4356 ;
  assign n4358 = x26 & ~n4357 ;
  assign n4359 = x26 & ~n4355 ;
  assign n4360 = ~n4354 & n4359 ;
  assign n4361 = ( ~n340 & n4358 ) | ( ~n340 & n4360 ) | ( n4358 & n4360 ) ;
  assign n4362 = ~x26 & n4357 ;
  assign n4363 = ~x26 & n4355 ;
  assign n4364 = ( ~x26 & n4354 ) | ( ~x26 & n4363 ) | ( n4354 & n4363 ) ;
  assign n4365 = ( n340 & n4362 ) | ( n340 & n4364 ) | ( n4362 & n4364 ) ;
  assign n4366 = n4361 | n4365 ;
  assign n4367 = ( n4102 & ~n4350 ) | ( n4102 & n4366 ) | ( ~n4350 & n4366 ) ;
  assign n4368 = ( ~n4102 & n4350 ) | ( ~n4102 & n4367 ) | ( n4350 & n4367 ) ;
  assign n4369 = x73 & n2429 ;
  assign n4370 = x72 & n2424 ;
  assign n4371 = x71 & ~n2423 ;
  assign n4372 = n2631 & n4371 ;
  assign n4373 = n4370 | n4372 ;
  assign n4374 = n4369 | n4373 ;
  assign n4375 = ( ~n610 & n2432 ) | ( ~n610 & n4374 ) | ( n2432 & n4374 ) ;
  assign n4376 = n2432 & n4369 ;
  assign n4377 = ( n2432 & n4373 ) | ( n2432 & n4376 ) | ( n4373 & n4376 ) ;
  assign n4378 = ( n598 & n4375 ) | ( n598 & n4377 ) | ( n4375 & n4377 ) ;
  assign n4379 = ( x23 & ~n4374 ) | ( x23 & n4378 ) | ( ~n4374 & n4378 ) ;
  assign n4380 = ~n4378 & n4379 ;
  assign n4381 = x23 | n4369 ;
  assign n4382 = n4373 | n4381 ;
  assign n4383 = n4378 | n4382 ;
  assign n4384 = ( ~x23 & n4380 ) | ( ~x23 & n4383 ) | ( n4380 & n4383 ) ;
  assign n4385 = ~n4350 & n4384 ;
  assign n4386 = n4366 & n4384 ;
  assign n4387 = ( n4102 & n4385 ) | ( n4102 & n4386 ) | ( n4385 & n4386 ) ;
  assign n4388 = ~n4366 & n4383 ;
  assign n4389 = x23 | n4366 ;
  assign n4390 = ( n4380 & n4388 ) | ( n4380 & ~n4389 ) | ( n4388 & ~n4389 ) ;
  assign n4391 = ( n4368 & n4387 ) | ( n4368 & n4390 ) | ( n4387 & n4390 ) ;
  assign n4392 = n4350 & ~n4384 ;
  assign n4393 = n4366 | n4384 ;
  assign n4394 = ( n4102 & ~n4392 ) | ( n4102 & n4393 ) | ( ~n4392 & n4393 ) ;
  assign n4395 = n4366 & ~n4383 ;
  assign n4396 = x23 & n4366 ;
  assign n4397 = ( ~n4380 & n4395 ) | ( ~n4380 & n4396 ) | ( n4395 & n4396 ) ;
  assign n4398 = ( n4368 & n4394 ) | ( n4368 & ~n4397 ) | ( n4394 & ~n4397 ) ;
  assign n4399 = ~n4391 & n4398 ;
  assign n4400 = n4122 | n4126 ;
  assign n4401 = ( n4122 & n4128 ) | ( n4122 & n4400 ) | ( n4128 & n4400 ) ;
  assign n4402 = n4399 & n4401 ;
  assign n4403 = n4399 | n4401 ;
  assign n4404 = ~n4402 & n4403 ;
  assign n4405 = x76 & n1859 ;
  assign n4406 = x75 & n1854 ;
  assign n4407 = x74 & ~n1853 ;
  assign n4408 = n2037 & n4407 ;
  assign n4409 = n4406 | n4408 ;
  assign n4410 = n4405 | n4409 ;
  assign n4411 = n1862 | n4405 ;
  assign n4412 = n4409 | n4411 ;
  assign n4413 = ( n923 & n4410 ) | ( n923 & n4412 ) | ( n4410 & n4412 ) ;
  assign n4414 = x20 & n4412 ;
  assign n4415 = x20 & n4405 ;
  assign n4416 = ( x20 & n4409 ) | ( x20 & n4415 ) | ( n4409 & n4415 ) ;
  assign n4417 = ( n923 & n4414 ) | ( n923 & n4416 ) | ( n4414 & n4416 ) ;
  assign n4418 = x20 & ~n4416 ;
  assign n4419 = x20 & ~n4412 ;
  assign n4420 = ( ~n923 & n4418 ) | ( ~n923 & n4419 ) | ( n4418 & n4419 ) ;
  assign n4421 = ( n4413 & ~n4417 ) | ( n4413 & n4420 ) | ( ~n4417 & n4420 ) ;
  assign n4422 = n4404 | n4421 ;
  assign n4423 = n4404 & n4421 ;
  assign n4424 = n4422 & ~n4423 ;
  assign n4425 = n4150 | n4151 ;
  assign n4426 = ( n4150 & n4153 ) | ( n4150 & n4425 ) | ( n4153 & n4425 ) ;
  assign n4427 = n4424 & n4426 ;
  assign n4428 = n4424 | n4426 ;
  assign n4429 = ~n4427 & n4428 ;
  assign n4430 = x79 & n1383 ;
  assign n4431 = x78 & n1378 ;
  assign n4432 = x77 & ~n1377 ;
  assign n4433 = n1542 & n4432 ;
  assign n4434 = n4431 | n4433 ;
  assign n4435 = n4430 | n4434 ;
  assign n4436 = n1386 | n4430 ;
  assign n4437 = n4434 | n4436 ;
  assign n4438 = ( n1332 & n4435 ) | ( n1332 & n4437 ) | ( n4435 & n4437 ) ;
  assign n4439 = x17 & n4437 ;
  assign n4440 = x17 & n4430 ;
  assign n4441 = ( x17 & n4434 ) | ( x17 & n4440 ) | ( n4434 & n4440 ) ;
  assign n4442 = ( n1332 & n4439 ) | ( n1332 & n4441 ) | ( n4439 & n4441 ) ;
  assign n4443 = x17 & ~n4441 ;
  assign n4444 = x17 & ~n4437 ;
  assign n4445 = ( ~n1332 & n4443 ) | ( ~n1332 & n4444 ) | ( n4443 & n4444 ) ;
  assign n4446 = ( n4438 & ~n4442 ) | ( n4438 & n4445 ) | ( ~n4442 & n4445 ) ;
  assign n4447 = n4429 & n4446 ;
  assign n4448 = n4429 & ~n4447 ;
  assign n4449 = ~n4429 & n4446 ;
  assign n4450 = n4448 | n4449 ;
  assign n4451 = n4174 | n4182 ;
  assign n4452 = n4450 | n4451 ;
  assign n4453 = n4450 & n4451 ;
  assign n4454 = n4452 & ~n4453 ;
  assign n4455 = x82 & n962 ;
  assign n4456 = x81 & n957 ;
  assign n4457 = x80 & ~n956 ;
  assign n4458 = n1105 & n4457 ;
  assign n4459 = n4456 | n4458 ;
  assign n4460 = n4455 | n4459 ;
  assign n4461 = n965 | n4455 ;
  assign n4462 = n4459 | n4461 ;
  assign n4463 = ( n1811 & n4460 ) | ( n1811 & n4462 ) | ( n4460 & n4462 ) ;
  assign n4464 = x14 & n4462 ;
  assign n4465 = x14 & n4455 ;
  assign n4466 = ( x14 & n4459 ) | ( x14 & n4465 ) | ( n4459 & n4465 ) ;
  assign n4467 = ( n1811 & n4464 ) | ( n1811 & n4466 ) | ( n4464 & n4466 ) ;
  assign n4468 = x14 & ~n4466 ;
  assign n4469 = x14 & ~n4462 ;
  assign n4470 = ( ~n1811 & n4468 ) | ( ~n1811 & n4469 ) | ( n4468 & n4469 ) ;
  assign n4471 = ( n4463 & ~n4467 ) | ( n4463 & n4470 ) | ( ~n4467 & n4470 ) ;
  assign n4472 = n4454 & n4471 ;
  assign n4473 = n4454 & ~n4472 ;
  assign n4474 = ~n4454 & n4471 ;
  assign n4475 = n4473 | n4474 ;
  assign n4476 = n4201 | n4205 ;
  assign n4477 = ( n4201 & n4204 ) | ( n4201 & n4476 ) | ( n4204 & n4476 ) ;
  assign n4478 = n4475 | n4477 ;
  assign n4479 = n4475 & n4477 ;
  assign n4480 = n4478 & ~n4479 ;
  assign n4481 = x85 & n636 ;
  assign n4482 = x84 & n631 ;
  assign n4483 = x83 & ~n630 ;
  assign n4484 = n764 & n4483 ;
  assign n4485 = n4482 | n4484 ;
  assign n4486 = n4481 | n4485 ;
  assign n4487 = n639 | n4481 ;
  assign n4488 = n4485 | n4487 ;
  assign n4489 = ( n2381 & n4486 ) | ( n2381 & n4488 ) | ( n4486 & n4488 ) ;
  assign n4490 = x11 & n4488 ;
  assign n4491 = x11 & n4481 ;
  assign n4492 = ( x11 & n4485 ) | ( x11 & n4491 ) | ( n4485 & n4491 ) ;
  assign n4493 = ( n2381 & n4490 ) | ( n2381 & n4492 ) | ( n4490 & n4492 ) ;
  assign n4494 = x11 & ~n4492 ;
  assign n4495 = x11 & ~n4488 ;
  assign n4496 = ( ~n2381 & n4494 ) | ( ~n2381 & n4495 ) | ( n4494 & n4495 ) ;
  assign n4497 = ( n4489 & ~n4493 ) | ( n4489 & n4496 ) | ( ~n4493 & n4496 ) ;
  assign n4498 = n4480 & n4497 ;
  assign n4499 = n4480 & ~n4498 ;
  assign n4500 = ~n4480 & n4497 ;
  assign n4501 = n4499 | n4500 ;
  assign n4502 = n4327 & ~n4501 ;
  assign n4503 = ~n4327 & n4501 ;
  assign n4504 = n4502 | n4503 ;
  assign n4505 = x88 & n389 ;
  assign n4506 = x87 & n384 ;
  assign n4507 = x86 & ~n383 ;
  assign n4508 = n463 & n4507 ;
  assign n4509 = n4506 | n4508 ;
  assign n4510 = n4505 | n4509 ;
  assign n4511 = n392 | n4505 ;
  assign n4512 = n4509 | n4511 ;
  assign n4513 = ( ~n3039 & n4510 ) | ( ~n3039 & n4512 ) | ( n4510 & n4512 ) ;
  assign n4514 = n4510 & n4512 ;
  assign n4515 = ( n3023 & n4513 ) | ( n3023 & n4514 ) | ( n4513 & n4514 ) ;
  assign n4516 = x8 & n4512 ;
  assign n4517 = x8 & n4505 ;
  assign n4518 = ( x8 & n4509 ) | ( x8 & n4517 ) | ( n4509 & n4517 ) ;
  assign n4519 = ( ~n3039 & n4516 ) | ( ~n3039 & n4518 ) | ( n4516 & n4518 ) ;
  assign n4520 = n4516 & n4518 ;
  assign n4521 = ( n3023 & n4519 ) | ( n3023 & n4520 ) | ( n4519 & n4520 ) ;
  assign n4522 = x8 & ~n4518 ;
  assign n4523 = x8 & ~n4512 ;
  assign n4524 = ( n3039 & n4522 ) | ( n3039 & n4523 ) | ( n4522 & n4523 ) ;
  assign n4525 = n4522 | n4523 ;
  assign n4526 = ( ~n3023 & n4524 ) | ( ~n3023 & n4525 ) | ( n4524 & n4525 ) ;
  assign n4527 = ( n4515 & ~n4521 ) | ( n4515 & n4526 ) | ( ~n4521 & n4526 ) ;
  assign n4528 = n4504 & n4527 ;
  assign n4529 = n4504 | n4527 ;
  assign n4530 = ~n4528 & n4529 ;
  assign n4531 = n4252 | n4258 ;
  assign n4532 = ( n4252 & n4256 ) | ( n4252 & n4531 ) | ( n4256 & n4531 ) ;
  assign n4533 = n4530 | n4532 ;
  assign n4534 = n4530 & n4532 ;
  assign n4535 = n4533 & ~n4534 ;
  assign n4536 = x91 & n212 ;
  assign n4537 = x90 & n207 ;
  assign n4538 = x89 & ~n206 ;
  assign n4539 = n267 & n4538 ;
  assign n4540 = n4537 | n4539 ;
  assign n4541 = n4536 | n4540 ;
  assign n4542 = n215 | n4536 ;
  assign n4543 = n4540 | n4542 ;
  assign n4544 = ( n3768 & n4541 ) | ( n3768 & n4543 ) | ( n4541 & n4543 ) ;
  assign n4545 = x5 & n4543 ;
  assign n4546 = x5 & n4536 ;
  assign n4547 = ( x5 & n4540 ) | ( x5 & n4546 ) | ( n4540 & n4546 ) ;
  assign n4548 = ( n3768 & n4545 ) | ( n3768 & n4547 ) | ( n4545 & n4547 ) ;
  assign n4549 = x5 & ~n4547 ;
  assign n4550 = x5 & ~n4543 ;
  assign n4551 = ( ~n3768 & n4549 ) | ( ~n3768 & n4550 ) | ( n4549 & n4550 ) ;
  assign n4552 = ( n4544 & ~n4548 ) | ( n4544 & n4551 ) | ( ~n4548 & n4551 ) ;
  assign n4553 = n4535 & n4552 ;
  assign n4554 = n4535 & ~n4553 ;
  assign n4555 = ~n4535 & n4552 ;
  assign n4556 = n4554 | n4555 ;
  assign n4557 = n4282 & n4283 ;
  assign n4558 = n4279 | n4557 ;
  assign n4559 = n4556 | n4558 ;
  assign n4560 = n4556 & n4558 ;
  assign n4561 = n4559 & ~n4560 ;
  assign n4562 = x93 | x94 ;
  assign n4563 = x93 & x94 ;
  assign n4564 = n4562 & ~n4563 ;
  assign n4565 = n4288 | n4290 ;
  assign n4566 = n4564 & n4565 ;
  assign n4567 = n4288 | n4289 ;
  assign n4568 = n4564 & n4567 ;
  assign n4569 = ( n4029 & n4566 ) | ( n4029 & n4568 ) | ( n4566 & n4568 ) ;
  assign n4570 = n4288 & n4564 ;
  assign n4571 = ( n4294 & n4564 ) | ( n4294 & n4570 ) | ( n4564 & n4570 ) ;
  assign n4572 = ( n3274 & n4569 ) | ( n3274 & n4571 ) | ( n4569 & n4571 ) ;
  assign n4573 = ( n3276 & n4569 ) | ( n3276 & n4571 ) | ( n4569 & n4571 ) ;
  assign n4574 = ( n1493 & n4572 ) | ( n1493 & n4573 ) | ( n4572 & n4573 ) ;
  assign n4575 = n4564 | n4565 ;
  assign n4576 = n4564 | n4567 ;
  assign n4577 = ( n4029 & n4575 ) | ( n4029 & n4576 ) | ( n4575 & n4576 ) ;
  assign n4578 = n4288 | n4564 ;
  assign n4579 = n4294 | n4578 ;
  assign n4580 = ( n3274 & n4577 ) | ( n3274 & n4579 ) | ( n4577 & n4579 ) ;
  assign n4581 = ( n3276 & n4577 ) | ( n3276 & n4579 ) | ( n4577 & n4579 ) ;
  assign n4582 = ( n1493 & n4580 ) | ( n1493 & n4581 ) | ( n4580 & n4581 ) ;
  assign n4583 = ~n4574 & n4582 ;
  assign n4584 = x93 & n133 ;
  assign n4585 = x92 & ~n162 ;
  assign n4586 = ( n137 & n4584 ) | ( n137 & n4585 ) | ( n4584 & n4585 ) ;
  assign n4587 = x0 & x94 ;
  assign n4588 = ( ~n137 & n4584 ) | ( ~n137 & n4587 ) | ( n4584 & n4587 ) ;
  assign n4589 = n4586 | n4588 ;
  assign n4590 = n141 | n4589 ;
  assign n4591 = ( n4583 & n4589 ) | ( n4583 & n4590 ) | ( n4589 & n4590 ) ;
  assign n4592 = x2 & n4589 ;
  assign n4593 = ( x2 & n523 ) | ( x2 & n4589 ) | ( n523 & n4589 ) ;
  assign n4594 = ( n4583 & n4592 ) | ( n4583 & n4593 ) | ( n4592 & n4593 ) ;
  assign n4595 = x2 & ~n4593 ;
  assign n4596 = x2 & ~n4589 ;
  assign n4597 = ( ~n4583 & n4595 ) | ( ~n4583 & n4596 ) | ( n4595 & n4596 ) ;
  assign n4598 = ( n4591 & ~n4594 ) | ( n4591 & n4597 ) | ( ~n4594 & n4597 ) ;
  assign n4599 = n4561 & n4598 ;
  assign n4600 = n4561 & ~n4599 ;
  assign n4601 = ~n4561 & n4598 ;
  assign n4602 = n4600 | n4601 ;
  assign n4603 = n4321 | n4324 ;
  assign n4604 = n4602 & n4603 ;
  assign n4605 = n4602 | n4603 ;
  assign n4606 = ~n4604 & n4605 ;
  assign n4607 = x70 & n3080 ;
  assign n4608 = x69 & ~n3079 ;
  assign n4609 = n3309 & n4608 ;
  assign n4610 = n4607 | n4609 ;
  assign n4611 = x71 & n3085 ;
  assign n4612 = n3088 | n4611 ;
  assign n4613 = n4610 | n4612 ;
  assign n4614 = x26 & ~n4613 ;
  assign n4615 = x26 & ~n4611 ;
  assign n4616 = ~n4610 & n4615 ;
  assign n4617 = ( ~n438 & n4614 ) | ( ~n438 & n4616 ) | ( n4614 & n4616 ) ;
  assign n4618 = ~x26 & n4613 ;
  assign n4619 = ~x26 & n4611 ;
  assign n4620 = ( ~x26 & n4610 ) | ( ~x26 & n4619 ) | ( n4610 & n4619 ) ;
  assign n4621 = ( n438 & n4618 ) | ( n438 & n4620 ) | ( n4618 & n4620 ) ;
  assign n4622 = n4617 | n4621 ;
  assign n4623 = ~x30 & x31 ;
  assign n4624 = x30 & ~x31 ;
  assign n4625 = n4623 | n4624 ;
  assign n4626 = ~n4330 & n4625 ;
  assign n4627 = x64 & n4626 ;
  assign n4628 = ~x31 & x32 ;
  assign n4629 = x31 & ~x32 ;
  assign n4630 = n4628 | n4629 ;
  assign n4631 = n4330 & ~n4630 ;
  assign n4632 = x65 & n4631 ;
  assign n4633 = n4627 | n4632 ;
  assign n4634 = n4330 & n4630 ;
  assign n4635 = x32 | n144 ;
  assign n4636 = ( x32 & n4634 ) | ( x32 & n4635 ) | ( n4634 & n4635 ) ;
  assign n4637 = ~x32 & n4636 ;
  assign n4638 = ( ~x32 & n4633 ) | ( ~x32 & n4637 ) | ( n4633 & n4637 ) ;
  assign n4639 = x32 & ~x64 ;
  assign n4640 = ( x32 & ~n4330 ) | ( x32 & n4639 ) | ( ~n4330 & n4639 ) ;
  assign n4641 = n4636 & n4640 ;
  assign n4642 = ( n4633 & n4640 ) | ( n4633 & n4641 ) | ( n4640 & n4641 ) ;
  assign n4643 = n144 & n4634 ;
  assign n4644 = n4640 & ~n4643 ;
  assign n4645 = ~n4633 & n4644 ;
  assign n4646 = ( n4638 & n4642 ) | ( n4638 & n4645 ) | ( n4642 & n4645 ) ;
  assign n4647 = n4636 | n4640 ;
  assign n4648 = n4633 | n4647 ;
  assign n4649 = ~n4640 & n4643 ;
  assign n4650 = ( n4633 & ~n4640 ) | ( n4633 & n4649 ) | ( ~n4640 & n4649 ) ;
  assign n4651 = ( n4638 & n4648 ) | ( n4638 & ~n4650 ) | ( n4648 & ~n4650 ) ;
  assign n4652 = ~n4646 & n4651 ;
  assign n4653 = n241 & n3819 ;
  assign n4654 = x68 & n3816 ;
  assign n4655 = x67 & n3811 ;
  assign n4656 = x66 & ~n3810 ;
  assign n4657 = n4067 & n4656 ;
  assign n4658 = n4655 | n4657 ;
  assign n4659 = n4654 | n4658 ;
  assign n4660 = n4653 | n4659 ;
  assign n4661 = x29 | n4654 ;
  assign n4662 = n4658 | n4661 ;
  assign n4663 = n4653 | n4662 ;
  assign n4664 = ~x29 & n4662 ;
  assign n4665 = ( ~x29 & n4653 ) | ( ~x29 & n4664 ) | ( n4653 & n4664 ) ;
  assign n4666 = ( ~n4660 & n4663 ) | ( ~n4660 & n4665 ) | ( n4663 & n4665 ) ;
  assign n4667 = n4652 & ~n4666 ;
  assign n4668 = ~n4652 & n4666 ;
  assign n4669 = n4667 | n4668 ;
  assign n4670 = ( n4081 & n4331 ) | ( n4081 & n4347 ) | ( n4331 & n4347 ) ;
  assign n4671 = n4669 | n4670 ;
  assign n4672 = n4669 & n4670 ;
  assign n4673 = n4671 & ~n4672 ;
  assign n4674 = n4622 & n4673 ;
  assign n4675 = n4622 | n4673 ;
  assign n4676 = ~n4674 & n4675 ;
  assign n4677 = n4350 & n4366 ;
  assign n4678 = n4350 & ~n4677 ;
  assign n4679 = ~n4350 & n4366 ;
  assign n4680 = n4102 & ~n4679 ;
  assign n4681 = ~n4678 & n4680 ;
  assign n4682 = ( n4102 & n4677 ) | ( n4102 & ~n4681 ) | ( n4677 & ~n4681 ) ;
  assign n4683 = n4676 & n4682 ;
  assign n4684 = n4676 | n4682 ;
  assign n4685 = ~n4683 & n4684 ;
  assign n4686 = x74 & n2429 ;
  assign n4687 = x73 & n2424 ;
  assign n4688 = x72 & ~n2423 ;
  assign n4689 = n2631 & n4688 ;
  assign n4690 = n4687 | n4689 ;
  assign n4691 = n4686 | n4690 ;
  assign n4692 = n2432 | n4686 ;
  assign n4693 = n4690 | n4692 ;
  assign n4694 = ( n710 & n4691 ) | ( n710 & n4693 ) | ( n4691 & n4693 ) ;
  assign n4695 = x23 & n4693 ;
  assign n4696 = x23 & n4686 ;
  assign n4697 = ( x23 & n4690 ) | ( x23 & n4696 ) | ( n4690 & n4696 ) ;
  assign n4698 = ( n710 & n4695 ) | ( n710 & n4697 ) | ( n4695 & n4697 ) ;
  assign n4699 = x23 & ~n4697 ;
  assign n4700 = x23 & ~n4693 ;
  assign n4701 = ( ~n710 & n4699 ) | ( ~n710 & n4700 ) | ( n4699 & n4700 ) ;
  assign n4702 = ( n4694 & ~n4698 ) | ( n4694 & n4701 ) | ( ~n4698 & n4701 ) ;
  assign n4703 = n4685 & n4702 ;
  assign n4704 = n4685 & ~n4703 ;
  assign n4705 = n4391 | n4399 ;
  assign n4706 = ( n4391 & n4401 ) | ( n4391 & n4705 ) | ( n4401 & n4705 ) ;
  assign n4707 = ~n4685 & n4702 ;
  assign n4708 = n4706 & n4707 ;
  assign n4709 = ( n4704 & n4706 ) | ( n4704 & n4708 ) | ( n4706 & n4708 ) ;
  assign n4710 = n4706 | n4707 ;
  assign n4711 = n4704 | n4710 ;
  assign n4712 = ~n4709 & n4711 ;
  assign n4713 = x77 & n1859 ;
  assign n4714 = x76 & n1854 ;
  assign n4715 = x75 & ~n1853 ;
  assign n4716 = n2037 & n4715 ;
  assign n4717 = n4714 | n4716 ;
  assign n4718 = n4713 | n4717 ;
  assign n4719 = n1862 | n4713 ;
  assign n4720 = n4717 | n4719 ;
  assign n4721 = ( n1059 & n4718 ) | ( n1059 & n4720 ) | ( n4718 & n4720 ) ;
  assign n4722 = x20 & n4720 ;
  assign n4723 = x20 & n4713 ;
  assign n4724 = ( x20 & n4717 ) | ( x20 & n4723 ) | ( n4717 & n4723 ) ;
  assign n4725 = ( n1059 & n4722 ) | ( n1059 & n4724 ) | ( n4722 & n4724 ) ;
  assign n4726 = x20 & ~n4724 ;
  assign n4727 = x20 & ~n4720 ;
  assign n4728 = ( ~n1059 & n4726 ) | ( ~n1059 & n4727 ) | ( n4726 & n4727 ) ;
  assign n4729 = ( n4721 & ~n4725 ) | ( n4721 & n4728 ) | ( ~n4725 & n4728 ) ;
  assign n4730 = n4712 | n4729 ;
  assign n4731 = n4712 & n4729 ;
  assign n4732 = n4730 & ~n4731 ;
  assign n4733 = n4423 | n4424 ;
  assign n4734 = ( n4423 & n4426 ) | ( n4423 & n4733 ) | ( n4426 & n4733 ) ;
  assign n4735 = n4732 & n4734 ;
  assign n4736 = n4732 | n4734 ;
  assign n4737 = ~n4735 & n4736 ;
  assign n4738 = x80 & n1383 ;
  assign n4739 = x79 & n1378 ;
  assign n4740 = x78 & ~n1377 ;
  assign n4741 = n1542 & n4740 ;
  assign n4742 = n4739 | n4741 ;
  assign n4743 = n4738 | n4742 ;
  assign n4744 = n1386 | n4738 ;
  assign n4745 = n4742 | n4744 ;
  assign n4746 = ( n1499 & n4743 ) | ( n1499 & n4745 ) | ( n4743 & n4745 ) ;
  assign n4747 = x17 & n4745 ;
  assign n4748 = x17 & n4738 ;
  assign n4749 = ( x17 & n4742 ) | ( x17 & n4748 ) | ( n4742 & n4748 ) ;
  assign n4750 = ( n1499 & n4747 ) | ( n1499 & n4749 ) | ( n4747 & n4749 ) ;
  assign n4751 = x17 & ~n4749 ;
  assign n4752 = x17 & ~n4745 ;
  assign n4753 = ( ~n1499 & n4751 ) | ( ~n1499 & n4752 ) | ( n4751 & n4752 ) ;
  assign n4754 = ( n4746 & ~n4750 ) | ( n4746 & n4753 ) | ( ~n4750 & n4753 ) ;
  assign n4755 = n4737 & n4754 ;
  assign n4756 = n4737 & ~n4755 ;
  assign n4757 = ~n4737 & n4754 ;
  assign n4758 = n4756 | n4757 ;
  assign n4759 = n4447 | n4449 ;
  assign n4760 = n4448 | n4759 ;
  assign n4761 = ( n4447 & n4451 ) | ( n4447 & n4760 ) | ( n4451 & n4760 ) ;
  assign n4762 = n4758 | n4761 ;
  assign n4763 = n4758 & n4761 ;
  assign n4764 = n4762 & ~n4763 ;
  assign n4765 = x83 & n962 ;
  assign n4766 = x82 & n957 ;
  assign n4767 = x81 & ~n956 ;
  assign n4768 = n1105 & n4767 ;
  assign n4769 = n4766 | n4768 ;
  assign n4770 = n4765 | n4769 ;
  assign n4771 = n965 | n4765 ;
  assign n4772 = n4769 | n4771 ;
  assign n4773 = ( n2009 & n4770 ) | ( n2009 & n4772 ) | ( n4770 & n4772 ) ;
  assign n4774 = x14 & n4772 ;
  assign n4775 = x14 & n4765 ;
  assign n4776 = ( x14 & n4769 ) | ( x14 & n4775 ) | ( n4769 & n4775 ) ;
  assign n4777 = ( n2009 & n4774 ) | ( n2009 & n4776 ) | ( n4774 & n4776 ) ;
  assign n4778 = x14 & ~n4776 ;
  assign n4779 = x14 & ~n4772 ;
  assign n4780 = ( ~n2009 & n4778 ) | ( ~n2009 & n4779 ) | ( n4778 & n4779 ) ;
  assign n4781 = ( n4773 & ~n4777 ) | ( n4773 & n4780 ) | ( ~n4777 & n4780 ) ;
  assign n4782 = n4764 & n4781 ;
  assign n4783 = n4764 & ~n4782 ;
  assign n4784 = ~n4764 & n4781 ;
  assign n4785 = n4783 | n4784 ;
  assign n4786 = n4472 | n4477 ;
  assign n4787 = ( n4472 & n4475 ) | ( n4472 & n4786 ) | ( n4475 & n4786 ) ;
  assign n4788 = n4785 | n4787 ;
  assign n4789 = n4785 & n4787 ;
  assign n4790 = n4788 & ~n4789 ;
  assign n4791 = x86 & n636 ;
  assign n4792 = x85 & n631 ;
  assign n4793 = x84 & ~n630 ;
  assign n4794 = n764 & n4793 ;
  assign n4795 = n4792 | n4794 ;
  assign n4796 = n4791 | n4795 ;
  assign n4797 = n639 | n4791 ;
  assign n4798 = n4795 | n4797 ;
  assign n4799 = ( n2606 & n4796 ) | ( n2606 & n4798 ) | ( n4796 & n4798 ) ;
  assign n4800 = x11 & n4798 ;
  assign n4801 = x11 & n4791 ;
  assign n4802 = ( x11 & n4795 ) | ( x11 & n4801 ) | ( n4795 & n4801 ) ;
  assign n4803 = ( n2606 & n4800 ) | ( n2606 & n4802 ) | ( n4800 & n4802 ) ;
  assign n4804 = x11 & ~n4802 ;
  assign n4805 = x11 & ~n4798 ;
  assign n4806 = ( ~n2606 & n4804 ) | ( ~n2606 & n4805 ) | ( n4804 & n4805 ) ;
  assign n4807 = ( n4799 & ~n4803 ) | ( n4799 & n4806 ) | ( ~n4803 & n4806 ) ;
  assign n4808 = n4790 & n4807 ;
  assign n4809 = n4790 & ~n4808 ;
  assign n4810 = ( n4227 & n4480 ) | ( n4227 & n4497 ) | ( n4480 & n4497 ) ;
  assign n4811 = n4480 | n4497 ;
  assign n4812 = ( n4231 & n4810 ) | ( n4231 & n4811 ) | ( n4810 & n4811 ) ;
  assign n4813 = ~n4790 & n4807 ;
  assign n4814 = n4812 & n4813 ;
  assign n4815 = ( n4809 & n4812 ) | ( n4809 & n4814 ) | ( n4812 & n4814 ) ;
  assign n4816 = n4812 | n4813 ;
  assign n4817 = n4809 | n4816 ;
  assign n4818 = ~n4815 & n4817 ;
  assign n4819 = x89 & n389 ;
  assign n4820 = x88 & n384 ;
  assign n4821 = x87 & ~n383 ;
  assign n4822 = n463 & n4821 ;
  assign n4823 = n4820 | n4822 ;
  assign n4824 = n4819 | n4823 ;
  assign n4825 = n392 | n4819 ;
  assign n4826 = n4823 | n4825 ;
  assign n4827 = ( n3282 & n4824 ) | ( n3282 & n4826 ) | ( n4824 & n4826 ) ;
  assign n4828 = x8 & n4826 ;
  assign n4829 = x8 & n4819 ;
  assign n4830 = ( x8 & n4823 ) | ( x8 & n4829 ) | ( n4823 & n4829 ) ;
  assign n4831 = ( n3282 & n4828 ) | ( n3282 & n4830 ) | ( n4828 & n4830 ) ;
  assign n4832 = x8 & ~n4830 ;
  assign n4833 = x8 & ~n4826 ;
  assign n4834 = ( ~n3282 & n4832 ) | ( ~n3282 & n4833 ) | ( n4832 & n4833 ) ;
  assign n4835 = ( n4827 & ~n4831 ) | ( n4827 & n4834 ) | ( ~n4831 & n4834 ) ;
  assign n4836 = n4818 & n4835 ;
  assign n4837 = n4818 & ~n4836 ;
  assign n4838 = ~n4818 & n4835 ;
  assign n4839 = n4837 | n4838 ;
  assign n4840 = n4528 | n4532 ;
  assign n4841 = ( n4528 & n4530 ) | ( n4528 & n4840 ) | ( n4530 & n4840 ) ;
  assign n4842 = n4839 | n4841 ;
  assign n4843 = n4839 & n4841 ;
  assign n4844 = n4842 & ~n4843 ;
  assign n4845 = x92 & n212 ;
  assign n4846 = x91 & n207 ;
  assign n4847 = x90 & ~n206 ;
  assign n4848 = n267 & n4847 ;
  assign n4849 = n4846 | n4848 ;
  assign n4850 = n4845 | n4849 ;
  assign n4851 = n215 | n4845 ;
  assign n4852 = n4849 | n4851 ;
  assign n4853 = ( n4040 & n4850 ) | ( n4040 & n4852 ) | ( n4850 & n4852 ) ;
  assign n4854 = x5 & n4852 ;
  assign n4855 = x5 & n4845 ;
  assign n4856 = ( x5 & n4849 ) | ( x5 & n4855 ) | ( n4849 & n4855 ) ;
  assign n4857 = ( n4040 & n4854 ) | ( n4040 & n4856 ) | ( n4854 & n4856 ) ;
  assign n4858 = x5 & ~n4856 ;
  assign n4859 = x5 & ~n4852 ;
  assign n4860 = ( ~n4040 & n4858 ) | ( ~n4040 & n4859 ) | ( n4858 & n4859 ) ;
  assign n4861 = ( n4853 & ~n4857 ) | ( n4853 & n4860 ) | ( ~n4857 & n4860 ) ;
  assign n4862 = n4844 & n4861 ;
  assign n4863 = n4844 & ~n4862 ;
  assign n4864 = ~n4844 & n4861 ;
  assign n4865 = n4863 | n4864 ;
  assign n4866 = n4553 | n4560 ;
  assign n4867 = n4865 | n4866 ;
  assign n4868 = n4865 & n4866 ;
  assign n4869 = n4867 & ~n4868 ;
  assign n4870 = x94 | x95 ;
  assign n4871 = x94 & x95 ;
  assign n4872 = n4870 & ~n4871 ;
  assign n4873 = n4563 | n4564 ;
  assign n4874 = n4872 & n4873 ;
  assign n4875 = n4563 & n4872 ;
  assign n4876 = ( n4565 & n4874 ) | ( n4565 & n4875 ) | ( n4874 & n4875 ) ;
  assign n4877 = ( n4567 & n4874 ) | ( n4567 & n4875 ) | ( n4874 & n4875 ) ;
  assign n4878 = ( n4029 & n4876 ) | ( n4029 & n4877 ) | ( n4876 & n4877 ) ;
  assign n4879 = ( n4288 & n4874 ) | ( n4288 & n4875 ) | ( n4874 & n4875 ) ;
  assign n4880 = n4874 | n4875 ;
  assign n4881 = ( n4294 & n4879 ) | ( n4294 & n4880 ) | ( n4879 & n4880 ) ;
  assign n4882 = ( n3274 & n4878 ) | ( n3274 & n4881 ) | ( n4878 & n4881 ) ;
  assign n4883 = ( n3276 & n4878 ) | ( n3276 & n4881 ) | ( n4878 & n4881 ) ;
  assign n4884 = ( n1493 & n4882 ) | ( n1493 & n4883 ) | ( n4882 & n4883 ) ;
  assign n4885 = ( n4563 & n4565 ) | ( n4563 & n4873 ) | ( n4565 & n4873 ) ;
  assign n4886 = ( n4563 & n4567 ) | ( n4563 & n4873 ) | ( n4567 & n4873 ) ;
  assign n4887 = ( n4029 & n4885 ) | ( n4029 & n4886 ) | ( n4885 & n4886 ) ;
  assign n4888 = n4872 | n4887 ;
  assign n4889 = n4563 | n4873 ;
  assign n4890 = n4872 | n4889 ;
  assign n4891 = ( n4288 & n4563 ) | ( n4288 & n4873 ) | ( n4563 & n4873 ) ;
  assign n4892 = n4872 | n4891 ;
  assign n4893 = ( n4294 & n4890 ) | ( n4294 & n4892 ) | ( n4890 & n4892 ) ;
  assign n4894 = ( n3274 & n4888 ) | ( n3274 & n4893 ) | ( n4888 & n4893 ) ;
  assign n4895 = ( n3276 & n4888 ) | ( n3276 & n4893 ) | ( n4888 & n4893 ) ;
  assign n4896 = ( n1493 & n4894 ) | ( n1493 & n4895 ) | ( n4894 & n4895 ) ;
  assign n4897 = ~n4884 & n4896 ;
  assign n4898 = x94 & n133 ;
  assign n4899 = x93 & ~n162 ;
  assign n4900 = ( n137 & n4898 ) | ( n137 & n4899 ) | ( n4898 & n4899 ) ;
  assign n4901 = x0 & x95 ;
  assign n4902 = ( ~n137 & n4898 ) | ( ~n137 & n4901 ) | ( n4898 & n4901 ) ;
  assign n4903 = n4900 | n4902 ;
  assign n4904 = n141 | n4903 ;
  assign n4905 = ( n4897 & n4903 ) | ( n4897 & n4904 ) | ( n4903 & n4904 ) ;
  assign n4906 = x2 & n4903 ;
  assign n4907 = ( x2 & n523 ) | ( x2 & n4903 ) | ( n523 & n4903 ) ;
  assign n4908 = ( n4897 & n4906 ) | ( n4897 & n4907 ) | ( n4906 & n4907 ) ;
  assign n4909 = x2 & ~n4907 ;
  assign n4910 = x2 & ~n4903 ;
  assign n4911 = ( ~n4897 & n4909 ) | ( ~n4897 & n4910 ) | ( n4909 & n4910 ) ;
  assign n4912 = ( n4905 & ~n4908 ) | ( n4905 & n4911 ) | ( ~n4908 & n4911 ) ;
  assign n4913 = n4869 & n4912 ;
  assign n4914 = n4869 & ~n4913 ;
  assign n4915 = ~n4869 & n4912 ;
  assign n4916 = n4914 | n4915 ;
  assign n4917 = n4599 | n4603 ;
  assign n4918 = ( n4599 & n4602 ) | ( n4599 & n4917 ) | ( n4602 & n4917 ) ;
  assign n4919 = n4916 & n4918 ;
  assign n4920 = n4916 | n4918 ;
  assign n4921 = ~n4919 & n4920 ;
  assign n4922 = x87 & n636 ;
  assign n4923 = x86 & n631 ;
  assign n4924 = x85 & ~n630 ;
  assign n4925 = n764 & n4924 ;
  assign n4926 = n4923 | n4925 ;
  assign n4927 = n4922 | n4926 ;
  assign n4928 = n639 | n4922 ;
  assign n4929 = n4926 | n4928 ;
  assign n4930 = ( n2816 & n4927 ) | ( n2816 & n4929 ) | ( n4927 & n4929 ) ;
  assign n4931 = x11 & n4929 ;
  assign n4932 = x11 & n4922 ;
  assign n4933 = ( x11 & n4926 ) | ( x11 & n4932 ) | ( n4926 & n4932 ) ;
  assign n4934 = ( n2816 & n4931 ) | ( n2816 & n4933 ) | ( n4931 & n4933 ) ;
  assign n4935 = x11 & ~n4933 ;
  assign n4936 = x11 & ~n4929 ;
  assign n4937 = ( ~n2816 & n4935 ) | ( ~n2816 & n4936 ) | ( n4935 & n4936 ) ;
  assign n4938 = ( n4930 & ~n4934 ) | ( n4930 & n4937 ) | ( ~n4934 & n4937 ) ;
  assign n4939 = n4731 | n4735 ;
  assign n4940 = n4703 | n4709 ;
  assign n4941 = x66 & n4631 ;
  assign n4942 = x65 & n4626 ;
  assign n4943 = ~n4330 & n4630 ;
  assign n4944 = x64 & ~n4625 ;
  assign n4945 = n4943 & n4944 ;
  assign n4946 = n4942 | n4945 ;
  assign n4947 = n4941 | n4946 ;
  assign n4948 = n159 & n4634 ;
  assign n4949 = n4947 | n4948 ;
  assign n4950 = x32 | n4634 ;
  assign n4951 = ( x32 & n159 ) | ( x32 & n4950 ) | ( n159 & n4950 ) ;
  assign n4952 = n4947 | n4951 ;
  assign n4953 = ~x32 & n4951 ;
  assign n4954 = ( ~x32 & n4947 ) | ( ~x32 & n4953 ) | ( n4947 & n4953 ) ;
  assign n4955 = ( ~n4949 & n4952 ) | ( ~n4949 & n4954 ) | ( n4952 & n4954 ) ;
  assign n4956 = n4646 | n4955 ;
  assign n4957 = n4646 & n4955 ;
  assign n4958 = n4956 & ~n4957 ;
  assign n4959 = n293 & n3819 ;
  assign n4960 = x69 & n3816 ;
  assign n4961 = x68 & n3811 ;
  assign n4962 = x67 & ~n3810 ;
  assign n4963 = n4067 & n4962 ;
  assign n4964 = n4961 | n4963 ;
  assign n4965 = n4960 | n4964 ;
  assign n4966 = n4959 | n4965 ;
  assign n4967 = x29 | n4960 ;
  assign n4968 = n4964 | n4967 ;
  assign n4969 = n4959 | n4968 ;
  assign n4970 = ~x29 & n4968 ;
  assign n4971 = ( ~x29 & n4959 ) | ( ~x29 & n4970 ) | ( n4959 & n4970 ) ;
  assign n4972 = ( ~n4966 & n4969 ) | ( ~n4966 & n4971 ) | ( n4969 & n4971 ) ;
  assign n4973 = n4958 | n4972 ;
  assign n4974 = n4958 & n4972 ;
  assign n4975 = n4973 & ~n4974 ;
  assign n4976 = ( n4652 & n4666 ) | ( n4652 & n4670 ) | ( n4666 & n4670 ) ;
  assign n4977 = n4974 | n4976 ;
  assign n4978 = ( n4974 & n4975 ) | ( n4974 & n4977 ) | ( n4975 & n4977 ) ;
  assign n4979 = n4973 & ~n4978 ;
  assign n4980 = ~n4975 & n4976 ;
  assign n4981 = n4979 | n4980 ;
  assign n4982 = x72 & n3085 ;
  assign n4983 = x71 & n3080 ;
  assign n4984 = x70 & ~n3079 ;
  assign n4985 = n3309 & n4984 ;
  assign n4986 = n4983 | n4985 ;
  assign n4987 = n4982 | n4986 ;
  assign n4988 = ( n513 & n3088 ) | ( n513 & n4987 ) | ( n3088 & n4987 ) ;
  assign n4989 = ( x26 & n3088 ) | ( x26 & ~n4982 ) | ( n3088 & ~n4982 ) ;
  assign n4990 = x26 & n3088 ;
  assign n4991 = ( ~n4986 & n4989 ) | ( ~n4986 & n4990 ) | ( n4989 & n4990 ) ;
  assign n4992 = ( x26 & n513 ) | ( x26 & n4991 ) | ( n513 & n4991 ) ;
  assign n4993 = ~n4988 & n4992 ;
  assign n4994 = n4987 | n4991 ;
  assign n4995 = x26 | n4987 ;
  assign n4996 = ( n513 & n4994 ) | ( n513 & n4995 ) | ( n4994 & n4995 ) ;
  assign n4997 = ( ~x26 & n4993 ) | ( ~x26 & n4996 ) | ( n4993 & n4996 ) ;
  assign n4998 = n4976 & n4997 ;
  assign n4999 = ~n4975 & n4998 ;
  assign n5000 = ( n4979 & n4997 ) | ( n4979 & n4999 ) | ( n4997 & n4999 ) ;
  assign n5001 = n4981 & ~n5000 ;
  assign n5002 = ~n4976 & n4997 ;
  assign n5003 = ( n4975 & n4997 ) | ( n4975 & n5002 ) | ( n4997 & n5002 ) ;
  assign n5004 = ~n4979 & n5003 ;
  assign n5005 = n5001 | n5004 ;
  assign n5006 = n4674 | n4676 ;
  assign n5007 = ( n4674 & n4682 ) | ( n4674 & n5006 ) | ( n4682 & n5006 ) ;
  assign n5008 = n5005 | n5007 ;
  assign n5009 = n5005 & n5007 ;
  assign n5010 = n5008 & ~n5009 ;
  assign n5011 = x75 & n2429 ;
  assign n5012 = x74 & n2424 ;
  assign n5013 = x73 & ~n2423 ;
  assign n5014 = n2631 & n5013 ;
  assign n5015 = n5012 | n5014 ;
  assign n5016 = n5011 | n5015 ;
  assign n5017 = n2432 | n5011 ;
  assign n5018 = n5015 | n5017 ;
  assign n5019 = ( n746 & n5016 ) | ( n746 & n5018 ) | ( n5016 & n5018 ) ;
  assign n5020 = x23 & n5018 ;
  assign n5021 = x23 & n5011 ;
  assign n5022 = ( x23 & n5015 ) | ( x23 & n5021 ) | ( n5015 & n5021 ) ;
  assign n5023 = ( n746 & n5020 ) | ( n746 & n5022 ) | ( n5020 & n5022 ) ;
  assign n5024 = x23 & ~n5022 ;
  assign n5025 = x23 & ~n5018 ;
  assign n5026 = ( ~n746 & n5024 ) | ( ~n746 & n5025 ) | ( n5024 & n5025 ) ;
  assign n5027 = ( n5019 & ~n5023 ) | ( n5019 & n5026 ) | ( ~n5023 & n5026 ) ;
  assign n5028 = n5010 & n5027 ;
  assign n5029 = n5010 | n5027 ;
  assign n5030 = ~n5028 & n5029 ;
  assign n5031 = n4940 & n5030 ;
  assign n5032 = n4940 & ~n5031 ;
  assign n5033 = x78 & n1859 ;
  assign n5034 = x77 & n1854 ;
  assign n5035 = x76 & ~n1853 ;
  assign n5036 = n2037 & n5035 ;
  assign n5037 = n5034 | n5036 ;
  assign n5038 = n5033 | n5037 ;
  assign n5039 = n1862 | n5033 ;
  assign n5040 = n5037 | n5039 ;
  assign n5041 = ( n1192 & n5038 ) | ( n1192 & n5040 ) | ( n5038 & n5040 ) ;
  assign n5042 = x20 & n5040 ;
  assign n5043 = x20 & n5033 ;
  assign n5044 = ( x20 & n5037 ) | ( x20 & n5043 ) | ( n5037 & n5043 ) ;
  assign n5045 = ( n1192 & n5042 ) | ( n1192 & n5044 ) | ( n5042 & n5044 ) ;
  assign n5046 = x20 & ~n5044 ;
  assign n5047 = x20 & ~n5040 ;
  assign n5048 = ( ~n1192 & n5046 ) | ( ~n1192 & n5047 ) | ( n5046 & n5047 ) ;
  assign n5049 = ( n5041 & ~n5045 ) | ( n5041 & n5048 ) | ( ~n5045 & n5048 ) ;
  assign n5050 = n5030 & n5049 ;
  assign n5051 = ~n5030 & n5049 ;
  assign n5052 = ( ~n4940 & n5049 ) | ( ~n4940 & n5051 ) | ( n5049 & n5051 ) ;
  assign n5053 = ( n5032 & n5050 ) | ( n5032 & n5052 ) | ( n5050 & n5052 ) ;
  assign n5054 = n5030 | n5049 ;
  assign n5055 = n5030 & ~n5049 ;
  assign n5056 = n4940 & n5055 ;
  assign n5057 = ( n5032 & n5054 ) | ( n5032 & ~n5056 ) | ( n5054 & ~n5056 ) ;
  assign n5058 = ~n5053 & n5057 ;
  assign n5059 = n4939 & n5058 ;
  assign n5060 = n4939 | n5058 ;
  assign n5061 = ~n5059 & n5060 ;
  assign n5062 = x81 & n1383 ;
  assign n5063 = x80 & n1378 ;
  assign n5064 = x79 & ~n1377 ;
  assign n5065 = n1542 & n5064 ;
  assign n5066 = n5063 | n5065 ;
  assign n5067 = n5062 | n5066 ;
  assign n5068 = n1386 | n5062 ;
  assign n5069 = n5066 | n5068 ;
  assign n5070 = ( n1651 & n5067 ) | ( n1651 & n5069 ) | ( n5067 & n5069 ) ;
  assign n5071 = x17 & n5069 ;
  assign n5072 = x17 & n5062 ;
  assign n5073 = ( x17 & n5066 ) | ( x17 & n5072 ) | ( n5066 & n5072 ) ;
  assign n5074 = ( n1651 & n5071 ) | ( n1651 & n5073 ) | ( n5071 & n5073 ) ;
  assign n5075 = x17 & ~n5073 ;
  assign n5076 = x17 & ~n5069 ;
  assign n5077 = ( ~n1651 & n5075 ) | ( ~n1651 & n5076 ) | ( n5075 & n5076 ) ;
  assign n5078 = ( n5070 & ~n5074 ) | ( n5070 & n5077 ) | ( ~n5074 & n5077 ) ;
  assign n5079 = n5061 & n5078 ;
  assign n5080 = n5061 & ~n5079 ;
  assign n5081 = ~n5061 & n5078 ;
  assign n5082 = n5080 | n5081 ;
  assign n5083 = n4755 | n4757 ;
  assign n5084 = n4756 | n5083 ;
  assign n5085 = ( n4755 & n4761 ) | ( n4755 & n5084 ) | ( n4761 & n5084 ) ;
  assign n5086 = n5082 | n5085 ;
  assign n5087 = n5082 & n5085 ;
  assign n5088 = n5086 & ~n5087 ;
  assign n5089 = x84 & n962 ;
  assign n5090 = x83 & n957 ;
  assign n5091 = x82 & ~n956 ;
  assign n5092 = n1105 & n5091 ;
  assign n5093 = n5090 | n5092 ;
  assign n5094 = n5089 | n5093 ;
  assign n5095 = n965 | n5089 ;
  assign n5096 = n5093 | n5095 ;
  assign n5097 = ( n2194 & n5094 ) | ( n2194 & n5096 ) | ( n5094 & n5096 ) ;
  assign n5098 = x14 & n5096 ;
  assign n5099 = x14 & n5089 ;
  assign n5100 = ( x14 & n5093 ) | ( x14 & n5099 ) | ( n5093 & n5099 ) ;
  assign n5101 = ( n2194 & n5098 ) | ( n2194 & n5100 ) | ( n5098 & n5100 ) ;
  assign n5102 = x14 & ~n5100 ;
  assign n5103 = x14 & ~n5096 ;
  assign n5104 = ( ~n2194 & n5102 ) | ( ~n2194 & n5103 ) | ( n5102 & n5103 ) ;
  assign n5105 = ( n5097 & ~n5101 ) | ( n5097 & n5104 ) | ( ~n5101 & n5104 ) ;
  assign n5106 = n5088 | n5105 ;
  assign n5107 = n5088 & n5105 ;
  assign n5108 = n5106 & ~n5107 ;
  assign n5109 = n4782 & n5108 ;
  assign n5110 = ( n4789 & n5108 ) | ( n4789 & n5109 ) | ( n5108 & n5109 ) ;
  assign n5111 = n5108 & ~n5110 ;
  assign n5112 = n4782 & ~n5108 ;
  assign n5113 = ( n4789 & ~n5108 ) | ( n4789 & n5112 ) | ( ~n5108 & n5112 ) ;
  assign n5114 = n4938 & n5113 ;
  assign n5115 = ( n4938 & n5111 ) | ( n4938 & n5114 ) | ( n5111 & n5114 ) ;
  assign n5116 = n4938 | n5113 ;
  assign n5117 = n5111 | n5116 ;
  assign n5118 = ~n5115 & n5117 ;
  assign n5119 = n4808 | n4815 ;
  assign n5120 = n5118 & n5119 ;
  assign n5121 = n5118 | n5119 ;
  assign n5122 = ~n5120 & n5121 ;
  assign n5123 = x90 & n389 ;
  assign n5124 = x89 & n384 ;
  assign n5125 = x88 & ~n383 ;
  assign n5126 = n463 & n5125 ;
  assign n5127 = n5124 | n5126 ;
  assign n5128 = n5123 | n5127 ;
  assign n5129 = n392 | n5123 ;
  assign n5130 = n5127 | n5129 ;
  assign n5131 = ( n3519 & n5128 ) | ( n3519 & n5130 ) | ( n5128 & n5130 ) ;
  assign n5132 = x8 & n5130 ;
  assign n5133 = x8 & n5123 ;
  assign n5134 = ( x8 & n5127 ) | ( x8 & n5133 ) | ( n5127 & n5133 ) ;
  assign n5135 = ( n3519 & n5132 ) | ( n3519 & n5134 ) | ( n5132 & n5134 ) ;
  assign n5136 = x8 & ~n5134 ;
  assign n5137 = x8 & ~n5130 ;
  assign n5138 = ( ~n3519 & n5136 ) | ( ~n3519 & n5137 ) | ( n5136 & n5137 ) ;
  assign n5139 = ( n5131 & ~n5135 ) | ( n5131 & n5138 ) | ( ~n5135 & n5138 ) ;
  assign n5140 = n5122 & n5139 ;
  assign n5141 = n5122 & ~n5140 ;
  assign n5142 = ~n5122 & n5139 ;
  assign n5143 = n5141 | n5142 ;
  assign n5144 = n4836 | n4843 ;
  assign n5145 = n5143 | n5144 ;
  assign n5146 = n5143 & n5144 ;
  assign n5147 = n5145 & ~n5146 ;
  assign n5148 = x93 & n212 ;
  assign n5149 = x92 & n207 ;
  assign n5150 = x91 & ~n206 ;
  assign n5151 = n267 & n5150 ;
  assign n5152 = n5149 | n5151 ;
  assign n5153 = n5148 | n5152 ;
  assign n5154 = n215 | n5148 ;
  assign n5155 = n5152 | n5154 ;
  assign n5156 = ( n4305 & n5153 ) | ( n4305 & n5155 ) | ( n5153 & n5155 ) ;
  assign n5157 = x5 & n5155 ;
  assign n5158 = x5 & n5148 ;
  assign n5159 = ( x5 & n5152 ) | ( x5 & n5158 ) | ( n5152 & n5158 ) ;
  assign n5160 = ( n4305 & n5157 ) | ( n4305 & n5159 ) | ( n5157 & n5159 ) ;
  assign n5161 = x5 & ~n5159 ;
  assign n5162 = x5 & ~n5155 ;
  assign n5163 = ( ~n4305 & n5161 ) | ( ~n4305 & n5162 ) | ( n5161 & n5162 ) ;
  assign n5164 = ( n5156 & ~n5160 ) | ( n5156 & n5163 ) | ( ~n5160 & n5163 ) ;
  assign n5165 = n5147 & n5164 ;
  assign n5166 = n5147 | n5164 ;
  assign n5167 = ~n5165 & n5166 ;
  assign n5168 = n4862 & n5167 ;
  assign n5169 = ( n4868 & n5167 ) | ( n4868 & n5168 ) | ( n5167 & n5168 ) ;
  assign n5170 = n4862 | n4864 ;
  assign n5171 = n4863 | n5170 ;
  assign n5172 = ( n4862 & n4866 ) | ( n4862 & n5171 ) | ( n4866 & n5171 ) ;
  assign n5173 = n5167 | n5172 ;
  assign n5174 = ~n5169 & n5173 ;
  assign n5175 = x95 | x96 ;
  assign n5176 = x95 & x96 ;
  assign n5177 = n5175 & ~n5176 ;
  assign n5178 = n4871 | n4872 ;
  assign n5179 = ( n4871 & n4873 ) | ( n4871 & n5178 ) | ( n4873 & n5178 ) ;
  assign n5180 = n5177 & n5179 ;
  assign n5181 = n4563 | n4871 ;
  assign n5182 = ( n4871 & n4872 ) | ( n4871 & n5181 ) | ( n4872 & n5181 ) ;
  assign n5183 = n5177 & n5182 ;
  assign n5184 = ( n4029 & n4565 ) | ( n4029 & n4567 ) | ( n4565 & n4567 ) ;
  assign n5185 = ( n5180 & n5183 ) | ( n5180 & n5184 ) | ( n5183 & n5184 ) ;
  assign n5186 = n4288 | n4294 ;
  assign n5187 = ( n5180 & n5183 ) | ( n5180 & n5186 ) | ( n5183 & n5186 ) ;
  assign n5188 = ( n3274 & n5185 ) | ( n3274 & n5187 ) | ( n5185 & n5187 ) ;
  assign n5189 = ( n3276 & n5185 ) | ( n3276 & n5187 ) | ( n5185 & n5187 ) ;
  assign n5190 = ( n1493 & n5188 ) | ( n1493 & n5189 ) | ( n5188 & n5189 ) ;
  assign n5191 = ( n4565 & n5179 ) | ( n4565 & n5182 ) | ( n5179 & n5182 ) ;
  assign n5192 = ( n4567 & n5179 ) | ( n4567 & n5182 ) | ( n5179 & n5182 ) ;
  assign n5193 = ( n4029 & n5191 ) | ( n4029 & n5192 ) | ( n5191 & n5192 ) ;
  assign n5194 = n5177 | n5193 ;
  assign n5195 = ( n4288 & n5179 ) | ( n4288 & n5182 ) | ( n5179 & n5182 ) ;
  assign n5196 = n5179 | n5182 ;
  assign n5197 = ( n4294 & n5195 ) | ( n4294 & n5196 ) | ( n5195 & n5196 ) ;
  assign n5198 = n5177 | n5197 ;
  assign n5199 = ( n3274 & n5194 ) | ( n3274 & n5198 ) | ( n5194 & n5198 ) ;
  assign n5200 = ( n3276 & n5194 ) | ( n3276 & n5198 ) | ( n5194 & n5198 ) ;
  assign n5201 = ( n1493 & n5199 ) | ( n1493 & n5200 ) | ( n5199 & n5200 ) ;
  assign n5202 = ~n5190 & n5201 ;
  assign n5203 = x95 & n133 ;
  assign n5204 = x94 & ~n162 ;
  assign n5205 = ( n137 & n5203 ) | ( n137 & n5204 ) | ( n5203 & n5204 ) ;
  assign n5206 = x0 & x96 ;
  assign n5207 = ( ~n137 & n5203 ) | ( ~n137 & n5206 ) | ( n5203 & n5206 ) ;
  assign n5208 = n5205 | n5207 ;
  assign n5209 = n141 | n5208 ;
  assign n5210 = ( n5202 & n5208 ) | ( n5202 & n5209 ) | ( n5208 & n5209 ) ;
  assign n5211 = x2 & n5208 ;
  assign n5212 = ( x2 & n523 ) | ( x2 & n5208 ) | ( n523 & n5208 ) ;
  assign n5213 = ( n5202 & n5211 ) | ( n5202 & n5212 ) | ( n5211 & n5212 ) ;
  assign n5214 = x2 & ~n5212 ;
  assign n5215 = x2 & ~n5208 ;
  assign n5216 = ( ~n5202 & n5214 ) | ( ~n5202 & n5215 ) | ( n5214 & n5215 ) ;
  assign n5217 = ( n5210 & ~n5213 ) | ( n5210 & n5216 ) | ( ~n5213 & n5216 ) ;
  assign n5218 = n5174 & ~n5217 ;
  assign n5219 = ~n5174 & n5217 ;
  assign n5220 = n5218 | n5219 ;
  assign n5221 = n4913 | n4918 ;
  assign n5222 = ( n4913 & n4916 ) | ( n4913 & n5221 ) | ( n4916 & n5221 ) ;
  assign n5223 = n5220 & n5222 ;
  assign n5224 = n5220 | n5222 ;
  assign n5225 = ~n5223 & n5224 ;
  assign n5226 = n5165 | n5169 ;
  assign n5227 = n5107 | n5110 ;
  assign n5228 = n5079 | n5087 ;
  assign n5229 = n5053 | n5059 ;
  assign n5230 = x32 & ~x33 ;
  assign n5231 = ~x32 & x33 ;
  assign n5232 = n5230 | n5231 ;
  assign n5233 = x64 & n5232 ;
  assign n5234 = ~n4646 & n5233 ;
  assign n5235 = ( ~n4955 & n5233 ) | ( ~n4955 & n5234 ) | ( n5233 & n5234 ) ;
  assign n5236 = n4646 & ~n5233 ;
  assign n5237 = n4955 & n5236 ;
  assign n5238 = n5235 | n5237 ;
  assign n5239 = x67 & n4631 ;
  assign n5240 = x66 & n4626 ;
  assign n5241 = x65 & ~n4625 ;
  assign n5242 = n4943 & n5241 ;
  assign n5243 = n5240 | n5242 ;
  assign n5244 = n5239 | n5243 ;
  assign n5245 = n186 & n4634 ;
  assign n5246 = n5244 | n5245 ;
  assign n5247 = x32 & ~n5246 ;
  assign n5248 = ~x32 & n5246 ;
  assign n5249 = n5247 | n5248 ;
  assign n5250 = n5238 & n5249 ;
  assign n5251 = n5238 | n5249 ;
  assign n5252 = ~n5250 & n5251 ;
  assign n5253 = x69 & n3811 ;
  assign n5254 = x68 & ~n3810 ;
  assign n5255 = n4067 & n5254 ;
  assign n5256 = n5253 | n5255 ;
  assign n5257 = x70 & n3816 ;
  assign n5258 = n3819 | n5257 ;
  assign n5259 = n5256 | n5258 ;
  assign n5260 = x29 & ~n5259 ;
  assign n5261 = x29 & ~n5257 ;
  assign n5262 = ~n5256 & n5261 ;
  assign n5263 = ( ~n340 & n5260 ) | ( ~n340 & n5262 ) | ( n5260 & n5262 ) ;
  assign n5264 = ~x29 & n5259 ;
  assign n5265 = ~x29 & n5257 ;
  assign n5266 = ( ~x29 & n5256 ) | ( ~x29 & n5265 ) | ( n5256 & n5265 ) ;
  assign n5267 = ( n340 & n5264 ) | ( n340 & n5266 ) | ( n5264 & n5266 ) ;
  assign n5268 = n5263 | n5267 ;
  assign n5269 = ( n4978 & ~n5252 ) | ( n4978 & n5268 ) | ( ~n5252 & n5268 ) ;
  assign n5270 = ( ~n4978 & n5252 ) | ( ~n4978 & n5269 ) | ( n5252 & n5269 ) ;
  assign n5271 = x73 & n3085 ;
  assign n5272 = x72 & n3080 ;
  assign n5273 = x71 & ~n3079 ;
  assign n5274 = n3309 & n5273 ;
  assign n5275 = n5272 | n5274 ;
  assign n5276 = n5271 | n5275 ;
  assign n5277 = ( ~n610 & n3088 ) | ( ~n610 & n5276 ) | ( n3088 & n5276 ) ;
  assign n5278 = n3088 & n5271 ;
  assign n5279 = ( n3088 & n5275 ) | ( n3088 & n5278 ) | ( n5275 & n5278 ) ;
  assign n5280 = ( n598 & n5277 ) | ( n598 & n5279 ) | ( n5277 & n5279 ) ;
  assign n5281 = ( x26 & ~n5276 ) | ( x26 & n5280 ) | ( ~n5276 & n5280 ) ;
  assign n5282 = ~n5280 & n5281 ;
  assign n5283 = x26 | n5271 ;
  assign n5284 = n5275 | n5283 ;
  assign n5285 = n5280 | n5284 ;
  assign n5286 = ( ~x26 & n5282 ) | ( ~x26 & n5285 ) | ( n5282 & n5285 ) ;
  assign n5287 = ~n5252 & n5286 ;
  assign n5288 = n5268 & n5286 ;
  assign n5289 = ( n4978 & n5287 ) | ( n4978 & n5288 ) | ( n5287 & n5288 ) ;
  assign n5290 = ~n5268 & n5285 ;
  assign n5291 = x26 | n5268 ;
  assign n5292 = ( n5282 & n5290 ) | ( n5282 & ~n5291 ) | ( n5290 & ~n5291 ) ;
  assign n5293 = ( n5270 & n5289 ) | ( n5270 & n5292 ) | ( n5289 & n5292 ) ;
  assign n5294 = n5252 & ~n5286 ;
  assign n5295 = n5268 | n5286 ;
  assign n5296 = ( n4978 & ~n5294 ) | ( n4978 & n5295 ) | ( ~n5294 & n5295 ) ;
  assign n5297 = n5268 & ~n5285 ;
  assign n5298 = x26 & n5268 ;
  assign n5299 = ( ~n5282 & n5297 ) | ( ~n5282 & n5298 ) | ( n5297 & n5298 ) ;
  assign n5300 = ( n5270 & n5296 ) | ( n5270 & ~n5299 ) | ( n5296 & ~n5299 ) ;
  assign n5301 = ~n5293 & n5300 ;
  assign n5302 = n5000 & n5301 ;
  assign n5303 = ( n5009 & n5301 ) | ( n5009 & n5302 ) | ( n5301 & n5302 ) ;
  assign n5304 = n5000 | n5301 ;
  assign n5305 = n5009 | n5304 ;
  assign n5306 = ~n5303 & n5305 ;
  assign n5307 = x76 & n2429 ;
  assign n5308 = x75 & n2424 ;
  assign n5309 = x74 & ~n2423 ;
  assign n5310 = n2631 & n5309 ;
  assign n5311 = n5308 | n5310 ;
  assign n5312 = n5307 | n5311 ;
  assign n5313 = n2432 | n5307 ;
  assign n5314 = n5311 | n5313 ;
  assign n5315 = ( n923 & n5312 ) | ( n923 & n5314 ) | ( n5312 & n5314 ) ;
  assign n5316 = x23 & n5314 ;
  assign n5317 = x23 & n5307 ;
  assign n5318 = ( x23 & n5311 ) | ( x23 & n5317 ) | ( n5311 & n5317 ) ;
  assign n5319 = ( n923 & n5316 ) | ( n923 & n5318 ) | ( n5316 & n5318 ) ;
  assign n5320 = x23 & ~n5318 ;
  assign n5321 = x23 & ~n5314 ;
  assign n5322 = ( ~n923 & n5320 ) | ( ~n923 & n5321 ) | ( n5320 & n5321 ) ;
  assign n5323 = ( n5315 & ~n5319 ) | ( n5315 & n5322 ) | ( ~n5319 & n5322 ) ;
  assign n5324 = n5306 | n5323 ;
  assign n5325 = n5306 & n5323 ;
  assign n5326 = n5324 & ~n5325 ;
  assign n5327 = n5028 | n5030 ;
  assign n5328 = ( n4940 & n5028 ) | ( n4940 & n5327 ) | ( n5028 & n5327 ) ;
  assign n5329 = n5326 & n5328 ;
  assign n5330 = n5326 | n5328 ;
  assign n5331 = ~n5329 & n5330 ;
  assign n5332 = x79 & n1859 ;
  assign n5333 = x78 & n1854 ;
  assign n5334 = x77 & ~n1853 ;
  assign n5335 = n2037 & n5334 ;
  assign n5336 = n5333 | n5335 ;
  assign n5337 = n5332 | n5336 ;
  assign n5338 = n1862 | n5332 ;
  assign n5339 = n5336 | n5338 ;
  assign n5340 = ( n1332 & n5337 ) | ( n1332 & n5339 ) | ( n5337 & n5339 ) ;
  assign n5341 = x20 & n5339 ;
  assign n5342 = x20 & n5332 ;
  assign n5343 = ( x20 & n5336 ) | ( x20 & n5342 ) | ( n5336 & n5342 ) ;
  assign n5344 = ( n1332 & n5341 ) | ( n1332 & n5343 ) | ( n5341 & n5343 ) ;
  assign n5345 = x20 & ~n5343 ;
  assign n5346 = x20 & ~n5339 ;
  assign n5347 = ( ~n1332 & n5345 ) | ( ~n1332 & n5346 ) | ( n5345 & n5346 ) ;
  assign n5348 = ( n5340 & ~n5344 ) | ( n5340 & n5347 ) | ( ~n5344 & n5347 ) ;
  assign n5349 = n5331 & n5348 ;
  assign n5350 = n5331 & ~n5349 ;
  assign n5351 = ~n5331 & n5348 ;
  assign n5352 = n5350 | n5351 ;
  assign n5353 = n5229 & ~n5352 ;
  assign n5354 = ~n5229 & n5352 ;
  assign n5355 = n5353 | n5354 ;
  assign n5356 = x82 & n1383 ;
  assign n5357 = x81 & n1378 ;
  assign n5358 = x80 & ~n1377 ;
  assign n5359 = n1542 & n5358 ;
  assign n5360 = n5357 | n5359 ;
  assign n5361 = n5356 | n5360 ;
  assign n5362 = n1386 | n5356 ;
  assign n5363 = n5360 | n5362 ;
  assign n5364 = ( n1811 & n5361 ) | ( n1811 & n5363 ) | ( n5361 & n5363 ) ;
  assign n5365 = x17 & n5363 ;
  assign n5366 = x17 & n5356 ;
  assign n5367 = ( x17 & n5360 ) | ( x17 & n5366 ) | ( n5360 & n5366 ) ;
  assign n5368 = ( n1811 & n5365 ) | ( n1811 & n5367 ) | ( n5365 & n5367 ) ;
  assign n5369 = x17 & ~n5367 ;
  assign n5370 = x17 & ~n5363 ;
  assign n5371 = ( ~n1811 & n5369 ) | ( ~n1811 & n5370 ) | ( n5369 & n5370 ) ;
  assign n5372 = ( n5364 & ~n5368 ) | ( n5364 & n5371 ) | ( ~n5368 & n5371 ) ;
  assign n5373 = n5355 & n5372 ;
  assign n5374 = n5355 | n5372 ;
  assign n5375 = ~n5373 & n5374 ;
  assign n5376 = n5228 | n5375 ;
  assign n5377 = n5228 & n5375 ;
  assign n5378 = n5376 & ~n5377 ;
  assign n5379 = x85 & n962 ;
  assign n5380 = x84 & n957 ;
  assign n5381 = x83 & ~n956 ;
  assign n5382 = n1105 & n5381 ;
  assign n5383 = n5380 | n5382 ;
  assign n5384 = n5379 | n5383 ;
  assign n5385 = n965 | n5379 ;
  assign n5386 = n5383 | n5385 ;
  assign n5387 = ( n2381 & n5384 ) | ( n2381 & n5386 ) | ( n5384 & n5386 ) ;
  assign n5388 = x14 & n5386 ;
  assign n5389 = x14 & n5379 ;
  assign n5390 = ( x14 & n5383 ) | ( x14 & n5389 ) | ( n5383 & n5389 ) ;
  assign n5391 = ( n2381 & n5388 ) | ( n2381 & n5390 ) | ( n5388 & n5390 ) ;
  assign n5392 = x14 & ~n5390 ;
  assign n5393 = x14 & ~n5386 ;
  assign n5394 = ( ~n2381 & n5392 ) | ( ~n2381 & n5393 ) | ( n5392 & n5393 ) ;
  assign n5395 = ( n5387 & ~n5391 ) | ( n5387 & n5394 ) | ( ~n5391 & n5394 ) ;
  assign n5396 = n5378 & n5395 ;
  assign n5397 = n5378 & ~n5396 ;
  assign n5398 = ~n5378 & n5395 ;
  assign n5399 = n5397 | n5398 ;
  assign n5400 = n5227 & ~n5399 ;
  assign n5401 = ~n5227 & n5399 ;
  assign n5402 = n5400 | n5401 ;
  assign n5403 = x88 & n636 ;
  assign n5404 = x87 & n631 ;
  assign n5405 = x86 & ~n630 ;
  assign n5406 = n764 & n5405 ;
  assign n5407 = n5404 | n5406 ;
  assign n5408 = n5403 | n5407 ;
  assign n5409 = n639 | n5403 ;
  assign n5410 = n5407 | n5409 ;
  assign n5411 = ( ~n3039 & n5408 ) | ( ~n3039 & n5410 ) | ( n5408 & n5410 ) ;
  assign n5412 = n5408 & n5410 ;
  assign n5413 = ( n3023 & n5411 ) | ( n3023 & n5412 ) | ( n5411 & n5412 ) ;
  assign n5414 = x11 & n5410 ;
  assign n5415 = x11 & n5403 ;
  assign n5416 = ( x11 & n5407 ) | ( x11 & n5415 ) | ( n5407 & n5415 ) ;
  assign n5417 = ( ~n3039 & n5414 ) | ( ~n3039 & n5416 ) | ( n5414 & n5416 ) ;
  assign n5418 = n5414 & n5416 ;
  assign n5419 = ( n3023 & n5417 ) | ( n3023 & n5418 ) | ( n5417 & n5418 ) ;
  assign n5420 = x11 & ~n5416 ;
  assign n5421 = x11 & ~n5410 ;
  assign n5422 = ( n3039 & n5420 ) | ( n3039 & n5421 ) | ( n5420 & n5421 ) ;
  assign n5423 = n5420 | n5421 ;
  assign n5424 = ( ~n3023 & n5422 ) | ( ~n3023 & n5423 ) | ( n5422 & n5423 ) ;
  assign n5425 = ( n5413 & ~n5419 ) | ( n5413 & n5424 ) | ( ~n5419 & n5424 ) ;
  assign n5426 = n5402 | n5425 ;
  assign n5427 = n5402 & n5425 ;
  assign n5428 = n5426 & ~n5427 ;
  assign n5429 = n5115 | n5118 ;
  assign n5430 = ( n5115 & n5119 ) | ( n5115 & n5429 ) | ( n5119 & n5429 ) ;
  assign n5431 = n5428 & n5430 ;
  assign n5432 = n5428 | n5430 ;
  assign n5433 = ~n5431 & n5432 ;
  assign n5434 = x91 & n389 ;
  assign n5435 = x90 & n384 ;
  assign n5436 = x89 & ~n383 ;
  assign n5437 = n463 & n5436 ;
  assign n5438 = n5435 | n5437 ;
  assign n5439 = n5434 | n5438 ;
  assign n5440 = n392 | n5434 ;
  assign n5441 = n5438 | n5440 ;
  assign n5442 = ( n3768 & n5439 ) | ( n3768 & n5441 ) | ( n5439 & n5441 ) ;
  assign n5443 = x8 & n5441 ;
  assign n5444 = x8 & n5434 ;
  assign n5445 = ( x8 & n5438 ) | ( x8 & n5444 ) | ( n5438 & n5444 ) ;
  assign n5446 = ( n3768 & n5443 ) | ( n3768 & n5445 ) | ( n5443 & n5445 ) ;
  assign n5447 = x8 & ~n5445 ;
  assign n5448 = x8 & ~n5441 ;
  assign n5449 = ( ~n3768 & n5447 ) | ( ~n3768 & n5448 ) | ( n5447 & n5448 ) ;
  assign n5450 = ( n5442 & ~n5446 ) | ( n5442 & n5449 ) | ( ~n5446 & n5449 ) ;
  assign n5451 = n5433 & n5450 ;
  assign n5452 = n5433 & ~n5451 ;
  assign n5453 = ~n5433 & n5450 ;
  assign n5454 = n5452 | n5453 ;
  assign n5455 = n5140 | n5146 ;
  assign n5456 = n5454 | n5455 ;
  assign n5457 = n5454 & n5455 ;
  assign n5458 = n5456 & ~n5457 ;
  assign n5459 = x94 & n212 ;
  assign n5460 = x93 & n207 ;
  assign n5461 = x92 & ~n206 ;
  assign n5462 = n267 & n5461 ;
  assign n5463 = n5460 | n5462 ;
  assign n5464 = n5459 | n5463 ;
  assign n5465 = n215 | n5459 ;
  assign n5466 = n5463 | n5465 ;
  assign n5467 = ( n4583 & n5464 ) | ( n4583 & n5466 ) | ( n5464 & n5466 ) ;
  assign n5468 = x5 & n5466 ;
  assign n5469 = x5 & n5459 ;
  assign n5470 = ( x5 & n5463 ) | ( x5 & n5469 ) | ( n5463 & n5469 ) ;
  assign n5471 = ( n4583 & n5468 ) | ( n4583 & n5470 ) | ( n5468 & n5470 ) ;
  assign n5472 = x5 & ~n5470 ;
  assign n5473 = x5 & ~n5466 ;
  assign n5474 = ( ~n4583 & n5472 ) | ( ~n4583 & n5473 ) | ( n5472 & n5473 ) ;
  assign n5475 = ( n5467 & ~n5471 ) | ( n5467 & n5474 ) | ( ~n5471 & n5474 ) ;
  assign n5476 = n5458 & n5475 ;
  assign n5477 = n5458 & ~n5476 ;
  assign n5478 = ~n5458 & n5475 ;
  assign n5479 = n5477 | n5478 ;
  assign n5480 = n5226 & ~n5479 ;
  assign n5481 = ~n5226 & n5479 ;
  assign n5482 = n5480 | n5481 ;
  assign n5483 = x96 | x97 ;
  assign n5484 = x96 & x97 ;
  assign n5485 = n5483 & ~n5484 ;
  assign n5486 = n5176 | n5177 ;
  assign n5487 = ( n5176 & n5182 ) | ( n5176 & n5486 ) | ( n5182 & n5486 ) ;
  assign n5488 = n5485 & n5487 ;
  assign n5489 = n5485 & n5486 ;
  assign n5490 = n5176 & n5485 ;
  assign n5491 = ( n5179 & n5489 ) | ( n5179 & n5490 ) | ( n5489 & n5490 ) ;
  assign n5492 = ( n5184 & n5488 ) | ( n5184 & n5491 ) | ( n5488 & n5491 ) ;
  assign n5493 = ( n5186 & n5488 ) | ( n5186 & n5491 ) | ( n5488 & n5491 ) ;
  assign n5494 = ( n3274 & n5492 ) | ( n3274 & n5493 ) | ( n5492 & n5493 ) ;
  assign n5495 = ( n3276 & n5492 ) | ( n3276 & n5493 ) | ( n5492 & n5493 ) ;
  assign n5496 = ( n1493 & n5494 ) | ( n1493 & n5495 ) | ( n5494 & n5495 ) ;
  assign n5497 = ( n5176 & n5179 ) | ( n5176 & n5486 ) | ( n5179 & n5486 ) ;
  assign n5498 = n5485 | n5497 ;
  assign n5499 = n5485 | n5487 ;
  assign n5500 = ( n5184 & n5498 ) | ( n5184 & n5499 ) | ( n5498 & n5499 ) ;
  assign n5501 = ( n5186 & n5498 ) | ( n5186 & n5499 ) | ( n5498 & n5499 ) ;
  assign n5502 = ( n3274 & n5500 ) | ( n3274 & n5501 ) | ( n5500 & n5501 ) ;
  assign n5503 = ( n3276 & n5500 ) | ( n3276 & n5501 ) | ( n5500 & n5501 ) ;
  assign n5504 = ( n1493 & n5502 ) | ( n1493 & n5503 ) | ( n5502 & n5503 ) ;
  assign n5505 = ~n5496 & n5504 ;
  assign n5506 = x96 & n133 ;
  assign n5507 = x95 & ~n162 ;
  assign n5508 = ( n137 & n5506 ) | ( n137 & n5507 ) | ( n5506 & n5507 ) ;
  assign n5509 = x0 & x97 ;
  assign n5510 = ( ~n137 & n5506 ) | ( ~n137 & n5509 ) | ( n5506 & n5509 ) ;
  assign n5511 = n5508 | n5510 ;
  assign n5512 = n141 | n5511 ;
  assign n5513 = ( n5505 & n5511 ) | ( n5505 & n5512 ) | ( n5511 & n5512 ) ;
  assign n5514 = x2 & n5511 ;
  assign n5515 = ( x2 & n523 ) | ( x2 & n5511 ) | ( n523 & n5511 ) ;
  assign n5516 = ( n5505 & n5514 ) | ( n5505 & n5515 ) | ( n5514 & n5515 ) ;
  assign n5517 = x2 & ~n5515 ;
  assign n5518 = x2 & ~n5511 ;
  assign n5519 = ( ~n5505 & n5517 ) | ( ~n5505 & n5518 ) | ( n5517 & n5518 ) ;
  assign n5520 = ( n5513 & ~n5516 ) | ( n5513 & n5519 ) | ( ~n5516 & n5519 ) ;
  assign n5521 = n5482 & n5520 ;
  assign n5522 = n5482 | n5520 ;
  assign n5523 = ~n5521 & n5522 ;
  assign n5524 = ( n5174 & n5217 ) | ( n5174 & n5222 ) | ( n5217 & n5222 ) ;
  assign n5525 = n5523 | n5524 ;
  assign n5526 = n5523 & n5524 ;
  assign n5527 = n5525 & ~n5526 ;
  assign n5528 = n5226 & n5479 ;
  assign n5529 = n5476 | n5528 ;
  assign n5530 = x70 & n3811 ;
  assign n5531 = x69 & ~n3810 ;
  assign n5532 = n4067 & n5531 ;
  assign n5533 = n5530 | n5532 ;
  assign n5534 = x71 & n3816 ;
  assign n5535 = n3819 | n5534 ;
  assign n5536 = n5533 | n5535 ;
  assign n5537 = x29 & ~n5536 ;
  assign n5538 = x29 & ~n5534 ;
  assign n5539 = ~n5533 & n5538 ;
  assign n5540 = ( ~n438 & n5537 ) | ( ~n438 & n5539 ) | ( n5537 & n5539 ) ;
  assign n5541 = ~x29 & n5536 ;
  assign n5542 = ~x29 & n5534 ;
  assign n5543 = ( ~x29 & n5533 ) | ( ~x29 & n5542 ) | ( n5533 & n5542 ) ;
  assign n5544 = ( n438 & n5541 ) | ( n438 & n5543 ) | ( n5541 & n5543 ) ;
  assign n5545 = n5540 | n5544 ;
  assign n5546 = ~x33 & x34 ;
  assign n5547 = x33 & ~x34 ;
  assign n5548 = n5546 | n5547 ;
  assign n5549 = ~n5232 & n5548 ;
  assign n5550 = x64 & n5549 ;
  assign n5551 = ~x34 & x35 ;
  assign n5552 = x34 & ~x35 ;
  assign n5553 = n5551 | n5552 ;
  assign n5554 = n5232 & ~n5553 ;
  assign n5555 = x65 & n5554 ;
  assign n5556 = n5550 | n5555 ;
  assign n5557 = n5232 & n5553 ;
  assign n5558 = x35 | n144 ;
  assign n5559 = ( x35 & n5557 ) | ( x35 & n5558 ) | ( n5557 & n5558 ) ;
  assign n5560 = ~x35 & n5559 ;
  assign n5561 = ( ~x35 & n5556 ) | ( ~x35 & n5560 ) | ( n5556 & n5560 ) ;
  assign n5562 = x35 & ~x64 ;
  assign n5563 = ( x35 & ~n5232 ) | ( x35 & n5562 ) | ( ~n5232 & n5562 ) ;
  assign n5564 = n5559 & n5563 ;
  assign n5565 = ( n5556 & n5563 ) | ( n5556 & n5564 ) | ( n5563 & n5564 ) ;
  assign n5566 = n144 & n5557 ;
  assign n5567 = n5563 & ~n5566 ;
  assign n5568 = ~n5556 & n5567 ;
  assign n5569 = ( n5561 & n5565 ) | ( n5561 & n5568 ) | ( n5565 & n5568 ) ;
  assign n5570 = n5559 | n5563 ;
  assign n5571 = n5556 | n5570 ;
  assign n5572 = ~n5563 & n5566 ;
  assign n5573 = ( n5556 & ~n5563 ) | ( n5556 & n5572 ) | ( ~n5563 & n5572 ) ;
  assign n5574 = ( n5561 & n5571 ) | ( n5561 & ~n5573 ) | ( n5571 & ~n5573 ) ;
  assign n5575 = ~n5569 & n5574 ;
  assign n5576 = n241 & n4634 ;
  assign n5577 = x68 & n4631 ;
  assign n5578 = x67 & n4626 ;
  assign n5579 = x66 & ~n4625 ;
  assign n5580 = n4943 & n5579 ;
  assign n5581 = n5578 | n5580 ;
  assign n5582 = n5577 | n5581 ;
  assign n5583 = n5576 | n5582 ;
  assign n5584 = x32 | n5577 ;
  assign n5585 = n5581 | n5584 ;
  assign n5586 = n5576 | n5585 ;
  assign n5587 = ~x32 & n5585 ;
  assign n5588 = ( ~x32 & n5576 ) | ( ~x32 & n5587 ) | ( n5576 & n5587 ) ;
  assign n5589 = ( ~n5583 & n5586 ) | ( ~n5583 & n5588 ) | ( n5586 & n5588 ) ;
  assign n5590 = n5575 | n5589 ;
  assign n5591 = n5575 & n5589 ;
  assign n5592 = n5590 & ~n5591 ;
  assign n5593 = ( n4957 & n5233 ) | ( n4957 & n5249 ) | ( n5233 & n5249 ) ;
  assign n5594 = n5592 | n5593 ;
  assign n5595 = n5592 & n5593 ;
  assign n5596 = n5594 & ~n5595 ;
  assign n5597 = n5545 | n5596 ;
  assign n5598 = n5545 & n5596 ;
  assign n5599 = n5597 & ~n5598 ;
  assign n5600 = n5252 & n5268 ;
  assign n5601 = n5252 & ~n5600 ;
  assign n5602 = ~n5252 & n5268 ;
  assign n5603 = n4978 & ~n5602 ;
  assign n5604 = ~n5601 & n5603 ;
  assign n5605 = ( n4978 & n5600 ) | ( n4978 & ~n5604 ) | ( n5600 & ~n5604 ) ;
  assign n5606 = n5599 & n5605 ;
  assign n5607 = n5599 | n5605 ;
  assign n5608 = ~n5606 & n5607 ;
  assign n5609 = x74 & n3085 ;
  assign n5610 = x73 & n3080 ;
  assign n5611 = x72 & ~n3079 ;
  assign n5612 = n3309 & n5611 ;
  assign n5613 = n5610 | n5612 ;
  assign n5614 = n5609 | n5613 ;
  assign n5615 = n3088 | n5609 ;
  assign n5616 = n5613 | n5615 ;
  assign n5617 = ( n710 & n5614 ) | ( n710 & n5616 ) | ( n5614 & n5616 ) ;
  assign n5618 = x26 & n5616 ;
  assign n5619 = x26 & n5609 ;
  assign n5620 = ( x26 & n5613 ) | ( x26 & n5619 ) | ( n5613 & n5619 ) ;
  assign n5621 = ( n710 & n5618 ) | ( n710 & n5620 ) | ( n5618 & n5620 ) ;
  assign n5622 = x26 & ~n5620 ;
  assign n5623 = x26 & ~n5616 ;
  assign n5624 = ( ~n710 & n5622 ) | ( ~n710 & n5623 ) | ( n5622 & n5623 ) ;
  assign n5625 = ( n5617 & ~n5621 ) | ( n5617 & n5624 ) | ( ~n5621 & n5624 ) ;
  assign n5626 = n5608 & n5625 ;
  assign n5627 = n5608 & ~n5626 ;
  assign n5628 = ~n5608 & n5625 ;
  assign n5629 = n5627 | n5628 ;
  assign n5630 = n5293 | n5303 ;
  assign n5631 = n5629 | n5630 ;
  assign n5632 = n5629 & n5630 ;
  assign n5633 = n5631 & ~n5632 ;
  assign n5634 = x77 & n2429 ;
  assign n5635 = x76 & n2424 ;
  assign n5636 = x75 & ~n2423 ;
  assign n5637 = n2631 & n5636 ;
  assign n5638 = n5635 | n5637 ;
  assign n5639 = n5634 | n5638 ;
  assign n5640 = n2432 | n5634 ;
  assign n5641 = n5638 | n5640 ;
  assign n5642 = ( n1059 & n5639 ) | ( n1059 & n5641 ) | ( n5639 & n5641 ) ;
  assign n5643 = x23 & n5641 ;
  assign n5644 = x23 & n5634 ;
  assign n5645 = ( x23 & n5638 ) | ( x23 & n5644 ) | ( n5638 & n5644 ) ;
  assign n5646 = ( n1059 & n5643 ) | ( n1059 & n5645 ) | ( n5643 & n5645 ) ;
  assign n5647 = x23 & ~n5645 ;
  assign n5648 = x23 & ~n5641 ;
  assign n5649 = ( ~n1059 & n5647 ) | ( ~n1059 & n5648 ) | ( n5647 & n5648 ) ;
  assign n5650 = ( n5642 & ~n5646 ) | ( n5642 & n5649 ) | ( ~n5646 & n5649 ) ;
  assign n5651 = n5633 & n5650 ;
  assign n5652 = n5633 | n5650 ;
  assign n5653 = ~n5651 & n5652 ;
  assign n5654 = n5325 | n5326 ;
  assign n5655 = ( n5325 & n5328 ) | ( n5325 & n5654 ) | ( n5328 & n5654 ) ;
  assign n5656 = n5653 & n5655 ;
  assign n5657 = ~n5653 & n5655 ;
  assign n5658 = ( n5653 & ~n5656 ) | ( n5653 & n5657 ) | ( ~n5656 & n5657 ) ;
  assign n5659 = x80 & n1859 ;
  assign n5660 = x79 & n1854 ;
  assign n5661 = x78 & ~n1853 ;
  assign n5662 = n2037 & n5661 ;
  assign n5663 = n5660 | n5662 ;
  assign n5664 = n5659 | n5663 ;
  assign n5665 = n1862 | n5659 ;
  assign n5666 = n5663 | n5665 ;
  assign n5667 = ( n1499 & n5664 ) | ( n1499 & n5666 ) | ( n5664 & n5666 ) ;
  assign n5668 = x20 & n5666 ;
  assign n5669 = x20 & n5659 ;
  assign n5670 = ( x20 & n5663 ) | ( x20 & n5669 ) | ( n5663 & n5669 ) ;
  assign n5671 = ( n1499 & n5668 ) | ( n1499 & n5670 ) | ( n5668 & n5670 ) ;
  assign n5672 = x20 & ~n5670 ;
  assign n5673 = x20 & ~n5666 ;
  assign n5674 = ( ~n1499 & n5672 ) | ( ~n1499 & n5673 ) | ( n5672 & n5673 ) ;
  assign n5675 = ( n5667 & ~n5671 ) | ( n5667 & n5674 ) | ( ~n5671 & n5674 ) ;
  assign n5676 = n5658 & n5675 ;
  assign n5677 = n5658 & ~n5676 ;
  assign n5678 = ( n5053 & n5331 ) | ( n5053 & n5348 ) | ( n5331 & n5348 ) ;
  assign n5679 = n5331 | n5348 ;
  assign n5680 = ( n5059 & n5678 ) | ( n5059 & n5679 ) | ( n5678 & n5679 ) ;
  assign n5681 = ~n5658 & n5675 ;
  assign n5682 = n5680 & n5681 ;
  assign n5683 = ( n5677 & n5680 ) | ( n5677 & n5682 ) | ( n5680 & n5682 ) ;
  assign n5684 = n5680 | n5681 ;
  assign n5685 = n5677 | n5684 ;
  assign n5686 = ~n5683 & n5685 ;
  assign n5687 = x83 & n1383 ;
  assign n5688 = x82 & n1378 ;
  assign n5689 = x81 & ~n1377 ;
  assign n5690 = n1542 & n5689 ;
  assign n5691 = n5688 | n5690 ;
  assign n5692 = n5687 | n5691 ;
  assign n5693 = n1386 | n5687 ;
  assign n5694 = n5691 | n5693 ;
  assign n5695 = ( n2009 & n5692 ) | ( n2009 & n5694 ) | ( n5692 & n5694 ) ;
  assign n5696 = x17 & n5694 ;
  assign n5697 = x17 & n5687 ;
  assign n5698 = ( x17 & n5691 ) | ( x17 & n5697 ) | ( n5691 & n5697 ) ;
  assign n5699 = ( n2009 & n5696 ) | ( n2009 & n5698 ) | ( n5696 & n5698 ) ;
  assign n5700 = x17 & ~n5698 ;
  assign n5701 = x17 & ~n5694 ;
  assign n5702 = ( ~n2009 & n5700 ) | ( ~n2009 & n5701 ) | ( n5700 & n5701 ) ;
  assign n5703 = ( n5695 & ~n5699 ) | ( n5695 & n5702 ) | ( ~n5699 & n5702 ) ;
  assign n5704 = n5686 & n5703 ;
  assign n5705 = n5686 & ~n5704 ;
  assign n5706 = ~n5686 & n5703 ;
  assign n5707 = n5705 | n5706 ;
  assign n5708 = n5373 | n5375 ;
  assign n5709 = ( n5228 & n5373 ) | ( n5228 & n5708 ) | ( n5373 & n5708 ) ;
  assign n5710 = n5707 | n5709 ;
  assign n5711 = n5707 & n5709 ;
  assign n5712 = n5710 & ~n5711 ;
  assign n5713 = x86 & n962 ;
  assign n5714 = x85 & n957 ;
  assign n5715 = x84 & ~n956 ;
  assign n5716 = n1105 & n5715 ;
  assign n5717 = n5714 | n5716 ;
  assign n5718 = n5713 | n5717 ;
  assign n5719 = n965 | n5713 ;
  assign n5720 = n5717 | n5719 ;
  assign n5721 = ( n2606 & n5718 ) | ( n2606 & n5720 ) | ( n5718 & n5720 ) ;
  assign n5722 = x14 & n5720 ;
  assign n5723 = x14 & n5713 ;
  assign n5724 = ( x14 & n5717 ) | ( x14 & n5723 ) | ( n5717 & n5723 ) ;
  assign n5725 = ( n2606 & n5722 ) | ( n2606 & n5724 ) | ( n5722 & n5724 ) ;
  assign n5726 = x14 & ~n5724 ;
  assign n5727 = x14 & ~n5720 ;
  assign n5728 = ( ~n2606 & n5726 ) | ( ~n2606 & n5727 ) | ( n5726 & n5727 ) ;
  assign n5729 = ( n5721 & ~n5725 ) | ( n5721 & n5728 ) | ( ~n5725 & n5728 ) ;
  assign n5730 = n5712 & n5729 ;
  assign n5731 = n5712 & ~n5730 ;
  assign n5732 = ~n5712 & n5729 ;
  assign n5733 = n5731 | n5732 ;
  assign n5734 = ( n5107 & n5378 ) | ( n5107 & n5395 ) | ( n5378 & n5395 ) ;
  assign n5735 = n5378 | n5395 ;
  assign n5736 = ( n5110 & n5734 ) | ( n5110 & n5735 ) | ( n5734 & n5735 ) ;
  assign n5737 = n5733 | n5736 ;
  assign n5738 = n5733 & n5736 ;
  assign n5739 = n5737 & ~n5738 ;
  assign n5740 = x89 & n636 ;
  assign n5741 = x88 & n631 ;
  assign n5742 = x87 & ~n630 ;
  assign n5743 = n764 & n5742 ;
  assign n5744 = n5741 | n5743 ;
  assign n5745 = n5740 | n5744 ;
  assign n5746 = n639 | n5740 ;
  assign n5747 = n5744 | n5746 ;
  assign n5748 = ( n3282 & n5745 ) | ( n3282 & n5747 ) | ( n5745 & n5747 ) ;
  assign n5749 = x11 & n5747 ;
  assign n5750 = x11 & n5740 ;
  assign n5751 = ( x11 & n5744 ) | ( x11 & n5750 ) | ( n5744 & n5750 ) ;
  assign n5752 = ( n3282 & n5749 ) | ( n3282 & n5751 ) | ( n5749 & n5751 ) ;
  assign n5753 = x11 & ~n5751 ;
  assign n5754 = x11 & ~n5747 ;
  assign n5755 = ( ~n3282 & n5753 ) | ( ~n3282 & n5754 ) | ( n5753 & n5754 ) ;
  assign n5756 = ( n5748 & ~n5752 ) | ( n5748 & n5755 ) | ( ~n5752 & n5755 ) ;
  assign n5757 = n5739 & n5756 ;
  assign n5758 = n5739 | n5756 ;
  assign n5759 = ~n5757 & n5758 ;
  assign n5760 = n5427 | n5431 ;
  assign n5761 = n5759 & n5760 ;
  assign n5762 = n5760 & ~n5761 ;
  assign n5763 = ( n5759 & ~n5761 ) | ( n5759 & n5762 ) | ( ~n5761 & n5762 ) ;
  assign n5764 = x92 & n389 ;
  assign n5765 = x91 & n384 ;
  assign n5766 = x90 & ~n383 ;
  assign n5767 = n463 & n5766 ;
  assign n5768 = n5765 | n5767 ;
  assign n5769 = n5764 | n5768 ;
  assign n5770 = n392 | n5764 ;
  assign n5771 = n5768 | n5770 ;
  assign n5772 = ( n4040 & n5769 ) | ( n4040 & n5771 ) | ( n5769 & n5771 ) ;
  assign n5773 = x8 & n5771 ;
  assign n5774 = x8 & n5764 ;
  assign n5775 = ( x8 & n5768 ) | ( x8 & n5774 ) | ( n5768 & n5774 ) ;
  assign n5776 = ( n4040 & n5773 ) | ( n4040 & n5775 ) | ( n5773 & n5775 ) ;
  assign n5777 = x8 & ~n5775 ;
  assign n5778 = x8 & ~n5771 ;
  assign n5779 = ( ~n4040 & n5777 ) | ( ~n4040 & n5778 ) | ( n5777 & n5778 ) ;
  assign n5780 = ( n5772 & ~n5776 ) | ( n5772 & n5779 ) | ( ~n5776 & n5779 ) ;
  assign n5781 = n5759 & n5780 ;
  assign n5782 = ~n5759 & n5780 ;
  assign n5783 = ( ~n5760 & n5780 ) | ( ~n5760 & n5782 ) | ( n5780 & n5782 ) ;
  assign n5784 = ( n5762 & n5781 ) | ( n5762 & n5783 ) | ( n5781 & n5783 ) ;
  assign n5785 = n5763 & ~n5784 ;
  assign n5786 = n5760 & n5781 ;
  assign n5787 = ( ~n5762 & n5782 ) | ( ~n5762 & n5786 ) | ( n5782 & n5786 ) ;
  assign n5788 = n5785 | n5787 ;
  assign n5789 = n5451 | n5453 ;
  assign n5790 = n5452 | n5789 ;
  assign n5791 = ( n5451 & n5455 ) | ( n5451 & n5790 ) | ( n5455 & n5790 ) ;
  assign n5792 = n5788 | n5791 ;
  assign n5793 = n5788 & n5791 ;
  assign n5794 = n5792 & ~n5793 ;
  assign n5795 = x95 & n212 ;
  assign n5796 = x94 & n207 ;
  assign n5797 = x93 & ~n206 ;
  assign n5798 = n267 & n5797 ;
  assign n5799 = n5796 | n5798 ;
  assign n5800 = n5795 | n5799 ;
  assign n5801 = n215 | n5795 ;
  assign n5802 = n5799 | n5801 ;
  assign n5803 = ( n4897 & n5800 ) | ( n4897 & n5802 ) | ( n5800 & n5802 ) ;
  assign n5804 = x5 & n5802 ;
  assign n5805 = x5 & n5795 ;
  assign n5806 = ( x5 & n5799 ) | ( x5 & n5805 ) | ( n5799 & n5805 ) ;
  assign n5807 = ( n4897 & n5804 ) | ( n4897 & n5806 ) | ( n5804 & n5806 ) ;
  assign n5808 = x5 & ~n5806 ;
  assign n5809 = x5 & ~n5802 ;
  assign n5810 = ( ~n4897 & n5808 ) | ( ~n4897 & n5809 ) | ( n5808 & n5809 ) ;
  assign n5811 = ( n5803 & ~n5807 ) | ( n5803 & n5810 ) | ( ~n5807 & n5810 ) ;
  assign n5812 = n5794 & n5811 ;
  assign n5813 = n5794 | n5811 ;
  assign n5814 = ~n5812 & n5813 ;
  assign n5815 = n5476 & n5813 ;
  assign n5816 = ~n5812 & n5815 ;
  assign n5817 = ( n5528 & n5814 ) | ( n5528 & n5816 ) | ( n5814 & n5816 ) ;
  assign n5818 = n5529 & ~n5817 ;
  assign n5819 = n5814 & ~n5815 ;
  assign n5820 = ~n5813 & n5814 ;
  assign n5821 = ( ~n5528 & n5819 ) | ( ~n5528 & n5820 ) | ( n5819 & n5820 ) ;
  assign n5822 = n5818 | n5821 ;
  assign n5823 = ( n1493 & n3274 ) | ( n1493 & n3276 ) | ( n3274 & n3276 ) ;
  assign n5824 = x97 | x98 ;
  assign n5825 = x97 & x98 ;
  assign n5826 = n5824 & ~n5825 ;
  assign n5827 = n5484 | n5491 ;
  assign n5828 = n5484 | n5485 ;
  assign n5829 = ( n5484 & n5487 ) | ( n5484 & n5828 ) | ( n5487 & n5828 ) ;
  assign n5830 = ( n5184 & n5827 ) | ( n5184 & n5829 ) | ( n5827 & n5829 ) ;
  assign n5831 = n5826 | n5830 ;
  assign n5832 = ( n5186 & n5827 ) | ( n5186 & n5829 ) | ( n5827 & n5829 ) ;
  assign n5833 = n5826 | n5832 ;
  assign n5834 = ( n5823 & n5831 ) | ( n5823 & n5833 ) | ( n5831 & n5833 ) ;
  assign n5835 = x97 & n133 ;
  assign n5836 = x96 & ~n162 ;
  assign n5837 = ( n137 & n5835 ) | ( n137 & n5836 ) | ( n5835 & n5836 ) ;
  assign n5838 = x0 & x98 ;
  assign n5839 = ( ~n137 & n5835 ) | ( ~n137 & n5838 ) | ( n5835 & n5838 ) ;
  assign n5840 = n5837 | n5839 ;
  assign n5841 = n141 | n5840 ;
  assign n5842 = n5484 & n5826 ;
  assign n5843 = ( n5491 & n5826 ) | ( n5491 & n5842 ) | ( n5826 & n5842 ) ;
  assign n5844 = n5826 & n5828 ;
  assign n5845 = ( n5487 & n5842 ) | ( n5487 & n5844 ) | ( n5842 & n5844 ) ;
  assign n5846 = ( n5184 & n5843 ) | ( n5184 & n5845 ) | ( n5843 & n5845 ) ;
  assign n5847 = ( n5186 & n5843 ) | ( n5186 & n5845 ) | ( n5843 & n5845 ) ;
  assign n5848 = ( n3274 & n5846 ) | ( n3274 & n5847 ) | ( n5846 & n5847 ) ;
  assign n5849 = ( n3276 & n5846 ) | ( n3276 & n5847 ) | ( n5846 & n5847 ) ;
  assign n5850 = ( n1493 & n5848 ) | ( n1493 & n5849 ) | ( n5848 & n5849 ) ;
  assign n5851 = ( n5840 & n5841 ) | ( n5840 & ~n5850 ) | ( n5841 & ~n5850 ) ;
  assign n5852 = n5840 & n5841 ;
  assign n5853 = ( n5834 & n5851 ) | ( n5834 & n5852 ) | ( n5851 & n5852 ) ;
  assign n5854 = x2 & n5840 ;
  assign n5855 = ( x2 & n523 ) | ( x2 & n5840 ) | ( n523 & n5840 ) ;
  assign n5856 = ( ~n5850 & n5854 ) | ( ~n5850 & n5855 ) | ( n5854 & n5855 ) ;
  assign n5857 = n5854 & n5855 ;
  assign n5858 = ( n5834 & n5856 ) | ( n5834 & n5857 ) | ( n5856 & n5857 ) ;
  assign n5859 = x2 & ~n5855 ;
  assign n5860 = x2 & ~n5840 ;
  assign n5861 = ( n5850 & n5859 ) | ( n5850 & n5860 ) | ( n5859 & n5860 ) ;
  assign n5862 = n5859 | n5860 ;
  assign n5863 = ( ~n5834 & n5861 ) | ( ~n5834 & n5862 ) | ( n5861 & n5862 ) ;
  assign n5864 = ( n5853 & ~n5858 ) | ( n5853 & n5863 ) | ( ~n5858 & n5863 ) ;
  assign n5865 = n5821 | n5864 ;
  assign n5866 = n5818 | n5865 ;
  assign n5867 = ~n5864 & n5866 ;
  assign n5868 = ( ~n5822 & n5866 ) | ( ~n5822 & n5867 ) | ( n5866 & n5867 ) ;
  assign n5869 = n5521 | n5526 ;
  assign n5870 = n5868 & n5869 ;
  assign n5871 = n5868 | n5869 ;
  assign n5872 = ~n5870 & n5871 ;
  assign n5873 = n5704 | n5711 ;
  assign n5874 = x78 & n2429 ;
  assign n5875 = x77 & n2424 ;
  assign n5876 = x76 & ~n2423 ;
  assign n5877 = n2631 & n5876 ;
  assign n5878 = n5875 | n5877 ;
  assign n5879 = n5874 | n5878 ;
  assign n5880 = n2432 | n5874 ;
  assign n5881 = n5878 | n5880 ;
  assign n5882 = ( n1192 & n5879 ) | ( n1192 & n5881 ) | ( n5879 & n5881 ) ;
  assign n5883 = x23 & n5881 ;
  assign n5884 = x23 & n5874 ;
  assign n5885 = ( x23 & n5878 ) | ( x23 & n5884 ) | ( n5878 & n5884 ) ;
  assign n5886 = ( n1192 & n5883 ) | ( n1192 & n5885 ) | ( n5883 & n5885 ) ;
  assign n5887 = x23 & ~n5885 ;
  assign n5888 = x23 & ~n5881 ;
  assign n5889 = ( ~n1192 & n5887 ) | ( ~n1192 & n5888 ) | ( n5887 & n5888 ) ;
  assign n5890 = ( n5882 & ~n5886 ) | ( n5882 & n5889 ) | ( ~n5886 & n5889 ) ;
  assign n5891 = x66 & n5554 ;
  assign n5892 = x65 & n5549 ;
  assign n5893 = ~n5232 & n5553 ;
  assign n5894 = x64 & ~n5548 ;
  assign n5895 = n5893 & n5894 ;
  assign n5896 = n5892 | n5895 ;
  assign n5897 = n5891 | n5896 ;
  assign n5898 = n159 & n5557 ;
  assign n5899 = n5897 | n5898 ;
  assign n5900 = x35 | n5557 ;
  assign n5901 = ( x35 & n159 ) | ( x35 & n5900 ) | ( n159 & n5900 ) ;
  assign n5902 = n5897 | n5901 ;
  assign n5903 = ~x35 & n5901 ;
  assign n5904 = ( ~x35 & n5897 ) | ( ~x35 & n5903 ) | ( n5897 & n5903 ) ;
  assign n5905 = ( ~n5899 & n5902 ) | ( ~n5899 & n5904 ) | ( n5902 & n5904 ) ;
  assign n5906 = n5569 | n5905 ;
  assign n5907 = n5569 & n5905 ;
  assign n5908 = n5906 & ~n5907 ;
  assign n5909 = n293 & n4634 ;
  assign n5910 = x69 & n4631 ;
  assign n5911 = x68 & n4626 ;
  assign n5912 = x67 & ~n4625 ;
  assign n5913 = n4943 & n5912 ;
  assign n5914 = n5911 | n5913 ;
  assign n5915 = n5910 | n5914 ;
  assign n5916 = n5909 | n5915 ;
  assign n5917 = x32 | n5910 ;
  assign n5918 = n5914 | n5917 ;
  assign n5919 = n5909 | n5918 ;
  assign n5920 = ~x32 & n5918 ;
  assign n5921 = ( ~x32 & n5909 ) | ( ~x32 & n5920 ) | ( n5909 & n5920 ) ;
  assign n5922 = ( ~n5916 & n5919 ) | ( ~n5916 & n5921 ) | ( n5919 & n5921 ) ;
  assign n5923 = n5908 | n5922 ;
  assign n5924 = n5908 & n5922 ;
  assign n5925 = n5923 & ~n5924 ;
  assign n5926 = n5591 | n5593 ;
  assign n5927 = ( n5591 & n5592 ) | ( n5591 & n5926 ) | ( n5592 & n5926 ) ;
  assign n5928 = ~n5925 & n5927 ;
  assign n5929 = n5925 & n5927 ;
  assign n5930 = n5925 & ~n5929 ;
  assign n5931 = n5928 | n5930 ;
  assign n5932 = x72 & n3816 ;
  assign n5933 = x71 & n3811 ;
  assign n5934 = x70 & ~n3810 ;
  assign n5935 = n4067 & n5934 ;
  assign n5936 = n5933 | n5935 ;
  assign n5937 = n5932 | n5936 ;
  assign n5938 = ( n513 & n3819 ) | ( n513 & n5937 ) | ( n3819 & n5937 ) ;
  assign n5939 = ( x29 & n3819 ) | ( x29 & ~n5932 ) | ( n3819 & ~n5932 ) ;
  assign n5940 = x29 & n3819 ;
  assign n5941 = ( ~n5936 & n5939 ) | ( ~n5936 & n5940 ) | ( n5939 & n5940 ) ;
  assign n5942 = ( x29 & n513 ) | ( x29 & n5941 ) | ( n513 & n5941 ) ;
  assign n5943 = ~n5938 & n5942 ;
  assign n5944 = n5937 | n5941 ;
  assign n5945 = x29 | n5937 ;
  assign n5946 = ( n513 & n5944 ) | ( n513 & n5945 ) | ( n5944 & n5945 ) ;
  assign n5947 = ( ~x29 & n5943 ) | ( ~x29 & n5946 ) | ( n5943 & n5946 ) ;
  assign n5948 = n5928 & n5947 ;
  assign n5949 = ( n5930 & n5947 ) | ( n5930 & n5948 ) | ( n5947 & n5948 ) ;
  assign n5950 = n5931 & ~n5949 ;
  assign n5951 = ~n5928 & n5947 ;
  assign n5952 = ~n5930 & n5951 ;
  assign n5953 = n5950 | n5952 ;
  assign n5954 = n5598 | n5599 ;
  assign n5955 = ( n5598 & n5605 ) | ( n5598 & n5954 ) | ( n5605 & n5954 ) ;
  assign n5956 = n5953 & n5955 ;
  assign n5957 = n5953 | n5955 ;
  assign n5958 = ~n5956 & n5957 ;
  assign n5959 = x75 & n3085 ;
  assign n5960 = x74 & n3080 ;
  assign n5961 = x73 & ~n3079 ;
  assign n5962 = n3309 & n5961 ;
  assign n5963 = n5960 | n5962 ;
  assign n5964 = n5959 | n5963 ;
  assign n5965 = n3088 | n5959 ;
  assign n5966 = n5963 | n5965 ;
  assign n5967 = ( n746 & n5964 ) | ( n746 & n5966 ) | ( n5964 & n5966 ) ;
  assign n5968 = x26 & n5966 ;
  assign n5969 = x26 & n5959 ;
  assign n5970 = ( x26 & n5963 ) | ( x26 & n5969 ) | ( n5963 & n5969 ) ;
  assign n5971 = ( n746 & n5968 ) | ( n746 & n5970 ) | ( n5968 & n5970 ) ;
  assign n5972 = x26 & ~n5970 ;
  assign n5973 = x26 & ~n5966 ;
  assign n5974 = ( ~n746 & n5972 ) | ( ~n746 & n5973 ) | ( n5972 & n5973 ) ;
  assign n5975 = ( n5967 & ~n5971 ) | ( n5967 & n5974 ) | ( ~n5971 & n5974 ) ;
  assign n5976 = n5958 & n5975 ;
  assign n5977 = n5958 & ~n5976 ;
  assign n5978 = ~n5958 & n5975 ;
  assign n5979 = n5977 | n5978 ;
  assign n5980 = n5626 | n5630 ;
  assign n5981 = ( n5626 & n5629 ) | ( n5626 & n5980 ) | ( n5629 & n5980 ) ;
  assign n5982 = ~n5979 & n5981 ;
  assign n5983 = n5890 & n5982 ;
  assign n5984 = n5979 & ~n5981 ;
  assign n5985 = ( n5890 & n5983 ) | ( n5890 & n5984 ) | ( n5983 & n5984 ) ;
  assign n5986 = n5890 | n5982 ;
  assign n5987 = n5984 | n5986 ;
  assign n5988 = ~n5985 & n5987 ;
  assign n5989 = n5651 | n5655 ;
  assign n5990 = ( n5651 & n5653 ) | ( n5651 & n5989 ) | ( n5653 & n5989 ) ;
  assign n5991 = n5988 & n5990 ;
  assign n5992 = n5988 | n5990 ;
  assign n5993 = ~n5991 & n5992 ;
  assign n5994 = x81 & n1859 ;
  assign n5995 = x80 & n1854 ;
  assign n5996 = x79 & ~n1853 ;
  assign n5997 = n2037 & n5996 ;
  assign n5998 = n5995 | n5997 ;
  assign n5999 = n5994 | n5998 ;
  assign n6000 = n1862 | n5994 ;
  assign n6001 = n5998 | n6000 ;
  assign n6002 = ( n1651 & n5999 ) | ( n1651 & n6001 ) | ( n5999 & n6001 ) ;
  assign n6003 = x20 & n6001 ;
  assign n6004 = x20 & n5994 ;
  assign n6005 = ( x20 & n5998 ) | ( x20 & n6004 ) | ( n5998 & n6004 ) ;
  assign n6006 = ( n1651 & n6003 ) | ( n1651 & n6005 ) | ( n6003 & n6005 ) ;
  assign n6007 = x20 & ~n6005 ;
  assign n6008 = x20 & ~n6001 ;
  assign n6009 = ( ~n1651 & n6007 ) | ( ~n1651 & n6008 ) | ( n6007 & n6008 ) ;
  assign n6010 = ( n6002 & ~n6006 ) | ( n6002 & n6009 ) | ( ~n6006 & n6009 ) ;
  assign n6011 = n5993 & n6010 ;
  assign n6012 = n5993 & ~n6011 ;
  assign n6013 = ~n5993 & n6010 ;
  assign n6014 = n6012 | n6013 ;
  assign n6015 = n5676 | n5683 ;
  assign n6016 = n6014 | n6015 ;
  assign n6017 = n6014 & n6015 ;
  assign n6018 = n6016 & ~n6017 ;
  assign n6019 = x84 & n1383 ;
  assign n6020 = x83 & n1378 ;
  assign n6021 = x82 & ~n1377 ;
  assign n6022 = n1542 & n6021 ;
  assign n6023 = n6020 | n6022 ;
  assign n6024 = n6019 | n6023 ;
  assign n6025 = n1386 | n6019 ;
  assign n6026 = n6023 | n6025 ;
  assign n6027 = ( n2194 & n6024 ) | ( n2194 & n6026 ) | ( n6024 & n6026 ) ;
  assign n6028 = x17 & n6026 ;
  assign n6029 = x17 & n6019 ;
  assign n6030 = ( x17 & n6023 ) | ( x17 & n6029 ) | ( n6023 & n6029 ) ;
  assign n6031 = ( n2194 & n6028 ) | ( n2194 & n6030 ) | ( n6028 & n6030 ) ;
  assign n6032 = x17 & ~n6030 ;
  assign n6033 = x17 & ~n6026 ;
  assign n6034 = ( ~n2194 & n6032 ) | ( ~n2194 & n6033 ) | ( n6032 & n6033 ) ;
  assign n6035 = ( n6027 & ~n6031 ) | ( n6027 & n6034 ) | ( ~n6031 & n6034 ) ;
  assign n6036 = n6018 & n6035 ;
  assign n6037 = n6018 | n6035 ;
  assign n6038 = ~n6036 & n6037 ;
  assign n6039 = n5873 & n6038 ;
  assign n6040 = n5873 & ~n6039 ;
  assign n6041 = x87 & n962 ;
  assign n6042 = x86 & n957 ;
  assign n6043 = x85 & ~n956 ;
  assign n6044 = n1105 & n6043 ;
  assign n6045 = n6042 | n6044 ;
  assign n6046 = n6041 | n6045 ;
  assign n6047 = n965 | n6041 ;
  assign n6048 = n6045 | n6047 ;
  assign n6049 = ( n2816 & n6046 ) | ( n2816 & n6048 ) | ( n6046 & n6048 ) ;
  assign n6050 = x14 & n6048 ;
  assign n6051 = x14 & n6041 ;
  assign n6052 = ( x14 & n6045 ) | ( x14 & n6051 ) | ( n6045 & n6051 ) ;
  assign n6053 = ( n2816 & n6050 ) | ( n2816 & n6052 ) | ( n6050 & n6052 ) ;
  assign n6054 = x14 & ~n6052 ;
  assign n6055 = x14 & ~n6048 ;
  assign n6056 = ( ~n2816 & n6054 ) | ( ~n2816 & n6055 ) | ( n6054 & n6055 ) ;
  assign n6057 = ( n6049 & ~n6053 ) | ( n6049 & n6056 ) | ( ~n6053 & n6056 ) ;
  assign n6058 = n6038 & n6057 ;
  assign n6059 = ~n6038 & n6057 ;
  assign n6060 = ( ~n5873 & n6057 ) | ( ~n5873 & n6059 ) | ( n6057 & n6059 ) ;
  assign n6061 = ( n6040 & n6058 ) | ( n6040 & n6060 ) | ( n6058 & n6060 ) ;
  assign n6062 = n6038 | n6057 ;
  assign n6063 = n6038 & ~n6057 ;
  assign n6064 = n5873 & n6063 ;
  assign n6065 = ( n6040 & n6062 ) | ( n6040 & ~n6064 ) | ( n6062 & ~n6064 ) ;
  assign n6066 = ~n6061 & n6065 ;
  assign n6067 = n5730 | n5736 ;
  assign n6068 = ( n5730 & n5733 ) | ( n5730 & n6067 ) | ( n5733 & n6067 ) ;
  assign n6069 = n6066 & n6068 ;
  assign n6070 = n6066 | n6068 ;
  assign n6071 = ~n6069 & n6070 ;
  assign n6072 = x90 & n636 ;
  assign n6073 = x89 & n631 ;
  assign n6074 = x88 & ~n630 ;
  assign n6075 = n764 & n6074 ;
  assign n6076 = n6073 | n6075 ;
  assign n6077 = n6072 | n6076 ;
  assign n6078 = n639 | n6072 ;
  assign n6079 = n6076 | n6078 ;
  assign n6080 = ( n3519 & n6077 ) | ( n3519 & n6079 ) | ( n6077 & n6079 ) ;
  assign n6081 = x11 & n6079 ;
  assign n6082 = x11 & n6072 ;
  assign n6083 = ( x11 & n6076 ) | ( x11 & n6082 ) | ( n6076 & n6082 ) ;
  assign n6084 = ( n3519 & n6081 ) | ( n3519 & n6083 ) | ( n6081 & n6083 ) ;
  assign n6085 = x11 & ~n6083 ;
  assign n6086 = x11 & ~n6079 ;
  assign n6087 = ( ~n3519 & n6085 ) | ( ~n3519 & n6086 ) | ( n6085 & n6086 ) ;
  assign n6088 = ( n6080 & ~n6084 ) | ( n6080 & n6087 ) | ( ~n6084 & n6087 ) ;
  assign n6089 = n6071 | n6088 ;
  assign n6090 = n6071 & n6088 ;
  assign n6091 = n6089 & ~n6090 ;
  assign n6092 = n5757 | n5759 ;
  assign n6093 = ( n5757 & n5760 ) | ( n5757 & n6092 ) | ( n5760 & n6092 ) ;
  assign n6094 = n6091 & n6093 ;
  assign n6095 = n6091 | n6093 ;
  assign n6096 = ~n6094 & n6095 ;
  assign n6097 = x93 & n389 ;
  assign n6098 = x92 & n384 ;
  assign n6099 = x91 & ~n383 ;
  assign n6100 = n463 & n6099 ;
  assign n6101 = n6098 | n6100 ;
  assign n6102 = n6097 | n6101 ;
  assign n6103 = n392 | n6097 ;
  assign n6104 = n6101 | n6103 ;
  assign n6105 = ( n4305 & n6102 ) | ( n4305 & n6104 ) | ( n6102 & n6104 ) ;
  assign n6106 = x8 & n6104 ;
  assign n6107 = x8 & n6097 ;
  assign n6108 = ( x8 & n6101 ) | ( x8 & n6107 ) | ( n6101 & n6107 ) ;
  assign n6109 = ( n4305 & n6106 ) | ( n4305 & n6108 ) | ( n6106 & n6108 ) ;
  assign n6110 = x8 & ~n6108 ;
  assign n6111 = x8 & ~n6104 ;
  assign n6112 = ( ~n4305 & n6110 ) | ( ~n4305 & n6111 ) | ( n6110 & n6111 ) ;
  assign n6113 = ( n6105 & ~n6109 ) | ( n6105 & n6112 ) | ( ~n6109 & n6112 ) ;
  assign n6114 = n6096 & n6113 ;
  assign n6115 = n6096 & ~n6114 ;
  assign n6116 = ~n6096 & n6113 ;
  assign n6117 = n6115 | n6116 ;
  assign n6118 = n5784 | n5793 ;
  assign n6119 = n6117 | n6118 ;
  assign n6120 = n6117 & n6118 ;
  assign n6121 = n6119 & ~n6120 ;
  assign n6122 = x96 & n212 ;
  assign n6123 = x95 & n207 ;
  assign n6124 = x94 & ~n206 ;
  assign n6125 = n267 & n6124 ;
  assign n6126 = n6123 | n6125 ;
  assign n6127 = n6122 | n6126 ;
  assign n6128 = n215 | n6122 ;
  assign n6129 = n6126 | n6128 ;
  assign n6130 = ( n5202 & n6127 ) | ( n5202 & n6129 ) | ( n6127 & n6129 ) ;
  assign n6131 = x5 & n6129 ;
  assign n6132 = x5 & n6122 ;
  assign n6133 = ( x5 & n6126 ) | ( x5 & n6132 ) | ( n6126 & n6132 ) ;
  assign n6134 = ( n5202 & n6131 ) | ( n5202 & n6133 ) | ( n6131 & n6133 ) ;
  assign n6135 = x5 & ~n6133 ;
  assign n6136 = x5 & ~n6129 ;
  assign n6137 = ( ~n5202 & n6135 ) | ( ~n5202 & n6136 ) | ( n6135 & n6136 ) ;
  assign n6138 = ( n6130 & ~n6134 ) | ( n6130 & n6137 ) | ( ~n6134 & n6137 ) ;
  assign n6139 = n6121 & n6138 ;
  assign n6140 = n6121 | n6138 ;
  assign n6141 = ~n6139 & n6140 ;
  assign n6142 = n5812 | n5815 ;
  assign n6143 = n5812 | n5813 ;
  assign n6144 = ( n5528 & n6142 ) | ( n5528 & n6143 ) | ( n6142 & n6143 ) ;
  assign n6145 = n6141 & n6144 ;
  assign n6146 = n6144 & ~n6145 ;
  assign n6147 = ( n6141 & ~n6145 ) | ( n6141 & n6146 ) | ( ~n6145 & n6146 ) ;
  assign n6148 = x98 | x99 ;
  assign n6149 = x98 & x99 ;
  assign n6150 = n6148 & ~n6149 ;
  assign n6151 = n5825 | n5845 ;
  assign n6152 = n5825 | n5826 ;
  assign n6153 = n5484 | n5825 ;
  assign n6154 = ( n5825 & n5826 ) | ( n5825 & n6153 ) | ( n5826 & n6153 ) ;
  assign n6155 = ( n5491 & n6152 ) | ( n5491 & n6154 ) | ( n6152 & n6154 ) ;
  assign n6156 = ( n5184 & n6151 ) | ( n5184 & n6155 ) | ( n6151 & n6155 ) ;
  assign n6157 = n6150 & n6156 ;
  assign n6158 = ( n5186 & n6151 ) | ( n5186 & n6155 ) | ( n6151 & n6155 ) ;
  assign n6159 = n6150 & n6158 ;
  assign n6160 = ( n5823 & n6157 ) | ( n5823 & n6159 ) | ( n6157 & n6159 ) ;
  assign n6161 = n6150 | n6156 ;
  assign n6162 = n6150 | n6158 ;
  assign n6163 = ( n5823 & n6161 ) | ( n5823 & n6162 ) | ( n6161 & n6162 ) ;
  assign n6164 = ~n6160 & n6163 ;
  assign n6165 = x98 & n133 ;
  assign n6166 = x97 & ~n162 ;
  assign n6167 = ( n137 & n6165 ) | ( n137 & n6166 ) | ( n6165 & n6166 ) ;
  assign n6168 = x0 & x99 ;
  assign n6169 = ( ~n137 & n6165 ) | ( ~n137 & n6168 ) | ( n6165 & n6168 ) ;
  assign n6170 = n6167 | n6169 ;
  assign n6171 = n141 | n6170 ;
  assign n6172 = ( n6164 & n6170 ) | ( n6164 & n6171 ) | ( n6170 & n6171 ) ;
  assign n6173 = x2 & n6170 ;
  assign n6174 = ( x2 & n523 ) | ( x2 & n6170 ) | ( n523 & n6170 ) ;
  assign n6175 = ( n6164 & n6173 ) | ( n6164 & n6174 ) | ( n6173 & n6174 ) ;
  assign n6176 = x2 & ~n6174 ;
  assign n6177 = x2 & ~n6170 ;
  assign n6178 = ( ~n6164 & n6176 ) | ( ~n6164 & n6177 ) | ( n6176 & n6177 ) ;
  assign n6179 = ( n6172 & ~n6175 ) | ( n6172 & n6178 ) | ( ~n6175 & n6178 ) ;
  assign n6180 = n6147 & ~n6179 ;
  assign n6181 = ~n6147 & n6179 ;
  assign n6182 = n6180 | n6181 ;
  assign n6183 = ~n5821 & n5864 ;
  assign n6184 = ~n5818 & n6183 ;
  assign n6185 = ( n5864 & n5870 ) | ( n5864 & ~n6184 ) | ( n5870 & ~n6184 ) ;
  assign n6186 = n6182 & n6185 ;
  assign n6187 = n6182 | n6185 ;
  assign n6188 = ~n6186 & n6187 ;
  assign n6189 = n6139 | n6145 ;
  assign n6190 = n6061 | n6069 ;
  assign n6191 = n5985 | n5991 ;
  assign n6192 = n5924 | n5929 ;
  assign n6193 = x35 & ~x36 ;
  assign n6194 = ~x35 & x36 ;
  assign n6195 = n6193 | n6194 ;
  assign n6196 = x64 & n6195 ;
  assign n6197 = ~n5569 & n6196 ;
  assign n6198 = ( ~n5905 & n6196 ) | ( ~n5905 & n6197 ) | ( n6196 & n6197 ) ;
  assign n6199 = n5569 & ~n6196 ;
  assign n6200 = n5905 & n6199 ;
  assign n6201 = n6198 | n6200 ;
  assign n6202 = x67 & n5554 ;
  assign n6203 = x66 & n5549 ;
  assign n6204 = x65 & ~n5548 ;
  assign n6205 = n5893 & n6204 ;
  assign n6206 = n6203 | n6205 ;
  assign n6207 = n6202 | n6206 ;
  assign n6208 = n186 & n5557 ;
  assign n6209 = n6207 | n6208 ;
  assign n6210 = x35 & ~n6209 ;
  assign n6211 = ~x35 & n6209 ;
  assign n6212 = n6210 | n6211 ;
  assign n6213 = n6201 & n6212 ;
  assign n6214 = n6201 | n6212 ;
  assign n6215 = ~n6213 & n6214 ;
  assign n6216 = x69 & n4626 ;
  assign n6217 = x68 & ~n4625 ;
  assign n6218 = n4943 & n6217 ;
  assign n6219 = n6216 | n6218 ;
  assign n6220 = x70 & n4631 ;
  assign n6221 = n4634 | n6220 ;
  assign n6222 = n6219 | n6221 ;
  assign n6223 = x32 & ~n6222 ;
  assign n6224 = x32 & ~n6220 ;
  assign n6225 = ~n6219 & n6224 ;
  assign n6226 = ( ~n340 & n6223 ) | ( ~n340 & n6225 ) | ( n6223 & n6225 ) ;
  assign n6227 = ~x32 & n6222 ;
  assign n6228 = ~x32 & n6220 ;
  assign n6229 = ( ~x32 & n6219 ) | ( ~x32 & n6228 ) | ( n6219 & n6228 ) ;
  assign n6230 = ( n340 & n6227 ) | ( n340 & n6229 ) | ( n6227 & n6229 ) ;
  assign n6231 = n6226 | n6230 ;
  assign n6232 = ( n5924 & ~n6215 ) | ( n5924 & n6231 ) | ( ~n6215 & n6231 ) ;
  assign n6233 = n6215 & ~n6231 ;
  assign n6234 = ( n5929 & n6232 ) | ( n5929 & ~n6233 ) | ( n6232 & ~n6233 ) ;
  assign n6235 = ( ~n6192 & n6215 ) | ( ~n6192 & n6234 ) | ( n6215 & n6234 ) ;
  assign n6236 = x73 & n3816 ;
  assign n6237 = x72 & n3811 ;
  assign n6238 = x71 & ~n3810 ;
  assign n6239 = n4067 & n6238 ;
  assign n6240 = n6237 | n6239 ;
  assign n6241 = n6236 | n6240 ;
  assign n6242 = ( ~n610 & n3819 ) | ( ~n610 & n6241 ) | ( n3819 & n6241 ) ;
  assign n6243 = n3819 & n6236 ;
  assign n6244 = ( n3819 & n6240 ) | ( n3819 & n6243 ) | ( n6240 & n6243 ) ;
  assign n6245 = ( n598 & n6242 ) | ( n598 & n6244 ) | ( n6242 & n6244 ) ;
  assign n6246 = ( x29 & ~n6241 ) | ( x29 & n6245 ) | ( ~n6241 & n6245 ) ;
  assign n6247 = ~n6245 & n6246 ;
  assign n6248 = x29 | n6236 ;
  assign n6249 = n6240 | n6248 ;
  assign n6250 = n6245 | n6249 ;
  assign n6251 = ( ~x29 & n6247 ) | ( ~x29 & n6250 ) | ( n6247 & n6250 ) ;
  assign n6252 = n6234 & n6251 ;
  assign n6253 = ~n6231 & n6250 ;
  assign n6254 = x29 | n6231 ;
  assign n6255 = ( n6247 & n6253 ) | ( n6247 & ~n6254 ) | ( n6253 & ~n6254 ) ;
  assign n6256 = ( n6235 & n6252 ) | ( n6235 & n6255 ) | ( n6252 & n6255 ) ;
  assign n6257 = n6234 | n6251 ;
  assign n6258 = n6231 & ~n6250 ;
  assign n6259 = x29 & n6231 ;
  assign n6260 = ( ~n6247 & n6258 ) | ( ~n6247 & n6259 ) | ( n6258 & n6259 ) ;
  assign n6261 = ( n6235 & n6257 ) | ( n6235 & ~n6260 ) | ( n6257 & ~n6260 ) ;
  assign n6262 = ~n6256 & n6261 ;
  assign n6263 = n5949 & n6262 ;
  assign n6264 = ( n5956 & n6262 ) | ( n5956 & n6263 ) | ( n6262 & n6263 ) ;
  assign n6265 = n5949 | n6262 ;
  assign n6266 = n5956 | n6265 ;
  assign n6267 = ~n6264 & n6266 ;
  assign n6268 = x76 & n3085 ;
  assign n6269 = x75 & n3080 ;
  assign n6270 = x74 & ~n3079 ;
  assign n6271 = n3309 & n6270 ;
  assign n6272 = n6269 | n6271 ;
  assign n6273 = n6268 | n6272 ;
  assign n6274 = n3088 | n6268 ;
  assign n6275 = n6272 | n6274 ;
  assign n6276 = ( n923 & n6273 ) | ( n923 & n6275 ) | ( n6273 & n6275 ) ;
  assign n6277 = x26 & n6275 ;
  assign n6278 = x26 & n6268 ;
  assign n6279 = ( x26 & n6272 ) | ( x26 & n6278 ) | ( n6272 & n6278 ) ;
  assign n6280 = ( n923 & n6277 ) | ( n923 & n6279 ) | ( n6277 & n6279 ) ;
  assign n6281 = x26 & ~n6279 ;
  assign n6282 = x26 & ~n6275 ;
  assign n6283 = ( ~n923 & n6281 ) | ( ~n923 & n6282 ) | ( n6281 & n6282 ) ;
  assign n6284 = ( n6276 & ~n6280 ) | ( n6276 & n6283 ) | ( ~n6280 & n6283 ) ;
  assign n6285 = n6267 | n6284 ;
  assign n6286 = n6267 & n6284 ;
  assign n6287 = n6285 & ~n6286 ;
  assign n6288 = n5979 & n5981 ;
  assign n6289 = n5976 & n6287 ;
  assign n6290 = ( n6287 & n6288 ) | ( n6287 & n6289 ) | ( n6288 & n6289 ) ;
  assign n6291 = n5976 | n6287 ;
  assign n6292 = n6288 | n6291 ;
  assign n6293 = ~n6290 & n6292 ;
  assign n6294 = x79 & n2429 ;
  assign n6295 = x78 & n2424 ;
  assign n6296 = x77 & ~n2423 ;
  assign n6297 = n2631 & n6296 ;
  assign n6298 = n6295 | n6297 ;
  assign n6299 = n6294 | n6298 ;
  assign n6300 = n2432 | n6294 ;
  assign n6301 = n6298 | n6300 ;
  assign n6302 = ( n1332 & n6299 ) | ( n1332 & n6301 ) | ( n6299 & n6301 ) ;
  assign n6303 = x23 & n6301 ;
  assign n6304 = x23 & n6294 ;
  assign n6305 = ( x23 & n6298 ) | ( x23 & n6304 ) | ( n6298 & n6304 ) ;
  assign n6306 = ( n1332 & n6303 ) | ( n1332 & n6305 ) | ( n6303 & n6305 ) ;
  assign n6307 = x23 & ~n6305 ;
  assign n6308 = x23 & ~n6301 ;
  assign n6309 = ( ~n1332 & n6307 ) | ( ~n1332 & n6308 ) | ( n6307 & n6308 ) ;
  assign n6310 = ( n6302 & ~n6306 ) | ( n6302 & n6309 ) | ( ~n6306 & n6309 ) ;
  assign n6311 = n6293 & n6310 ;
  assign n6312 = n6293 & ~n6311 ;
  assign n6313 = ~n6293 & n6310 ;
  assign n6314 = n6312 | n6313 ;
  assign n6315 = n6191 & ~n6314 ;
  assign n6316 = ~n6191 & n6314 ;
  assign n6317 = n6315 | n6316 ;
  assign n6318 = x82 & n1859 ;
  assign n6319 = x81 & n1854 ;
  assign n6320 = x80 & ~n1853 ;
  assign n6321 = n2037 & n6320 ;
  assign n6322 = n6319 | n6321 ;
  assign n6323 = n6318 | n6322 ;
  assign n6324 = n1862 | n6318 ;
  assign n6325 = n6322 | n6324 ;
  assign n6326 = ( n1811 & n6323 ) | ( n1811 & n6325 ) | ( n6323 & n6325 ) ;
  assign n6327 = x20 & n6325 ;
  assign n6328 = x20 & n6318 ;
  assign n6329 = ( x20 & n6322 ) | ( x20 & n6328 ) | ( n6322 & n6328 ) ;
  assign n6330 = ( n1811 & n6327 ) | ( n1811 & n6329 ) | ( n6327 & n6329 ) ;
  assign n6331 = x20 & ~n6329 ;
  assign n6332 = x20 & ~n6325 ;
  assign n6333 = ( ~n1811 & n6331 ) | ( ~n1811 & n6332 ) | ( n6331 & n6332 ) ;
  assign n6334 = ( n6326 & ~n6330 ) | ( n6326 & n6333 ) | ( ~n6330 & n6333 ) ;
  assign n6335 = n6317 & n6334 ;
  assign n6336 = n6317 | n6334 ;
  assign n6337 = ~n6335 & n6336 ;
  assign n6338 = n6011 | n6017 ;
  assign n6339 = n6337 | n6338 ;
  assign n6340 = n6337 & n6338 ;
  assign n6341 = n6339 & ~n6340 ;
  assign n6342 = x85 & n1383 ;
  assign n6343 = x84 & n1378 ;
  assign n6344 = x83 & ~n1377 ;
  assign n6345 = n1542 & n6344 ;
  assign n6346 = n6343 | n6345 ;
  assign n6347 = n6342 | n6346 ;
  assign n6348 = n1386 | n6342 ;
  assign n6349 = n6346 | n6348 ;
  assign n6350 = ( n2381 & n6347 ) | ( n2381 & n6349 ) | ( n6347 & n6349 ) ;
  assign n6351 = x17 & n6349 ;
  assign n6352 = x17 & n6342 ;
  assign n6353 = ( x17 & n6346 ) | ( x17 & n6352 ) | ( n6346 & n6352 ) ;
  assign n6354 = ( n2381 & n6351 ) | ( n2381 & n6353 ) | ( n6351 & n6353 ) ;
  assign n6355 = x17 & ~n6353 ;
  assign n6356 = x17 & ~n6349 ;
  assign n6357 = ( ~n2381 & n6355 ) | ( ~n2381 & n6356 ) | ( n6355 & n6356 ) ;
  assign n6358 = ( n6350 & ~n6354 ) | ( n6350 & n6357 ) | ( ~n6354 & n6357 ) ;
  assign n6359 = n6341 & n6358 ;
  assign n6360 = n6341 & ~n6359 ;
  assign n6361 = ~n6341 & n6358 ;
  assign n6362 = n6360 | n6361 ;
  assign n6363 = n6036 | n6038 ;
  assign n6364 = ( n5873 & n6036 ) | ( n5873 & n6363 ) | ( n6036 & n6363 ) ;
  assign n6365 = ~n6362 & n6364 ;
  assign n6366 = n6362 & ~n6364 ;
  assign n6367 = n6365 | n6366 ;
  assign n6368 = x88 & n962 ;
  assign n6369 = x87 & n957 ;
  assign n6370 = x86 & ~n956 ;
  assign n6371 = n1105 & n6370 ;
  assign n6372 = n6369 | n6371 ;
  assign n6373 = n6368 | n6372 ;
  assign n6374 = n965 | n6368 ;
  assign n6375 = n6372 | n6374 ;
  assign n6376 = ( ~n3039 & n6373 ) | ( ~n3039 & n6375 ) | ( n6373 & n6375 ) ;
  assign n6377 = n6373 & n6375 ;
  assign n6378 = ( n3023 & n6376 ) | ( n3023 & n6377 ) | ( n6376 & n6377 ) ;
  assign n6379 = x14 & n6375 ;
  assign n6380 = x14 & n6368 ;
  assign n6381 = ( x14 & n6372 ) | ( x14 & n6380 ) | ( n6372 & n6380 ) ;
  assign n6382 = ( ~n3039 & n6379 ) | ( ~n3039 & n6381 ) | ( n6379 & n6381 ) ;
  assign n6383 = n6379 & n6381 ;
  assign n6384 = ( n3023 & n6382 ) | ( n3023 & n6383 ) | ( n6382 & n6383 ) ;
  assign n6385 = x14 & ~n6381 ;
  assign n6386 = x14 & ~n6375 ;
  assign n6387 = ( n3039 & n6385 ) | ( n3039 & n6386 ) | ( n6385 & n6386 ) ;
  assign n6388 = n6385 | n6386 ;
  assign n6389 = ( ~n3023 & n6387 ) | ( ~n3023 & n6388 ) | ( n6387 & n6388 ) ;
  assign n6390 = ( n6378 & ~n6384 ) | ( n6378 & n6389 ) | ( ~n6384 & n6389 ) ;
  assign n6391 = n6367 | n6390 ;
  assign n6392 = n6367 & n6390 ;
  assign n6393 = n6391 & ~n6392 ;
  assign n6394 = n6190 & n6393 ;
  assign n6395 = n6190 | n6393 ;
  assign n6396 = ~n6394 & n6395 ;
  assign n6397 = x91 & n636 ;
  assign n6398 = x90 & n631 ;
  assign n6399 = x89 & ~n630 ;
  assign n6400 = n764 & n6399 ;
  assign n6401 = n6398 | n6400 ;
  assign n6402 = n6397 | n6401 ;
  assign n6403 = n639 | n6397 ;
  assign n6404 = n6401 | n6403 ;
  assign n6405 = ( n3768 & n6402 ) | ( n3768 & n6404 ) | ( n6402 & n6404 ) ;
  assign n6406 = x11 & n6404 ;
  assign n6407 = x11 & n6397 ;
  assign n6408 = ( x11 & n6401 ) | ( x11 & n6407 ) | ( n6401 & n6407 ) ;
  assign n6409 = ( n3768 & n6406 ) | ( n3768 & n6408 ) | ( n6406 & n6408 ) ;
  assign n6410 = x11 & ~n6408 ;
  assign n6411 = x11 & ~n6404 ;
  assign n6412 = ( ~n3768 & n6410 ) | ( ~n3768 & n6411 ) | ( n6410 & n6411 ) ;
  assign n6413 = ( n6405 & ~n6409 ) | ( n6405 & n6412 ) | ( ~n6409 & n6412 ) ;
  assign n6414 = n6396 & n6413 ;
  assign n6415 = n6396 & ~n6414 ;
  assign n6416 = ~n6396 & n6413 ;
  assign n6417 = n6415 | n6416 ;
  assign n6418 = n6090 | n6091 ;
  assign n6419 = ( n6090 & n6093 ) | ( n6090 & n6418 ) | ( n6093 & n6418 ) ;
  assign n6420 = ~n6417 & n6419 ;
  assign n6421 = n6417 & ~n6419 ;
  assign n6422 = n6420 | n6421 ;
  assign n6423 = x94 & n389 ;
  assign n6424 = x93 & n384 ;
  assign n6425 = x92 & ~n383 ;
  assign n6426 = n463 & n6425 ;
  assign n6427 = n6424 | n6426 ;
  assign n6428 = n6423 | n6427 ;
  assign n6429 = n392 | n6423 ;
  assign n6430 = n6427 | n6429 ;
  assign n6431 = ( n4583 & n6428 ) | ( n4583 & n6430 ) | ( n6428 & n6430 ) ;
  assign n6432 = x8 & n6430 ;
  assign n6433 = x8 & n6423 ;
  assign n6434 = ( x8 & n6427 ) | ( x8 & n6433 ) | ( n6427 & n6433 ) ;
  assign n6435 = ( n4583 & n6432 ) | ( n4583 & n6434 ) | ( n6432 & n6434 ) ;
  assign n6436 = x8 & ~n6434 ;
  assign n6437 = x8 & ~n6430 ;
  assign n6438 = ( ~n4583 & n6436 ) | ( ~n4583 & n6437 ) | ( n6436 & n6437 ) ;
  assign n6439 = ( n6431 & ~n6435 ) | ( n6431 & n6438 ) | ( ~n6435 & n6438 ) ;
  assign n6440 = n6422 | n6439 ;
  assign n6441 = n6422 & n6439 ;
  assign n6442 = n6440 & ~n6441 ;
  assign n6443 = n6114 | n6116 ;
  assign n6444 = n6115 | n6443 ;
  assign n6445 = ( n6114 & n6118 ) | ( n6114 & n6444 ) | ( n6118 & n6444 ) ;
  assign n6446 = n6442 & n6445 ;
  assign n6447 = n6442 | n6445 ;
  assign n6448 = ~n6446 & n6447 ;
  assign n6449 = x97 & n212 ;
  assign n6450 = x96 & n207 ;
  assign n6451 = x95 & ~n206 ;
  assign n6452 = n267 & n6451 ;
  assign n6453 = n6450 | n6452 ;
  assign n6454 = n6449 | n6453 ;
  assign n6455 = n215 | n6449 ;
  assign n6456 = n6453 | n6455 ;
  assign n6457 = ( n5505 & n6454 ) | ( n5505 & n6456 ) | ( n6454 & n6456 ) ;
  assign n6458 = x5 & n6456 ;
  assign n6459 = x5 & n6449 ;
  assign n6460 = ( x5 & n6453 ) | ( x5 & n6459 ) | ( n6453 & n6459 ) ;
  assign n6461 = ( n5505 & n6458 ) | ( n5505 & n6460 ) | ( n6458 & n6460 ) ;
  assign n6462 = x5 & ~n6460 ;
  assign n6463 = x5 & ~n6456 ;
  assign n6464 = ( ~n5505 & n6462 ) | ( ~n5505 & n6463 ) | ( n6462 & n6463 ) ;
  assign n6465 = ( n6457 & ~n6461 ) | ( n6457 & n6464 ) | ( ~n6461 & n6464 ) ;
  assign n6466 = n6448 & n6465 ;
  assign n6467 = n6448 | n6465 ;
  assign n6468 = ~n6466 & n6467 ;
  assign n6469 = n6189 & n6468 ;
  assign n6470 = n6189 | n6468 ;
  assign n6471 = ~n6469 & n6470 ;
  assign n6472 = x99 | x100 ;
  assign n6473 = x99 & x100 ;
  assign n6474 = n6472 & ~n6473 ;
  assign n6475 = n6149 & n6474 ;
  assign n6476 = ( n6159 & n6474 ) | ( n6159 & n6475 ) | ( n6474 & n6475 ) ;
  assign n6477 = ( n6157 & n6474 ) | ( n6157 & n6475 ) | ( n6474 & n6475 ) ;
  assign n6478 = ( n5823 & n6476 ) | ( n5823 & n6477 ) | ( n6476 & n6477 ) ;
  assign n6479 = n6149 | n6474 ;
  assign n6480 = n6159 | n6479 ;
  assign n6481 = n6157 | n6479 ;
  assign n6482 = ( n5823 & n6480 ) | ( n5823 & n6481 ) | ( n6480 & n6481 ) ;
  assign n6483 = ~n6478 & n6482 ;
  assign n6484 = x99 & n133 ;
  assign n6485 = x98 & ~n162 ;
  assign n6486 = ( n137 & n6484 ) | ( n137 & n6485 ) | ( n6484 & n6485 ) ;
  assign n6487 = x0 & x100 ;
  assign n6488 = ( ~n137 & n6484 ) | ( ~n137 & n6487 ) | ( n6484 & n6487 ) ;
  assign n6489 = n6486 | n6488 ;
  assign n6490 = n141 | n6489 ;
  assign n6491 = ( n6483 & n6489 ) | ( n6483 & n6490 ) | ( n6489 & n6490 ) ;
  assign n6492 = x2 & n6489 ;
  assign n6493 = ( x2 & n523 ) | ( x2 & n6489 ) | ( n523 & n6489 ) ;
  assign n6494 = ( n6483 & n6492 ) | ( n6483 & n6493 ) | ( n6492 & n6493 ) ;
  assign n6495 = x2 & ~n6493 ;
  assign n6496 = x2 & ~n6489 ;
  assign n6497 = ( ~n6483 & n6495 ) | ( ~n6483 & n6496 ) | ( n6495 & n6496 ) ;
  assign n6498 = ( n6491 & ~n6494 ) | ( n6491 & n6497 ) | ( ~n6494 & n6497 ) ;
  assign n6499 = n6471 & n6498 ;
  assign n6500 = n6471 & ~n6499 ;
  assign n6501 = ~n6471 & n6498 ;
  assign n6502 = n6500 | n6501 ;
  assign n6503 = ( n6147 & n6179 ) | ( n6147 & ~n6184 ) | ( n6179 & ~n6184 ) ;
  assign n6504 = ( n5864 & ~n6145 ) | ( n5864 & n6179 ) | ( ~n6145 & n6179 ) ;
  assign n6505 = ( n5864 & n6141 ) | ( n5864 & n6179 ) | ( n6141 & n6179 ) ;
  assign n6506 = ( n6146 & n6504 ) | ( n6146 & n6505 ) | ( n6504 & n6505 ) ;
  assign n6507 = ( n5870 & n6503 ) | ( n5870 & n6506 ) | ( n6503 & n6506 ) ;
  assign n6508 = n6502 | n6507 ;
  assign n6509 = n6502 & n6507 ;
  assign n6510 = n6508 & ~n6509 ;
  assign n6511 = n6392 | n6394 ;
  assign n6512 = x70 & n4626 ;
  assign n6513 = x69 & ~n4625 ;
  assign n6514 = n4943 & n6513 ;
  assign n6515 = n6512 | n6514 ;
  assign n6516 = x71 & n4631 ;
  assign n6517 = n4634 | n6516 ;
  assign n6518 = n6515 | n6517 ;
  assign n6519 = x32 & ~n6518 ;
  assign n6520 = x32 & ~n6516 ;
  assign n6521 = ~n6515 & n6520 ;
  assign n6522 = ( ~n438 & n6519 ) | ( ~n438 & n6521 ) | ( n6519 & n6521 ) ;
  assign n6523 = ~x32 & n6518 ;
  assign n6524 = ~x32 & n6516 ;
  assign n6525 = ( ~x32 & n6515 ) | ( ~x32 & n6524 ) | ( n6515 & n6524 ) ;
  assign n6526 = ( n438 & n6523 ) | ( n438 & n6525 ) | ( n6523 & n6525 ) ;
  assign n6527 = n6522 | n6526 ;
  assign n6528 = ~x36 & x37 ;
  assign n6529 = x36 & ~x37 ;
  assign n6530 = n6528 | n6529 ;
  assign n6531 = ~n6195 & n6530 ;
  assign n6532 = x64 & n6531 ;
  assign n6533 = ~x37 & x38 ;
  assign n6534 = x37 & ~x38 ;
  assign n6535 = n6533 | n6534 ;
  assign n6536 = n6195 & ~n6535 ;
  assign n6537 = x65 & n6536 ;
  assign n6538 = n6532 | n6537 ;
  assign n6539 = n6195 & n6535 ;
  assign n6540 = x38 | n144 ;
  assign n6541 = ( x38 & n6539 ) | ( x38 & n6540 ) | ( n6539 & n6540 ) ;
  assign n6542 = ~x38 & n6541 ;
  assign n6543 = ( ~x38 & n6538 ) | ( ~x38 & n6542 ) | ( n6538 & n6542 ) ;
  assign n6544 = x38 & ~x64 ;
  assign n6545 = ( x38 & ~n6195 ) | ( x38 & n6544 ) | ( ~n6195 & n6544 ) ;
  assign n6546 = n6541 & n6545 ;
  assign n6547 = ( n6538 & n6545 ) | ( n6538 & n6546 ) | ( n6545 & n6546 ) ;
  assign n6548 = n144 & n6539 ;
  assign n6549 = n6545 & ~n6548 ;
  assign n6550 = ~n6538 & n6549 ;
  assign n6551 = ( n6543 & n6547 ) | ( n6543 & n6550 ) | ( n6547 & n6550 ) ;
  assign n6552 = n6541 | n6545 ;
  assign n6553 = n6538 | n6552 ;
  assign n6554 = ~n6545 & n6548 ;
  assign n6555 = ( n6538 & ~n6545 ) | ( n6538 & n6554 ) | ( ~n6545 & n6554 ) ;
  assign n6556 = ( n6543 & n6553 ) | ( n6543 & ~n6555 ) | ( n6553 & ~n6555 ) ;
  assign n6557 = ~n6551 & n6556 ;
  assign n6558 = n241 & n5557 ;
  assign n6559 = x68 & n5554 ;
  assign n6560 = x67 & n5549 ;
  assign n6561 = x66 & ~n5548 ;
  assign n6562 = n5893 & n6561 ;
  assign n6563 = n6560 | n6562 ;
  assign n6564 = n6559 | n6563 ;
  assign n6565 = n6558 | n6564 ;
  assign n6566 = x35 | n6559 ;
  assign n6567 = n6563 | n6566 ;
  assign n6568 = n6558 | n6567 ;
  assign n6569 = ~x35 & n6567 ;
  assign n6570 = ( ~x35 & n6558 ) | ( ~x35 & n6569 ) | ( n6558 & n6569 ) ;
  assign n6571 = ( ~n6565 & n6568 ) | ( ~n6565 & n6570 ) | ( n6568 & n6570 ) ;
  assign n6572 = n6557 | n6571 ;
  assign n6573 = n6557 & n6571 ;
  assign n6574 = n6572 & ~n6573 ;
  assign n6575 = ( n5907 & n6196 ) | ( n5907 & n6212 ) | ( n6196 & n6212 ) ;
  assign n6576 = n6574 | n6575 ;
  assign n6577 = n6574 & n6575 ;
  assign n6578 = n6576 & ~n6577 ;
  assign n6579 = n6527 | n6578 ;
  assign n6580 = n6527 & n6578 ;
  assign n6581 = n6579 & ~n6580 ;
  assign n6582 = ~n6215 & n6231 ;
  assign n6583 = n6192 & ~n6582 ;
  assign n6584 = n6215 & n6231 ;
  assign n6585 = n6215 & ~n6584 ;
  assign n6586 = ( n6192 & n6584 ) | ( n6192 & n6585 ) | ( n6584 & n6585 ) ;
  assign n6587 = n6192 | n6584 ;
  assign n6588 = ( ~n6583 & n6586 ) | ( ~n6583 & n6587 ) | ( n6586 & n6587 ) ;
  assign n6589 = n6581 & n6588 ;
  assign n6590 = n6581 | n6588 ;
  assign n6591 = ~n6589 & n6590 ;
  assign n6592 = x74 & n3816 ;
  assign n6593 = x73 & n3811 ;
  assign n6594 = x72 & ~n3810 ;
  assign n6595 = n4067 & n6594 ;
  assign n6596 = n6593 | n6595 ;
  assign n6597 = n6592 | n6596 ;
  assign n6598 = n3819 | n6592 ;
  assign n6599 = n6596 | n6598 ;
  assign n6600 = ( n710 & n6597 ) | ( n710 & n6599 ) | ( n6597 & n6599 ) ;
  assign n6601 = x29 & n6599 ;
  assign n6602 = x29 & n6592 ;
  assign n6603 = ( x29 & n6596 ) | ( x29 & n6602 ) | ( n6596 & n6602 ) ;
  assign n6604 = ( n710 & n6601 ) | ( n710 & n6603 ) | ( n6601 & n6603 ) ;
  assign n6605 = x29 & ~n6603 ;
  assign n6606 = x29 & ~n6599 ;
  assign n6607 = ( ~n710 & n6605 ) | ( ~n710 & n6606 ) | ( n6605 & n6606 ) ;
  assign n6608 = ( n6600 & ~n6604 ) | ( n6600 & n6607 ) | ( ~n6604 & n6607 ) ;
  assign n6609 = n6591 | n6608 ;
  assign n6610 = n6591 & n6608 ;
  assign n6611 = n6609 & ~n6610 ;
  assign n6612 = n6256 | n6264 ;
  assign n6613 = n6611 & n6612 ;
  assign n6614 = n6611 | n6612 ;
  assign n6615 = ~n6613 & n6614 ;
  assign n6616 = x77 & n3085 ;
  assign n6617 = x76 & n3080 ;
  assign n6618 = x75 & ~n3079 ;
  assign n6619 = n3309 & n6618 ;
  assign n6620 = n6617 | n6619 ;
  assign n6621 = n6616 | n6620 ;
  assign n6622 = n3088 | n6616 ;
  assign n6623 = n6620 | n6622 ;
  assign n6624 = ( n1059 & n6621 ) | ( n1059 & n6623 ) | ( n6621 & n6623 ) ;
  assign n6625 = x26 & n6623 ;
  assign n6626 = x26 & n6616 ;
  assign n6627 = ( x26 & n6620 ) | ( x26 & n6626 ) | ( n6620 & n6626 ) ;
  assign n6628 = ( n1059 & n6625 ) | ( n1059 & n6627 ) | ( n6625 & n6627 ) ;
  assign n6629 = x26 & ~n6627 ;
  assign n6630 = x26 & ~n6623 ;
  assign n6631 = ( ~n1059 & n6629 ) | ( ~n1059 & n6630 ) | ( n6629 & n6630 ) ;
  assign n6632 = ( n6624 & ~n6628 ) | ( n6624 & n6631 ) | ( ~n6628 & n6631 ) ;
  assign n6633 = n6615 | n6632 ;
  assign n6634 = n6615 & n6632 ;
  assign n6635 = n6633 & ~n6634 ;
  assign n6636 = n6286 | n6290 ;
  assign n6637 = n6635 & n6636 ;
  assign n6638 = n6635 | n6636 ;
  assign n6639 = ~n6637 & n6638 ;
  assign n6640 = x80 & n2429 ;
  assign n6641 = x79 & n2424 ;
  assign n6642 = x78 & ~n2423 ;
  assign n6643 = n2631 & n6642 ;
  assign n6644 = n6641 | n6643 ;
  assign n6645 = n6640 | n6644 ;
  assign n6646 = n2432 | n6640 ;
  assign n6647 = n6644 | n6646 ;
  assign n6648 = ( n1499 & n6645 ) | ( n1499 & n6647 ) | ( n6645 & n6647 ) ;
  assign n6649 = x23 & n6647 ;
  assign n6650 = x23 & n6640 ;
  assign n6651 = ( x23 & n6644 ) | ( x23 & n6650 ) | ( n6644 & n6650 ) ;
  assign n6652 = ( n1499 & n6649 ) | ( n1499 & n6651 ) | ( n6649 & n6651 ) ;
  assign n6653 = x23 & ~n6651 ;
  assign n6654 = x23 & ~n6647 ;
  assign n6655 = ( ~n1499 & n6653 ) | ( ~n1499 & n6654 ) | ( n6653 & n6654 ) ;
  assign n6656 = ( n6648 & ~n6652 ) | ( n6648 & n6655 ) | ( ~n6652 & n6655 ) ;
  assign n6657 = n6639 & n6656 ;
  assign n6658 = n6639 & ~n6657 ;
  assign n6659 = ( n5985 & n6293 ) | ( n5985 & n6310 ) | ( n6293 & n6310 ) ;
  assign n6660 = n6293 | n6310 ;
  assign n6661 = ( n5991 & n6659 ) | ( n5991 & n6660 ) | ( n6659 & n6660 ) ;
  assign n6662 = ~n6639 & n6656 ;
  assign n6663 = n6661 & n6662 ;
  assign n6664 = ( n6658 & n6661 ) | ( n6658 & n6663 ) | ( n6661 & n6663 ) ;
  assign n6665 = n6661 | n6662 ;
  assign n6666 = n6658 | n6665 ;
  assign n6667 = ~n6664 & n6666 ;
  assign n6668 = x83 & n1859 ;
  assign n6669 = x82 & n1854 ;
  assign n6670 = x81 & ~n1853 ;
  assign n6671 = n2037 & n6670 ;
  assign n6672 = n6669 | n6671 ;
  assign n6673 = n6668 | n6672 ;
  assign n6674 = n1862 | n6668 ;
  assign n6675 = n6672 | n6674 ;
  assign n6676 = ( n2009 & n6673 ) | ( n2009 & n6675 ) | ( n6673 & n6675 ) ;
  assign n6677 = x20 & n6675 ;
  assign n6678 = x20 & n6668 ;
  assign n6679 = ( x20 & n6672 ) | ( x20 & n6678 ) | ( n6672 & n6678 ) ;
  assign n6680 = ( n2009 & n6677 ) | ( n2009 & n6679 ) | ( n6677 & n6679 ) ;
  assign n6681 = x20 & ~n6679 ;
  assign n6682 = x20 & ~n6675 ;
  assign n6683 = ( ~n2009 & n6681 ) | ( ~n2009 & n6682 ) | ( n6681 & n6682 ) ;
  assign n6684 = ( n6676 & ~n6680 ) | ( n6676 & n6683 ) | ( ~n6680 & n6683 ) ;
  assign n6685 = n6667 & n6684 ;
  assign n6686 = n6667 & ~n6685 ;
  assign n6687 = ~n6667 & n6684 ;
  assign n6688 = n6686 | n6687 ;
  assign n6689 = n6335 | n6337 ;
  assign n6690 = ( n6335 & n6338 ) | ( n6335 & n6689 ) | ( n6338 & n6689 ) ;
  assign n6691 = n6688 | n6690 ;
  assign n6692 = n6688 & n6690 ;
  assign n6693 = n6691 & ~n6692 ;
  assign n6694 = x86 & n1383 ;
  assign n6695 = x85 & n1378 ;
  assign n6696 = x84 & ~n1377 ;
  assign n6697 = n1542 & n6696 ;
  assign n6698 = n6695 | n6697 ;
  assign n6699 = n6694 | n6698 ;
  assign n6700 = n1386 | n6694 ;
  assign n6701 = n6698 | n6700 ;
  assign n6702 = ( n2606 & n6699 ) | ( n2606 & n6701 ) | ( n6699 & n6701 ) ;
  assign n6703 = x17 & n6701 ;
  assign n6704 = x17 & n6694 ;
  assign n6705 = ( x17 & n6698 ) | ( x17 & n6704 ) | ( n6698 & n6704 ) ;
  assign n6706 = ( n2606 & n6703 ) | ( n2606 & n6705 ) | ( n6703 & n6705 ) ;
  assign n6707 = x17 & ~n6705 ;
  assign n6708 = x17 & ~n6701 ;
  assign n6709 = ( ~n2606 & n6707 ) | ( ~n2606 & n6708 ) | ( n6707 & n6708 ) ;
  assign n6710 = ( n6702 & ~n6706 ) | ( n6702 & n6709 ) | ( ~n6706 & n6709 ) ;
  assign n6711 = n6693 & n6710 ;
  assign n6712 = n6693 & ~n6711 ;
  assign n6713 = ~n6693 & n6710 ;
  assign n6714 = n6712 | n6713 ;
  assign n6715 = ( n6341 & n6358 ) | ( n6341 & n6364 ) | ( n6358 & n6364 ) ;
  assign n6716 = n6714 | n6715 ;
  assign n6717 = n6714 & n6715 ;
  assign n6718 = n6716 & ~n6717 ;
  assign n6719 = x89 & n962 ;
  assign n6720 = x88 & n957 ;
  assign n6721 = x87 & ~n956 ;
  assign n6722 = n1105 & n6721 ;
  assign n6723 = n6720 | n6722 ;
  assign n6724 = n6719 | n6723 ;
  assign n6725 = n965 | n6719 ;
  assign n6726 = n6723 | n6725 ;
  assign n6727 = ( n3282 & n6724 ) | ( n3282 & n6726 ) | ( n6724 & n6726 ) ;
  assign n6728 = x14 & n6726 ;
  assign n6729 = x14 & n6719 ;
  assign n6730 = ( x14 & n6723 ) | ( x14 & n6729 ) | ( n6723 & n6729 ) ;
  assign n6731 = ( n3282 & n6728 ) | ( n3282 & n6730 ) | ( n6728 & n6730 ) ;
  assign n6732 = x14 & ~n6730 ;
  assign n6733 = x14 & ~n6726 ;
  assign n6734 = ( ~n3282 & n6732 ) | ( ~n3282 & n6733 ) | ( n6732 & n6733 ) ;
  assign n6735 = ( n6727 & ~n6731 ) | ( n6727 & n6734 ) | ( ~n6731 & n6734 ) ;
  assign n6736 = n6718 & n6735 ;
  assign n6737 = n6718 | n6735 ;
  assign n6738 = ~n6736 & n6737 ;
  assign n6739 = n6511 & n6738 ;
  assign n6740 = n6511 & ~n6739 ;
  assign n6741 = x92 & n636 ;
  assign n6742 = x91 & n631 ;
  assign n6743 = x90 & ~n630 ;
  assign n6744 = n764 & n6743 ;
  assign n6745 = n6742 | n6744 ;
  assign n6746 = n6741 | n6745 ;
  assign n6747 = n639 | n6741 ;
  assign n6748 = n6745 | n6747 ;
  assign n6749 = ( n4040 & n6746 ) | ( n4040 & n6748 ) | ( n6746 & n6748 ) ;
  assign n6750 = x11 & n6748 ;
  assign n6751 = x11 & n6741 ;
  assign n6752 = ( x11 & n6745 ) | ( x11 & n6751 ) | ( n6745 & n6751 ) ;
  assign n6753 = ( n4040 & n6750 ) | ( n4040 & n6752 ) | ( n6750 & n6752 ) ;
  assign n6754 = x11 & ~n6752 ;
  assign n6755 = x11 & ~n6748 ;
  assign n6756 = ( ~n4040 & n6754 ) | ( ~n4040 & n6755 ) | ( n6754 & n6755 ) ;
  assign n6757 = ( n6749 & ~n6753 ) | ( n6749 & n6756 ) | ( ~n6753 & n6756 ) ;
  assign n6758 = n6738 & n6757 ;
  assign n6759 = ~n6738 & n6757 ;
  assign n6760 = ( ~n6511 & n6757 ) | ( ~n6511 & n6759 ) | ( n6757 & n6759 ) ;
  assign n6761 = ( n6740 & n6758 ) | ( n6740 & n6760 ) | ( n6758 & n6760 ) ;
  assign n6762 = n6738 | n6757 ;
  assign n6763 = n6738 & ~n6757 ;
  assign n6764 = n6511 & n6763 ;
  assign n6765 = ( n6740 & n6762 ) | ( n6740 & ~n6764 ) | ( n6762 & ~n6764 ) ;
  assign n6766 = ~n6761 & n6765 ;
  assign n6767 = ( n6396 & n6413 ) | ( n6396 & n6419 ) | ( n6413 & n6419 ) ;
  assign n6768 = n6766 | n6767 ;
  assign n6769 = n6766 & n6767 ;
  assign n6770 = n6768 & ~n6769 ;
  assign n6771 = x95 & n389 ;
  assign n6772 = x94 & n384 ;
  assign n6773 = x93 & ~n383 ;
  assign n6774 = n463 & n6773 ;
  assign n6775 = n6772 | n6774 ;
  assign n6776 = n6771 | n6775 ;
  assign n6777 = n392 | n6771 ;
  assign n6778 = n6775 | n6777 ;
  assign n6779 = ( n4897 & n6776 ) | ( n4897 & n6778 ) | ( n6776 & n6778 ) ;
  assign n6780 = x8 & n6778 ;
  assign n6781 = x8 & n6771 ;
  assign n6782 = ( x8 & n6775 ) | ( x8 & n6781 ) | ( n6775 & n6781 ) ;
  assign n6783 = ( n4897 & n6780 ) | ( n4897 & n6782 ) | ( n6780 & n6782 ) ;
  assign n6784 = x8 & ~n6782 ;
  assign n6785 = x8 & ~n6778 ;
  assign n6786 = ( ~n4897 & n6784 ) | ( ~n4897 & n6785 ) | ( n6784 & n6785 ) ;
  assign n6787 = ( n6779 & ~n6783 ) | ( n6779 & n6786 ) | ( ~n6783 & n6786 ) ;
  assign n6788 = n6770 | n6787 ;
  assign n6789 = n6770 & n6787 ;
  assign n6790 = n6788 & ~n6789 ;
  assign n6791 = n6441 | n6442 ;
  assign n6792 = ( n6441 & n6445 ) | ( n6441 & n6791 ) | ( n6445 & n6791 ) ;
  assign n6793 = n6790 & n6792 ;
  assign n6794 = n6790 | n6792 ;
  assign n6795 = ~n6793 & n6794 ;
  assign n6796 = x98 & n212 ;
  assign n6797 = x97 & n207 ;
  assign n6798 = x96 & ~n206 ;
  assign n6799 = n267 & n6798 ;
  assign n6800 = n6797 | n6799 ;
  assign n6801 = n6796 | n6800 ;
  assign n6802 = n215 | n6796 ;
  assign n6803 = n6800 | n6802 ;
  assign n6804 = ( ~n5850 & n6801 ) | ( ~n5850 & n6803 ) | ( n6801 & n6803 ) ;
  assign n6805 = n6801 & n6803 ;
  assign n6806 = ( n5834 & n6804 ) | ( n5834 & n6805 ) | ( n6804 & n6805 ) ;
  assign n6807 = x5 & n6803 ;
  assign n6808 = x5 & n6796 ;
  assign n6809 = ( x5 & n6800 ) | ( x5 & n6808 ) | ( n6800 & n6808 ) ;
  assign n6810 = ( ~n5850 & n6807 ) | ( ~n5850 & n6809 ) | ( n6807 & n6809 ) ;
  assign n6811 = n6807 & n6809 ;
  assign n6812 = ( n5834 & n6810 ) | ( n5834 & n6811 ) | ( n6810 & n6811 ) ;
  assign n6813 = x5 & ~n6809 ;
  assign n6814 = x5 & ~n6803 ;
  assign n6815 = ( n5850 & n6813 ) | ( n5850 & n6814 ) | ( n6813 & n6814 ) ;
  assign n6816 = n6813 | n6814 ;
  assign n6817 = ( ~n5834 & n6815 ) | ( ~n5834 & n6816 ) | ( n6815 & n6816 ) ;
  assign n6818 = ( n6806 & ~n6812 ) | ( n6806 & n6817 ) | ( ~n6812 & n6817 ) ;
  assign n6819 = n6795 & n6818 ;
  assign n6820 = n6795 & ~n6819 ;
  assign n6821 = ~n6795 & n6818 ;
  assign n6822 = n6820 | n6821 ;
  assign n6823 = n6466 | n6468 ;
  assign n6824 = ( n6189 & n6466 ) | ( n6189 & n6823 ) | ( n6466 & n6823 ) ;
  assign n6825 = n6822 | n6824 ;
  assign n6826 = n6822 & n6824 ;
  assign n6827 = n6825 & ~n6826 ;
  assign n6828 = x100 | x101 ;
  assign n6829 = x100 & x101 ;
  assign n6830 = n6828 & ~n6829 ;
  assign n6831 = n6149 | n6473 ;
  assign n6832 = ( n6473 & n6474 ) | ( n6473 & n6831 ) | ( n6474 & n6831 ) ;
  assign n6833 = n6830 & n6832 ;
  assign n6834 = n6473 | n6474 ;
  assign n6835 = n6830 & n6834 ;
  assign n6836 = ( n6159 & n6833 ) | ( n6159 & n6835 ) | ( n6833 & n6835 ) ;
  assign n6837 = ( n6157 & n6833 ) | ( n6157 & n6835 ) | ( n6833 & n6835 ) ;
  assign n6838 = ( n5823 & n6836 ) | ( n5823 & n6837 ) | ( n6836 & n6837 ) ;
  assign n6839 = n6830 | n6832 ;
  assign n6840 = n6830 | n6834 ;
  assign n6841 = ( n6159 & n6839 ) | ( n6159 & n6840 ) | ( n6839 & n6840 ) ;
  assign n6842 = ( n6157 & n6839 ) | ( n6157 & n6840 ) | ( n6839 & n6840 ) ;
  assign n6843 = ( n5823 & n6841 ) | ( n5823 & n6842 ) | ( n6841 & n6842 ) ;
  assign n6844 = ~n6838 & n6843 ;
  assign n6845 = x100 & n133 ;
  assign n6846 = x99 & ~n162 ;
  assign n6847 = ( n137 & n6845 ) | ( n137 & n6846 ) | ( n6845 & n6846 ) ;
  assign n6848 = x0 & x101 ;
  assign n6849 = ( ~n137 & n6845 ) | ( ~n137 & n6848 ) | ( n6845 & n6848 ) ;
  assign n6850 = n6847 | n6849 ;
  assign n6851 = n141 | n6850 ;
  assign n6852 = ( n6844 & n6850 ) | ( n6844 & n6851 ) | ( n6850 & n6851 ) ;
  assign n6853 = x2 & n6850 ;
  assign n6854 = ( x2 & n523 ) | ( x2 & n6850 ) | ( n523 & n6850 ) ;
  assign n6855 = ( n6844 & n6853 ) | ( n6844 & n6854 ) | ( n6853 & n6854 ) ;
  assign n6856 = x2 & ~n6854 ;
  assign n6857 = x2 & ~n6850 ;
  assign n6858 = ( ~n6844 & n6856 ) | ( ~n6844 & n6857 ) | ( n6856 & n6857 ) ;
  assign n6859 = ( n6852 & ~n6855 ) | ( n6852 & n6858 ) | ( ~n6855 & n6858 ) ;
  assign n6860 = n6827 | n6859 ;
  assign n6861 = n6827 & n6859 ;
  assign n6862 = n6860 & ~n6861 ;
  assign n6863 = n6499 | n6507 ;
  assign n6864 = ( n6499 & n6502 ) | ( n6499 & n6863 ) | ( n6502 & n6863 ) ;
  assign n6865 = n6862 | n6864 ;
  assign n6866 = n6862 & n6864 ;
  assign n6867 = n6865 & ~n6866 ;
  assign n6868 = n6610 | n6613 ;
  assign n6869 = x66 & n6536 ;
  assign n6870 = x65 & n6531 ;
  assign n6871 = ~n6195 & n6535 ;
  assign n6872 = x64 & ~n6530 ;
  assign n6873 = n6871 & n6872 ;
  assign n6874 = n6870 | n6873 ;
  assign n6875 = n6869 | n6874 ;
  assign n6876 = n159 & n6539 ;
  assign n6877 = n6875 | n6876 ;
  assign n6878 = x38 | n6539 ;
  assign n6879 = ( x38 & n159 ) | ( x38 & n6878 ) | ( n159 & n6878 ) ;
  assign n6880 = n6875 | n6879 ;
  assign n6881 = ~x38 & n6879 ;
  assign n6882 = ( ~x38 & n6875 ) | ( ~x38 & n6881 ) | ( n6875 & n6881 ) ;
  assign n6883 = ( ~n6877 & n6880 ) | ( ~n6877 & n6882 ) | ( n6880 & n6882 ) ;
  assign n6884 = n6551 | n6883 ;
  assign n6885 = n6551 & n6883 ;
  assign n6886 = n6884 & ~n6885 ;
  assign n6887 = n293 & n5557 ;
  assign n6888 = x69 & n5554 ;
  assign n6889 = x68 & n5549 ;
  assign n6890 = x67 & ~n5548 ;
  assign n6891 = n5893 & n6890 ;
  assign n6892 = n6889 | n6891 ;
  assign n6893 = n6888 | n6892 ;
  assign n6894 = n6887 | n6893 ;
  assign n6895 = x35 | n6888 ;
  assign n6896 = n6892 | n6895 ;
  assign n6897 = n6887 | n6896 ;
  assign n6898 = ~x35 & n6896 ;
  assign n6899 = ( ~x35 & n6887 ) | ( ~x35 & n6898 ) | ( n6887 & n6898 ) ;
  assign n6900 = ( ~n6894 & n6897 ) | ( ~n6894 & n6899 ) | ( n6897 & n6899 ) ;
  assign n6901 = n6886 & n6900 ;
  assign n6902 = n6886 & ~n6901 ;
  assign n6903 = ~n6886 & n6900 ;
  assign n6904 = n6902 | n6903 ;
  assign n6905 = n6573 | n6575 ;
  assign n6906 = ( n6573 & n6574 ) | ( n6573 & n6905 ) | ( n6574 & n6905 ) ;
  assign n6907 = ~n6904 & n6906 ;
  assign n6908 = n6904 & ~n6906 ;
  assign n6909 = n6907 | n6908 ;
  assign n6910 = x72 & n4631 ;
  assign n6911 = x71 & n4626 ;
  assign n6912 = x70 & ~n4625 ;
  assign n6913 = n4943 & n6912 ;
  assign n6914 = n6911 | n6913 ;
  assign n6915 = n6910 | n6914 ;
  assign n6916 = ( n513 & n4634 ) | ( n513 & n6915 ) | ( n4634 & n6915 ) ;
  assign n6917 = ( x32 & n4634 ) | ( x32 & ~n6910 ) | ( n4634 & ~n6910 ) ;
  assign n6918 = x32 & n4634 ;
  assign n6919 = ( ~n6914 & n6917 ) | ( ~n6914 & n6918 ) | ( n6917 & n6918 ) ;
  assign n6920 = ( x32 & n513 ) | ( x32 & n6919 ) | ( n513 & n6919 ) ;
  assign n6921 = ~n6916 & n6920 ;
  assign n6922 = n6915 | n6919 ;
  assign n6923 = x32 | n6915 ;
  assign n6924 = ( n513 & n6922 ) | ( n513 & n6923 ) | ( n6922 & n6923 ) ;
  assign n6925 = ( ~x32 & n6921 ) | ( ~x32 & n6924 ) | ( n6921 & n6924 ) ;
  assign n6926 = n6909 & n6925 ;
  assign n6927 = n6909 | n6925 ;
  assign n6928 = ~n6926 & n6927 ;
  assign n6929 = n6580 | n6581 ;
  assign n6930 = ( n6580 & n6588 ) | ( n6580 & n6929 ) | ( n6588 & n6929 ) ;
  assign n6931 = n6928 & n6930 ;
  assign n6932 = n6928 | n6930 ;
  assign n6933 = ~n6931 & n6932 ;
  assign n6934 = x75 & n3816 ;
  assign n6935 = x74 & n3811 ;
  assign n6936 = x73 & ~n3810 ;
  assign n6937 = n4067 & n6936 ;
  assign n6938 = n6935 | n6937 ;
  assign n6939 = n6934 | n6938 ;
  assign n6940 = n3819 | n6934 ;
  assign n6941 = n6938 | n6940 ;
  assign n6942 = ( n746 & n6939 ) | ( n746 & n6941 ) | ( n6939 & n6941 ) ;
  assign n6943 = x29 & n6941 ;
  assign n6944 = x29 & n6934 ;
  assign n6945 = ( x29 & n6938 ) | ( x29 & n6944 ) | ( n6938 & n6944 ) ;
  assign n6946 = ( n746 & n6943 ) | ( n746 & n6945 ) | ( n6943 & n6945 ) ;
  assign n6947 = x29 & ~n6945 ;
  assign n6948 = x29 & ~n6941 ;
  assign n6949 = ( ~n746 & n6947 ) | ( ~n746 & n6948 ) | ( n6947 & n6948 ) ;
  assign n6950 = ( n6942 & ~n6946 ) | ( n6942 & n6949 ) | ( ~n6946 & n6949 ) ;
  assign n6951 = n6933 & n6950 ;
  assign n6952 = n6933 & ~n6951 ;
  assign n6953 = ~n6933 & n6950 ;
  assign n6954 = n6952 | n6953 ;
  assign n6955 = n6868 & n6954 ;
  assign n6956 = n6868 & ~n6955 ;
  assign n6957 = n6954 & ~n6955 ;
  assign n6958 = n6956 | n6957 ;
  assign n6959 = x78 & n3085 ;
  assign n6960 = x77 & n3080 ;
  assign n6961 = x76 & ~n3079 ;
  assign n6962 = n3309 & n6961 ;
  assign n6963 = n6960 | n6962 ;
  assign n6964 = n6959 | n6963 ;
  assign n6965 = n3088 | n6959 ;
  assign n6966 = n6963 | n6965 ;
  assign n6967 = ( n1192 & n6964 ) | ( n1192 & n6966 ) | ( n6964 & n6966 ) ;
  assign n6968 = x26 & n6966 ;
  assign n6969 = x26 & n6959 ;
  assign n6970 = ( x26 & n6963 ) | ( x26 & n6969 ) | ( n6963 & n6969 ) ;
  assign n6971 = ( n1192 & n6968 ) | ( n1192 & n6970 ) | ( n6968 & n6970 ) ;
  assign n6972 = x26 & ~n6970 ;
  assign n6973 = x26 & ~n6966 ;
  assign n6974 = ( ~n1192 & n6972 ) | ( ~n1192 & n6973 ) | ( n6972 & n6973 ) ;
  assign n6975 = ( n6967 & ~n6971 ) | ( n6967 & n6974 ) | ( ~n6971 & n6974 ) ;
  assign n6976 = n6958 | n6975 ;
  assign n6977 = n6958 & n6975 ;
  assign n6978 = n6976 & ~n6977 ;
  assign n6979 = n6634 | n6635 ;
  assign n6980 = ( n6634 & n6636 ) | ( n6634 & n6979 ) | ( n6636 & n6979 ) ;
  assign n6981 = n6978 & n6980 ;
  assign n6982 = n6978 | n6980 ;
  assign n6983 = ~n6981 & n6982 ;
  assign n6984 = x81 & n2429 ;
  assign n6985 = x80 & n2424 ;
  assign n6986 = x79 & ~n2423 ;
  assign n6987 = n2631 & n6986 ;
  assign n6988 = n6985 | n6987 ;
  assign n6989 = n6984 | n6988 ;
  assign n6990 = n2432 | n6984 ;
  assign n6991 = n6988 | n6990 ;
  assign n6992 = ( n1651 & n6989 ) | ( n1651 & n6991 ) | ( n6989 & n6991 ) ;
  assign n6993 = x23 & n6991 ;
  assign n6994 = x23 & n6984 ;
  assign n6995 = ( x23 & n6988 ) | ( x23 & n6994 ) | ( n6988 & n6994 ) ;
  assign n6996 = ( n1651 & n6993 ) | ( n1651 & n6995 ) | ( n6993 & n6995 ) ;
  assign n6997 = x23 & ~n6995 ;
  assign n6998 = x23 & ~n6991 ;
  assign n6999 = ( ~n1651 & n6997 ) | ( ~n1651 & n6998 ) | ( n6997 & n6998 ) ;
  assign n7000 = ( n6992 & ~n6996 ) | ( n6992 & n6999 ) | ( ~n6996 & n6999 ) ;
  assign n7001 = n6983 & n7000 ;
  assign n7002 = n6983 & ~n7001 ;
  assign n7003 = ~n6983 & n7000 ;
  assign n7004 = n7002 | n7003 ;
  assign n7005 = n6657 | n6664 ;
  assign n7006 = n7004 | n7005 ;
  assign n7007 = n7004 & n7005 ;
  assign n7008 = n7006 & ~n7007 ;
  assign n7009 = x84 & n1859 ;
  assign n7010 = x83 & n1854 ;
  assign n7011 = x82 & ~n1853 ;
  assign n7012 = n2037 & n7011 ;
  assign n7013 = n7010 | n7012 ;
  assign n7014 = n7009 | n7013 ;
  assign n7015 = n1862 | n7009 ;
  assign n7016 = n7013 | n7015 ;
  assign n7017 = ( n2194 & n7014 ) | ( n2194 & n7016 ) | ( n7014 & n7016 ) ;
  assign n7018 = x20 & n7016 ;
  assign n7019 = x20 & n7009 ;
  assign n7020 = ( x20 & n7013 ) | ( x20 & n7019 ) | ( n7013 & n7019 ) ;
  assign n7021 = ( n2194 & n7018 ) | ( n2194 & n7020 ) | ( n7018 & n7020 ) ;
  assign n7022 = x20 & ~n7020 ;
  assign n7023 = x20 & ~n7016 ;
  assign n7024 = ( ~n2194 & n7022 ) | ( ~n2194 & n7023 ) | ( n7022 & n7023 ) ;
  assign n7025 = ( n7017 & ~n7021 ) | ( n7017 & n7024 ) | ( ~n7021 & n7024 ) ;
  assign n7026 = n7008 & n7025 ;
  assign n7027 = n7008 & ~n7026 ;
  assign n7028 = ~n7008 & n7025 ;
  assign n7029 = n7027 | n7028 ;
  assign n7030 = n6685 | n6692 ;
  assign n7031 = n7029 | n7030 ;
  assign n7032 = n7029 & n7030 ;
  assign n7033 = n7031 & ~n7032 ;
  assign n7034 = x87 & n1383 ;
  assign n7035 = x86 & n1378 ;
  assign n7036 = x85 & ~n1377 ;
  assign n7037 = n1542 & n7036 ;
  assign n7038 = n7035 | n7037 ;
  assign n7039 = n7034 | n7038 ;
  assign n7040 = n1386 | n7034 ;
  assign n7041 = n7038 | n7040 ;
  assign n7042 = ( n2816 & n7039 ) | ( n2816 & n7041 ) | ( n7039 & n7041 ) ;
  assign n7043 = x17 & n7041 ;
  assign n7044 = x17 & n7034 ;
  assign n7045 = ( x17 & n7038 ) | ( x17 & n7044 ) | ( n7038 & n7044 ) ;
  assign n7046 = ( n2816 & n7043 ) | ( n2816 & n7045 ) | ( n7043 & n7045 ) ;
  assign n7047 = x17 & ~n7045 ;
  assign n7048 = x17 & ~n7041 ;
  assign n7049 = ( ~n2816 & n7047 ) | ( ~n2816 & n7048 ) | ( n7047 & n7048 ) ;
  assign n7050 = ( n7042 & ~n7046 ) | ( n7042 & n7049 ) | ( ~n7046 & n7049 ) ;
  assign n7051 = n7033 & n7050 ;
  assign n7052 = n7033 | n7050 ;
  assign n7053 = ~n7051 & n7052 ;
  assign n7054 = n6711 & n7053 ;
  assign n7055 = ( n6717 & n7053 ) | ( n6717 & n7054 ) | ( n7053 & n7054 ) ;
  assign n7056 = x90 & n962 ;
  assign n7057 = x89 & n957 ;
  assign n7058 = x88 & ~n956 ;
  assign n7059 = n1105 & n7058 ;
  assign n7060 = n7057 | n7059 ;
  assign n7061 = n7056 | n7060 ;
  assign n7062 = n965 | n7056 ;
  assign n7063 = n7060 | n7062 ;
  assign n7064 = ( n3519 & n7061 ) | ( n3519 & n7063 ) | ( n7061 & n7063 ) ;
  assign n7065 = x14 & n7063 ;
  assign n7066 = x14 & n7056 ;
  assign n7067 = ( x14 & n7060 ) | ( x14 & n7066 ) | ( n7060 & n7066 ) ;
  assign n7068 = ( n3519 & n7065 ) | ( n3519 & n7067 ) | ( n7065 & n7067 ) ;
  assign n7069 = x14 & ~n7067 ;
  assign n7070 = x14 & ~n7063 ;
  assign n7071 = ( ~n3519 & n7069 ) | ( ~n3519 & n7070 ) | ( n7069 & n7070 ) ;
  assign n7072 = ( n7064 & ~n7068 ) | ( n7064 & n7071 ) | ( ~n7068 & n7071 ) ;
  assign n7073 = n6711 | n6715 ;
  assign n7074 = ( n6711 & n6714 ) | ( n6711 & n7073 ) | ( n6714 & n7073 ) ;
  assign n7075 = n7072 & n7074 ;
  assign n7076 = ( n7053 & n7072 ) | ( n7053 & n7075 ) | ( n7072 & n7075 ) ;
  assign n7077 = ~n7055 & n7076 ;
  assign n7078 = n7072 | n7074 ;
  assign n7079 = n7053 | n7078 ;
  assign n7080 = ( ~n7055 & n7072 ) | ( ~n7055 & n7079 ) | ( n7072 & n7079 ) ;
  assign n7081 = ~n7077 & n7080 ;
  assign n7082 = n6736 | n6738 ;
  assign n7083 = ( n6511 & n6736 ) | ( n6511 & n7082 ) | ( n6736 & n7082 ) ;
  assign n7084 = n7081 & n7083 ;
  assign n7085 = n7081 | n7083 ;
  assign n7086 = ~n7084 & n7085 ;
  assign n7087 = x93 & n636 ;
  assign n7088 = x92 & n631 ;
  assign n7089 = x91 & ~n630 ;
  assign n7090 = n764 & n7089 ;
  assign n7091 = n7088 | n7090 ;
  assign n7092 = n7087 | n7091 ;
  assign n7093 = n639 | n7087 ;
  assign n7094 = n7091 | n7093 ;
  assign n7095 = ( n4305 & n7092 ) | ( n4305 & n7094 ) | ( n7092 & n7094 ) ;
  assign n7096 = x11 & n7094 ;
  assign n7097 = x11 & n7087 ;
  assign n7098 = ( x11 & n7091 ) | ( x11 & n7097 ) | ( n7091 & n7097 ) ;
  assign n7099 = ( n4305 & n7096 ) | ( n4305 & n7098 ) | ( n7096 & n7098 ) ;
  assign n7100 = x11 & ~n7098 ;
  assign n7101 = x11 & ~n7094 ;
  assign n7102 = ( ~n4305 & n7100 ) | ( ~n4305 & n7101 ) | ( n7100 & n7101 ) ;
  assign n7103 = ( n7095 & ~n7099 ) | ( n7095 & n7102 ) | ( ~n7099 & n7102 ) ;
  assign n7104 = n7086 | n7103 ;
  assign n7105 = n7086 & n7103 ;
  assign n7106 = n7104 & ~n7105 ;
  assign n7107 = n6761 | n6767 ;
  assign n7108 = ( n6761 & n6766 ) | ( n6761 & n7107 ) | ( n6766 & n7107 ) ;
  assign n7109 = n7106 & n7108 ;
  assign n7110 = n7106 | n7108 ;
  assign n7111 = ~n7109 & n7110 ;
  assign n7112 = x96 & n389 ;
  assign n7113 = x95 & n384 ;
  assign n7114 = x94 & ~n383 ;
  assign n7115 = n463 & n7114 ;
  assign n7116 = n7113 | n7115 ;
  assign n7117 = n7112 | n7116 ;
  assign n7118 = n392 | n7112 ;
  assign n7119 = n7116 | n7118 ;
  assign n7120 = ( n5202 & n7117 ) | ( n5202 & n7119 ) | ( n7117 & n7119 ) ;
  assign n7121 = x8 & n7119 ;
  assign n7122 = x8 & n7112 ;
  assign n7123 = ( x8 & n7116 ) | ( x8 & n7122 ) | ( n7116 & n7122 ) ;
  assign n7124 = ( n5202 & n7121 ) | ( n5202 & n7123 ) | ( n7121 & n7123 ) ;
  assign n7125 = x8 & ~n7123 ;
  assign n7126 = x8 & ~n7119 ;
  assign n7127 = ( ~n5202 & n7125 ) | ( ~n5202 & n7126 ) | ( n7125 & n7126 ) ;
  assign n7128 = ( n7120 & ~n7124 ) | ( n7120 & n7127 ) | ( ~n7124 & n7127 ) ;
  assign n7129 = n7111 | n7128 ;
  assign n7130 = n7111 & n7128 ;
  assign n7131 = n7129 & ~n7130 ;
  assign n7132 = n6789 | n6790 ;
  assign n7133 = ( n6789 & n6792 ) | ( n6789 & n7132 ) | ( n6792 & n7132 ) ;
  assign n7134 = n7131 & n7133 ;
  assign n7135 = n7131 | n7133 ;
  assign n7136 = ~n7134 & n7135 ;
  assign n7137 = x99 & n212 ;
  assign n7138 = x98 & n207 ;
  assign n7139 = x97 & ~n206 ;
  assign n7140 = n267 & n7139 ;
  assign n7141 = n7138 | n7140 ;
  assign n7142 = n7137 | n7141 ;
  assign n7143 = n215 | n7137 ;
  assign n7144 = n7141 | n7143 ;
  assign n7145 = ( n6164 & n7142 ) | ( n6164 & n7144 ) | ( n7142 & n7144 ) ;
  assign n7146 = x5 & n7144 ;
  assign n7147 = x5 & n7137 ;
  assign n7148 = ( x5 & n7141 ) | ( x5 & n7147 ) | ( n7141 & n7147 ) ;
  assign n7149 = ( n6164 & n7146 ) | ( n6164 & n7148 ) | ( n7146 & n7148 ) ;
  assign n7150 = x5 & ~n7148 ;
  assign n7151 = x5 & ~n7144 ;
  assign n7152 = ( ~n6164 & n7150 ) | ( ~n6164 & n7151 ) | ( n7150 & n7151 ) ;
  assign n7153 = ( n7145 & ~n7149 ) | ( n7145 & n7152 ) | ( ~n7149 & n7152 ) ;
  assign n7154 = n7136 | n7153 ;
  assign n7155 = n7136 & n7153 ;
  assign n7156 = n7154 & ~n7155 ;
  assign n7157 = n6819 & n7156 ;
  assign n7158 = ( n6826 & n7156 ) | ( n6826 & n7157 ) | ( n7156 & n7157 ) ;
  assign n7159 = n6819 | n7156 ;
  assign n7160 = n6826 | n7159 ;
  assign n7161 = ~n7158 & n7160 ;
  assign n7162 = x101 | x102 ;
  assign n7163 = x101 & x102 ;
  assign n7164 = n7162 & ~n7163 ;
  assign n7165 = n6829 | n6830 ;
  assign n7166 = ( n6829 & n6832 ) | ( n6829 & n7165 ) | ( n6832 & n7165 ) ;
  assign n7167 = n7164 & n7166 ;
  assign n7168 = ( n6829 & n6834 ) | ( n6829 & n7165 ) | ( n6834 & n7165 ) ;
  assign n7169 = n7164 & n7168 ;
  assign n7170 = ( n6159 & n7167 ) | ( n6159 & n7169 ) | ( n7167 & n7169 ) ;
  assign n7171 = ( n6157 & n7167 ) | ( n6157 & n7169 ) | ( n7167 & n7169 ) ;
  assign n7172 = ( n5823 & n7170 ) | ( n5823 & n7171 ) | ( n7170 & n7171 ) ;
  assign n7173 = n7164 | n7168 ;
  assign n7174 = n7164 | n7166 ;
  assign n7175 = ( n6159 & n7173 ) | ( n6159 & n7174 ) | ( n7173 & n7174 ) ;
  assign n7176 = ( n6157 & n7173 ) | ( n6157 & n7174 ) | ( n7173 & n7174 ) ;
  assign n7177 = ( n5823 & n7175 ) | ( n5823 & n7176 ) | ( n7175 & n7176 ) ;
  assign n7178 = ~n7172 & n7177 ;
  assign n7179 = x101 & n133 ;
  assign n7180 = x100 & ~n162 ;
  assign n7181 = ( n137 & n7179 ) | ( n137 & n7180 ) | ( n7179 & n7180 ) ;
  assign n7182 = x0 & x102 ;
  assign n7183 = ( ~n137 & n7179 ) | ( ~n137 & n7182 ) | ( n7179 & n7182 ) ;
  assign n7184 = n7181 | n7183 ;
  assign n7185 = n141 | n7184 ;
  assign n7186 = ( n7178 & n7184 ) | ( n7178 & n7185 ) | ( n7184 & n7185 ) ;
  assign n7187 = x2 & n7184 ;
  assign n7188 = ( x2 & n523 ) | ( x2 & n7184 ) | ( n523 & n7184 ) ;
  assign n7189 = ( n7178 & n7187 ) | ( n7178 & n7188 ) | ( n7187 & n7188 ) ;
  assign n7190 = x2 & ~n7188 ;
  assign n7191 = x2 & ~n7184 ;
  assign n7192 = ( ~n7178 & n7190 ) | ( ~n7178 & n7191 ) | ( n7190 & n7191 ) ;
  assign n7193 = ( n7186 & ~n7189 ) | ( n7186 & n7192 ) | ( ~n7189 & n7192 ) ;
  assign n7194 = n7161 & n7193 ;
  assign n7195 = n7161 & ~n7194 ;
  assign n7196 = ~n7161 & n7193 ;
  assign n7197 = n7195 | n7196 ;
  assign n7198 = n6861 | n6862 ;
  assign n7199 = ( n6861 & n6864 ) | ( n6861 & n7198 ) | ( n6864 & n7198 ) ;
  assign n7200 = n7197 & n7199 ;
  assign n7201 = n7197 | n7199 ;
  assign n7202 = ~n7200 & n7201 ;
  assign n7203 = n7155 | n7158 ;
  assign n7204 = n7077 | n7084 ;
  assign n7205 = x38 & ~x39 ;
  assign n7206 = ~x38 & x39 ;
  assign n7207 = n7205 | n7206 ;
  assign n7208 = x64 & n7207 ;
  assign n7209 = ~n6551 & n7208 ;
  assign n7210 = ( ~n6883 & n7208 ) | ( ~n6883 & n7209 ) | ( n7208 & n7209 ) ;
  assign n7211 = n6551 & ~n7208 ;
  assign n7212 = n6883 & n7211 ;
  assign n7213 = n7210 | n7212 ;
  assign n7214 = x67 & n6536 ;
  assign n7215 = x66 & n6531 ;
  assign n7216 = x65 & ~n6530 ;
  assign n7217 = n6871 & n7216 ;
  assign n7218 = n7215 | n7217 ;
  assign n7219 = n7214 | n7218 ;
  assign n7220 = n186 & n6539 ;
  assign n7221 = n7219 | n7220 ;
  assign n7222 = x38 & ~n7221 ;
  assign n7223 = ~x38 & n7221 ;
  assign n7224 = n7222 | n7223 ;
  assign n7225 = n7213 & n7224 ;
  assign n7226 = n7213 | n7224 ;
  assign n7227 = ~n7225 & n7226 ;
  assign n7228 = x69 & n5549 ;
  assign n7229 = x68 & ~n5548 ;
  assign n7230 = n5893 & n7229 ;
  assign n7231 = n7228 | n7230 ;
  assign n7232 = x70 & n5554 ;
  assign n7233 = n5557 | n7232 ;
  assign n7234 = n7231 | n7233 ;
  assign n7235 = x35 & ~n7234 ;
  assign n7236 = x35 & ~n7232 ;
  assign n7237 = ~n7231 & n7236 ;
  assign n7238 = ( ~n340 & n7235 ) | ( ~n340 & n7237 ) | ( n7235 & n7237 ) ;
  assign n7239 = ~x35 & n7234 ;
  assign n7240 = ~x35 & n7232 ;
  assign n7241 = ( ~x35 & n7231 ) | ( ~x35 & n7240 ) | ( n7231 & n7240 ) ;
  assign n7242 = ( n340 & n7239 ) | ( n340 & n7241 ) | ( n7239 & n7241 ) ;
  assign n7243 = n7238 | n7242 ;
  assign n7244 = n7227 & n7243 ;
  assign n7245 = n7227 & ~n7244 ;
  assign n7246 = ( n6886 & n6900 ) | ( n6886 & n6906 ) | ( n6900 & n6906 ) ;
  assign n7247 = ~n7227 & n7243 ;
  assign n7248 = n7246 & n7247 ;
  assign n7249 = ( n7245 & n7246 ) | ( n7245 & n7248 ) | ( n7246 & n7248 ) ;
  assign n7250 = n7246 | n7247 ;
  assign n7251 = n7245 | n7250 ;
  assign n7252 = ~n7249 & n7251 ;
  assign n7253 = x73 & n4631 ;
  assign n7254 = x72 & n4626 ;
  assign n7255 = x71 & ~n4625 ;
  assign n7256 = n4943 & n7255 ;
  assign n7257 = n7254 | n7256 ;
  assign n7258 = n7253 | n7257 ;
  assign n7259 = ( ~n610 & n4634 ) | ( ~n610 & n7258 ) | ( n4634 & n7258 ) ;
  assign n7260 = n4634 & n7253 ;
  assign n7261 = ( n4634 & n7257 ) | ( n4634 & n7260 ) | ( n7257 & n7260 ) ;
  assign n7262 = ( n598 & n7259 ) | ( n598 & n7261 ) | ( n7259 & n7261 ) ;
  assign n7263 = ( x32 & ~n7258 ) | ( x32 & n7262 ) | ( ~n7258 & n7262 ) ;
  assign n7264 = ~n7262 & n7263 ;
  assign n7265 = x32 | n7253 ;
  assign n7266 = n7257 | n7265 ;
  assign n7267 = n7262 | n7266 ;
  assign n7268 = ( ~x32 & n7264 ) | ( ~x32 & n7267 ) | ( n7264 & n7267 ) ;
  assign n7269 = n7252 & n7268 ;
  assign n7270 = n7252 & ~n7269 ;
  assign n7271 = n6926 | n6931 ;
  assign n7272 = ~n7252 & n7268 ;
  assign n7273 = n6926 & n7272 ;
  assign n7274 = ( n6931 & n7272 ) | ( n6931 & n7273 ) | ( n7272 & n7273 ) ;
  assign n7275 = ( n7270 & n7271 ) | ( n7270 & n7274 ) | ( n7271 & n7274 ) ;
  assign n7276 = n6926 | n7272 ;
  assign n7277 = n6931 | n7276 ;
  assign n7278 = n7270 | n7277 ;
  assign n7279 = ~n7275 & n7278 ;
  assign n7280 = x76 & n3816 ;
  assign n7281 = x75 & n3811 ;
  assign n7282 = x74 & ~n3810 ;
  assign n7283 = n4067 & n7282 ;
  assign n7284 = n7281 | n7283 ;
  assign n7285 = n7280 | n7284 ;
  assign n7286 = n3819 | n7280 ;
  assign n7287 = n7284 | n7286 ;
  assign n7288 = ( n923 & n7285 ) | ( n923 & n7287 ) | ( n7285 & n7287 ) ;
  assign n7289 = x29 & n7287 ;
  assign n7290 = x29 & n7280 ;
  assign n7291 = ( x29 & n7284 ) | ( x29 & n7290 ) | ( n7284 & n7290 ) ;
  assign n7292 = ( n923 & n7289 ) | ( n923 & n7291 ) | ( n7289 & n7291 ) ;
  assign n7293 = x29 & ~n7291 ;
  assign n7294 = x29 & ~n7287 ;
  assign n7295 = ( ~n923 & n7293 ) | ( ~n923 & n7294 ) | ( n7293 & n7294 ) ;
  assign n7296 = ( n7288 & ~n7292 ) | ( n7288 & n7295 ) | ( ~n7292 & n7295 ) ;
  assign n7297 = n7279 | n7296 ;
  assign n7298 = n7279 & n7296 ;
  assign n7299 = n7297 & ~n7298 ;
  assign n7300 = n6951 | n6955 ;
  assign n7301 = n7299 & n7300 ;
  assign n7302 = n7299 | n7300 ;
  assign n7303 = ~n7301 & n7302 ;
  assign n7304 = x79 & n3085 ;
  assign n7305 = x78 & n3080 ;
  assign n7306 = x77 & ~n3079 ;
  assign n7307 = n3309 & n7306 ;
  assign n7308 = n7305 | n7307 ;
  assign n7309 = n7304 | n7308 ;
  assign n7310 = n3088 | n7304 ;
  assign n7311 = n7308 | n7310 ;
  assign n7312 = ( n1332 & n7309 ) | ( n1332 & n7311 ) | ( n7309 & n7311 ) ;
  assign n7313 = x26 & n7311 ;
  assign n7314 = x26 & n7304 ;
  assign n7315 = ( x26 & n7308 ) | ( x26 & n7314 ) | ( n7308 & n7314 ) ;
  assign n7316 = ( n1332 & n7313 ) | ( n1332 & n7315 ) | ( n7313 & n7315 ) ;
  assign n7317 = x26 & ~n7315 ;
  assign n7318 = x26 & ~n7311 ;
  assign n7319 = ( ~n1332 & n7317 ) | ( ~n1332 & n7318 ) | ( n7317 & n7318 ) ;
  assign n7320 = ( n7312 & ~n7316 ) | ( n7312 & n7319 ) | ( ~n7316 & n7319 ) ;
  assign n7321 = n7303 & n7320 ;
  assign n7322 = n7303 & ~n7321 ;
  assign n7323 = ~n7303 & n7320 ;
  assign n7324 = n7322 | n7323 ;
  assign n7325 = n6977 | n6980 ;
  assign n7326 = ( n6977 & n6978 ) | ( n6977 & n7325 ) | ( n6978 & n7325 ) ;
  assign n7327 = ~n7324 & n7326 ;
  assign n7328 = n7324 & ~n7326 ;
  assign n7329 = n7327 | n7328 ;
  assign n7330 = x82 & n2429 ;
  assign n7331 = x81 & n2424 ;
  assign n7332 = x80 & ~n2423 ;
  assign n7333 = n2631 & n7332 ;
  assign n7334 = n7331 | n7333 ;
  assign n7335 = n7330 | n7334 ;
  assign n7336 = n2432 | n7330 ;
  assign n7337 = n7334 | n7336 ;
  assign n7338 = ( n1811 & n7335 ) | ( n1811 & n7337 ) | ( n7335 & n7337 ) ;
  assign n7339 = x23 & n7337 ;
  assign n7340 = x23 & n7330 ;
  assign n7341 = ( x23 & n7334 ) | ( x23 & n7340 ) | ( n7334 & n7340 ) ;
  assign n7342 = ( n1811 & n7339 ) | ( n1811 & n7341 ) | ( n7339 & n7341 ) ;
  assign n7343 = x23 & ~n7341 ;
  assign n7344 = x23 & ~n7337 ;
  assign n7345 = ( ~n1811 & n7343 ) | ( ~n1811 & n7344 ) | ( n7343 & n7344 ) ;
  assign n7346 = ( n7338 & ~n7342 ) | ( n7338 & n7345 ) | ( ~n7342 & n7345 ) ;
  assign n7347 = n7329 & n7346 ;
  assign n7348 = n7329 | n7346 ;
  assign n7349 = ~n7347 & n7348 ;
  assign n7350 = n7001 | n7005 ;
  assign n7351 = ( n7001 & n7004 ) | ( n7001 & n7350 ) | ( n7004 & n7350 ) ;
  assign n7352 = n7349 | n7351 ;
  assign n7353 = n7349 & n7351 ;
  assign n7354 = n7352 & ~n7353 ;
  assign n7355 = x85 & n1859 ;
  assign n7356 = x84 & n1854 ;
  assign n7357 = x83 & ~n1853 ;
  assign n7358 = n2037 & n7357 ;
  assign n7359 = n7356 | n7358 ;
  assign n7360 = n7355 | n7359 ;
  assign n7361 = n1862 | n7355 ;
  assign n7362 = n7359 | n7361 ;
  assign n7363 = ( n2381 & n7360 ) | ( n2381 & n7362 ) | ( n7360 & n7362 ) ;
  assign n7364 = x20 & n7362 ;
  assign n7365 = x20 & n7355 ;
  assign n7366 = ( x20 & n7359 ) | ( x20 & n7365 ) | ( n7359 & n7365 ) ;
  assign n7367 = ( n2381 & n7364 ) | ( n2381 & n7366 ) | ( n7364 & n7366 ) ;
  assign n7368 = x20 & ~n7366 ;
  assign n7369 = x20 & ~n7362 ;
  assign n7370 = ( ~n2381 & n7368 ) | ( ~n2381 & n7369 ) | ( n7368 & n7369 ) ;
  assign n7371 = ( n7363 & ~n7367 ) | ( n7363 & n7370 ) | ( ~n7367 & n7370 ) ;
  assign n7372 = n7354 & n7371 ;
  assign n7373 = n7354 & ~n7372 ;
  assign n7374 = ~n7354 & n7371 ;
  assign n7375 = n7373 | n7374 ;
  assign n7376 = n7026 | n7030 ;
  assign n7377 = ( n7026 & n7029 ) | ( n7026 & n7376 ) | ( n7029 & n7376 ) ;
  assign n7378 = n7375 | n7377 ;
  assign n7379 = n7375 & n7377 ;
  assign n7380 = n7378 & ~n7379 ;
  assign n7381 = x88 & n1383 ;
  assign n7382 = x87 & n1378 ;
  assign n7383 = x86 & ~n1377 ;
  assign n7384 = n1542 & n7383 ;
  assign n7385 = n7382 | n7384 ;
  assign n7386 = n7381 | n7385 ;
  assign n7387 = n1386 | n7381 ;
  assign n7388 = n7385 | n7387 ;
  assign n7389 = ( ~n3039 & n7386 ) | ( ~n3039 & n7388 ) | ( n7386 & n7388 ) ;
  assign n7390 = n7386 & n7388 ;
  assign n7391 = ( n3023 & n7389 ) | ( n3023 & n7390 ) | ( n7389 & n7390 ) ;
  assign n7392 = x17 & n7388 ;
  assign n7393 = x17 & n7381 ;
  assign n7394 = ( x17 & n7385 ) | ( x17 & n7393 ) | ( n7385 & n7393 ) ;
  assign n7395 = ( ~n3039 & n7392 ) | ( ~n3039 & n7394 ) | ( n7392 & n7394 ) ;
  assign n7396 = n7392 & n7394 ;
  assign n7397 = ( n3023 & n7395 ) | ( n3023 & n7396 ) | ( n7395 & n7396 ) ;
  assign n7398 = x17 & ~n7394 ;
  assign n7399 = x17 & ~n7388 ;
  assign n7400 = ( n3039 & n7398 ) | ( n3039 & n7399 ) | ( n7398 & n7399 ) ;
  assign n7401 = n7398 | n7399 ;
  assign n7402 = ( ~n3023 & n7400 ) | ( ~n3023 & n7401 ) | ( n7400 & n7401 ) ;
  assign n7403 = ( n7391 & ~n7397 ) | ( n7391 & n7402 ) | ( ~n7397 & n7402 ) ;
  assign n7404 = n7380 | n7403 ;
  assign n7405 = n7380 & n7403 ;
  assign n7406 = n7404 & ~n7405 ;
  assign n7407 = n7051 | n7053 ;
  assign n7408 = n6717 | n7051 ;
  assign n7409 = ( n7054 & n7407 ) | ( n7054 & n7408 ) | ( n7407 & n7408 ) ;
  assign n7410 = n7406 & n7409 ;
  assign n7411 = n7406 | n7409 ;
  assign n7412 = ~n7410 & n7411 ;
  assign n7413 = x91 & n962 ;
  assign n7414 = x90 & n957 ;
  assign n7415 = x89 & ~n956 ;
  assign n7416 = n1105 & n7415 ;
  assign n7417 = n7414 | n7416 ;
  assign n7418 = n7413 | n7417 ;
  assign n7419 = n965 | n7413 ;
  assign n7420 = n7417 | n7419 ;
  assign n7421 = ( n3768 & n7418 ) | ( n3768 & n7420 ) | ( n7418 & n7420 ) ;
  assign n7422 = x14 & n7420 ;
  assign n7423 = x14 & n7413 ;
  assign n7424 = ( x14 & n7417 ) | ( x14 & n7423 ) | ( n7417 & n7423 ) ;
  assign n7425 = ( n3768 & n7422 ) | ( n3768 & n7424 ) | ( n7422 & n7424 ) ;
  assign n7426 = x14 & ~n7424 ;
  assign n7427 = x14 & ~n7420 ;
  assign n7428 = ( ~n3768 & n7426 ) | ( ~n3768 & n7427 ) | ( n7426 & n7427 ) ;
  assign n7429 = ( n7421 & ~n7425 ) | ( n7421 & n7428 ) | ( ~n7425 & n7428 ) ;
  assign n7430 = n7412 & n7429 ;
  assign n7431 = n7412 & ~n7430 ;
  assign n7432 = ~n7412 & n7429 ;
  assign n7433 = n7431 | n7432 ;
  assign n7434 = n7204 & ~n7433 ;
  assign n7435 = ~n7204 & n7433 ;
  assign n7436 = n7434 | n7435 ;
  assign n7437 = x94 & n636 ;
  assign n7438 = x93 & n631 ;
  assign n7439 = x92 & ~n630 ;
  assign n7440 = n764 & n7439 ;
  assign n7441 = n7438 | n7440 ;
  assign n7442 = n7437 | n7441 ;
  assign n7443 = n639 | n7437 ;
  assign n7444 = n7441 | n7443 ;
  assign n7445 = ( n4583 & n7442 ) | ( n4583 & n7444 ) | ( n7442 & n7444 ) ;
  assign n7446 = x11 & n7444 ;
  assign n7447 = x11 & n7437 ;
  assign n7448 = ( x11 & n7441 ) | ( x11 & n7447 ) | ( n7441 & n7447 ) ;
  assign n7449 = ( n4583 & n7446 ) | ( n4583 & n7448 ) | ( n7446 & n7448 ) ;
  assign n7450 = x11 & ~n7448 ;
  assign n7451 = x11 & ~n7444 ;
  assign n7452 = ( ~n4583 & n7450 ) | ( ~n4583 & n7451 ) | ( n7450 & n7451 ) ;
  assign n7453 = ( n7445 & ~n7449 ) | ( n7445 & n7452 ) | ( ~n7449 & n7452 ) ;
  assign n7454 = n7436 & n7453 ;
  assign n7455 = n7436 | n7453 ;
  assign n7456 = ~n7454 & n7455 ;
  assign n7457 = n7105 | n7109 ;
  assign n7458 = n7456 & n7457 ;
  assign n7459 = n7456 | n7457 ;
  assign n7460 = ~n7458 & n7459 ;
  assign n7461 = x97 & n389 ;
  assign n7462 = x96 & n384 ;
  assign n7463 = x95 & ~n383 ;
  assign n7464 = n463 & n7463 ;
  assign n7465 = n7462 | n7464 ;
  assign n7466 = n7461 | n7465 ;
  assign n7467 = n392 | n7461 ;
  assign n7468 = n7465 | n7467 ;
  assign n7469 = ( n5505 & n7466 ) | ( n5505 & n7468 ) | ( n7466 & n7468 ) ;
  assign n7470 = x8 & n7468 ;
  assign n7471 = x8 & n7461 ;
  assign n7472 = ( x8 & n7465 ) | ( x8 & n7471 ) | ( n7465 & n7471 ) ;
  assign n7473 = ( n5505 & n7470 ) | ( n5505 & n7472 ) | ( n7470 & n7472 ) ;
  assign n7474 = x8 & ~n7472 ;
  assign n7475 = x8 & ~n7468 ;
  assign n7476 = ( ~n5505 & n7474 ) | ( ~n5505 & n7475 ) | ( n7474 & n7475 ) ;
  assign n7477 = ( n7469 & ~n7473 ) | ( n7469 & n7476 ) | ( ~n7473 & n7476 ) ;
  assign n7478 = n7460 & n7477 ;
  assign n7479 = n7460 & ~n7478 ;
  assign n7480 = ~n7460 & n7477 ;
  assign n7481 = n7130 | n7131 ;
  assign n7482 = ( n7130 & n7133 ) | ( n7130 & n7481 ) | ( n7133 & n7481 ) ;
  assign n7483 = ~n7480 & n7482 ;
  assign n7484 = ~n7479 & n7483 ;
  assign n7485 = n7480 & ~n7482 ;
  assign n7486 = ( n7479 & ~n7482 ) | ( n7479 & n7485 ) | ( ~n7482 & n7485 ) ;
  assign n7487 = n7484 | n7486 ;
  assign n7488 = x100 & n212 ;
  assign n7489 = x99 & n207 ;
  assign n7490 = x98 & ~n206 ;
  assign n7491 = n267 & n7490 ;
  assign n7492 = n7489 | n7491 ;
  assign n7493 = n7488 | n7492 ;
  assign n7494 = n215 | n7488 ;
  assign n7495 = n7492 | n7494 ;
  assign n7496 = ( n6483 & n7493 ) | ( n6483 & n7495 ) | ( n7493 & n7495 ) ;
  assign n7497 = x5 & n7495 ;
  assign n7498 = x5 & n7488 ;
  assign n7499 = ( x5 & n7492 ) | ( x5 & n7498 ) | ( n7492 & n7498 ) ;
  assign n7500 = ( n6483 & n7497 ) | ( n6483 & n7499 ) | ( n7497 & n7499 ) ;
  assign n7501 = x5 & ~n7499 ;
  assign n7502 = x5 & ~n7495 ;
  assign n7503 = ( ~n6483 & n7501 ) | ( ~n6483 & n7502 ) | ( n7501 & n7502 ) ;
  assign n7504 = ( n7496 & ~n7500 ) | ( n7496 & n7503 ) | ( ~n7500 & n7503 ) ;
  assign n7505 = n7487 | n7504 ;
  assign n7506 = n7487 & n7504 ;
  assign n7507 = n7505 & ~n7506 ;
  assign n7508 = n7203 & n7507 ;
  assign n7509 = n7203 | n7507 ;
  assign n7510 = ~n7508 & n7509 ;
  assign n7511 = x102 | x103 ;
  assign n7512 = x102 & x103 ;
  assign n7513 = n7511 & ~n7512 ;
  assign n7514 = n7163 | n7164 ;
  assign n7515 = n7513 & n7514 ;
  assign n7516 = n7163 & n7513 ;
  assign n7517 = ( n7166 & n7515 ) | ( n7166 & n7516 ) | ( n7515 & n7516 ) ;
  assign n7518 = ( n7168 & n7515 ) | ( n7168 & n7516 ) | ( n7515 & n7516 ) ;
  assign n7519 = ( n6159 & n7517 ) | ( n6159 & n7518 ) | ( n7517 & n7518 ) ;
  assign n7520 = ( n6157 & n7517 ) | ( n6157 & n7518 ) | ( n7517 & n7518 ) ;
  assign n7521 = ( n5823 & n7519 ) | ( n5823 & n7520 ) | ( n7519 & n7520 ) ;
  assign n7522 = n7513 | n7514 ;
  assign n7523 = n7163 | n7513 ;
  assign n7524 = ( n7168 & n7522 ) | ( n7168 & n7523 ) | ( n7522 & n7523 ) ;
  assign n7525 = ( n7166 & n7522 ) | ( n7166 & n7523 ) | ( n7522 & n7523 ) ;
  assign n7526 = ( n6159 & n7524 ) | ( n6159 & n7525 ) | ( n7524 & n7525 ) ;
  assign n7527 = ( n6157 & n7524 ) | ( n6157 & n7525 ) | ( n7524 & n7525 ) ;
  assign n7528 = ( n5823 & n7526 ) | ( n5823 & n7527 ) | ( n7526 & n7527 ) ;
  assign n7529 = ~n7521 & n7528 ;
  assign n7530 = x102 & n133 ;
  assign n7531 = x101 & ~n162 ;
  assign n7532 = ( n137 & n7530 ) | ( n137 & n7531 ) | ( n7530 & n7531 ) ;
  assign n7533 = x0 & x103 ;
  assign n7534 = ( ~n137 & n7530 ) | ( ~n137 & n7533 ) | ( n7530 & n7533 ) ;
  assign n7535 = n7532 | n7534 ;
  assign n7536 = n141 | n7535 ;
  assign n7537 = ( n7529 & n7535 ) | ( n7529 & n7536 ) | ( n7535 & n7536 ) ;
  assign n7538 = x2 & n7535 ;
  assign n7539 = ( x2 & n523 ) | ( x2 & n7535 ) | ( n523 & n7535 ) ;
  assign n7540 = ( n7529 & n7538 ) | ( n7529 & n7539 ) | ( n7538 & n7539 ) ;
  assign n7541 = x2 & ~n7539 ;
  assign n7542 = x2 & ~n7535 ;
  assign n7543 = ( ~n7529 & n7541 ) | ( ~n7529 & n7542 ) | ( n7541 & n7542 ) ;
  assign n7544 = ( n7537 & ~n7540 ) | ( n7537 & n7543 ) | ( ~n7540 & n7543 ) ;
  assign n7545 = n7510 & n7544 ;
  assign n7546 = n7510 & ~n7545 ;
  assign n7547 = ~n7510 & n7544 ;
  assign n7548 = n7546 | n7547 ;
  assign n7549 = n7194 | n7200 ;
  assign n7550 = n7548 & n7549 ;
  assign n7551 = n7548 | n7549 ;
  assign n7552 = ~n7550 & n7551 ;
  assign n7553 = n7545 | n7550 ;
  assign n7554 = ( n7077 & n7412 ) | ( n7077 & n7429 ) | ( n7412 & n7429 ) ;
  assign n7555 = n7412 | n7429 ;
  assign n7556 = ( n7084 & n7554 ) | ( n7084 & n7555 ) | ( n7554 & n7555 ) ;
  assign n7557 = n7269 | n7275 ;
  assign n7558 = ~x39 & x40 ;
  assign n7559 = x39 & ~x40 ;
  assign n7560 = n7558 | n7559 ;
  assign n7561 = ~n7207 & n7560 ;
  assign n7562 = x64 & n7561 ;
  assign n7563 = ~x40 & x41 ;
  assign n7564 = x40 & ~x41 ;
  assign n7565 = n7563 | n7564 ;
  assign n7566 = n7207 & ~n7565 ;
  assign n7567 = x65 & n7566 ;
  assign n7568 = n7562 | n7567 ;
  assign n7569 = n7207 & n7565 ;
  assign n7570 = x41 | n144 ;
  assign n7571 = ( x41 & n7569 ) | ( x41 & n7570 ) | ( n7569 & n7570 ) ;
  assign n7572 = ~x41 & n7571 ;
  assign n7573 = ( ~x41 & n7568 ) | ( ~x41 & n7572 ) | ( n7568 & n7572 ) ;
  assign n7574 = x41 & ~x64 ;
  assign n7575 = ( x41 & ~n7207 ) | ( x41 & n7574 ) | ( ~n7207 & n7574 ) ;
  assign n7576 = n7571 & n7575 ;
  assign n7577 = ( n7568 & n7575 ) | ( n7568 & n7576 ) | ( n7575 & n7576 ) ;
  assign n7578 = n144 & n7569 ;
  assign n7579 = n7575 & ~n7578 ;
  assign n7580 = ~n7568 & n7579 ;
  assign n7581 = ( n7573 & n7577 ) | ( n7573 & n7580 ) | ( n7577 & n7580 ) ;
  assign n7582 = n7571 | n7575 ;
  assign n7583 = n7568 | n7582 ;
  assign n7584 = ~n7575 & n7578 ;
  assign n7585 = ( n7568 & ~n7575 ) | ( n7568 & n7584 ) | ( ~n7575 & n7584 ) ;
  assign n7586 = ( n7573 & n7583 ) | ( n7573 & ~n7585 ) | ( n7583 & ~n7585 ) ;
  assign n7587 = ~n7581 & n7586 ;
  assign n7588 = n241 & n6539 ;
  assign n7589 = x68 & n6536 ;
  assign n7590 = x67 & n6531 ;
  assign n7591 = x66 & ~n6530 ;
  assign n7592 = n6871 & n7591 ;
  assign n7593 = n7590 | n7592 ;
  assign n7594 = n7589 | n7593 ;
  assign n7595 = n7588 | n7594 ;
  assign n7596 = x38 | n7589 ;
  assign n7597 = n7593 | n7596 ;
  assign n7598 = n7588 | n7597 ;
  assign n7599 = ~x38 & n7597 ;
  assign n7600 = ( ~x38 & n7588 ) | ( ~x38 & n7599 ) | ( n7588 & n7599 ) ;
  assign n7601 = ( ~n7595 & n7598 ) | ( ~n7595 & n7600 ) | ( n7598 & n7600 ) ;
  assign n7602 = n7587 | n7601 ;
  assign n7603 = n7587 & n7601 ;
  assign n7604 = n7602 & ~n7603 ;
  assign n7605 = ( n6885 & n7208 ) | ( n6885 & n7224 ) | ( n7208 & n7224 ) ;
  assign n7606 = n7604 | n7605 ;
  assign n7607 = n7604 & n7605 ;
  assign n7608 = n7606 & ~n7607 ;
  assign n7609 = x70 & n5549 ;
  assign n7610 = x69 & ~n5548 ;
  assign n7611 = n5893 & n7610 ;
  assign n7612 = n7609 | n7611 ;
  assign n7613 = x71 & n5554 ;
  assign n7614 = n5557 | n7613 ;
  assign n7615 = n7612 | n7614 ;
  assign n7616 = x35 & ~n7615 ;
  assign n7617 = x35 & ~n7613 ;
  assign n7618 = ~n7612 & n7617 ;
  assign n7619 = ( ~n438 & n7616 ) | ( ~n438 & n7618 ) | ( n7616 & n7618 ) ;
  assign n7620 = ~x35 & n7615 ;
  assign n7621 = ~x35 & n7613 ;
  assign n7622 = ( ~x35 & n7612 ) | ( ~x35 & n7621 ) | ( n7612 & n7621 ) ;
  assign n7623 = ( n438 & n7620 ) | ( n438 & n7622 ) | ( n7620 & n7622 ) ;
  assign n7624 = n7619 | n7623 ;
  assign n7625 = n7608 & n7624 ;
  assign n7626 = n7608 & ~n7625 ;
  assign n7627 = ~n7608 & n7624 ;
  assign n7628 = n7626 | n7627 ;
  assign n7629 = n7244 | n7249 ;
  assign n7630 = n7628 | n7629 ;
  assign n7631 = n7628 & n7629 ;
  assign n7632 = n7630 & ~n7631 ;
  assign n7633 = x74 & n4631 ;
  assign n7634 = x73 & n4626 ;
  assign n7635 = x72 & ~n4625 ;
  assign n7636 = n4943 & n7635 ;
  assign n7637 = n7634 | n7636 ;
  assign n7638 = n7633 | n7637 ;
  assign n7639 = n4634 | n7633 ;
  assign n7640 = n7637 | n7639 ;
  assign n7641 = ( n710 & n7638 ) | ( n710 & n7640 ) | ( n7638 & n7640 ) ;
  assign n7642 = x32 & n7640 ;
  assign n7643 = x32 & n7633 ;
  assign n7644 = ( x32 & n7637 ) | ( x32 & n7643 ) | ( n7637 & n7643 ) ;
  assign n7645 = ( n710 & n7642 ) | ( n710 & n7644 ) | ( n7642 & n7644 ) ;
  assign n7646 = x32 & ~n7644 ;
  assign n7647 = x32 & ~n7640 ;
  assign n7648 = ( ~n710 & n7646 ) | ( ~n710 & n7647 ) | ( n7646 & n7647 ) ;
  assign n7649 = ( n7641 & ~n7645 ) | ( n7641 & n7648 ) | ( ~n7645 & n7648 ) ;
  assign n7650 = n7632 & n7649 ;
  assign n7651 = n7632 | n7649 ;
  assign n7652 = ~n7650 & n7651 ;
  assign n7653 = n7269 & n7649 ;
  assign n7654 = ( n7269 & n7632 ) | ( n7269 & n7653 ) | ( n7632 & n7653 ) ;
  assign n7655 = ~n7650 & n7654 ;
  assign n7656 = ( n7275 & n7652 ) | ( n7275 & n7655 ) | ( n7652 & n7655 ) ;
  assign n7657 = n7557 & ~n7656 ;
  assign n7658 = x77 & n3816 ;
  assign n7659 = x76 & n3811 ;
  assign n7660 = x75 & ~n3810 ;
  assign n7661 = n4067 & n7660 ;
  assign n7662 = n7659 | n7661 ;
  assign n7663 = n7658 | n7662 ;
  assign n7664 = n3819 | n7658 ;
  assign n7665 = n7662 | n7664 ;
  assign n7666 = ( n1059 & n7663 ) | ( n1059 & n7665 ) | ( n7663 & n7665 ) ;
  assign n7667 = x29 & n7665 ;
  assign n7668 = x29 & n7658 ;
  assign n7669 = ( x29 & n7662 ) | ( x29 & n7668 ) | ( n7662 & n7668 ) ;
  assign n7670 = ( n1059 & n7667 ) | ( n1059 & n7669 ) | ( n7667 & n7669 ) ;
  assign n7671 = x29 & ~n7669 ;
  assign n7672 = x29 & ~n7665 ;
  assign n7673 = ( ~n1059 & n7671 ) | ( ~n1059 & n7672 ) | ( n7671 & n7672 ) ;
  assign n7674 = ( n7666 & ~n7670 ) | ( n7666 & n7673 ) | ( ~n7670 & n7673 ) ;
  assign n7675 = ( n7275 & n7651 ) | ( n7275 & n7654 ) | ( n7651 & n7654 ) ;
  assign n7676 = n7652 & n7674 ;
  assign n7677 = ~n7675 & n7676 ;
  assign n7678 = ( n7657 & n7674 ) | ( n7657 & n7677 ) | ( n7674 & n7677 ) ;
  assign n7679 = n7652 | n7674 ;
  assign n7680 = ( n7674 & ~n7675 ) | ( n7674 & n7679 ) | ( ~n7675 & n7679 ) ;
  assign n7681 = n7657 | n7680 ;
  assign n7682 = ~n7678 & n7681 ;
  assign n7683 = n7298 | n7299 ;
  assign n7684 = ( n7298 & n7300 ) | ( n7298 & n7683 ) | ( n7300 & n7683 ) ;
  assign n7685 = n7682 & n7684 ;
  assign n7686 = n7682 | n7684 ;
  assign n7687 = ~n7685 & n7686 ;
  assign n7688 = x80 & n3085 ;
  assign n7689 = x79 & n3080 ;
  assign n7690 = x78 & ~n3079 ;
  assign n7691 = n3309 & n7690 ;
  assign n7692 = n7689 | n7691 ;
  assign n7693 = n7688 | n7692 ;
  assign n7694 = n3088 | n7688 ;
  assign n7695 = n7692 | n7694 ;
  assign n7696 = ( n1499 & n7693 ) | ( n1499 & n7695 ) | ( n7693 & n7695 ) ;
  assign n7697 = x26 & n7695 ;
  assign n7698 = x26 & n7688 ;
  assign n7699 = ( x26 & n7692 ) | ( x26 & n7698 ) | ( n7692 & n7698 ) ;
  assign n7700 = ( n1499 & n7697 ) | ( n1499 & n7699 ) | ( n7697 & n7699 ) ;
  assign n7701 = x26 & ~n7699 ;
  assign n7702 = x26 & ~n7695 ;
  assign n7703 = ( ~n1499 & n7701 ) | ( ~n1499 & n7702 ) | ( n7701 & n7702 ) ;
  assign n7704 = ( n7696 & ~n7700 ) | ( n7696 & n7703 ) | ( ~n7700 & n7703 ) ;
  assign n7705 = n7687 & n7704 ;
  assign n7706 = n7687 & ~n7705 ;
  assign n7707 = ~n7687 & n7704 ;
  assign n7708 = n7706 | n7707 ;
  assign n7709 = ( n7303 & n7320 ) | ( n7303 & n7326 ) | ( n7320 & n7326 ) ;
  assign n7710 = n7708 | n7709 ;
  assign n7711 = n7708 & n7709 ;
  assign n7712 = n7710 & ~n7711 ;
  assign n7713 = x83 & n2429 ;
  assign n7714 = x82 & n2424 ;
  assign n7715 = x81 & ~n2423 ;
  assign n7716 = n2631 & n7715 ;
  assign n7717 = n7714 | n7716 ;
  assign n7718 = n7713 | n7717 ;
  assign n7719 = n2432 | n7713 ;
  assign n7720 = n7717 | n7719 ;
  assign n7721 = ( n2009 & n7718 ) | ( n2009 & n7720 ) | ( n7718 & n7720 ) ;
  assign n7722 = x23 & n7720 ;
  assign n7723 = x23 & n7713 ;
  assign n7724 = ( x23 & n7717 ) | ( x23 & n7723 ) | ( n7717 & n7723 ) ;
  assign n7725 = ( n2009 & n7722 ) | ( n2009 & n7724 ) | ( n7722 & n7724 ) ;
  assign n7726 = x23 & ~n7724 ;
  assign n7727 = x23 & ~n7720 ;
  assign n7728 = ( ~n2009 & n7726 ) | ( ~n2009 & n7727 ) | ( n7726 & n7727 ) ;
  assign n7729 = ( n7721 & ~n7725 ) | ( n7721 & n7728 ) | ( ~n7725 & n7728 ) ;
  assign n7730 = n7712 & n7729 ;
  assign n7731 = n7712 & ~n7730 ;
  assign n7732 = ~n7712 & n7729 ;
  assign n7733 = n7731 | n7732 ;
  assign n7734 = n7347 | n7353 ;
  assign n7735 = n7733 | n7734 ;
  assign n7736 = n7733 & n7734 ;
  assign n7737 = n7735 & ~n7736 ;
  assign n7738 = x86 & n1859 ;
  assign n7739 = x85 & n1854 ;
  assign n7740 = x84 & ~n1853 ;
  assign n7741 = n2037 & n7740 ;
  assign n7742 = n7739 | n7741 ;
  assign n7743 = n7738 | n7742 ;
  assign n7744 = n1862 | n7738 ;
  assign n7745 = n7742 | n7744 ;
  assign n7746 = ( n2606 & n7743 ) | ( n2606 & n7745 ) | ( n7743 & n7745 ) ;
  assign n7747 = x20 & n7745 ;
  assign n7748 = x20 & n7738 ;
  assign n7749 = ( x20 & n7742 ) | ( x20 & n7748 ) | ( n7742 & n7748 ) ;
  assign n7750 = ( n2606 & n7747 ) | ( n2606 & n7749 ) | ( n7747 & n7749 ) ;
  assign n7751 = x20 & ~n7749 ;
  assign n7752 = x20 & ~n7745 ;
  assign n7753 = ( ~n2606 & n7751 ) | ( ~n2606 & n7752 ) | ( n7751 & n7752 ) ;
  assign n7754 = ( n7746 & ~n7750 ) | ( n7746 & n7753 ) | ( ~n7750 & n7753 ) ;
  assign n7755 = n7737 & n7754 ;
  assign n7756 = n7737 & ~n7755 ;
  assign n7757 = ~n7737 & n7754 ;
  assign n7758 = n7756 | n7757 ;
  assign n7759 = n7372 | n7379 ;
  assign n7760 = n7758 | n7759 ;
  assign n7761 = n7758 & n7759 ;
  assign n7762 = n7760 & ~n7761 ;
  assign n7763 = x89 & n1383 ;
  assign n7764 = x88 & n1378 ;
  assign n7765 = x87 & ~n1377 ;
  assign n7766 = n1542 & n7765 ;
  assign n7767 = n7764 | n7766 ;
  assign n7768 = n7763 | n7767 ;
  assign n7769 = n1386 | n7763 ;
  assign n7770 = n7767 | n7769 ;
  assign n7771 = ( n3282 & n7768 ) | ( n3282 & n7770 ) | ( n7768 & n7770 ) ;
  assign n7772 = x17 & n7770 ;
  assign n7773 = x17 & n7763 ;
  assign n7774 = ( x17 & n7767 ) | ( x17 & n7773 ) | ( n7767 & n7773 ) ;
  assign n7775 = ( n3282 & n7772 ) | ( n3282 & n7774 ) | ( n7772 & n7774 ) ;
  assign n7776 = x17 & ~n7774 ;
  assign n7777 = x17 & ~n7770 ;
  assign n7778 = ( ~n3282 & n7776 ) | ( ~n3282 & n7777 ) | ( n7776 & n7777 ) ;
  assign n7779 = ( n7771 & ~n7775 ) | ( n7771 & n7778 ) | ( ~n7775 & n7778 ) ;
  assign n7780 = n7762 & n7779 ;
  assign n7781 = n7762 & ~n7780 ;
  assign n7782 = ~n7762 & n7779 ;
  assign n7783 = n7781 | n7782 ;
  assign n7784 = n7405 | n7406 ;
  assign n7785 = ( n7405 & n7409 ) | ( n7405 & n7784 ) | ( n7409 & n7784 ) ;
  assign n7786 = n7783 & n7785 ;
  assign n7787 = n7783 | n7785 ;
  assign n7788 = ~n7786 & n7787 ;
  assign n7789 = x92 & n962 ;
  assign n7790 = x91 & n957 ;
  assign n7791 = x90 & ~n956 ;
  assign n7792 = n1105 & n7791 ;
  assign n7793 = n7790 | n7792 ;
  assign n7794 = n7789 | n7793 ;
  assign n7795 = n965 | n7789 ;
  assign n7796 = n7793 | n7795 ;
  assign n7797 = ( n4040 & n7794 ) | ( n4040 & n7796 ) | ( n7794 & n7796 ) ;
  assign n7798 = x14 & n7796 ;
  assign n7799 = x14 & n7789 ;
  assign n7800 = ( x14 & n7793 ) | ( x14 & n7799 ) | ( n7793 & n7799 ) ;
  assign n7801 = ( n4040 & n7798 ) | ( n4040 & n7800 ) | ( n7798 & n7800 ) ;
  assign n7802 = x14 & ~n7800 ;
  assign n7803 = x14 & ~n7796 ;
  assign n7804 = ( ~n4040 & n7802 ) | ( ~n4040 & n7803 ) | ( n7802 & n7803 ) ;
  assign n7805 = ( n7797 & ~n7801 ) | ( n7797 & n7804 ) | ( ~n7801 & n7804 ) ;
  assign n7806 = n7788 & n7805 ;
  assign n7807 = n7788 & ~n7806 ;
  assign n7808 = ~n7788 & n7805 ;
  assign n7809 = n7556 & n7808 ;
  assign n7810 = ( n7556 & n7807 ) | ( n7556 & n7809 ) | ( n7807 & n7809 ) ;
  assign n7811 = n7556 & ~n7810 ;
  assign n7812 = n7807 | n7808 ;
  assign n7813 = ~n7810 & n7812 ;
  assign n7814 = n7811 | n7813 ;
  assign n7815 = x95 & n636 ;
  assign n7816 = x94 & n631 ;
  assign n7817 = x93 & ~n630 ;
  assign n7818 = n764 & n7817 ;
  assign n7819 = n7816 | n7818 ;
  assign n7820 = n7815 | n7819 ;
  assign n7821 = n639 | n7815 ;
  assign n7822 = n7819 | n7821 ;
  assign n7823 = ( n4897 & n7820 ) | ( n4897 & n7822 ) | ( n7820 & n7822 ) ;
  assign n7824 = x11 & n7822 ;
  assign n7825 = x11 & n7815 ;
  assign n7826 = ( x11 & n7819 ) | ( x11 & n7825 ) | ( n7819 & n7825 ) ;
  assign n7827 = ( n4897 & n7824 ) | ( n4897 & n7826 ) | ( n7824 & n7826 ) ;
  assign n7828 = x11 & ~n7826 ;
  assign n7829 = x11 & ~n7822 ;
  assign n7830 = ( ~n4897 & n7828 ) | ( ~n4897 & n7829 ) | ( n7828 & n7829 ) ;
  assign n7831 = ( n7823 & ~n7827 ) | ( n7823 & n7830 ) | ( ~n7827 & n7830 ) ;
  assign n7832 = n7814 | n7831 ;
  assign n7833 = n7814 & n7831 ;
  assign n7834 = n7832 & ~n7833 ;
  assign n7835 = n7454 | n7457 ;
  assign n7836 = ( n7454 & n7456 ) | ( n7454 & n7835 ) | ( n7456 & n7835 ) ;
  assign n7837 = n7834 & n7836 ;
  assign n7838 = n7834 | n7836 ;
  assign n7839 = ~n7837 & n7838 ;
  assign n7840 = x98 & n389 ;
  assign n7841 = x97 & n384 ;
  assign n7842 = x96 & ~n383 ;
  assign n7843 = n463 & n7842 ;
  assign n7844 = n7841 | n7843 ;
  assign n7845 = n7840 | n7844 ;
  assign n7846 = n392 | n7840 ;
  assign n7847 = n7844 | n7846 ;
  assign n7848 = ( ~n5850 & n7845 ) | ( ~n5850 & n7847 ) | ( n7845 & n7847 ) ;
  assign n7849 = n7845 & n7847 ;
  assign n7850 = ( n5834 & n7848 ) | ( n5834 & n7849 ) | ( n7848 & n7849 ) ;
  assign n7851 = x8 & n7847 ;
  assign n7852 = x8 & n7840 ;
  assign n7853 = ( x8 & n7844 ) | ( x8 & n7852 ) | ( n7844 & n7852 ) ;
  assign n7854 = ( ~n5850 & n7851 ) | ( ~n5850 & n7853 ) | ( n7851 & n7853 ) ;
  assign n7855 = n7851 & n7853 ;
  assign n7856 = ( n5834 & n7854 ) | ( n5834 & n7855 ) | ( n7854 & n7855 ) ;
  assign n7857 = x8 & ~n7853 ;
  assign n7858 = x8 & ~n7847 ;
  assign n7859 = ( n5850 & n7857 ) | ( n5850 & n7858 ) | ( n7857 & n7858 ) ;
  assign n7860 = n7857 | n7858 ;
  assign n7861 = ( ~n5834 & n7859 ) | ( ~n5834 & n7860 ) | ( n7859 & n7860 ) ;
  assign n7862 = ( n7850 & ~n7856 ) | ( n7850 & n7861 ) | ( ~n7856 & n7861 ) ;
  assign n7863 = n7839 | n7862 ;
  assign n7864 = n7839 & n7862 ;
  assign n7865 = n7863 & ~n7864 ;
  assign n7866 = ( n7460 & n7477 ) | ( n7460 & n7482 ) | ( n7477 & n7482 ) ;
  assign n7867 = n7865 | n7866 ;
  assign n7868 = n7865 & n7866 ;
  assign n7869 = n7867 & ~n7868 ;
  assign n7870 = x101 & n212 ;
  assign n7871 = x100 & n207 ;
  assign n7872 = x99 & ~n206 ;
  assign n7873 = n267 & n7872 ;
  assign n7874 = n7871 | n7873 ;
  assign n7875 = n7870 | n7874 ;
  assign n7876 = n215 | n7870 ;
  assign n7877 = n7874 | n7876 ;
  assign n7878 = ( n6844 & n7875 ) | ( n6844 & n7877 ) | ( n7875 & n7877 ) ;
  assign n7879 = x5 & n7877 ;
  assign n7880 = x5 & n7870 ;
  assign n7881 = ( x5 & n7874 ) | ( x5 & n7880 ) | ( n7874 & n7880 ) ;
  assign n7882 = ( n6844 & n7879 ) | ( n6844 & n7881 ) | ( n7879 & n7881 ) ;
  assign n7883 = x5 & ~n7881 ;
  assign n7884 = x5 & ~n7877 ;
  assign n7885 = ( ~n6844 & n7883 ) | ( ~n6844 & n7884 ) | ( n7883 & n7884 ) ;
  assign n7886 = ( n7878 & ~n7882 ) | ( n7878 & n7885 ) | ( ~n7882 & n7885 ) ;
  assign n7887 = n7869 & n7886 ;
  assign n7888 = n7869 & ~n7887 ;
  assign n7889 = ~n7869 & n7886 ;
  assign n7890 = n7888 | n7889 ;
  assign n7891 = n7506 | n7507 ;
  assign n7892 = ( n7203 & n7506 ) | ( n7203 & n7891 ) | ( n7506 & n7891 ) ;
  assign n7893 = ~n7890 & n7892 ;
  assign n7894 = n7890 & ~n7892 ;
  assign n7895 = n7893 | n7894 ;
  assign n7896 = x103 | x104 ;
  assign n7897 = x103 & x104 ;
  assign n7898 = n7896 & ~n7897 ;
  assign n7899 = n7512 & n7898 ;
  assign n7900 = ( n7517 & n7898 ) | ( n7517 & n7899 ) | ( n7898 & n7899 ) ;
  assign n7901 = ( n7518 & n7898 ) | ( n7518 & n7899 ) | ( n7898 & n7899 ) ;
  assign n7902 = ( n6159 & n7900 ) | ( n6159 & n7901 ) | ( n7900 & n7901 ) ;
  assign n7903 = ( n6157 & n7900 ) | ( n6157 & n7901 ) | ( n7900 & n7901 ) ;
  assign n7904 = ( n5823 & n7902 ) | ( n5823 & n7903 ) | ( n7902 & n7903 ) ;
  assign n7905 = n7512 | n7898 ;
  assign n7906 = n7518 | n7905 ;
  assign n7907 = n7517 | n7905 ;
  assign n7908 = ( n6159 & n7906 ) | ( n6159 & n7907 ) | ( n7906 & n7907 ) ;
  assign n7909 = ( n6157 & n7906 ) | ( n6157 & n7907 ) | ( n7906 & n7907 ) ;
  assign n7910 = ( n5823 & n7908 ) | ( n5823 & n7909 ) | ( n7908 & n7909 ) ;
  assign n7911 = ~n7904 & n7910 ;
  assign n7912 = x103 & n133 ;
  assign n7913 = x102 & ~n162 ;
  assign n7914 = ( n137 & n7912 ) | ( n137 & n7913 ) | ( n7912 & n7913 ) ;
  assign n7915 = x0 & x104 ;
  assign n7916 = ( ~n137 & n7912 ) | ( ~n137 & n7915 ) | ( n7912 & n7915 ) ;
  assign n7917 = n7914 | n7916 ;
  assign n7918 = n141 | n7917 ;
  assign n7919 = ( n7911 & n7917 ) | ( n7911 & n7918 ) | ( n7917 & n7918 ) ;
  assign n7920 = x2 & n7917 ;
  assign n7921 = ( x2 & n523 ) | ( x2 & n7917 ) | ( n523 & n7917 ) ;
  assign n7922 = ( n7911 & n7920 ) | ( n7911 & n7921 ) | ( n7920 & n7921 ) ;
  assign n7923 = x2 & ~n7921 ;
  assign n7924 = x2 & ~n7917 ;
  assign n7925 = ( ~n7911 & n7923 ) | ( ~n7911 & n7924 ) | ( n7923 & n7924 ) ;
  assign n7926 = ( n7919 & ~n7922 ) | ( n7919 & n7925 ) | ( ~n7922 & n7925 ) ;
  assign n7927 = n7895 & n7926 ;
  assign n7928 = n7895 | n7926 ;
  assign n7929 = ~n7927 & n7928 ;
  assign n7930 = n7553 & n7929 ;
  assign n7931 = n7553 | n7929 ;
  assign n7932 = ~n7930 & n7931 ;
  assign n7933 = x75 & n4631 ;
  assign n7934 = x74 & n4626 ;
  assign n7935 = x73 & ~n4625 ;
  assign n7936 = n4943 & n7935 ;
  assign n7937 = n7934 | n7936 ;
  assign n7938 = n7933 | n7937 ;
  assign n7939 = n4634 | n7933 ;
  assign n7940 = n7937 | n7939 ;
  assign n7941 = ( n746 & n7938 ) | ( n746 & n7940 ) | ( n7938 & n7940 ) ;
  assign n7942 = x32 & n7940 ;
  assign n7943 = x32 & n7933 ;
  assign n7944 = ( x32 & n7937 ) | ( x32 & n7943 ) | ( n7937 & n7943 ) ;
  assign n7945 = ( n746 & n7942 ) | ( n746 & n7944 ) | ( n7942 & n7944 ) ;
  assign n7946 = x32 & ~n7944 ;
  assign n7947 = x32 & ~n7940 ;
  assign n7948 = ( ~n746 & n7946 ) | ( ~n746 & n7947 ) | ( n7946 & n7947 ) ;
  assign n7949 = ( n7941 & ~n7945 ) | ( n7941 & n7948 ) | ( ~n7945 & n7948 ) ;
  assign n7950 = n7625 | n7631 ;
  assign n7951 = x66 & n7566 ;
  assign n7952 = x65 & n7561 ;
  assign n7953 = ~n7207 & n7565 ;
  assign n7954 = x64 & ~n7560 ;
  assign n7955 = n7953 & n7954 ;
  assign n7956 = n7952 | n7955 ;
  assign n7957 = n7951 | n7956 ;
  assign n7958 = n159 & n7569 ;
  assign n7959 = n7957 | n7958 ;
  assign n7960 = x41 | n7569 ;
  assign n7961 = ( x41 & n159 ) | ( x41 & n7960 ) | ( n159 & n7960 ) ;
  assign n7962 = n7957 | n7961 ;
  assign n7963 = ~x41 & n7961 ;
  assign n7964 = ( ~x41 & n7957 ) | ( ~x41 & n7963 ) | ( n7957 & n7963 ) ;
  assign n7965 = ( ~n7959 & n7962 ) | ( ~n7959 & n7964 ) | ( n7962 & n7964 ) ;
  assign n7966 = n7581 | n7965 ;
  assign n7967 = n7581 & n7965 ;
  assign n7968 = n7966 & ~n7967 ;
  assign n7969 = n293 & n6539 ;
  assign n7970 = x69 & n6536 ;
  assign n7971 = x68 & n6531 ;
  assign n7972 = x67 & ~n6530 ;
  assign n7973 = n6871 & n7972 ;
  assign n7974 = n7971 | n7973 ;
  assign n7975 = n7970 | n7974 ;
  assign n7976 = n7969 | n7975 ;
  assign n7977 = x38 | n7970 ;
  assign n7978 = n7974 | n7977 ;
  assign n7979 = n7969 | n7978 ;
  assign n7980 = ~x38 & n7978 ;
  assign n7981 = ( ~x38 & n7969 ) | ( ~x38 & n7980 ) | ( n7969 & n7980 ) ;
  assign n7982 = ( ~n7976 & n7979 ) | ( ~n7976 & n7981 ) | ( n7979 & n7981 ) ;
  assign n7983 = n7968 & n7982 ;
  assign n7984 = n7968 & ~n7983 ;
  assign n7985 = ~n7968 & n7982 ;
  assign n7986 = n7984 | n7985 ;
  assign n7987 = n7603 | n7605 ;
  assign n7988 = ( n7603 & n7604 ) | ( n7603 & n7987 ) | ( n7604 & n7987 ) ;
  assign n7989 = n7986 & n7988 ;
  assign n7990 = n7986 | n7988 ;
  assign n7991 = ~n7989 & n7990 ;
  assign n7992 = x72 & n5554 ;
  assign n7993 = x71 & n5549 ;
  assign n7994 = x70 & ~n5548 ;
  assign n7995 = n5893 & n7994 ;
  assign n7996 = n7993 | n7995 ;
  assign n7997 = n7992 | n7996 ;
  assign n7998 = ( n513 & n5557 ) | ( n513 & n7997 ) | ( n5557 & n7997 ) ;
  assign n7999 = ( x35 & n5557 ) | ( x35 & ~n7992 ) | ( n5557 & ~n7992 ) ;
  assign n8000 = x35 & n5557 ;
  assign n8001 = ( ~n7996 & n7999 ) | ( ~n7996 & n8000 ) | ( n7999 & n8000 ) ;
  assign n8002 = ( x35 & n513 ) | ( x35 & n8001 ) | ( n513 & n8001 ) ;
  assign n8003 = ~n7998 & n8002 ;
  assign n8004 = n7997 | n8001 ;
  assign n8005 = x35 | n7997 ;
  assign n8006 = ( n513 & n8004 ) | ( n513 & n8005 ) | ( n8004 & n8005 ) ;
  assign n8007 = ( ~x35 & n8003 ) | ( ~x35 & n8006 ) | ( n8003 & n8006 ) ;
  assign n8008 = n7991 & n8007 ;
  assign n8009 = n7991 & ~n8008 ;
  assign n8010 = ~n7991 & n8007 ;
  assign n8011 = n8009 | n8010 ;
  assign n8012 = ~n7950 & n8011 ;
  assign n8013 = n7949 & n8012 ;
  assign n8014 = n7950 & ~n8011 ;
  assign n8015 = ( n7949 & n8013 ) | ( n7949 & n8014 ) | ( n8013 & n8014 ) ;
  assign n8016 = n7949 | n8012 ;
  assign n8017 = n8014 | n8016 ;
  assign n8018 = ~n8015 & n8017 ;
  assign n8019 = n7650 | n7654 ;
  assign n8020 = n7650 | n7651 ;
  assign n8021 = ( n7275 & n8019 ) | ( n7275 & n8020 ) | ( n8019 & n8020 ) ;
  assign n8022 = n8018 & n8021 ;
  assign n8023 = n8018 | n8021 ;
  assign n8024 = ~n8022 & n8023 ;
  assign n8025 = x78 & n3816 ;
  assign n8026 = x77 & n3811 ;
  assign n8027 = x76 & ~n3810 ;
  assign n8028 = n4067 & n8027 ;
  assign n8029 = n8026 | n8028 ;
  assign n8030 = n8025 | n8029 ;
  assign n8031 = n3819 | n8025 ;
  assign n8032 = n8029 | n8031 ;
  assign n8033 = ( n1192 & n8030 ) | ( n1192 & n8032 ) | ( n8030 & n8032 ) ;
  assign n8034 = x29 & n8032 ;
  assign n8035 = x29 & n8025 ;
  assign n8036 = ( x29 & n8029 ) | ( x29 & n8035 ) | ( n8029 & n8035 ) ;
  assign n8037 = ( n1192 & n8034 ) | ( n1192 & n8036 ) | ( n8034 & n8036 ) ;
  assign n8038 = x29 & ~n8036 ;
  assign n8039 = x29 & ~n8032 ;
  assign n8040 = ( ~n1192 & n8038 ) | ( ~n1192 & n8039 ) | ( n8038 & n8039 ) ;
  assign n8041 = ( n8033 & ~n8037 ) | ( n8033 & n8040 ) | ( ~n8037 & n8040 ) ;
  assign n8042 = n8024 | n8041 ;
  assign n8043 = n8024 & n8041 ;
  assign n8044 = n8042 & ~n8043 ;
  assign n8045 = n7678 | n7682 ;
  assign n8046 = ( n7678 & n7684 ) | ( n7678 & n8045 ) | ( n7684 & n8045 ) ;
  assign n8047 = n8044 & n8046 ;
  assign n8048 = n8044 | n8046 ;
  assign n8049 = ~n8047 & n8048 ;
  assign n8050 = x81 & n3085 ;
  assign n8051 = x80 & n3080 ;
  assign n8052 = x79 & ~n3079 ;
  assign n8053 = n3309 & n8052 ;
  assign n8054 = n8051 | n8053 ;
  assign n8055 = n8050 | n8054 ;
  assign n8056 = n3088 | n8050 ;
  assign n8057 = n8054 | n8056 ;
  assign n8058 = ( n1651 & n8055 ) | ( n1651 & n8057 ) | ( n8055 & n8057 ) ;
  assign n8059 = x26 & n8057 ;
  assign n8060 = x26 & n8050 ;
  assign n8061 = ( x26 & n8054 ) | ( x26 & n8060 ) | ( n8054 & n8060 ) ;
  assign n8062 = ( n1651 & n8059 ) | ( n1651 & n8061 ) | ( n8059 & n8061 ) ;
  assign n8063 = x26 & ~n8061 ;
  assign n8064 = x26 & ~n8057 ;
  assign n8065 = ( ~n1651 & n8063 ) | ( ~n1651 & n8064 ) | ( n8063 & n8064 ) ;
  assign n8066 = ( n8058 & ~n8062 ) | ( n8058 & n8065 ) | ( ~n8062 & n8065 ) ;
  assign n8067 = n8049 | n8066 ;
  assign n8068 = n8049 & n8066 ;
  assign n8069 = n8067 & ~n8068 ;
  assign n8070 = n7705 | n7709 ;
  assign n8071 = ( n7705 & n7708 ) | ( n7705 & n8070 ) | ( n7708 & n8070 ) ;
  assign n8072 = n8069 & n8071 ;
  assign n8073 = n8069 | n8071 ;
  assign n8074 = ~n8072 & n8073 ;
  assign n8075 = x84 & n2429 ;
  assign n8076 = x83 & n2424 ;
  assign n8077 = x82 & ~n2423 ;
  assign n8078 = n2631 & n8077 ;
  assign n8079 = n8076 | n8078 ;
  assign n8080 = n8075 | n8079 ;
  assign n8081 = n2432 | n8075 ;
  assign n8082 = n8079 | n8081 ;
  assign n8083 = ( n2194 & n8080 ) | ( n2194 & n8082 ) | ( n8080 & n8082 ) ;
  assign n8084 = x23 & n8082 ;
  assign n8085 = x23 & n8075 ;
  assign n8086 = ( x23 & n8079 ) | ( x23 & n8085 ) | ( n8079 & n8085 ) ;
  assign n8087 = ( n2194 & n8084 ) | ( n2194 & n8086 ) | ( n8084 & n8086 ) ;
  assign n8088 = x23 & ~n8086 ;
  assign n8089 = x23 & ~n8082 ;
  assign n8090 = ( ~n2194 & n8088 ) | ( ~n2194 & n8089 ) | ( n8088 & n8089 ) ;
  assign n8091 = ( n8083 & ~n8087 ) | ( n8083 & n8090 ) | ( ~n8087 & n8090 ) ;
  assign n8092 = n8074 & n8091 ;
  assign n8093 = n8074 & ~n8092 ;
  assign n8094 = ~n8074 & n8091 ;
  assign n8095 = n8093 | n8094 ;
  assign n8096 = n7730 | n7736 ;
  assign n8097 = n8095 | n8096 ;
  assign n8098 = n8095 & n8096 ;
  assign n8099 = n8097 & ~n8098 ;
  assign n8100 = x87 & n1859 ;
  assign n8101 = x86 & n1854 ;
  assign n8102 = x85 & ~n1853 ;
  assign n8103 = n2037 & n8102 ;
  assign n8104 = n8101 | n8103 ;
  assign n8105 = n8100 | n8104 ;
  assign n8106 = n1862 | n8100 ;
  assign n8107 = n8104 | n8106 ;
  assign n8108 = ( n2816 & n8105 ) | ( n2816 & n8107 ) | ( n8105 & n8107 ) ;
  assign n8109 = x20 & n8107 ;
  assign n8110 = x20 & n8100 ;
  assign n8111 = ( x20 & n8104 ) | ( x20 & n8110 ) | ( n8104 & n8110 ) ;
  assign n8112 = ( n2816 & n8109 ) | ( n2816 & n8111 ) | ( n8109 & n8111 ) ;
  assign n8113 = x20 & ~n8111 ;
  assign n8114 = x20 & ~n8107 ;
  assign n8115 = ( ~n2816 & n8113 ) | ( ~n2816 & n8114 ) | ( n8113 & n8114 ) ;
  assign n8116 = ( n8108 & ~n8112 ) | ( n8108 & n8115 ) | ( ~n8112 & n8115 ) ;
  assign n8117 = n8099 | n8116 ;
  assign n8118 = n8099 & n8116 ;
  assign n8119 = n7755 | n7761 ;
  assign n8120 = n8117 & ~n8118 ;
  assign n8121 = n8118 | n8120 ;
  assign n8122 = ( n8118 & n8119 ) | ( n8118 & n8121 ) | ( n8119 & n8121 ) ;
  assign n8123 = n8117 & ~n8122 ;
  assign n8124 = x90 & n1383 ;
  assign n8125 = x89 & n1378 ;
  assign n8126 = x88 & ~n1377 ;
  assign n8127 = n1542 & n8126 ;
  assign n8128 = n8125 | n8127 ;
  assign n8129 = n8124 | n8128 ;
  assign n8130 = n1386 | n8124 ;
  assign n8131 = n8128 | n8130 ;
  assign n8132 = ( n3519 & n8129 ) | ( n3519 & n8131 ) | ( n8129 & n8131 ) ;
  assign n8133 = x17 & n8131 ;
  assign n8134 = x17 & n8124 ;
  assign n8135 = ( x17 & n8128 ) | ( x17 & n8134 ) | ( n8128 & n8134 ) ;
  assign n8136 = ( n3519 & n8133 ) | ( n3519 & n8135 ) | ( n8133 & n8135 ) ;
  assign n8137 = x17 & ~n8135 ;
  assign n8138 = x17 & ~n8131 ;
  assign n8139 = ( ~n3519 & n8137 ) | ( ~n3519 & n8138 ) | ( n8137 & n8138 ) ;
  assign n8140 = ( n8132 & ~n8136 ) | ( n8132 & n8139 ) | ( ~n8136 & n8139 ) ;
  assign n8141 = ~n8120 & n8140 ;
  assign n8142 = n8119 & n8141 ;
  assign n8143 = ( n8123 & n8140 ) | ( n8123 & n8142 ) | ( n8140 & n8142 ) ;
  assign n8144 = n8120 & ~n8140 ;
  assign n8145 = ( n8119 & n8140 ) | ( n8119 & ~n8144 ) | ( n8140 & ~n8144 ) ;
  assign n8146 = n8123 | n8145 ;
  assign n8147 = ~n8143 & n8146 ;
  assign n8148 = n7780 | n7785 ;
  assign n8149 = ( n7780 & n7783 ) | ( n7780 & n8148 ) | ( n7783 & n8148 ) ;
  assign n8150 = n8147 & n8149 ;
  assign n8151 = n8147 | n8149 ;
  assign n8152 = ~n8150 & n8151 ;
  assign n8153 = x93 & n962 ;
  assign n8154 = x92 & n957 ;
  assign n8155 = x91 & ~n956 ;
  assign n8156 = n1105 & n8155 ;
  assign n8157 = n8154 | n8156 ;
  assign n8158 = n8153 | n8157 ;
  assign n8159 = n965 | n8153 ;
  assign n8160 = n8157 | n8159 ;
  assign n8161 = ( n4305 & n8158 ) | ( n4305 & n8160 ) | ( n8158 & n8160 ) ;
  assign n8162 = x14 & n8160 ;
  assign n8163 = x14 & n8153 ;
  assign n8164 = ( x14 & n8157 ) | ( x14 & n8163 ) | ( n8157 & n8163 ) ;
  assign n8165 = ( n4305 & n8162 ) | ( n4305 & n8164 ) | ( n8162 & n8164 ) ;
  assign n8166 = x14 & ~n8164 ;
  assign n8167 = x14 & ~n8160 ;
  assign n8168 = ( ~n4305 & n8166 ) | ( ~n4305 & n8167 ) | ( n8166 & n8167 ) ;
  assign n8169 = ( n8161 & ~n8165 ) | ( n8161 & n8168 ) | ( ~n8165 & n8168 ) ;
  assign n8170 = n8152 | n8169 ;
  assign n8171 = n8152 & n8169 ;
  assign n8172 = n8170 & ~n8171 ;
  assign n8173 = n7806 & n8172 ;
  assign n8174 = ( n7810 & n8172 ) | ( n7810 & n8173 ) | ( n8172 & n8173 ) ;
  assign n8175 = n7806 | n8172 ;
  assign n8176 = n7810 | n8175 ;
  assign n8177 = ~n8174 & n8176 ;
  assign n8178 = x96 & n636 ;
  assign n8179 = x95 & n631 ;
  assign n8180 = x94 & ~n630 ;
  assign n8181 = n764 & n8180 ;
  assign n8182 = n8179 | n8181 ;
  assign n8183 = n8178 | n8182 ;
  assign n8184 = n639 | n8178 ;
  assign n8185 = n8182 | n8184 ;
  assign n8186 = ( n5202 & n8183 ) | ( n5202 & n8185 ) | ( n8183 & n8185 ) ;
  assign n8187 = x11 & n8185 ;
  assign n8188 = x11 & n8178 ;
  assign n8189 = ( x11 & n8182 ) | ( x11 & n8188 ) | ( n8182 & n8188 ) ;
  assign n8190 = ( n5202 & n8187 ) | ( n5202 & n8189 ) | ( n8187 & n8189 ) ;
  assign n8191 = x11 & ~n8189 ;
  assign n8192 = x11 & ~n8185 ;
  assign n8193 = ( ~n5202 & n8191 ) | ( ~n5202 & n8192 ) | ( n8191 & n8192 ) ;
  assign n8194 = ( n8186 & ~n8190 ) | ( n8186 & n8193 ) | ( ~n8190 & n8193 ) ;
  assign n8195 = n8177 | n8194 ;
  assign n8196 = n8177 & n8194 ;
  assign n8197 = n8195 & ~n8196 ;
  assign n8198 = n7833 | n7836 ;
  assign n8199 = ( n7833 & n7834 ) | ( n7833 & n8198 ) | ( n7834 & n8198 ) ;
  assign n8200 = n8197 & n8199 ;
  assign n8201 = n8197 | n8199 ;
  assign n8202 = ~n8200 & n8201 ;
  assign n8203 = x99 & n389 ;
  assign n8204 = x98 & n384 ;
  assign n8205 = x97 & ~n383 ;
  assign n8206 = n463 & n8205 ;
  assign n8207 = n8204 | n8206 ;
  assign n8208 = n8203 | n8207 ;
  assign n8209 = n392 | n8203 ;
  assign n8210 = n8207 | n8209 ;
  assign n8211 = ( n6164 & n8208 ) | ( n6164 & n8210 ) | ( n8208 & n8210 ) ;
  assign n8212 = x8 & n8210 ;
  assign n8213 = x8 & n8203 ;
  assign n8214 = ( x8 & n8207 ) | ( x8 & n8213 ) | ( n8207 & n8213 ) ;
  assign n8215 = ( n6164 & n8212 ) | ( n6164 & n8214 ) | ( n8212 & n8214 ) ;
  assign n8216 = x8 & ~n8214 ;
  assign n8217 = x8 & ~n8210 ;
  assign n8218 = ( ~n6164 & n8216 ) | ( ~n6164 & n8217 ) | ( n8216 & n8217 ) ;
  assign n8219 = ( n8211 & ~n8215 ) | ( n8211 & n8218 ) | ( ~n8215 & n8218 ) ;
  assign n8220 = n8202 & n8219 ;
  assign n8221 = n8202 & ~n8220 ;
  assign n8222 = ~n8202 & n8219 ;
  assign n8223 = n8221 | n8222 ;
  assign n8224 = n7864 | n7866 ;
  assign n8225 = ( n7864 & n7865 ) | ( n7864 & n8224 ) | ( n7865 & n8224 ) ;
  assign n8226 = ~n8223 & n8225 ;
  assign n8227 = n8223 & ~n8225 ;
  assign n8228 = n8226 | n8227 ;
  assign n8229 = x102 & n212 ;
  assign n8230 = x101 & n207 ;
  assign n8231 = x100 & ~n206 ;
  assign n8232 = n267 & n8231 ;
  assign n8233 = n8230 | n8232 ;
  assign n8234 = n8229 | n8233 ;
  assign n8235 = n215 | n8229 ;
  assign n8236 = n8233 | n8235 ;
  assign n8237 = ( n7178 & n8234 ) | ( n7178 & n8236 ) | ( n8234 & n8236 ) ;
  assign n8238 = x5 & n8236 ;
  assign n8239 = x5 & n8229 ;
  assign n8240 = ( x5 & n8233 ) | ( x5 & n8239 ) | ( n8233 & n8239 ) ;
  assign n8241 = ( n7178 & n8238 ) | ( n7178 & n8240 ) | ( n8238 & n8240 ) ;
  assign n8242 = x5 & ~n8240 ;
  assign n8243 = x5 & ~n8236 ;
  assign n8244 = ( ~n7178 & n8242 ) | ( ~n7178 & n8243 ) | ( n8242 & n8243 ) ;
  assign n8245 = ( n8237 & ~n8241 ) | ( n8237 & n8244 ) | ( ~n8241 & n8244 ) ;
  assign n8246 = n8228 & n8245 ;
  assign n8247 = n8228 | n8245 ;
  assign n8248 = ~n8246 & n8247 ;
  assign n8249 = ( n7869 & n7886 ) | ( n7869 & n7892 ) | ( n7886 & n7892 ) ;
  assign n8250 = n8248 | n8249 ;
  assign n8251 = n8248 & n8249 ;
  assign n8252 = n8250 & ~n8251 ;
  assign n8253 = x104 | x105 ;
  assign n8254 = x104 & x105 ;
  assign n8255 = n8253 & ~n8254 ;
  assign n8256 = n7512 | n7897 ;
  assign n8257 = ( n7897 & n7898 ) | ( n7897 & n8256 ) | ( n7898 & n8256 ) ;
  assign n8258 = n8255 & n8257 ;
  assign n8259 = n7897 | n7898 ;
  assign n8260 = n8255 & n8259 ;
  assign n8261 = ( n7517 & n8258 ) | ( n7517 & n8260 ) | ( n8258 & n8260 ) ;
  assign n8262 = ( n7518 & n8258 ) | ( n7518 & n8260 ) | ( n8258 & n8260 ) ;
  assign n8263 = ( n6159 & n8261 ) | ( n6159 & n8262 ) | ( n8261 & n8262 ) ;
  assign n8264 = ( n6157 & n8261 ) | ( n6157 & n8262 ) | ( n8261 & n8262 ) ;
  assign n8265 = ( n5823 & n8263 ) | ( n5823 & n8264 ) | ( n8263 & n8264 ) ;
  assign n8266 = n8255 | n8257 ;
  assign n8267 = n8255 | n8259 ;
  assign n8268 = ( n7518 & n8266 ) | ( n7518 & n8267 ) | ( n8266 & n8267 ) ;
  assign n8269 = ( n7517 & n8266 ) | ( n7517 & n8267 ) | ( n8266 & n8267 ) ;
  assign n8270 = ( n6159 & n8268 ) | ( n6159 & n8269 ) | ( n8268 & n8269 ) ;
  assign n8271 = ( n6157 & n8268 ) | ( n6157 & n8269 ) | ( n8268 & n8269 ) ;
  assign n8272 = ( n5823 & n8270 ) | ( n5823 & n8271 ) | ( n8270 & n8271 ) ;
  assign n8273 = ~n8265 & n8272 ;
  assign n8274 = x104 & n133 ;
  assign n8275 = x103 & ~n162 ;
  assign n8276 = ( n137 & n8274 ) | ( n137 & n8275 ) | ( n8274 & n8275 ) ;
  assign n8277 = x0 & x105 ;
  assign n8278 = ( ~n137 & n8274 ) | ( ~n137 & n8277 ) | ( n8274 & n8277 ) ;
  assign n8279 = n8276 | n8278 ;
  assign n8280 = n141 | n8279 ;
  assign n8281 = ( n8273 & n8279 ) | ( n8273 & n8280 ) | ( n8279 & n8280 ) ;
  assign n8282 = x2 & n8279 ;
  assign n8283 = ( x2 & n523 ) | ( x2 & n8279 ) | ( n523 & n8279 ) ;
  assign n8284 = ( n8273 & n8282 ) | ( n8273 & n8283 ) | ( n8282 & n8283 ) ;
  assign n8285 = x2 & ~n8283 ;
  assign n8286 = x2 & ~n8279 ;
  assign n8287 = ( ~n8273 & n8285 ) | ( ~n8273 & n8286 ) | ( n8285 & n8286 ) ;
  assign n8288 = ( n8281 & ~n8284 ) | ( n8281 & n8287 ) | ( ~n8284 & n8287 ) ;
  assign n8289 = n8252 | n8288 ;
  assign n8290 = n8252 & n8288 ;
  assign n8291 = n8289 & ~n8290 ;
  assign n8292 = n7927 | n7929 ;
  assign n8293 = ( n7553 & n7927 ) | ( n7553 & n8292 ) | ( n7927 & n8292 ) ;
  assign n8294 = n8291 & n8293 ;
  assign n8295 = n8291 | n8293 ;
  assign n8296 = ~n8294 & n8295 ;
  assign n8297 = n8143 | n8150 ;
  assign n8298 = x41 & ~x42 ;
  assign n8299 = ~x41 & x42 ;
  assign n8300 = n8298 | n8299 ;
  assign n8301 = x64 & n8300 ;
  assign n8302 = ~n7581 & n8301 ;
  assign n8303 = ( ~n7965 & n8301 ) | ( ~n7965 & n8302 ) | ( n8301 & n8302 ) ;
  assign n8304 = n7581 & ~n8301 ;
  assign n8305 = n7965 & n8304 ;
  assign n8306 = n8303 | n8305 ;
  assign n8307 = x67 & n7566 ;
  assign n8308 = x66 & n7561 ;
  assign n8309 = x65 & ~n7560 ;
  assign n8310 = n7953 & n8309 ;
  assign n8311 = n8308 | n8310 ;
  assign n8312 = n8307 | n8311 ;
  assign n8313 = n186 & n7569 ;
  assign n8314 = n8312 | n8313 ;
  assign n8315 = x41 & ~n8314 ;
  assign n8316 = ~x41 & n8314 ;
  assign n8317 = n8315 | n8316 ;
  assign n8318 = n8306 & n8317 ;
  assign n8319 = n8306 | n8317 ;
  assign n8320 = ~n8318 & n8319 ;
  assign n8321 = x69 & n6531 ;
  assign n8322 = x68 & ~n6530 ;
  assign n8323 = n6871 & n8322 ;
  assign n8324 = n8321 | n8323 ;
  assign n8325 = x70 & n6536 ;
  assign n8326 = n6539 | n8325 ;
  assign n8327 = n8324 | n8326 ;
  assign n8328 = x38 & ~n8327 ;
  assign n8329 = x38 & ~n8325 ;
  assign n8330 = ~n8324 & n8329 ;
  assign n8331 = ( ~n340 & n8328 ) | ( ~n340 & n8330 ) | ( n8328 & n8330 ) ;
  assign n8332 = ~x38 & n8327 ;
  assign n8333 = ~x38 & n8325 ;
  assign n8334 = ( ~x38 & n8324 ) | ( ~x38 & n8333 ) | ( n8324 & n8333 ) ;
  assign n8335 = ( n340 & n8332 ) | ( n340 & n8334 ) | ( n8332 & n8334 ) ;
  assign n8336 = n8331 | n8335 ;
  assign n8337 = n8320 & n8336 ;
  assign n8338 = n8320 & ~n8337 ;
  assign n8339 = ~n8320 & n8336 ;
  assign n8340 = n8338 | n8339 ;
  assign n8341 = n7983 | n7988 ;
  assign n8342 = ( n7983 & n7986 ) | ( n7983 & n8341 ) | ( n7986 & n8341 ) ;
  assign n8343 = n8340 | n8342 ;
  assign n8344 = n8340 & n8342 ;
  assign n8345 = n8343 & ~n8344 ;
  assign n8346 = x73 & n5554 ;
  assign n8347 = x72 & n5549 ;
  assign n8348 = x71 & ~n5548 ;
  assign n8349 = n5893 & n8348 ;
  assign n8350 = n8347 | n8349 ;
  assign n8351 = n8346 | n8350 ;
  assign n8352 = ( ~n610 & n5557 ) | ( ~n610 & n8351 ) | ( n5557 & n8351 ) ;
  assign n8353 = n5557 & n8346 ;
  assign n8354 = ( n5557 & n8350 ) | ( n5557 & n8353 ) | ( n8350 & n8353 ) ;
  assign n8355 = ( n598 & n8352 ) | ( n598 & n8354 ) | ( n8352 & n8354 ) ;
  assign n8356 = ( x35 & ~n8351 ) | ( x35 & n8355 ) | ( ~n8351 & n8355 ) ;
  assign n8357 = ~n8355 & n8356 ;
  assign n8358 = x35 | n8346 ;
  assign n8359 = n8350 | n8358 ;
  assign n8360 = n8355 | n8359 ;
  assign n8361 = ( ~x35 & n8357 ) | ( ~x35 & n8360 ) | ( n8357 & n8360 ) ;
  assign n8362 = n8345 | n8361 ;
  assign n8363 = n8345 & n8361 ;
  assign n8364 = n8362 & ~n8363 ;
  assign n8365 = n7950 & n8011 ;
  assign n8366 = n8008 | n8365 ;
  assign n8367 = n8364 & n8366 ;
  assign n8368 = n8364 | n8366 ;
  assign n8369 = ~n8367 & n8368 ;
  assign n8370 = x76 & n4631 ;
  assign n8371 = x75 & n4626 ;
  assign n8372 = x74 & ~n4625 ;
  assign n8373 = n4943 & n8372 ;
  assign n8374 = n8371 | n8373 ;
  assign n8375 = n8370 | n8374 ;
  assign n8376 = n4634 | n8370 ;
  assign n8377 = n8374 | n8376 ;
  assign n8378 = ( n923 & n8375 ) | ( n923 & n8377 ) | ( n8375 & n8377 ) ;
  assign n8379 = x32 & n8377 ;
  assign n8380 = x32 & n8370 ;
  assign n8381 = ( x32 & n8374 ) | ( x32 & n8380 ) | ( n8374 & n8380 ) ;
  assign n8382 = ( n923 & n8379 ) | ( n923 & n8381 ) | ( n8379 & n8381 ) ;
  assign n8383 = x32 & ~n8381 ;
  assign n8384 = x32 & ~n8377 ;
  assign n8385 = ( ~n923 & n8383 ) | ( ~n923 & n8384 ) | ( n8383 & n8384 ) ;
  assign n8386 = ( n8378 & ~n8382 ) | ( n8378 & n8385 ) | ( ~n8382 & n8385 ) ;
  assign n8387 = n8369 & n8386 ;
  assign n8388 = n8369 & ~n8387 ;
  assign n8389 = ~n8369 & n8386 ;
  assign n8390 = n8388 | n8389 ;
  assign n8391 = n8015 | n8021 ;
  assign n8392 = ( n8015 & n8018 ) | ( n8015 & n8391 ) | ( n8018 & n8391 ) ;
  assign n8393 = n8389 & n8392 ;
  assign n8394 = ( n8388 & n8392 ) | ( n8388 & n8393 ) | ( n8392 & n8393 ) ;
  assign n8395 = n8390 & ~n8394 ;
  assign n8396 = ~n8389 & n8392 ;
  assign n8397 = ~n8388 & n8396 ;
  assign n8398 = n8395 | n8397 ;
  assign n8399 = x79 & n3816 ;
  assign n8400 = x78 & n3811 ;
  assign n8401 = x77 & ~n3810 ;
  assign n8402 = n4067 & n8401 ;
  assign n8403 = n8400 | n8402 ;
  assign n8404 = n8399 | n8403 ;
  assign n8405 = n3819 | n8399 ;
  assign n8406 = n8403 | n8405 ;
  assign n8407 = ( n1332 & n8404 ) | ( n1332 & n8406 ) | ( n8404 & n8406 ) ;
  assign n8408 = x29 & n8406 ;
  assign n8409 = x29 & n8399 ;
  assign n8410 = ( x29 & n8403 ) | ( x29 & n8409 ) | ( n8403 & n8409 ) ;
  assign n8411 = ( n1332 & n8408 ) | ( n1332 & n8410 ) | ( n8408 & n8410 ) ;
  assign n8412 = x29 & ~n8410 ;
  assign n8413 = x29 & ~n8406 ;
  assign n8414 = ( ~n1332 & n8412 ) | ( ~n1332 & n8413 ) | ( n8412 & n8413 ) ;
  assign n8415 = ( n8407 & ~n8411 ) | ( n8407 & n8414 ) | ( ~n8411 & n8414 ) ;
  assign n8416 = n8043 | n8044 ;
  assign n8417 = ( n8043 & n8046 ) | ( n8043 & n8416 ) | ( n8046 & n8416 ) ;
  assign n8418 = ( ~n8398 & n8415 ) | ( ~n8398 & n8417 ) | ( n8415 & n8417 ) ;
  assign n8419 = x82 & n3085 ;
  assign n8420 = x81 & n3080 ;
  assign n8421 = x80 & ~n3079 ;
  assign n8422 = n3309 & n8421 ;
  assign n8423 = n8420 | n8422 ;
  assign n8424 = n8419 | n8423 ;
  assign n8425 = n3088 | n8419 ;
  assign n8426 = n8423 | n8425 ;
  assign n8427 = ( n1811 & n8424 ) | ( n1811 & n8426 ) | ( n8424 & n8426 ) ;
  assign n8428 = x26 & n8426 ;
  assign n8429 = x26 & n8419 ;
  assign n8430 = ( x26 & n8423 ) | ( x26 & n8429 ) | ( n8423 & n8429 ) ;
  assign n8431 = ( n1811 & n8428 ) | ( n1811 & n8430 ) | ( n8428 & n8430 ) ;
  assign n8432 = x26 & ~n8430 ;
  assign n8433 = x26 & ~n8426 ;
  assign n8434 = ( ~n1811 & n8432 ) | ( ~n1811 & n8433 ) | ( n8432 & n8433 ) ;
  assign n8435 = ( n8427 & ~n8431 ) | ( n8427 & n8434 ) | ( ~n8431 & n8434 ) ;
  assign n8436 = n8398 & n8435 ;
  assign n8437 = ~n8415 & n8435 ;
  assign n8438 = ( n8417 & n8436 ) | ( n8417 & n8437 ) | ( n8436 & n8437 ) ;
  assign n8439 = ~n8046 & n8435 ;
  assign n8440 = ~n8043 & n8435 ;
  assign n8441 = ( ~n8416 & n8439 ) | ( ~n8416 & n8440 ) | ( n8439 & n8440 ) ;
  assign n8442 = ( n8418 & n8438 ) | ( n8418 & n8441 ) | ( n8438 & n8441 ) ;
  assign n8443 = n8398 | n8435 ;
  assign n8444 = n8415 & ~n8435 ;
  assign n8445 = ( n8417 & n8443 ) | ( n8417 & ~n8444 ) | ( n8443 & ~n8444 ) ;
  assign n8446 = n8046 & ~n8435 ;
  assign n8447 = n8043 & ~n8435 ;
  assign n8448 = ( n8416 & n8446 ) | ( n8416 & n8447 ) | ( n8446 & n8447 ) ;
  assign n8449 = ( n8418 & n8445 ) | ( n8418 & ~n8448 ) | ( n8445 & ~n8448 ) ;
  assign n8450 = ~n8442 & n8449 ;
  assign n8451 = n8068 | n8069 ;
  assign n8452 = ( n8068 & n8071 ) | ( n8068 & n8451 ) | ( n8071 & n8451 ) ;
  assign n8453 = n8450 & n8452 ;
  assign n8454 = n8450 | n8452 ;
  assign n8455 = ~n8453 & n8454 ;
  assign n8456 = x85 & n2429 ;
  assign n8457 = x84 & n2424 ;
  assign n8458 = x83 & ~n2423 ;
  assign n8459 = n2631 & n8458 ;
  assign n8460 = n8457 | n8459 ;
  assign n8461 = n8456 | n8460 ;
  assign n8462 = n2432 | n8456 ;
  assign n8463 = n8460 | n8462 ;
  assign n8464 = ( n2381 & n8461 ) | ( n2381 & n8463 ) | ( n8461 & n8463 ) ;
  assign n8465 = x23 & n8463 ;
  assign n8466 = x23 & n8456 ;
  assign n8467 = ( x23 & n8460 ) | ( x23 & n8466 ) | ( n8460 & n8466 ) ;
  assign n8468 = ( n2381 & n8465 ) | ( n2381 & n8467 ) | ( n8465 & n8467 ) ;
  assign n8469 = x23 & ~n8467 ;
  assign n8470 = x23 & ~n8463 ;
  assign n8471 = ( ~n2381 & n8469 ) | ( ~n2381 & n8470 ) | ( n8469 & n8470 ) ;
  assign n8472 = ( n8464 & ~n8468 ) | ( n8464 & n8471 ) | ( ~n8468 & n8471 ) ;
  assign n8473 = n8455 & n8472 ;
  assign n8474 = n8455 & ~n8473 ;
  assign n8475 = ~n8455 & n8472 ;
  assign n8476 = n8474 | n8475 ;
  assign n8477 = n8092 | n8094 ;
  assign n8478 = n8093 | n8477 ;
  assign n8479 = ( n8092 & n8096 ) | ( n8092 & n8478 ) | ( n8096 & n8478 ) ;
  assign n8480 = n8476 | n8479 ;
  assign n8481 = n8476 & n8479 ;
  assign n8482 = n8480 & ~n8481 ;
  assign n8483 = x88 & n1859 ;
  assign n8484 = x87 & n1854 ;
  assign n8485 = x86 & ~n1853 ;
  assign n8486 = n2037 & n8485 ;
  assign n8487 = n8484 | n8486 ;
  assign n8488 = n8483 | n8487 ;
  assign n8489 = n1862 | n8483 ;
  assign n8490 = n8487 | n8489 ;
  assign n8491 = ( ~n3039 & n8488 ) | ( ~n3039 & n8490 ) | ( n8488 & n8490 ) ;
  assign n8492 = n8488 & n8490 ;
  assign n8493 = ( n3023 & n8491 ) | ( n3023 & n8492 ) | ( n8491 & n8492 ) ;
  assign n8494 = x20 & n8490 ;
  assign n8495 = x20 & n8483 ;
  assign n8496 = ( x20 & n8487 ) | ( x20 & n8495 ) | ( n8487 & n8495 ) ;
  assign n8497 = ( ~n3039 & n8494 ) | ( ~n3039 & n8496 ) | ( n8494 & n8496 ) ;
  assign n8498 = n8494 & n8496 ;
  assign n8499 = ( n3023 & n8497 ) | ( n3023 & n8498 ) | ( n8497 & n8498 ) ;
  assign n8500 = x20 & ~n8496 ;
  assign n8501 = x20 & ~n8490 ;
  assign n8502 = ( n3039 & n8500 ) | ( n3039 & n8501 ) | ( n8500 & n8501 ) ;
  assign n8503 = n8500 | n8501 ;
  assign n8504 = ( ~n3023 & n8502 ) | ( ~n3023 & n8503 ) | ( n8502 & n8503 ) ;
  assign n8505 = ( n8493 & ~n8499 ) | ( n8493 & n8504 ) | ( ~n8499 & n8504 ) ;
  assign n8506 = n8482 | n8505 ;
  assign n8507 = n8482 & n8505 ;
  assign n8508 = n8506 & ~n8507 ;
  assign n8509 = n8122 & n8508 ;
  assign n8510 = n8122 | n8508 ;
  assign n8511 = ~n8509 & n8510 ;
  assign n8512 = x91 & n1383 ;
  assign n8513 = x90 & n1378 ;
  assign n8514 = x89 & ~n1377 ;
  assign n8515 = n1542 & n8514 ;
  assign n8516 = n8513 | n8515 ;
  assign n8517 = n8512 | n8516 ;
  assign n8518 = n1386 | n8512 ;
  assign n8519 = n8516 | n8518 ;
  assign n8520 = ( n3768 & n8517 ) | ( n3768 & n8519 ) | ( n8517 & n8519 ) ;
  assign n8521 = x17 & n8519 ;
  assign n8522 = x17 & n8512 ;
  assign n8523 = ( x17 & n8516 ) | ( x17 & n8522 ) | ( n8516 & n8522 ) ;
  assign n8524 = ( n3768 & n8521 ) | ( n3768 & n8523 ) | ( n8521 & n8523 ) ;
  assign n8525 = x17 & ~n8523 ;
  assign n8526 = x17 & ~n8519 ;
  assign n8527 = ( ~n3768 & n8525 ) | ( ~n3768 & n8526 ) | ( n8525 & n8526 ) ;
  assign n8528 = ( n8520 & ~n8524 ) | ( n8520 & n8527 ) | ( ~n8524 & n8527 ) ;
  assign n8529 = n8511 & n8528 ;
  assign n8530 = n8511 & ~n8529 ;
  assign n8531 = ~n8511 & n8528 ;
  assign n8532 = n8530 | n8531 ;
  assign n8533 = n8297 & ~n8532 ;
  assign n8534 = ~n8297 & n8532 ;
  assign n8535 = n8533 | n8534 ;
  assign n8536 = x94 & n962 ;
  assign n8537 = x93 & n957 ;
  assign n8538 = x92 & ~n956 ;
  assign n8539 = n1105 & n8538 ;
  assign n8540 = n8537 | n8539 ;
  assign n8541 = n8536 | n8540 ;
  assign n8542 = n965 | n8536 ;
  assign n8543 = n8540 | n8542 ;
  assign n8544 = ( n4583 & n8541 ) | ( n4583 & n8543 ) | ( n8541 & n8543 ) ;
  assign n8545 = x14 & n8543 ;
  assign n8546 = x14 & n8536 ;
  assign n8547 = ( x14 & n8540 ) | ( x14 & n8546 ) | ( n8540 & n8546 ) ;
  assign n8548 = ( n4583 & n8545 ) | ( n4583 & n8547 ) | ( n8545 & n8547 ) ;
  assign n8549 = x14 & ~n8547 ;
  assign n8550 = x14 & ~n8543 ;
  assign n8551 = ( ~n4583 & n8549 ) | ( ~n4583 & n8550 ) | ( n8549 & n8550 ) ;
  assign n8552 = ( n8544 & ~n8548 ) | ( n8544 & n8551 ) | ( ~n8548 & n8551 ) ;
  assign n8553 = n8535 & n8552 ;
  assign n8554 = n8535 | n8552 ;
  assign n8555 = ~n8553 & n8554 ;
  assign n8556 = n7810 | n8171 ;
  assign n8557 = n8171 | n8172 ;
  assign n8558 = ( n8173 & n8556 ) | ( n8173 & n8557 ) | ( n8556 & n8557 ) ;
  assign n8559 = n8555 & n8558 ;
  assign n8560 = n8555 | n8558 ;
  assign n8561 = ~n8559 & n8560 ;
  assign n8562 = x97 & n636 ;
  assign n8563 = x96 & n631 ;
  assign n8564 = x95 & ~n630 ;
  assign n8565 = n764 & n8564 ;
  assign n8566 = n8563 | n8565 ;
  assign n8567 = n8562 | n8566 ;
  assign n8568 = n639 | n8562 ;
  assign n8569 = n8566 | n8568 ;
  assign n8570 = ( n5505 & n8567 ) | ( n5505 & n8569 ) | ( n8567 & n8569 ) ;
  assign n8571 = x11 & n8569 ;
  assign n8572 = x11 & n8562 ;
  assign n8573 = ( x11 & n8566 ) | ( x11 & n8572 ) | ( n8566 & n8572 ) ;
  assign n8574 = ( n5505 & n8571 ) | ( n5505 & n8573 ) | ( n8571 & n8573 ) ;
  assign n8575 = x11 & ~n8573 ;
  assign n8576 = x11 & ~n8569 ;
  assign n8577 = ( ~n5505 & n8575 ) | ( ~n5505 & n8576 ) | ( n8575 & n8576 ) ;
  assign n8578 = ( n8570 & ~n8574 ) | ( n8570 & n8577 ) | ( ~n8574 & n8577 ) ;
  assign n8579 = n8561 & n8578 ;
  assign n8580 = n8561 & ~n8579 ;
  assign n8581 = ~n8561 & n8578 ;
  assign n8582 = n8580 | n8581 ;
  assign n8583 = n8196 | n8200 ;
  assign n8584 = ~n8582 & n8583 ;
  assign n8585 = n8582 & ~n8583 ;
  assign n8586 = n8584 | n8585 ;
  assign n8587 = x100 & n389 ;
  assign n8588 = x99 & n384 ;
  assign n8589 = x98 & ~n383 ;
  assign n8590 = n463 & n8589 ;
  assign n8591 = n8588 | n8590 ;
  assign n8592 = n8587 | n8591 ;
  assign n8593 = n392 | n8587 ;
  assign n8594 = n8591 | n8593 ;
  assign n8595 = ( n6483 & n8592 ) | ( n6483 & n8594 ) | ( n8592 & n8594 ) ;
  assign n8596 = x8 & n8594 ;
  assign n8597 = x8 & n8587 ;
  assign n8598 = ( x8 & n8591 ) | ( x8 & n8597 ) | ( n8591 & n8597 ) ;
  assign n8599 = ( n6483 & n8596 ) | ( n6483 & n8598 ) | ( n8596 & n8598 ) ;
  assign n8600 = x8 & ~n8598 ;
  assign n8601 = x8 & ~n8594 ;
  assign n8602 = ( ~n6483 & n8600 ) | ( ~n6483 & n8601 ) | ( n8600 & n8601 ) ;
  assign n8603 = ( n8595 & ~n8599 ) | ( n8595 & n8602 ) | ( ~n8599 & n8602 ) ;
  assign n8604 = n8586 | n8603 ;
  assign n8605 = n8586 & n8603 ;
  assign n8606 = n8604 & ~n8605 ;
  assign n8607 = ( n8202 & n8219 ) | ( n8202 & n8225 ) | ( n8219 & n8225 ) ;
  assign n8608 = n8606 | n8607 ;
  assign n8609 = n8606 & n8607 ;
  assign n8610 = n8608 & ~n8609 ;
  assign n8611 = x103 & n212 ;
  assign n8612 = x102 & n207 ;
  assign n8613 = x101 & ~n206 ;
  assign n8614 = n267 & n8613 ;
  assign n8615 = n8612 | n8614 ;
  assign n8616 = n8611 | n8615 ;
  assign n8617 = n215 | n8611 ;
  assign n8618 = n8615 | n8617 ;
  assign n8619 = ( n7529 & n8616 ) | ( n7529 & n8618 ) | ( n8616 & n8618 ) ;
  assign n8620 = x5 & n8618 ;
  assign n8621 = x5 & n8611 ;
  assign n8622 = ( x5 & n8615 ) | ( x5 & n8621 ) | ( n8615 & n8621 ) ;
  assign n8623 = ( n7529 & n8620 ) | ( n7529 & n8622 ) | ( n8620 & n8622 ) ;
  assign n8624 = x5 & ~n8622 ;
  assign n8625 = x5 & ~n8618 ;
  assign n8626 = ( ~n7529 & n8624 ) | ( ~n7529 & n8625 ) | ( n8624 & n8625 ) ;
  assign n8627 = ( n8619 & ~n8623 ) | ( n8619 & n8626 ) | ( ~n8623 & n8626 ) ;
  assign n8628 = n8610 & n8627 ;
  assign n8629 = n8610 & ~n8628 ;
  assign n8630 = ~n8610 & n8627 ;
  assign n8631 = n8629 | n8630 ;
  assign n8632 = n8246 | n8249 ;
  assign n8633 = ( n8246 & n8248 ) | ( n8246 & n8632 ) | ( n8248 & n8632 ) ;
  assign n8634 = ~n8631 & n8633 ;
  assign n8635 = n8631 & ~n8633 ;
  assign n8636 = n8634 | n8635 ;
  assign n8637 = x105 | x106 ;
  assign n8638 = x105 & x106 ;
  assign n8639 = n8637 & ~n8638 ;
  assign n8640 = n8254 & n8639 ;
  assign n8641 = ( n8260 & n8639 ) | ( n8260 & n8640 ) | ( n8639 & n8640 ) ;
  assign n8642 = ( n8258 & n8639 ) | ( n8258 & n8640 ) | ( n8639 & n8640 ) ;
  assign n8643 = ( n7517 & n8641 ) | ( n7517 & n8642 ) | ( n8641 & n8642 ) ;
  assign n8644 = ( n7518 & n8641 ) | ( n7518 & n8642 ) | ( n8641 & n8642 ) ;
  assign n8645 = ( n6159 & n8643 ) | ( n6159 & n8644 ) | ( n8643 & n8644 ) ;
  assign n8646 = ( n6157 & n8643 ) | ( n6157 & n8644 ) | ( n8643 & n8644 ) ;
  assign n8647 = ( n5823 & n8645 ) | ( n5823 & n8646 ) | ( n8645 & n8646 ) ;
  assign n8648 = n8254 | n8639 ;
  assign n8649 = n8260 | n8648 ;
  assign n8650 = n8258 | n8648 ;
  assign n8651 = ( n7517 & n8649 ) | ( n7517 & n8650 ) | ( n8649 & n8650 ) ;
  assign n8652 = ( n7518 & n8649 ) | ( n7518 & n8650 ) | ( n8649 & n8650 ) ;
  assign n8653 = ( n6159 & n8651 ) | ( n6159 & n8652 ) | ( n8651 & n8652 ) ;
  assign n8654 = ( n6157 & n8651 ) | ( n6157 & n8652 ) | ( n8651 & n8652 ) ;
  assign n8655 = ( n5823 & n8653 ) | ( n5823 & n8654 ) | ( n8653 & n8654 ) ;
  assign n8656 = ~n8647 & n8655 ;
  assign n8657 = x105 & n133 ;
  assign n8658 = x104 & ~n162 ;
  assign n8659 = ( n137 & n8657 ) | ( n137 & n8658 ) | ( n8657 & n8658 ) ;
  assign n8660 = x0 & x106 ;
  assign n8661 = ( ~n137 & n8657 ) | ( ~n137 & n8660 ) | ( n8657 & n8660 ) ;
  assign n8662 = n8659 | n8661 ;
  assign n8663 = n141 | n8662 ;
  assign n8664 = ( n8656 & n8662 ) | ( n8656 & n8663 ) | ( n8662 & n8663 ) ;
  assign n8665 = x2 & n8662 ;
  assign n8666 = ( x2 & n523 ) | ( x2 & n8662 ) | ( n523 & n8662 ) ;
  assign n8667 = ( n8656 & n8665 ) | ( n8656 & n8666 ) | ( n8665 & n8666 ) ;
  assign n8668 = x2 & ~n8666 ;
  assign n8669 = x2 & ~n8662 ;
  assign n8670 = ( ~n8656 & n8668 ) | ( ~n8656 & n8669 ) | ( n8668 & n8669 ) ;
  assign n8671 = ( n8664 & ~n8667 ) | ( n8664 & n8670 ) | ( ~n8667 & n8670 ) ;
  assign n8672 = n8636 & n8671 ;
  assign n8673 = n8636 | n8671 ;
  assign n8674 = ~n8672 & n8673 ;
  assign n8675 = n8290 | n8291 ;
  assign n8676 = ( n8290 & n8293 ) | ( n8290 & n8675 ) | ( n8293 & n8675 ) ;
  assign n8677 = n8674 & n8676 ;
  assign n8678 = n8674 | n8676 ;
  assign n8679 = ~n8677 & n8678 ;
  assign n8680 = x104 & n212 ;
  assign n8681 = x103 & n207 ;
  assign n8682 = x102 & ~n206 ;
  assign n8683 = n267 & n8682 ;
  assign n8684 = n8681 | n8683 ;
  assign n8685 = n8680 | n8684 ;
  assign n8686 = n215 | n8680 ;
  assign n8687 = n8684 | n8686 ;
  assign n8688 = ( n7911 & n8685 ) | ( n7911 & n8687 ) | ( n8685 & n8687 ) ;
  assign n8689 = x5 & n8687 ;
  assign n8690 = x5 & n8680 ;
  assign n8691 = ( x5 & n8684 ) | ( x5 & n8690 ) | ( n8684 & n8690 ) ;
  assign n8692 = ( n7911 & n8689 ) | ( n7911 & n8691 ) | ( n8689 & n8691 ) ;
  assign n8693 = x5 & ~n8691 ;
  assign n8694 = x5 & ~n8687 ;
  assign n8695 = ( ~n7911 & n8693 ) | ( ~n7911 & n8694 ) | ( n8693 & n8694 ) ;
  assign n8696 = ( n8688 & ~n8692 ) | ( n8688 & n8695 ) | ( ~n8692 & n8695 ) ;
  assign n8697 = x95 & n962 ;
  assign n8698 = x94 & n957 ;
  assign n8699 = x93 & ~n956 ;
  assign n8700 = n1105 & n8699 ;
  assign n8701 = n8698 | n8700 ;
  assign n8702 = n8697 | n8701 ;
  assign n8703 = n965 | n8697 ;
  assign n8704 = n8701 | n8703 ;
  assign n8705 = ( n4897 & n8702 ) | ( n4897 & n8704 ) | ( n8702 & n8704 ) ;
  assign n8706 = x14 & n8704 ;
  assign n8707 = x14 & n8697 ;
  assign n8708 = ( x14 & n8701 ) | ( x14 & n8707 ) | ( n8701 & n8707 ) ;
  assign n8709 = ( n4897 & n8706 ) | ( n4897 & n8708 ) | ( n8706 & n8708 ) ;
  assign n8710 = x14 & ~n8708 ;
  assign n8711 = x14 & ~n8704 ;
  assign n8712 = ( ~n4897 & n8710 ) | ( ~n4897 & n8711 ) | ( n8710 & n8711 ) ;
  assign n8713 = ( n8705 & ~n8709 ) | ( n8705 & n8712 ) | ( ~n8709 & n8712 ) ;
  assign n8714 = n8363 | n8364 ;
  assign n8715 = ( n8363 & n8366 ) | ( n8363 & n8714 ) | ( n8366 & n8714 ) ;
  assign n8716 = ~x42 & x43 ;
  assign n8717 = x42 & ~x43 ;
  assign n8718 = n8716 | n8717 ;
  assign n8719 = ~n8300 & n8718 ;
  assign n8720 = x64 & n8719 ;
  assign n8721 = ~x43 & x44 ;
  assign n8722 = x43 & ~x44 ;
  assign n8723 = n8721 | n8722 ;
  assign n8724 = n8300 & ~n8723 ;
  assign n8725 = x65 & n8724 ;
  assign n8726 = n8720 | n8725 ;
  assign n8727 = n8300 & n8723 ;
  assign n8728 = x44 | n144 ;
  assign n8729 = ( x44 & n8727 ) | ( x44 & n8728 ) | ( n8727 & n8728 ) ;
  assign n8730 = ~x44 & n8729 ;
  assign n8731 = ( ~x44 & n8726 ) | ( ~x44 & n8730 ) | ( n8726 & n8730 ) ;
  assign n8732 = x44 & ~x64 ;
  assign n8733 = ( x44 & ~n8300 ) | ( x44 & n8732 ) | ( ~n8300 & n8732 ) ;
  assign n8734 = n8729 & n8733 ;
  assign n8735 = ( n8726 & n8733 ) | ( n8726 & n8734 ) | ( n8733 & n8734 ) ;
  assign n8736 = n144 & n8727 ;
  assign n8737 = n8733 & ~n8736 ;
  assign n8738 = ~n8726 & n8737 ;
  assign n8739 = ( n8731 & n8735 ) | ( n8731 & n8738 ) | ( n8735 & n8738 ) ;
  assign n8740 = n8729 | n8733 ;
  assign n8741 = n8726 | n8740 ;
  assign n8742 = ~n8733 & n8736 ;
  assign n8743 = ( n8726 & ~n8733 ) | ( n8726 & n8742 ) | ( ~n8733 & n8742 ) ;
  assign n8744 = ( n8731 & n8741 ) | ( n8731 & ~n8743 ) | ( n8741 & ~n8743 ) ;
  assign n8745 = ~n8739 & n8744 ;
  assign n8746 = n241 & n7569 ;
  assign n8747 = x68 & n7566 ;
  assign n8748 = x67 & n7561 ;
  assign n8749 = x66 & ~n7560 ;
  assign n8750 = n7953 & n8749 ;
  assign n8751 = n8748 | n8750 ;
  assign n8752 = n8747 | n8751 ;
  assign n8753 = n8746 | n8752 ;
  assign n8754 = x41 | n8747 ;
  assign n8755 = n8751 | n8754 ;
  assign n8756 = n8746 | n8755 ;
  assign n8757 = ~x41 & n8755 ;
  assign n8758 = ( ~x41 & n8746 ) | ( ~x41 & n8757 ) | ( n8746 & n8757 ) ;
  assign n8759 = ( ~n8753 & n8756 ) | ( ~n8753 & n8758 ) | ( n8756 & n8758 ) ;
  assign n8760 = n8745 | n8759 ;
  assign n8761 = n8745 & n8759 ;
  assign n8762 = n8760 & ~n8761 ;
  assign n8763 = ( n7967 & n8301 ) | ( n7967 & n8317 ) | ( n8301 & n8317 ) ;
  assign n8764 = n8762 | n8763 ;
  assign n8765 = n8762 & n8763 ;
  assign n8766 = n8764 & ~n8765 ;
  assign n8767 = x70 & n6531 ;
  assign n8768 = x69 & ~n6530 ;
  assign n8769 = n6871 & n8768 ;
  assign n8770 = n8767 | n8769 ;
  assign n8771 = x71 & n6536 ;
  assign n8772 = n6539 | n8771 ;
  assign n8773 = n8770 | n8772 ;
  assign n8774 = x38 & ~n8773 ;
  assign n8775 = x38 & ~n8771 ;
  assign n8776 = ~n8770 & n8775 ;
  assign n8777 = ( ~n438 & n8774 ) | ( ~n438 & n8776 ) | ( n8774 & n8776 ) ;
  assign n8778 = ~x38 & n8773 ;
  assign n8779 = ~x38 & n8771 ;
  assign n8780 = ( ~x38 & n8770 ) | ( ~x38 & n8779 ) | ( n8770 & n8779 ) ;
  assign n8781 = ( n438 & n8778 ) | ( n438 & n8780 ) | ( n8778 & n8780 ) ;
  assign n8782 = n8777 | n8781 ;
  assign n8783 = n8766 & n8782 ;
  assign n8784 = n8766 & ~n8783 ;
  assign n8785 = ~n8766 & n8782 ;
  assign n8786 = n8784 | n8785 ;
  assign n8787 = n8337 | n8342 ;
  assign n8788 = ( n8337 & n8340 ) | ( n8337 & n8787 ) | ( n8340 & n8787 ) ;
  assign n8789 = n8786 | n8788 ;
  assign n8790 = n8786 & n8788 ;
  assign n8791 = n8789 & ~n8790 ;
  assign n8792 = x74 & n5554 ;
  assign n8793 = x73 & n5549 ;
  assign n8794 = x72 & ~n5548 ;
  assign n8795 = n5893 & n8794 ;
  assign n8796 = n8793 | n8795 ;
  assign n8797 = n8792 | n8796 ;
  assign n8798 = n5557 | n8792 ;
  assign n8799 = n8796 | n8798 ;
  assign n8800 = ( n710 & n8797 ) | ( n710 & n8799 ) | ( n8797 & n8799 ) ;
  assign n8801 = x35 & n8799 ;
  assign n8802 = x35 & n8792 ;
  assign n8803 = ( x35 & n8796 ) | ( x35 & n8802 ) | ( n8796 & n8802 ) ;
  assign n8804 = ( n710 & n8801 ) | ( n710 & n8803 ) | ( n8801 & n8803 ) ;
  assign n8805 = x35 & ~n8803 ;
  assign n8806 = x35 & ~n8799 ;
  assign n8807 = ( ~n710 & n8805 ) | ( ~n710 & n8806 ) | ( n8805 & n8806 ) ;
  assign n8808 = ( n8800 & ~n8804 ) | ( n8800 & n8807 ) | ( ~n8804 & n8807 ) ;
  assign n8809 = n8791 & n8808 ;
  assign n8810 = n8791 | n8808 ;
  assign n8811 = ~n8809 & n8810 ;
  assign n8812 = n8715 & n8811 ;
  assign n8813 = n8715 & ~n8812 ;
  assign n8814 = x77 & n4631 ;
  assign n8815 = x76 & n4626 ;
  assign n8816 = x75 & ~n4625 ;
  assign n8817 = n4943 & n8816 ;
  assign n8818 = n8815 | n8817 ;
  assign n8819 = n8814 | n8818 ;
  assign n8820 = n4634 | n8814 ;
  assign n8821 = n8818 | n8820 ;
  assign n8822 = ( n1059 & n8819 ) | ( n1059 & n8821 ) | ( n8819 & n8821 ) ;
  assign n8823 = x32 & n8821 ;
  assign n8824 = x32 & n8814 ;
  assign n8825 = ( x32 & n8818 ) | ( x32 & n8824 ) | ( n8818 & n8824 ) ;
  assign n8826 = ( n1059 & n8823 ) | ( n1059 & n8825 ) | ( n8823 & n8825 ) ;
  assign n8827 = x32 & ~n8825 ;
  assign n8828 = x32 & ~n8821 ;
  assign n8829 = ( ~n1059 & n8827 ) | ( ~n1059 & n8828 ) | ( n8827 & n8828 ) ;
  assign n8830 = ( n8822 & ~n8826 ) | ( n8822 & n8829 ) | ( ~n8826 & n8829 ) ;
  assign n8831 = ~n8810 & n8811 ;
  assign n8832 = ( ~n8715 & n8811 ) | ( ~n8715 & n8831 ) | ( n8811 & n8831 ) ;
  assign n8833 = n8830 & n8832 ;
  assign n8834 = ( n8813 & n8830 ) | ( n8813 & n8833 ) | ( n8830 & n8833 ) ;
  assign n8835 = n8830 | n8832 ;
  assign n8836 = n8813 | n8835 ;
  assign n8837 = ~n8834 & n8836 ;
  assign n8838 = n8387 | n8392 ;
  assign n8839 = ( n8387 & n8390 ) | ( n8387 & n8838 ) | ( n8390 & n8838 ) ;
  assign n8840 = n8837 & n8839 ;
  assign n8841 = n8837 | n8839 ;
  assign n8842 = ~n8840 & n8841 ;
  assign n8843 = x80 & n3816 ;
  assign n8844 = x79 & n3811 ;
  assign n8845 = x78 & ~n3810 ;
  assign n8846 = n4067 & n8845 ;
  assign n8847 = n8844 | n8846 ;
  assign n8848 = n8843 | n8847 ;
  assign n8849 = n3819 | n8843 ;
  assign n8850 = n8847 | n8849 ;
  assign n8851 = ( n1499 & n8848 ) | ( n1499 & n8850 ) | ( n8848 & n8850 ) ;
  assign n8852 = x29 & n8850 ;
  assign n8853 = x29 & n8843 ;
  assign n8854 = ( x29 & n8847 ) | ( x29 & n8853 ) | ( n8847 & n8853 ) ;
  assign n8855 = ( n1499 & n8852 ) | ( n1499 & n8854 ) | ( n8852 & n8854 ) ;
  assign n8856 = x29 & ~n8854 ;
  assign n8857 = x29 & ~n8850 ;
  assign n8858 = ( ~n1499 & n8856 ) | ( ~n1499 & n8857 ) | ( n8856 & n8857 ) ;
  assign n8859 = ( n8851 & ~n8855 ) | ( n8851 & n8858 ) | ( ~n8855 & n8858 ) ;
  assign n8860 = n8842 & n8859 ;
  assign n8861 = n8842 & ~n8860 ;
  assign n8862 = ~n8842 & n8859 ;
  assign n8863 = n8861 | n8862 ;
  assign n8864 = ~n8397 & n8415 ;
  assign n8865 = ~n8395 & n8864 ;
  assign n8866 = n8417 & ~n8865 ;
  assign n8867 = n8397 & n8415 ;
  assign n8868 = ( n8395 & n8415 ) | ( n8395 & n8867 ) | ( n8415 & n8867 ) ;
  assign n8869 = n8398 & ~n8868 ;
  assign n8870 = ( n8417 & n8868 ) | ( n8417 & n8869 ) | ( n8868 & n8869 ) ;
  assign n8871 = n8417 | n8868 ;
  assign n8872 = ( ~n8866 & n8870 ) | ( ~n8866 & n8871 ) | ( n8870 & n8871 ) ;
  assign n8873 = n8863 | n8872 ;
  assign n8874 = n8863 & n8872 ;
  assign n8875 = n8873 & ~n8874 ;
  assign n8876 = x83 & n3085 ;
  assign n8877 = x82 & n3080 ;
  assign n8878 = x81 & ~n3079 ;
  assign n8879 = n3309 & n8878 ;
  assign n8880 = n8877 | n8879 ;
  assign n8881 = n8876 | n8880 ;
  assign n8882 = n3088 | n8876 ;
  assign n8883 = n8880 | n8882 ;
  assign n8884 = ( n2009 & n8881 ) | ( n2009 & n8883 ) | ( n8881 & n8883 ) ;
  assign n8885 = x26 & n8883 ;
  assign n8886 = x26 & n8876 ;
  assign n8887 = ( x26 & n8880 ) | ( x26 & n8886 ) | ( n8880 & n8886 ) ;
  assign n8888 = ( n2009 & n8885 ) | ( n2009 & n8887 ) | ( n8885 & n8887 ) ;
  assign n8889 = x26 & ~n8887 ;
  assign n8890 = x26 & ~n8883 ;
  assign n8891 = ( ~n2009 & n8889 ) | ( ~n2009 & n8890 ) | ( n8889 & n8890 ) ;
  assign n8892 = ( n8884 & ~n8888 ) | ( n8884 & n8891 ) | ( ~n8888 & n8891 ) ;
  assign n8893 = n8875 & n8892 ;
  assign n8894 = n8875 & ~n8893 ;
  assign n8895 = n8442 | n8450 ;
  assign n8896 = ( n8442 & n8452 ) | ( n8442 & n8895 ) | ( n8452 & n8895 ) ;
  assign n8897 = ~n8875 & n8892 ;
  assign n8898 = n8896 & n8897 ;
  assign n8899 = ( n8894 & n8896 ) | ( n8894 & n8898 ) | ( n8896 & n8898 ) ;
  assign n8900 = n8896 | n8897 ;
  assign n8901 = n8894 | n8900 ;
  assign n8902 = ~n8899 & n8901 ;
  assign n8903 = x86 & n2429 ;
  assign n8904 = x85 & n2424 ;
  assign n8905 = x84 & ~n2423 ;
  assign n8906 = n2631 & n8905 ;
  assign n8907 = n8904 | n8906 ;
  assign n8908 = n8903 | n8907 ;
  assign n8909 = n2432 | n8903 ;
  assign n8910 = n8907 | n8909 ;
  assign n8911 = ( n2606 & n8908 ) | ( n2606 & n8910 ) | ( n8908 & n8910 ) ;
  assign n8912 = x23 & n8910 ;
  assign n8913 = x23 & n8903 ;
  assign n8914 = ( x23 & n8907 ) | ( x23 & n8913 ) | ( n8907 & n8913 ) ;
  assign n8915 = ( n2606 & n8912 ) | ( n2606 & n8914 ) | ( n8912 & n8914 ) ;
  assign n8916 = x23 & ~n8914 ;
  assign n8917 = x23 & ~n8910 ;
  assign n8918 = ( ~n2606 & n8916 ) | ( ~n2606 & n8917 ) | ( n8916 & n8917 ) ;
  assign n8919 = ( n8911 & ~n8915 ) | ( n8911 & n8918 ) | ( ~n8915 & n8918 ) ;
  assign n8920 = n8902 & n8919 ;
  assign n8921 = n8902 & ~n8920 ;
  assign n8922 = ~n8902 & n8919 ;
  assign n8923 = n8921 | n8922 ;
  assign n8924 = n8473 | n8476 ;
  assign n8925 = ( n8473 & n8479 ) | ( n8473 & n8924 ) | ( n8479 & n8924 ) ;
  assign n8926 = n8923 | n8925 ;
  assign n8927 = n8923 & n8925 ;
  assign n8928 = n8926 & ~n8927 ;
  assign n8929 = x89 & n1859 ;
  assign n8930 = x88 & n1854 ;
  assign n8931 = x87 & ~n1853 ;
  assign n8932 = n2037 & n8931 ;
  assign n8933 = n8930 | n8932 ;
  assign n8934 = n8929 | n8933 ;
  assign n8935 = n1862 | n8929 ;
  assign n8936 = n8933 | n8935 ;
  assign n8937 = ( n3282 & n8934 ) | ( n3282 & n8936 ) | ( n8934 & n8936 ) ;
  assign n8938 = x20 & n8936 ;
  assign n8939 = x20 & n8929 ;
  assign n8940 = ( x20 & n8933 ) | ( x20 & n8939 ) | ( n8933 & n8939 ) ;
  assign n8941 = ( n3282 & n8938 ) | ( n3282 & n8940 ) | ( n8938 & n8940 ) ;
  assign n8942 = x20 & ~n8940 ;
  assign n8943 = x20 & ~n8936 ;
  assign n8944 = ( ~n3282 & n8942 ) | ( ~n3282 & n8943 ) | ( n8942 & n8943 ) ;
  assign n8945 = ( n8937 & ~n8941 ) | ( n8937 & n8944 ) | ( ~n8941 & n8944 ) ;
  assign n8946 = n8928 & n8945 ;
  assign n8947 = n8928 & ~n8946 ;
  assign n8948 = ~n8928 & n8945 ;
  assign n8949 = n8947 | n8948 ;
  assign n8950 = n8507 | n8508 ;
  assign n8951 = ( n8122 & n8507 ) | ( n8122 & n8950 ) | ( n8507 & n8950 ) ;
  assign n8952 = n8949 & n8951 ;
  assign n8953 = n8949 | n8951 ;
  assign n8954 = ~n8952 & n8953 ;
  assign n8955 = x92 & n1383 ;
  assign n8956 = x91 & n1378 ;
  assign n8957 = x90 & ~n1377 ;
  assign n8958 = n1542 & n8957 ;
  assign n8959 = n8956 | n8958 ;
  assign n8960 = n8955 | n8959 ;
  assign n8961 = n1386 | n8955 ;
  assign n8962 = n8959 | n8961 ;
  assign n8963 = ( n4040 & n8960 ) | ( n4040 & n8962 ) | ( n8960 & n8962 ) ;
  assign n8964 = x17 & n8962 ;
  assign n8965 = x17 & n8955 ;
  assign n8966 = ( x17 & n8959 ) | ( x17 & n8965 ) | ( n8959 & n8965 ) ;
  assign n8967 = ( n4040 & n8964 ) | ( n4040 & n8966 ) | ( n8964 & n8966 ) ;
  assign n8968 = x17 & ~n8966 ;
  assign n8969 = x17 & ~n8962 ;
  assign n8970 = ( ~n4040 & n8968 ) | ( ~n4040 & n8969 ) | ( n8968 & n8969 ) ;
  assign n8971 = ( n8963 & ~n8967 ) | ( n8963 & n8970 ) | ( ~n8967 & n8970 ) ;
  assign n8972 = n8954 & n8971 ;
  assign n8973 = n8954 & ~n8972 ;
  assign n8974 = ~n8954 & n8971 ;
  assign n8975 = ( n8143 & n8511 ) | ( n8143 & n8528 ) | ( n8511 & n8528 ) ;
  assign n8976 = n8511 | n8528 ;
  assign n8977 = ( n8150 & n8975 ) | ( n8150 & n8976 ) | ( n8975 & n8976 ) ;
  assign n8978 = ~n8974 & n8977 ;
  assign n8979 = ~n8973 & n8978 ;
  assign n8980 = n8713 & n8979 ;
  assign n8981 = n8974 & ~n8977 ;
  assign n8982 = ( n8973 & ~n8977 ) | ( n8973 & n8981 ) | ( ~n8977 & n8981 ) ;
  assign n8983 = ( n8713 & n8980 ) | ( n8713 & n8982 ) | ( n8980 & n8982 ) ;
  assign n8984 = n8713 | n8979 ;
  assign n8985 = n8982 | n8984 ;
  assign n8986 = ~n8983 & n8985 ;
  assign n8987 = n8553 | n8559 ;
  assign n8988 = n8986 & n8987 ;
  assign n8989 = n8986 | n8987 ;
  assign n8990 = ~n8988 & n8989 ;
  assign n8991 = x98 & n636 ;
  assign n8992 = x97 & n631 ;
  assign n8993 = x96 & ~n630 ;
  assign n8994 = n764 & n8993 ;
  assign n8995 = n8992 | n8994 ;
  assign n8996 = n8991 | n8995 ;
  assign n8997 = n639 | n8991 ;
  assign n8998 = n8995 | n8997 ;
  assign n8999 = ( ~n5850 & n8996 ) | ( ~n5850 & n8998 ) | ( n8996 & n8998 ) ;
  assign n9000 = n8996 & n8998 ;
  assign n9001 = ( n5834 & n8999 ) | ( n5834 & n9000 ) | ( n8999 & n9000 ) ;
  assign n9002 = x11 & n8998 ;
  assign n9003 = x11 & n8991 ;
  assign n9004 = ( x11 & n8995 ) | ( x11 & n9003 ) | ( n8995 & n9003 ) ;
  assign n9005 = ( ~n5850 & n9002 ) | ( ~n5850 & n9004 ) | ( n9002 & n9004 ) ;
  assign n9006 = n9002 & n9004 ;
  assign n9007 = ( n5834 & n9005 ) | ( n5834 & n9006 ) | ( n9005 & n9006 ) ;
  assign n9008 = x11 & ~n9004 ;
  assign n9009 = x11 & ~n8998 ;
  assign n9010 = ( n5850 & n9008 ) | ( n5850 & n9009 ) | ( n9008 & n9009 ) ;
  assign n9011 = n9008 | n9009 ;
  assign n9012 = ( ~n5834 & n9010 ) | ( ~n5834 & n9011 ) | ( n9010 & n9011 ) ;
  assign n9013 = ( n9001 & ~n9007 ) | ( n9001 & n9012 ) | ( ~n9007 & n9012 ) ;
  assign n9014 = n8990 & n9013 ;
  assign n9015 = n8990 & ~n9014 ;
  assign n9016 = ( n8196 & n8561 ) | ( n8196 & n8578 ) | ( n8561 & n8578 ) ;
  assign n9017 = n8561 | n8578 ;
  assign n9018 = ( n8200 & n9016 ) | ( n8200 & n9017 ) | ( n9016 & n9017 ) ;
  assign n9019 = ~n8990 & n9013 ;
  assign n9020 = n9018 & n9019 ;
  assign n9021 = ( n9015 & n9018 ) | ( n9015 & n9020 ) | ( n9018 & n9020 ) ;
  assign n9022 = n9018 | n9019 ;
  assign n9023 = n9015 | n9022 ;
  assign n9024 = ~n9021 & n9023 ;
  assign n9025 = x101 & n389 ;
  assign n9026 = x100 & n384 ;
  assign n9027 = x99 & ~n383 ;
  assign n9028 = n463 & n9027 ;
  assign n9029 = n9026 | n9028 ;
  assign n9030 = n9025 | n9029 ;
  assign n9031 = n392 | n9025 ;
  assign n9032 = n9029 | n9031 ;
  assign n9033 = ( n6844 & n9030 ) | ( n6844 & n9032 ) | ( n9030 & n9032 ) ;
  assign n9034 = x8 & n9032 ;
  assign n9035 = x8 & n9025 ;
  assign n9036 = ( x8 & n9029 ) | ( x8 & n9035 ) | ( n9029 & n9035 ) ;
  assign n9037 = ( n6844 & n9034 ) | ( n6844 & n9036 ) | ( n9034 & n9036 ) ;
  assign n9038 = x8 & ~n9036 ;
  assign n9039 = x8 & ~n9032 ;
  assign n9040 = ( ~n6844 & n9038 ) | ( ~n6844 & n9039 ) | ( n9038 & n9039 ) ;
  assign n9041 = ( n9033 & ~n9037 ) | ( n9033 & n9040 ) | ( ~n9037 & n9040 ) ;
  assign n9042 = n9024 | n9041 ;
  assign n9043 = n9024 & n9041 ;
  assign n9044 = n9042 & ~n9043 ;
  assign n9045 = n8605 | n8607 ;
  assign n9046 = ( n8605 & n8606 ) | ( n8605 & n9045 ) | ( n8606 & n9045 ) ;
  assign n9047 = n9044 & n9046 ;
  assign n9048 = n9044 & ~n9047 ;
  assign n9049 = ~n9044 & n9046 ;
  assign n9050 = n8696 & n9049 ;
  assign n9051 = ( n8696 & n9048 ) | ( n8696 & n9050 ) | ( n9048 & n9050 ) ;
  assign n9052 = n8696 | n9049 ;
  assign n9053 = n9048 | n9052 ;
  assign n9054 = ~n9051 & n9053 ;
  assign n9055 = n8628 | n8633 ;
  assign n9056 = ( n8628 & n8631 ) | ( n8628 & n9055 ) | ( n8631 & n9055 ) ;
  assign n9057 = n9054 & n9056 ;
  assign n9058 = n9054 | n9056 ;
  assign n9059 = ~n9057 & n9058 ;
  assign n9060 = x106 | x107 ;
  assign n9061 = x106 & x107 ;
  assign n9062 = n9060 & ~n9061 ;
  assign n9063 = n8254 | n8638 ;
  assign n9064 = ( n8638 & n8639 ) | ( n8638 & n9063 ) | ( n8639 & n9063 ) ;
  assign n9065 = n9062 & n9064 ;
  assign n9066 = n8638 | n8639 ;
  assign n9067 = n9062 & n9066 ;
  assign n9068 = ( n8260 & n9065 ) | ( n8260 & n9067 ) | ( n9065 & n9067 ) ;
  assign n9069 = ( n8258 & n9065 ) | ( n8258 & n9067 ) | ( n9065 & n9067 ) ;
  assign n9070 = ( n7517 & n9068 ) | ( n7517 & n9069 ) | ( n9068 & n9069 ) ;
  assign n9071 = ( n7518 & n9068 ) | ( n7518 & n9069 ) | ( n9068 & n9069 ) ;
  assign n9072 = ( n6159 & n9070 ) | ( n6159 & n9071 ) | ( n9070 & n9071 ) ;
  assign n9073 = ( n6157 & n9070 ) | ( n6157 & n9071 ) | ( n9070 & n9071 ) ;
  assign n9074 = ( n5823 & n9072 ) | ( n5823 & n9073 ) | ( n9072 & n9073 ) ;
  assign n9075 = ( n8260 & n9064 ) | ( n8260 & n9066 ) | ( n9064 & n9066 ) ;
  assign n9076 = ( n8258 & n9064 ) | ( n8258 & n9066 ) | ( n9064 & n9066 ) ;
  assign n9077 = ( n7518 & n9075 ) | ( n7518 & n9076 ) | ( n9075 & n9076 ) ;
  assign n9078 = n9062 | n9077 ;
  assign n9079 = ( n7517 & n9075 ) | ( n7517 & n9076 ) | ( n9075 & n9076 ) ;
  assign n9080 = n9062 | n9079 ;
  assign n9081 = ( n6159 & n9078 ) | ( n6159 & n9080 ) | ( n9078 & n9080 ) ;
  assign n9082 = ( n6157 & n9078 ) | ( n6157 & n9080 ) | ( n9078 & n9080 ) ;
  assign n9083 = ( n5823 & n9081 ) | ( n5823 & n9082 ) | ( n9081 & n9082 ) ;
  assign n9084 = ~n9074 & n9083 ;
  assign n9085 = x106 & n133 ;
  assign n9086 = x105 & ~n162 ;
  assign n9087 = ( n137 & n9085 ) | ( n137 & n9086 ) | ( n9085 & n9086 ) ;
  assign n9088 = x0 & x107 ;
  assign n9089 = ( ~n137 & n9085 ) | ( ~n137 & n9088 ) | ( n9085 & n9088 ) ;
  assign n9090 = n9087 | n9089 ;
  assign n9091 = n141 | n9090 ;
  assign n9092 = ( n9084 & n9090 ) | ( n9084 & n9091 ) | ( n9090 & n9091 ) ;
  assign n9093 = x2 & n9090 ;
  assign n9094 = ( x2 & n523 ) | ( x2 & n9090 ) | ( n523 & n9090 ) ;
  assign n9095 = ( n9084 & n9093 ) | ( n9084 & n9094 ) | ( n9093 & n9094 ) ;
  assign n9096 = x2 & ~n9094 ;
  assign n9097 = x2 & ~n9090 ;
  assign n9098 = ( ~n9084 & n9096 ) | ( ~n9084 & n9097 ) | ( n9096 & n9097 ) ;
  assign n9099 = ( n9092 & ~n9095 ) | ( n9092 & n9098 ) | ( ~n9095 & n9098 ) ;
  assign n9100 = n9059 & n9099 ;
  assign n9101 = n9059 & ~n9100 ;
  assign n9102 = ~n9059 & n9099 ;
  assign n9103 = n9101 | n9102 ;
  assign n9104 = n8672 | n8677 ;
  assign n9105 = n9103 & n9104 ;
  assign n9106 = n9103 | n9104 ;
  assign n9107 = ~n9105 & n9106 ;
  assign n9108 = n9100 | n9105 ;
  assign n9109 = n9051 | n9054 ;
  assign n9110 = ( n9051 & n9056 ) | ( n9051 & n9109 ) | ( n9056 & n9109 ) ;
  assign n9111 = n9043 | n9047 ;
  assign n9112 = x90 & n1859 ;
  assign n9113 = x89 & n1854 ;
  assign n9114 = x88 & ~n1853 ;
  assign n9115 = n2037 & n9114 ;
  assign n9116 = n9113 | n9115 ;
  assign n9117 = n9112 | n9116 ;
  assign n9118 = n1862 | n9112 ;
  assign n9119 = n9116 | n9118 ;
  assign n9120 = ( n3519 & n9117 ) | ( n3519 & n9119 ) | ( n9117 & n9119 ) ;
  assign n9121 = x20 & n9119 ;
  assign n9122 = x20 & n9112 ;
  assign n9123 = ( x20 & n9116 ) | ( x20 & n9122 ) | ( n9116 & n9122 ) ;
  assign n9124 = ( n3519 & n9121 ) | ( n3519 & n9123 ) | ( n9121 & n9123 ) ;
  assign n9125 = x20 & ~n9123 ;
  assign n9126 = x20 & ~n9119 ;
  assign n9127 = ( ~n3519 & n9125 ) | ( ~n3519 & n9126 ) | ( n9125 & n9126 ) ;
  assign n9128 = ( n9120 & ~n9124 ) | ( n9120 & n9127 ) | ( ~n9124 & n9127 ) ;
  assign n9129 = x75 & n5554 ;
  assign n9130 = x74 & n5549 ;
  assign n9131 = x73 & ~n5548 ;
  assign n9132 = n5893 & n9131 ;
  assign n9133 = n9130 | n9132 ;
  assign n9134 = n9129 | n9133 ;
  assign n9135 = n5557 | n9129 ;
  assign n9136 = n9133 | n9135 ;
  assign n9137 = ( n746 & n9134 ) | ( n746 & n9136 ) | ( n9134 & n9136 ) ;
  assign n9138 = x35 & n9136 ;
  assign n9139 = x35 & n9129 ;
  assign n9140 = ( x35 & n9133 ) | ( x35 & n9139 ) | ( n9133 & n9139 ) ;
  assign n9141 = ( n746 & n9138 ) | ( n746 & n9140 ) | ( n9138 & n9140 ) ;
  assign n9142 = x35 & ~n9140 ;
  assign n9143 = x35 & ~n9136 ;
  assign n9144 = ( ~n746 & n9142 ) | ( ~n746 & n9143 ) | ( n9142 & n9143 ) ;
  assign n9145 = ( n9137 & ~n9141 ) | ( n9137 & n9144 ) | ( ~n9141 & n9144 ) ;
  assign n9146 = n8783 | n8790 ;
  assign n9147 = x66 & n8724 ;
  assign n9148 = x65 & n8719 ;
  assign n9149 = ~n8300 & n8723 ;
  assign n9150 = x64 & ~n8718 ;
  assign n9151 = n9149 & n9150 ;
  assign n9152 = n9148 | n9151 ;
  assign n9153 = n9147 | n9152 ;
  assign n9154 = n159 & n8727 ;
  assign n9155 = n9153 | n9154 ;
  assign n9156 = x44 | n8727 ;
  assign n9157 = ( x44 & n159 ) | ( x44 & n9156 ) | ( n159 & n9156 ) ;
  assign n9158 = n9153 | n9157 ;
  assign n9159 = ~x44 & n9157 ;
  assign n9160 = ( ~x44 & n9153 ) | ( ~x44 & n9159 ) | ( n9153 & n9159 ) ;
  assign n9161 = ( ~n9155 & n9158 ) | ( ~n9155 & n9160 ) | ( n9158 & n9160 ) ;
  assign n9162 = n8739 | n9161 ;
  assign n9163 = n8739 & n9161 ;
  assign n9164 = n9162 & ~n9163 ;
  assign n9165 = n293 & n7569 ;
  assign n9166 = x69 & n7566 ;
  assign n9167 = x68 & n7561 ;
  assign n9168 = x67 & ~n7560 ;
  assign n9169 = n7953 & n9168 ;
  assign n9170 = n9167 | n9169 ;
  assign n9171 = n9166 | n9170 ;
  assign n9172 = n9165 | n9171 ;
  assign n9173 = x41 | n9166 ;
  assign n9174 = n9170 | n9173 ;
  assign n9175 = n9165 | n9174 ;
  assign n9176 = ~x41 & n9174 ;
  assign n9177 = ( ~x41 & n9165 ) | ( ~x41 & n9176 ) | ( n9165 & n9176 ) ;
  assign n9178 = ( ~n9172 & n9175 ) | ( ~n9172 & n9177 ) | ( n9175 & n9177 ) ;
  assign n9179 = n9164 & n9178 ;
  assign n9180 = n9164 & ~n9179 ;
  assign n9181 = ~n9164 & n9178 ;
  assign n9182 = n9180 | n9181 ;
  assign n9183 = n8761 | n8763 ;
  assign n9184 = ( n8761 & n8762 ) | ( n8761 & n9183 ) | ( n8762 & n9183 ) ;
  assign n9185 = n9182 & n9184 ;
  assign n9186 = n9182 | n9184 ;
  assign n9187 = ~n9185 & n9186 ;
  assign n9188 = x72 & n6536 ;
  assign n9189 = x71 & n6531 ;
  assign n9190 = x70 & ~n6530 ;
  assign n9191 = n6871 & n9190 ;
  assign n9192 = n9189 | n9191 ;
  assign n9193 = n9188 | n9192 ;
  assign n9194 = ( n513 & n6539 ) | ( n513 & n9193 ) | ( n6539 & n9193 ) ;
  assign n9195 = ( x38 & n6539 ) | ( x38 & ~n9188 ) | ( n6539 & ~n9188 ) ;
  assign n9196 = x38 & n6539 ;
  assign n9197 = ( ~n9192 & n9195 ) | ( ~n9192 & n9196 ) | ( n9195 & n9196 ) ;
  assign n9198 = ( x38 & n513 ) | ( x38 & n9197 ) | ( n513 & n9197 ) ;
  assign n9199 = ~n9194 & n9198 ;
  assign n9200 = n9193 | n9197 ;
  assign n9201 = x38 | n9193 ;
  assign n9202 = ( n513 & n9200 ) | ( n513 & n9201 ) | ( n9200 & n9201 ) ;
  assign n9203 = ( ~x38 & n9199 ) | ( ~x38 & n9202 ) | ( n9199 & n9202 ) ;
  assign n9204 = n9187 & n9203 ;
  assign n9205 = n9187 & ~n9204 ;
  assign n9206 = ~n9187 & n9203 ;
  assign n9207 = n9205 | n9206 ;
  assign n9208 = ~n9146 & n9207 ;
  assign n9209 = n9145 & n9208 ;
  assign n9210 = n9146 & ~n9207 ;
  assign n9211 = ( n9145 & n9209 ) | ( n9145 & n9210 ) | ( n9209 & n9210 ) ;
  assign n9212 = n9145 | n9208 ;
  assign n9213 = n9210 | n9212 ;
  assign n9214 = ~n9211 & n9213 ;
  assign n9215 = n8809 | n8810 ;
  assign n9216 = ( n8715 & n8809 ) | ( n8715 & n9215 ) | ( n8809 & n9215 ) ;
  assign n9217 = n9214 & n9216 ;
  assign n9218 = n9214 | n9216 ;
  assign n9219 = ~n9217 & n9218 ;
  assign n9220 = x78 & n4631 ;
  assign n9221 = x77 & n4626 ;
  assign n9222 = x76 & ~n4625 ;
  assign n9223 = n4943 & n9222 ;
  assign n9224 = n9221 | n9223 ;
  assign n9225 = n9220 | n9224 ;
  assign n9226 = n4634 | n9220 ;
  assign n9227 = n9224 | n9226 ;
  assign n9228 = ( n1192 & n9225 ) | ( n1192 & n9227 ) | ( n9225 & n9227 ) ;
  assign n9229 = x32 & n9227 ;
  assign n9230 = x32 & n9220 ;
  assign n9231 = ( x32 & n9224 ) | ( x32 & n9230 ) | ( n9224 & n9230 ) ;
  assign n9232 = ( n1192 & n9229 ) | ( n1192 & n9231 ) | ( n9229 & n9231 ) ;
  assign n9233 = x32 & ~n9231 ;
  assign n9234 = x32 & ~n9227 ;
  assign n9235 = ( ~n1192 & n9233 ) | ( ~n1192 & n9234 ) | ( n9233 & n9234 ) ;
  assign n9236 = ( n9228 & ~n9232 ) | ( n9228 & n9235 ) | ( ~n9232 & n9235 ) ;
  assign n9237 = n9219 | n9236 ;
  assign n9238 = n9219 & n9236 ;
  assign n9239 = n9237 & ~n9238 ;
  assign n9240 = n8834 | n8837 ;
  assign n9241 = ( n8834 & n8839 ) | ( n8834 & n9240 ) | ( n8839 & n9240 ) ;
  assign n9242 = n9239 & n9241 ;
  assign n9243 = n9239 | n9241 ;
  assign n9244 = ~n9242 & n9243 ;
  assign n9245 = x81 & n3816 ;
  assign n9246 = x80 & n3811 ;
  assign n9247 = x79 & ~n3810 ;
  assign n9248 = n4067 & n9247 ;
  assign n9249 = n9246 | n9248 ;
  assign n9250 = n9245 | n9249 ;
  assign n9251 = n3819 | n9245 ;
  assign n9252 = n9249 | n9251 ;
  assign n9253 = ( n1651 & n9250 ) | ( n1651 & n9252 ) | ( n9250 & n9252 ) ;
  assign n9254 = x29 & n9252 ;
  assign n9255 = x29 & n9245 ;
  assign n9256 = ( x29 & n9249 ) | ( x29 & n9255 ) | ( n9249 & n9255 ) ;
  assign n9257 = ( n1651 & n9254 ) | ( n1651 & n9256 ) | ( n9254 & n9256 ) ;
  assign n9258 = x29 & ~n9256 ;
  assign n9259 = x29 & ~n9252 ;
  assign n9260 = ( ~n1651 & n9258 ) | ( ~n1651 & n9259 ) | ( n9258 & n9259 ) ;
  assign n9261 = ( n9253 & ~n9257 ) | ( n9253 & n9260 ) | ( ~n9257 & n9260 ) ;
  assign n9262 = n9244 | n9261 ;
  assign n9263 = n9244 & n9261 ;
  assign n9264 = n9262 & ~n9263 ;
  assign n9265 = n8860 & n9264 ;
  assign n9266 = ( n8874 & n9264 ) | ( n8874 & n9265 ) | ( n9264 & n9265 ) ;
  assign n9267 = n8860 | n9264 ;
  assign n9268 = n8874 | n9267 ;
  assign n9269 = ~n9266 & n9268 ;
  assign n9270 = x84 & n3085 ;
  assign n9271 = x83 & n3080 ;
  assign n9272 = x82 & ~n3079 ;
  assign n9273 = n3309 & n9272 ;
  assign n9274 = n9271 | n9273 ;
  assign n9275 = n9270 | n9274 ;
  assign n9276 = n3088 | n9270 ;
  assign n9277 = n9274 | n9276 ;
  assign n9278 = ( n2194 & n9275 ) | ( n2194 & n9277 ) | ( n9275 & n9277 ) ;
  assign n9279 = x26 & n9277 ;
  assign n9280 = x26 & n9270 ;
  assign n9281 = ( x26 & n9274 ) | ( x26 & n9280 ) | ( n9274 & n9280 ) ;
  assign n9282 = ( n2194 & n9279 ) | ( n2194 & n9281 ) | ( n9279 & n9281 ) ;
  assign n9283 = x26 & ~n9281 ;
  assign n9284 = x26 & ~n9277 ;
  assign n9285 = ( ~n2194 & n9283 ) | ( ~n2194 & n9284 ) | ( n9283 & n9284 ) ;
  assign n9286 = ( n9278 & ~n9282 ) | ( n9278 & n9285 ) | ( ~n9282 & n9285 ) ;
  assign n9287 = n9269 & n9286 ;
  assign n9288 = n9269 & ~n9287 ;
  assign n9289 = ~n9269 & n9286 ;
  assign n9290 = n9288 | n9289 ;
  assign n9291 = n8893 | n8899 ;
  assign n9292 = n9290 | n9291 ;
  assign n9293 = n9290 & n9291 ;
  assign n9294 = n9292 & ~n9293 ;
  assign n9295 = x87 & n2429 ;
  assign n9296 = x86 & n2424 ;
  assign n9297 = x85 & ~n2423 ;
  assign n9298 = n2631 & n9297 ;
  assign n9299 = n9296 | n9298 ;
  assign n9300 = n9295 | n9299 ;
  assign n9301 = n2432 | n9295 ;
  assign n9302 = n9299 | n9301 ;
  assign n9303 = ( n2816 & n9300 ) | ( n2816 & n9302 ) | ( n9300 & n9302 ) ;
  assign n9304 = x23 & n9302 ;
  assign n9305 = x23 & n9295 ;
  assign n9306 = ( x23 & n9299 ) | ( x23 & n9305 ) | ( n9299 & n9305 ) ;
  assign n9307 = ( n2816 & n9304 ) | ( n2816 & n9306 ) | ( n9304 & n9306 ) ;
  assign n9308 = x23 & ~n9306 ;
  assign n9309 = x23 & ~n9302 ;
  assign n9310 = ( ~n2816 & n9308 ) | ( ~n2816 & n9309 ) | ( n9308 & n9309 ) ;
  assign n9311 = ( n9303 & ~n9307 ) | ( n9303 & n9310 ) | ( ~n9307 & n9310 ) ;
  assign n9312 = n9294 | n9311 ;
  assign n9313 = n9294 & n9311 ;
  assign n9314 = n9312 & ~n9313 ;
  assign n9315 = n8920 | n8925 ;
  assign n9316 = ( n8920 & n8923 ) | ( n8920 & n9315 ) | ( n8923 & n9315 ) ;
  assign n9317 = ~n9314 & n9316 ;
  assign n9318 = n9128 & n9317 ;
  assign n9319 = n9313 | n9314 ;
  assign n9320 = n9312 & ~n9316 ;
  assign n9321 = ( n9314 & ~n9319 ) | ( n9314 & n9320 ) | ( ~n9319 & n9320 ) ;
  assign n9322 = ( n9128 & n9318 ) | ( n9128 & n9321 ) | ( n9318 & n9321 ) ;
  assign n9323 = n9128 | n9317 ;
  assign n9324 = n9321 | n9323 ;
  assign n9325 = ~n9322 & n9324 ;
  assign n9326 = n8946 | n8951 ;
  assign n9327 = ( n8946 & n8949 ) | ( n8946 & n9326 ) | ( n8949 & n9326 ) ;
  assign n9328 = n9325 & n9327 ;
  assign n9329 = n9325 | n9327 ;
  assign n9330 = ~n9328 & n9329 ;
  assign n9331 = x93 & n1383 ;
  assign n9332 = x92 & n1378 ;
  assign n9333 = x91 & ~n1377 ;
  assign n9334 = n1542 & n9333 ;
  assign n9335 = n9332 | n9334 ;
  assign n9336 = n9331 | n9335 ;
  assign n9337 = n1386 | n9331 ;
  assign n9338 = n9335 | n9337 ;
  assign n9339 = ( n4305 & n9336 ) | ( n4305 & n9338 ) | ( n9336 & n9338 ) ;
  assign n9340 = x17 & n9338 ;
  assign n9341 = x17 & n9331 ;
  assign n9342 = ( x17 & n9335 ) | ( x17 & n9341 ) | ( n9335 & n9341 ) ;
  assign n9343 = ( n4305 & n9340 ) | ( n4305 & n9342 ) | ( n9340 & n9342 ) ;
  assign n9344 = x17 & ~n9342 ;
  assign n9345 = x17 & ~n9338 ;
  assign n9346 = ( ~n4305 & n9344 ) | ( ~n4305 & n9345 ) | ( n9344 & n9345 ) ;
  assign n9347 = ( n9339 & ~n9343 ) | ( n9339 & n9346 ) | ( ~n9343 & n9346 ) ;
  assign n9348 = n9330 | n9347 ;
  assign n9349 = n9330 & n9347 ;
  assign n9350 = n9348 & ~n9349 ;
  assign n9351 = n8974 & n8977 ;
  assign n9352 = ( n8973 & n8977 ) | ( n8973 & n9351 ) | ( n8977 & n9351 ) ;
  assign n9353 = n8972 | n9352 ;
  assign n9354 = n9350 & n9353 ;
  assign n9355 = n9350 | n9353 ;
  assign n9356 = ~n9354 & n9355 ;
  assign n9357 = x96 & n962 ;
  assign n9358 = x95 & n957 ;
  assign n9359 = x94 & ~n956 ;
  assign n9360 = n1105 & n9359 ;
  assign n9361 = n9358 | n9360 ;
  assign n9362 = n9357 | n9361 ;
  assign n9363 = n965 | n9357 ;
  assign n9364 = n9361 | n9363 ;
  assign n9365 = ( n5202 & n9362 ) | ( n5202 & n9364 ) | ( n9362 & n9364 ) ;
  assign n9366 = x14 & n9364 ;
  assign n9367 = x14 & n9357 ;
  assign n9368 = ( x14 & n9361 ) | ( x14 & n9367 ) | ( n9361 & n9367 ) ;
  assign n9369 = ( n5202 & n9366 ) | ( n5202 & n9368 ) | ( n9366 & n9368 ) ;
  assign n9370 = x14 & ~n9368 ;
  assign n9371 = x14 & ~n9364 ;
  assign n9372 = ( ~n5202 & n9370 ) | ( ~n5202 & n9371 ) | ( n9370 & n9371 ) ;
  assign n9373 = ( n9365 & ~n9369 ) | ( n9365 & n9372 ) | ( ~n9369 & n9372 ) ;
  assign n9374 = n9356 | n9373 ;
  assign n9375 = n9356 & n9373 ;
  assign n9376 = n9374 & ~n9375 ;
  assign n9377 = n8983 | n8986 ;
  assign n9378 = ( n8983 & n8987 ) | ( n8983 & n9377 ) | ( n8987 & n9377 ) ;
  assign n9379 = n9376 & n9378 ;
  assign n9380 = n9376 | n9378 ;
  assign n9381 = ~n9379 & n9380 ;
  assign n9382 = x99 & n636 ;
  assign n9383 = x98 & n631 ;
  assign n9384 = x97 & ~n630 ;
  assign n9385 = n764 & n9384 ;
  assign n9386 = n9383 | n9385 ;
  assign n9387 = n9382 | n9386 ;
  assign n9388 = n639 | n9382 ;
  assign n9389 = n9386 | n9388 ;
  assign n9390 = ( n6164 & n9387 ) | ( n6164 & n9389 ) | ( n9387 & n9389 ) ;
  assign n9391 = x11 & n9389 ;
  assign n9392 = x11 & n9382 ;
  assign n9393 = ( x11 & n9386 ) | ( x11 & n9392 ) | ( n9386 & n9392 ) ;
  assign n9394 = ( n6164 & n9391 ) | ( n6164 & n9393 ) | ( n9391 & n9393 ) ;
  assign n9395 = x11 & ~n9393 ;
  assign n9396 = x11 & ~n9389 ;
  assign n9397 = ( ~n6164 & n9395 ) | ( ~n6164 & n9396 ) | ( n9395 & n9396 ) ;
  assign n9398 = ( n9390 & ~n9394 ) | ( n9390 & n9397 ) | ( ~n9394 & n9397 ) ;
  assign n9399 = n9381 & n9398 ;
  assign n9400 = n9381 & ~n9399 ;
  assign n9401 = ~n9381 & n9398 ;
  assign n9402 = n9400 | n9401 ;
  assign n9403 = n9014 | n9021 ;
  assign n9404 = n9402 | n9403 ;
  assign n9405 = n9402 & n9403 ;
  assign n9406 = n9404 & ~n9405 ;
  assign n9407 = x102 & n389 ;
  assign n9408 = x101 & n384 ;
  assign n9409 = x100 & ~n383 ;
  assign n9410 = n463 & n9409 ;
  assign n9411 = n9408 | n9410 ;
  assign n9412 = n9407 | n9411 ;
  assign n9413 = n392 | n9407 ;
  assign n9414 = n9411 | n9413 ;
  assign n9415 = ( n7178 & n9412 ) | ( n7178 & n9414 ) | ( n9412 & n9414 ) ;
  assign n9416 = x8 & n9414 ;
  assign n9417 = x8 & n9407 ;
  assign n9418 = ( x8 & n9411 ) | ( x8 & n9417 ) | ( n9411 & n9417 ) ;
  assign n9419 = ( n7178 & n9416 ) | ( n7178 & n9418 ) | ( n9416 & n9418 ) ;
  assign n9420 = x8 & ~n9418 ;
  assign n9421 = x8 & ~n9414 ;
  assign n9422 = ( ~n7178 & n9420 ) | ( ~n7178 & n9421 ) | ( n9420 & n9421 ) ;
  assign n9423 = ( n9415 & ~n9419 ) | ( n9415 & n9422 ) | ( ~n9419 & n9422 ) ;
  assign n9424 = n9406 & n9423 ;
  assign n9425 = n9406 & ~n9424 ;
  assign n9426 = ~n9406 & n9423 ;
  assign n9427 = n9425 | n9426 ;
  assign n9428 = n9111 & n9427 ;
  assign n9429 = n9111 | n9427 ;
  assign n9430 = ~n9428 & n9429 ;
  assign n9431 = x105 & n212 ;
  assign n9432 = x104 & n207 ;
  assign n9433 = x103 & ~n206 ;
  assign n9434 = n267 & n9433 ;
  assign n9435 = n9432 | n9434 ;
  assign n9436 = n9431 | n9435 ;
  assign n9437 = n215 | n9431 ;
  assign n9438 = n9435 | n9437 ;
  assign n9439 = ( n8273 & n9436 ) | ( n8273 & n9438 ) | ( n9436 & n9438 ) ;
  assign n9440 = x5 & n9438 ;
  assign n9441 = x5 & n9431 ;
  assign n9442 = ( x5 & n9435 ) | ( x5 & n9441 ) | ( n9435 & n9441 ) ;
  assign n9443 = ( n8273 & n9440 ) | ( n8273 & n9442 ) | ( n9440 & n9442 ) ;
  assign n9444 = x5 & ~n9442 ;
  assign n9445 = x5 & ~n9438 ;
  assign n9446 = ( ~n8273 & n9444 ) | ( ~n8273 & n9445 ) | ( n9444 & n9445 ) ;
  assign n9447 = ( n9439 & ~n9443 ) | ( n9439 & n9446 ) | ( ~n9443 & n9446 ) ;
  assign n9448 = n9430 & n9447 ;
  assign n9449 = n9430 & ~n9448 ;
  assign n9450 = ~n9430 & n9447 ;
  assign n9451 = n9110 & n9450 ;
  assign n9452 = ( n9110 & n9449 ) | ( n9110 & n9451 ) | ( n9449 & n9451 ) ;
  assign n9453 = n9110 & ~n9452 ;
  assign n9454 = n9449 | n9450 ;
  assign n9455 = ~n9452 & n9454 ;
  assign n9456 = n9453 | n9455 ;
  assign n9457 = x107 | x108 ;
  assign n9458 = x107 & x108 ;
  assign n9459 = n9457 & ~n9458 ;
  assign n9460 = n9061 | n9062 ;
  assign n9461 = ( n9061 & n9064 ) | ( n9061 & n9460 ) | ( n9064 & n9460 ) ;
  assign n9462 = n9459 & n9461 ;
  assign n9463 = ( n9061 & n9066 ) | ( n9061 & n9460 ) | ( n9066 & n9460 ) ;
  assign n9464 = n9459 & n9463 ;
  assign n9465 = ( n8261 & n9462 ) | ( n8261 & n9464 ) | ( n9462 & n9464 ) ;
  assign n9466 = ( n8262 & n9462 ) | ( n8262 & n9464 ) | ( n9462 & n9464 ) ;
  assign n9467 = ( n6159 & n9465 ) | ( n6159 & n9466 ) | ( n9465 & n9466 ) ;
  assign n9468 = ( n6157 & n9465 ) | ( n6157 & n9466 ) | ( n9465 & n9466 ) ;
  assign n9469 = ( n5823 & n9467 ) | ( n5823 & n9468 ) | ( n9467 & n9468 ) ;
  assign n9470 = ( n8260 & n9461 ) | ( n8260 & n9463 ) | ( n9461 & n9463 ) ;
  assign n9471 = ( n8258 & n9461 ) | ( n8258 & n9463 ) | ( n9461 & n9463 ) ;
  assign n9472 = ( n7518 & n9470 ) | ( n7518 & n9471 ) | ( n9470 & n9471 ) ;
  assign n9473 = n9459 | n9472 ;
  assign n9474 = ( n7517 & n9470 ) | ( n7517 & n9471 ) | ( n9470 & n9471 ) ;
  assign n9475 = n9459 | n9474 ;
  assign n9476 = ( n6159 & n9473 ) | ( n6159 & n9475 ) | ( n9473 & n9475 ) ;
  assign n9477 = ( n6157 & n9473 ) | ( n6157 & n9475 ) | ( n9473 & n9475 ) ;
  assign n9478 = ( n5823 & n9476 ) | ( n5823 & n9477 ) | ( n9476 & n9477 ) ;
  assign n9479 = ~n9469 & n9478 ;
  assign n9480 = x107 & n133 ;
  assign n9481 = x106 & ~n162 ;
  assign n9482 = ( n137 & n9480 ) | ( n137 & n9481 ) | ( n9480 & n9481 ) ;
  assign n9483 = x0 & x108 ;
  assign n9484 = ( ~n137 & n9480 ) | ( ~n137 & n9483 ) | ( n9480 & n9483 ) ;
  assign n9485 = n9482 | n9484 ;
  assign n9486 = n141 | n9485 ;
  assign n9487 = ( n9479 & n9485 ) | ( n9479 & n9486 ) | ( n9485 & n9486 ) ;
  assign n9488 = x2 & n9485 ;
  assign n9489 = ( x2 & n523 ) | ( x2 & n9485 ) | ( n523 & n9485 ) ;
  assign n9490 = ( n9479 & n9488 ) | ( n9479 & n9489 ) | ( n9488 & n9489 ) ;
  assign n9491 = x2 & ~n9489 ;
  assign n9492 = x2 & ~n9485 ;
  assign n9493 = ( ~n9479 & n9491 ) | ( ~n9479 & n9492 ) | ( n9491 & n9492 ) ;
  assign n9494 = ( n9487 & ~n9490 ) | ( n9487 & n9493 ) | ( ~n9490 & n9493 ) ;
  assign n9495 = n9456 & ~n9494 ;
  assign n9496 = ~n9456 & n9494 ;
  assign n9497 = n9495 | n9496 ;
  assign n9498 = n9108 & n9497 ;
  assign n9499 = n9108 | n9497 ;
  assign n9500 = ~n9498 & n9499 ;
  assign n9501 = x44 & ~x45 ;
  assign n9502 = ~x44 & x45 ;
  assign n9503 = n9501 | n9502 ;
  assign n9504 = x64 & n9503 ;
  assign n9505 = ~n8739 & n9504 ;
  assign n9506 = ( ~n9161 & n9504 ) | ( ~n9161 & n9505 ) | ( n9504 & n9505 ) ;
  assign n9507 = n8739 & ~n9504 ;
  assign n9508 = n9161 & n9507 ;
  assign n9509 = n9506 | n9508 ;
  assign n9510 = x67 & n8724 ;
  assign n9511 = x66 & n8719 ;
  assign n9512 = x65 & ~n8718 ;
  assign n9513 = n9149 & n9512 ;
  assign n9514 = n9511 | n9513 ;
  assign n9515 = n9510 | n9514 ;
  assign n9516 = n186 & n8727 ;
  assign n9517 = n9515 | n9516 ;
  assign n9518 = x44 & ~n9517 ;
  assign n9519 = ~x44 & n9517 ;
  assign n9520 = n9518 | n9519 ;
  assign n9521 = n9509 & n9520 ;
  assign n9522 = n9509 | n9520 ;
  assign n9523 = ~n9521 & n9522 ;
  assign n9524 = x69 & n7561 ;
  assign n9525 = x68 & ~n7560 ;
  assign n9526 = n7953 & n9525 ;
  assign n9527 = n9524 | n9526 ;
  assign n9528 = x70 & n7566 ;
  assign n9529 = n7569 | n9528 ;
  assign n9530 = n9527 | n9529 ;
  assign n9531 = x41 & ~n9530 ;
  assign n9532 = x41 & ~n9528 ;
  assign n9533 = ~n9527 & n9532 ;
  assign n9534 = ( ~n340 & n9531 ) | ( ~n340 & n9533 ) | ( n9531 & n9533 ) ;
  assign n9535 = ~x41 & n9530 ;
  assign n9536 = ~x41 & n9528 ;
  assign n9537 = ( ~x41 & n9527 ) | ( ~x41 & n9536 ) | ( n9527 & n9536 ) ;
  assign n9538 = ( n340 & n9535 ) | ( n340 & n9537 ) | ( n9535 & n9537 ) ;
  assign n9539 = n9534 | n9538 ;
  assign n9540 = n9523 & n9539 ;
  assign n9541 = n9523 & ~n9540 ;
  assign n9542 = ~n9523 & n9539 ;
  assign n9543 = n9541 | n9542 ;
  assign n9544 = n9179 | n9184 ;
  assign n9545 = ( n9179 & n9182 ) | ( n9179 & n9544 ) | ( n9182 & n9544 ) ;
  assign n9546 = n9543 | n9545 ;
  assign n9547 = n9543 & n9545 ;
  assign n9548 = n9546 & ~n9547 ;
  assign n9549 = x73 & n6536 ;
  assign n9550 = x72 & n6531 ;
  assign n9551 = x71 & ~n6530 ;
  assign n9552 = n6871 & n9551 ;
  assign n9553 = n9550 | n9552 ;
  assign n9554 = n9549 | n9553 ;
  assign n9555 = ( ~n610 & n6539 ) | ( ~n610 & n9554 ) | ( n6539 & n9554 ) ;
  assign n9556 = n6539 & n9549 ;
  assign n9557 = ( n6539 & n9553 ) | ( n6539 & n9556 ) | ( n9553 & n9556 ) ;
  assign n9558 = ( n598 & n9555 ) | ( n598 & n9557 ) | ( n9555 & n9557 ) ;
  assign n9559 = ( x38 & ~n9554 ) | ( x38 & n9558 ) | ( ~n9554 & n9558 ) ;
  assign n9560 = ~n9558 & n9559 ;
  assign n9561 = x38 | n9549 ;
  assign n9562 = n9553 | n9561 ;
  assign n9563 = n9558 | n9562 ;
  assign n9564 = ( ~x38 & n9560 ) | ( ~x38 & n9563 ) | ( n9560 & n9563 ) ;
  assign n9565 = n9548 | n9564 ;
  assign n9566 = n9548 & n9564 ;
  assign n9567 = n9565 & ~n9566 ;
  assign n9568 = n9146 & n9207 ;
  assign n9569 = n9204 | n9568 ;
  assign n9570 = n9567 & n9569 ;
  assign n9571 = n9567 | n9569 ;
  assign n9572 = ~n9570 & n9571 ;
  assign n9573 = x76 & n5554 ;
  assign n9574 = x75 & n5549 ;
  assign n9575 = x74 & ~n5548 ;
  assign n9576 = n5893 & n9575 ;
  assign n9577 = n9574 | n9576 ;
  assign n9578 = n9573 | n9577 ;
  assign n9579 = n5557 | n9573 ;
  assign n9580 = n9577 | n9579 ;
  assign n9581 = ( n923 & n9578 ) | ( n923 & n9580 ) | ( n9578 & n9580 ) ;
  assign n9582 = x35 & n9580 ;
  assign n9583 = x35 & n9573 ;
  assign n9584 = ( x35 & n9577 ) | ( x35 & n9583 ) | ( n9577 & n9583 ) ;
  assign n9585 = ( n923 & n9582 ) | ( n923 & n9584 ) | ( n9582 & n9584 ) ;
  assign n9586 = x35 & ~n9584 ;
  assign n9587 = x35 & ~n9580 ;
  assign n9588 = ( ~n923 & n9586 ) | ( ~n923 & n9587 ) | ( n9586 & n9587 ) ;
  assign n9589 = ( n9581 & ~n9585 ) | ( n9581 & n9588 ) | ( ~n9585 & n9588 ) ;
  assign n9590 = n9572 & n9589 ;
  assign n9591 = n9572 & ~n9590 ;
  assign n9592 = ~n9572 & n9589 ;
  assign n9593 = n9591 | n9592 ;
  assign n9594 = n9211 | n9217 ;
  assign n9595 = n9593 & n9594 ;
  assign n9596 = n9593 & ~n9595 ;
  assign n9597 = ~n9593 & n9594 ;
  assign n9598 = n9596 | n9597 ;
  assign n9599 = x79 & n4631 ;
  assign n9600 = x78 & n4626 ;
  assign n9601 = x77 & ~n4625 ;
  assign n9602 = n4943 & n9601 ;
  assign n9603 = n9600 | n9602 ;
  assign n9604 = n9599 | n9603 ;
  assign n9605 = n4634 | n9599 ;
  assign n9606 = n9603 | n9605 ;
  assign n9607 = ( n1332 & n9604 ) | ( n1332 & n9606 ) | ( n9604 & n9606 ) ;
  assign n9608 = x32 & n9606 ;
  assign n9609 = x32 & n9599 ;
  assign n9610 = ( x32 & n9603 ) | ( x32 & n9609 ) | ( n9603 & n9609 ) ;
  assign n9611 = ( n1332 & n9608 ) | ( n1332 & n9610 ) | ( n9608 & n9610 ) ;
  assign n9612 = x32 & ~n9610 ;
  assign n9613 = x32 & ~n9606 ;
  assign n9614 = ( ~n1332 & n9612 ) | ( ~n1332 & n9613 ) | ( n9612 & n9613 ) ;
  assign n9615 = ( n9607 & ~n9611 ) | ( n9607 & n9614 ) | ( ~n9611 & n9614 ) ;
  assign n9616 = n9238 | n9239 ;
  assign n9617 = ( n9238 & n9241 ) | ( n9238 & n9616 ) | ( n9241 & n9616 ) ;
  assign n9618 = ( n9598 & ~n9615 ) | ( n9598 & n9617 ) | ( ~n9615 & n9617 ) ;
  assign n9619 = ( ~n9598 & n9615 ) | ( ~n9598 & n9618 ) | ( n9615 & n9618 ) ;
  assign n9620 = x82 & n3816 ;
  assign n9621 = x81 & n3811 ;
  assign n9622 = x80 & ~n3810 ;
  assign n9623 = n4067 & n9622 ;
  assign n9624 = n9621 | n9623 ;
  assign n9625 = n9620 | n9624 ;
  assign n9626 = n3819 | n9620 ;
  assign n9627 = n9624 | n9626 ;
  assign n9628 = ( n1811 & n9625 ) | ( n1811 & n9627 ) | ( n9625 & n9627 ) ;
  assign n9629 = x29 & n9627 ;
  assign n9630 = x29 & n9620 ;
  assign n9631 = ( x29 & n9624 ) | ( x29 & n9630 ) | ( n9624 & n9630 ) ;
  assign n9632 = ( n1811 & n9629 ) | ( n1811 & n9631 ) | ( n9629 & n9631 ) ;
  assign n9633 = x29 & ~n9631 ;
  assign n9634 = x29 & ~n9627 ;
  assign n9635 = ( ~n1811 & n9633 ) | ( ~n1811 & n9634 ) | ( n9633 & n9634 ) ;
  assign n9636 = ( n9628 & ~n9632 ) | ( n9628 & n9635 ) | ( ~n9632 & n9635 ) ;
  assign n9637 = n9618 & n9636 ;
  assign n9638 = ~n9617 & n9636 ;
  assign n9639 = ( n9619 & n9637 ) | ( n9619 & n9638 ) | ( n9637 & n9638 ) ;
  assign n9640 = n9618 | n9636 ;
  assign n9641 = n9617 & ~n9636 ;
  assign n9642 = ( n9619 & n9640 ) | ( n9619 & ~n9641 ) | ( n9640 & ~n9641 ) ;
  assign n9643 = ~n9639 & n9642 ;
  assign n9644 = n9263 & n9643 ;
  assign n9645 = ( n9266 & n9643 ) | ( n9266 & n9644 ) | ( n9643 & n9644 ) ;
  assign n9646 = n9263 | n9643 ;
  assign n9647 = n9266 | n9646 ;
  assign n9648 = ~n9645 & n9647 ;
  assign n9649 = x85 & n3085 ;
  assign n9650 = x84 & n3080 ;
  assign n9651 = x83 & ~n3079 ;
  assign n9652 = n3309 & n9651 ;
  assign n9653 = n9650 | n9652 ;
  assign n9654 = n9649 | n9653 ;
  assign n9655 = n3088 | n9649 ;
  assign n9656 = n9653 | n9655 ;
  assign n9657 = ( n2381 & n9654 ) | ( n2381 & n9656 ) | ( n9654 & n9656 ) ;
  assign n9658 = x26 & n9656 ;
  assign n9659 = x26 & n9649 ;
  assign n9660 = ( x26 & n9653 ) | ( x26 & n9659 ) | ( n9653 & n9659 ) ;
  assign n9661 = ( n2381 & n9658 ) | ( n2381 & n9660 ) | ( n9658 & n9660 ) ;
  assign n9662 = x26 & ~n9660 ;
  assign n9663 = x26 & ~n9656 ;
  assign n9664 = ( ~n2381 & n9662 ) | ( ~n2381 & n9663 ) | ( n9662 & n9663 ) ;
  assign n9665 = ( n9657 & ~n9661 ) | ( n9657 & n9664 ) | ( ~n9661 & n9664 ) ;
  assign n9666 = n9648 & n9665 ;
  assign n9667 = n9648 & ~n9666 ;
  assign n9668 = ~n9648 & n9665 ;
  assign n9669 = n9667 | n9668 ;
  assign n9670 = n9287 | n9293 ;
  assign n9671 = n9669 | n9670 ;
  assign n9672 = n9669 & n9670 ;
  assign n9673 = n9671 & ~n9672 ;
  assign n9674 = x88 & n2429 ;
  assign n9675 = x87 & n2424 ;
  assign n9676 = x86 & ~n2423 ;
  assign n9677 = n2631 & n9676 ;
  assign n9678 = n9675 | n9677 ;
  assign n9679 = n9674 | n9678 ;
  assign n9680 = n2432 | n9674 ;
  assign n9681 = n9678 | n9680 ;
  assign n9682 = ( ~n3039 & n9679 ) | ( ~n3039 & n9681 ) | ( n9679 & n9681 ) ;
  assign n9683 = n9679 & n9681 ;
  assign n9684 = ( n3023 & n9682 ) | ( n3023 & n9683 ) | ( n9682 & n9683 ) ;
  assign n9685 = x23 & n9681 ;
  assign n9686 = x23 & n9674 ;
  assign n9687 = ( x23 & n9678 ) | ( x23 & n9686 ) | ( n9678 & n9686 ) ;
  assign n9688 = ( ~n3039 & n9685 ) | ( ~n3039 & n9687 ) | ( n9685 & n9687 ) ;
  assign n9689 = n9685 & n9687 ;
  assign n9690 = ( n3023 & n9688 ) | ( n3023 & n9689 ) | ( n9688 & n9689 ) ;
  assign n9691 = x23 & ~n9687 ;
  assign n9692 = x23 & ~n9681 ;
  assign n9693 = ( n3039 & n9691 ) | ( n3039 & n9692 ) | ( n9691 & n9692 ) ;
  assign n9694 = n9691 | n9692 ;
  assign n9695 = ( ~n3023 & n9693 ) | ( ~n3023 & n9694 ) | ( n9693 & n9694 ) ;
  assign n9696 = ( n9684 & ~n9690 ) | ( n9684 & n9695 ) | ( ~n9690 & n9695 ) ;
  assign n9697 = n9673 | n9696 ;
  assign n9698 = n9673 & n9696 ;
  assign n9699 = n9697 & ~n9698 ;
  assign n9700 = ( n9313 & n9316 ) | ( n9313 & n9319 ) | ( n9316 & n9319 ) ;
  assign n9701 = n9699 & n9700 ;
  assign n9702 = n9699 | n9700 ;
  assign n9703 = ~n9701 & n9702 ;
  assign n9704 = x91 & n1859 ;
  assign n9705 = x90 & n1854 ;
  assign n9706 = x89 & ~n1853 ;
  assign n9707 = n2037 & n9706 ;
  assign n9708 = n9705 | n9707 ;
  assign n9709 = n9704 | n9708 ;
  assign n9710 = n1862 | n9704 ;
  assign n9711 = n9708 | n9710 ;
  assign n9712 = ( n3768 & n9709 ) | ( n3768 & n9711 ) | ( n9709 & n9711 ) ;
  assign n9713 = x20 & n9711 ;
  assign n9714 = x20 & n9704 ;
  assign n9715 = ( x20 & n9708 ) | ( x20 & n9714 ) | ( n9708 & n9714 ) ;
  assign n9716 = ( n3768 & n9713 ) | ( n3768 & n9715 ) | ( n9713 & n9715 ) ;
  assign n9717 = x20 & ~n9715 ;
  assign n9718 = x20 & ~n9711 ;
  assign n9719 = ( ~n3768 & n9717 ) | ( ~n3768 & n9718 ) | ( n9717 & n9718 ) ;
  assign n9720 = ( n9712 & ~n9716 ) | ( n9712 & n9719 ) | ( ~n9716 & n9719 ) ;
  assign n9721 = n9703 & n9720 ;
  assign n9722 = n9703 & ~n9721 ;
  assign n9723 = ~n9703 & n9720 ;
  assign n9724 = n9722 | n9723 ;
  assign n9725 = n9322 | n9325 ;
  assign n9726 = ( n9322 & n9327 ) | ( n9322 & n9725 ) | ( n9327 & n9725 ) ;
  assign n9727 = ~n9724 & n9726 ;
  assign n9728 = n9724 & ~n9726 ;
  assign n9729 = n9727 | n9728 ;
  assign n9730 = x94 & n1383 ;
  assign n9731 = x93 & n1378 ;
  assign n9732 = x92 & ~n1377 ;
  assign n9733 = n1542 & n9732 ;
  assign n9734 = n9731 | n9733 ;
  assign n9735 = n9730 | n9734 ;
  assign n9736 = n1386 | n9730 ;
  assign n9737 = n9734 | n9736 ;
  assign n9738 = ( n4583 & n9735 ) | ( n4583 & n9737 ) | ( n9735 & n9737 ) ;
  assign n9739 = x17 & n9737 ;
  assign n9740 = x17 & n9730 ;
  assign n9741 = ( x17 & n9734 ) | ( x17 & n9740 ) | ( n9734 & n9740 ) ;
  assign n9742 = ( n4583 & n9739 ) | ( n4583 & n9741 ) | ( n9739 & n9741 ) ;
  assign n9743 = x17 & ~n9741 ;
  assign n9744 = x17 & ~n9737 ;
  assign n9745 = ( ~n4583 & n9743 ) | ( ~n4583 & n9744 ) | ( n9743 & n9744 ) ;
  assign n9746 = ( n9738 & ~n9742 ) | ( n9738 & n9745 ) | ( ~n9742 & n9745 ) ;
  assign n9747 = n9729 & n9746 ;
  assign n9748 = n9729 | n9746 ;
  assign n9749 = ~n9747 & n9748 ;
  assign n9750 = n9349 | n9350 ;
  assign n9751 = ( n9349 & n9353 ) | ( n9349 & n9750 ) | ( n9353 & n9750 ) ;
  assign n9752 = n9749 & n9751 ;
  assign n9753 = n9749 | n9751 ;
  assign n9754 = ~n9752 & n9753 ;
  assign n9755 = x97 & n962 ;
  assign n9756 = x96 & n957 ;
  assign n9757 = x95 & ~n956 ;
  assign n9758 = n1105 & n9757 ;
  assign n9759 = n9756 | n9758 ;
  assign n9760 = n9755 | n9759 ;
  assign n9761 = n965 | n9755 ;
  assign n9762 = n9759 | n9761 ;
  assign n9763 = ( n5505 & n9760 ) | ( n5505 & n9762 ) | ( n9760 & n9762 ) ;
  assign n9764 = x14 & n9762 ;
  assign n9765 = x14 & n9755 ;
  assign n9766 = ( x14 & n9759 ) | ( x14 & n9765 ) | ( n9759 & n9765 ) ;
  assign n9767 = ( n5505 & n9764 ) | ( n5505 & n9766 ) | ( n9764 & n9766 ) ;
  assign n9768 = x14 & ~n9766 ;
  assign n9769 = x14 & ~n9762 ;
  assign n9770 = ( ~n5505 & n9768 ) | ( ~n5505 & n9769 ) | ( n9768 & n9769 ) ;
  assign n9771 = ( n9763 & ~n9767 ) | ( n9763 & n9770 ) | ( ~n9767 & n9770 ) ;
  assign n9772 = n9754 & n9771 ;
  assign n9773 = n9754 & ~n9772 ;
  assign n9774 = ~n9754 & n9771 ;
  assign n9775 = n9773 | n9774 ;
  assign n9776 = n9375 | n9379 ;
  assign n9777 = ~n9775 & n9776 ;
  assign n9778 = n9775 & ~n9776 ;
  assign n9779 = n9777 | n9778 ;
  assign n9780 = x100 & n636 ;
  assign n9781 = x99 & n631 ;
  assign n9782 = x98 & ~n630 ;
  assign n9783 = n764 & n9782 ;
  assign n9784 = n9781 | n9783 ;
  assign n9785 = n9780 | n9784 ;
  assign n9786 = n639 | n9780 ;
  assign n9787 = n9784 | n9786 ;
  assign n9788 = ( n6483 & n9785 ) | ( n6483 & n9787 ) | ( n9785 & n9787 ) ;
  assign n9789 = x11 & n9787 ;
  assign n9790 = x11 & n9780 ;
  assign n9791 = ( x11 & n9784 ) | ( x11 & n9790 ) | ( n9784 & n9790 ) ;
  assign n9792 = ( n6483 & n9789 ) | ( n6483 & n9791 ) | ( n9789 & n9791 ) ;
  assign n9793 = x11 & ~n9791 ;
  assign n9794 = x11 & ~n9787 ;
  assign n9795 = ( ~n6483 & n9793 ) | ( ~n6483 & n9794 ) | ( n9793 & n9794 ) ;
  assign n9796 = ( n9788 & ~n9792 ) | ( n9788 & n9795 ) | ( ~n9792 & n9795 ) ;
  assign n9797 = n9779 & n9796 ;
  assign n9798 = n9779 | n9796 ;
  assign n9799 = ~n9797 & n9798 ;
  assign n9800 = n9399 & n9799 ;
  assign n9801 = ( n9405 & n9799 ) | ( n9405 & n9800 ) | ( n9799 & n9800 ) ;
  assign n9802 = n9399 | n9799 ;
  assign n9803 = n9405 | n9802 ;
  assign n9804 = ~n9801 & n9803 ;
  assign n9805 = x103 & n389 ;
  assign n9806 = x102 & n384 ;
  assign n9807 = x101 & ~n383 ;
  assign n9808 = n463 & n9807 ;
  assign n9809 = n9806 | n9808 ;
  assign n9810 = n9805 | n9809 ;
  assign n9811 = n392 | n9805 ;
  assign n9812 = n9809 | n9811 ;
  assign n9813 = ( n7529 & n9810 ) | ( n7529 & n9812 ) | ( n9810 & n9812 ) ;
  assign n9814 = x8 & n9812 ;
  assign n9815 = x8 & n9805 ;
  assign n9816 = ( x8 & n9809 ) | ( x8 & n9815 ) | ( n9809 & n9815 ) ;
  assign n9817 = ( n7529 & n9814 ) | ( n7529 & n9816 ) | ( n9814 & n9816 ) ;
  assign n9818 = x8 & ~n9816 ;
  assign n9819 = x8 & ~n9812 ;
  assign n9820 = ( ~n7529 & n9818 ) | ( ~n7529 & n9819 ) | ( n9818 & n9819 ) ;
  assign n9821 = ( n9813 & ~n9817 ) | ( n9813 & n9820 ) | ( ~n9817 & n9820 ) ;
  assign n9822 = n9804 & n9821 ;
  assign n9823 = n9804 & ~n9822 ;
  assign n9824 = ~n9804 & n9821 ;
  assign n9825 = n9823 | n9824 ;
  assign n9826 = n9111 | n9424 ;
  assign n9827 = ( n9424 & n9427 ) | ( n9424 & n9826 ) | ( n9427 & n9826 ) ;
  assign n9828 = n9825 | n9827 ;
  assign n9829 = n9825 & n9827 ;
  assign n9830 = n9828 & ~n9829 ;
  assign n9831 = x106 & n212 ;
  assign n9832 = x105 & n207 ;
  assign n9833 = x104 & ~n206 ;
  assign n9834 = n267 & n9833 ;
  assign n9835 = n9832 | n9834 ;
  assign n9836 = n9831 | n9835 ;
  assign n9837 = n215 | n9831 ;
  assign n9838 = n9835 | n9837 ;
  assign n9839 = ( n8656 & n9836 ) | ( n8656 & n9838 ) | ( n9836 & n9838 ) ;
  assign n9840 = x5 & n9838 ;
  assign n9841 = x5 & n9831 ;
  assign n9842 = ( x5 & n9835 ) | ( x5 & n9841 ) | ( n9835 & n9841 ) ;
  assign n9843 = ( n8656 & n9840 ) | ( n8656 & n9842 ) | ( n9840 & n9842 ) ;
  assign n9844 = x5 & ~n9842 ;
  assign n9845 = x5 & ~n9838 ;
  assign n9846 = ( ~n8656 & n9844 ) | ( ~n8656 & n9845 ) | ( n9844 & n9845 ) ;
  assign n9847 = ( n9839 & ~n9843 ) | ( n9839 & n9846 ) | ( ~n9843 & n9846 ) ;
  assign n9848 = n9830 & n9847 ;
  assign n9849 = n9830 & ~n9848 ;
  assign n9850 = ~n9830 & n9847 ;
  assign n9851 = n9849 | n9850 ;
  assign n9852 = n9448 | n9452 ;
  assign n9853 = n9851 | n9852 ;
  assign n9854 = n9851 & n9852 ;
  assign n9855 = n9853 & ~n9854 ;
  assign n9856 = x108 | x109 ;
  assign n9857 = x108 & x109 ;
  assign n9858 = n9856 & ~n9857 ;
  assign n9859 = n9458 | n9459 ;
  assign n9860 = n9858 & n9859 ;
  assign n9861 = n9458 & n9858 ;
  assign n9862 = ( n9461 & n9860 ) | ( n9461 & n9861 ) | ( n9860 & n9861 ) ;
  assign n9863 = ( n9463 & n9860 ) | ( n9463 & n9861 ) | ( n9860 & n9861 ) ;
  assign n9864 = ( n8261 & n9862 ) | ( n8261 & n9863 ) | ( n9862 & n9863 ) ;
  assign n9865 = ( n8262 & n9862 ) | ( n8262 & n9863 ) | ( n9862 & n9863 ) ;
  assign n9866 = ( n6159 & n9864 ) | ( n6159 & n9865 ) | ( n9864 & n9865 ) ;
  assign n9867 = ( n6157 & n9864 ) | ( n6157 & n9865 ) | ( n9864 & n9865 ) ;
  assign n9868 = ( n5823 & n9866 ) | ( n5823 & n9867 ) | ( n9866 & n9867 ) ;
  assign n9869 = ( n9458 & n9463 ) | ( n9458 & n9859 ) | ( n9463 & n9859 ) ;
  assign n9870 = n9858 | n9869 ;
  assign n9871 = ( n9458 & n9461 ) | ( n9458 & n9859 ) | ( n9461 & n9859 ) ;
  assign n9872 = n9858 | n9871 ;
  assign n9873 = ( n8262 & n9870 ) | ( n8262 & n9872 ) | ( n9870 & n9872 ) ;
  assign n9874 = ( n8261 & n9870 ) | ( n8261 & n9872 ) | ( n9870 & n9872 ) ;
  assign n9875 = ( n6159 & n9873 ) | ( n6159 & n9874 ) | ( n9873 & n9874 ) ;
  assign n9876 = ( n6157 & n9873 ) | ( n6157 & n9874 ) | ( n9873 & n9874 ) ;
  assign n9877 = ( n5823 & n9875 ) | ( n5823 & n9876 ) | ( n9875 & n9876 ) ;
  assign n9878 = ~n9868 & n9877 ;
  assign n9879 = x108 & n133 ;
  assign n9880 = x107 & ~n162 ;
  assign n9881 = ( n137 & n9879 ) | ( n137 & n9880 ) | ( n9879 & n9880 ) ;
  assign n9882 = x0 & x109 ;
  assign n9883 = ( ~n137 & n9879 ) | ( ~n137 & n9882 ) | ( n9879 & n9882 ) ;
  assign n9884 = n9881 | n9883 ;
  assign n9885 = n141 | n9884 ;
  assign n9886 = ( n9878 & n9884 ) | ( n9878 & n9885 ) | ( n9884 & n9885 ) ;
  assign n9887 = x2 & n9884 ;
  assign n9888 = ( x2 & n523 ) | ( x2 & n9884 ) | ( n523 & n9884 ) ;
  assign n9889 = ( n9878 & n9887 ) | ( n9878 & n9888 ) | ( n9887 & n9888 ) ;
  assign n9890 = x2 & ~n9888 ;
  assign n9891 = x2 & ~n9884 ;
  assign n9892 = ( ~n9878 & n9890 ) | ( ~n9878 & n9891 ) | ( n9890 & n9891 ) ;
  assign n9893 = ( n9886 & ~n9889 ) | ( n9886 & n9892 ) | ( ~n9889 & n9892 ) ;
  assign n9894 = n9855 | n9893 ;
  assign n9895 = n9855 & n9893 ;
  assign n9896 = n9894 & ~n9895 ;
  assign n9897 = ( n9100 & n9456 ) | ( n9100 & n9494 ) | ( n9456 & n9494 ) ;
  assign n9898 = n9456 | n9494 ;
  assign n9899 = ( n9105 & n9897 ) | ( n9105 & n9898 ) | ( n9897 & n9898 ) ;
  assign n9900 = n9896 | n9899 ;
  assign n9901 = n9896 & n9899 ;
  assign n9902 = n9900 & ~n9901 ;
  assign n9903 = n9822 | n9827 ;
  assign n9904 = ( n9822 & n9825 ) | ( n9822 & n9903 ) | ( n9825 & n9903 ) ;
  assign n9905 = n9747 | n9752 ;
  assign n9906 = x95 & n1383 ;
  assign n9907 = x94 & n1378 ;
  assign n9908 = x93 & ~n1377 ;
  assign n9909 = n1542 & n9908 ;
  assign n9910 = n9907 | n9909 ;
  assign n9911 = n9906 | n9910 ;
  assign n9912 = n1386 | n9906 ;
  assign n9913 = n9910 | n9912 ;
  assign n9914 = ( n4897 & n9911 ) | ( n4897 & n9913 ) | ( n9911 & n9913 ) ;
  assign n9915 = x17 & n9913 ;
  assign n9916 = x17 & n9906 ;
  assign n9917 = ( x17 & n9910 ) | ( x17 & n9916 ) | ( n9910 & n9916 ) ;
  assign n9918 = ( n4897 & n9915 ) | ( n4897 & n9917 ) | ( n9915 & n9917 ) ;
  assign n9919 = x17 & ~n9917 ;
  assign n9920 = x17 & ~n9913 ;
  assign n9921 = ( ~n4897 & n9919 ) | ( ~n4897 & n9920 ) | ( n9919 & n9920 ) ;
  assign n9922 = ( n9914 & ~n9918 ) | ( n9914 & n9921 ) | ( ~n9918 & n9921 ) ;
  assign n9923 = n9566 | n9567 ;
  assign n9924 = ( n9566 & n9569 ) | ( n9566 & n9923 ) | ( n9569 & n9923 ) ;
  assign n9925 = ~x45 & x46 ;
  assign n9926 = x45 & ~x46 ;
  assign n9927 = n9925 | n9926 ;
  assign n9928 = ~n9503 & n9927 ;
  assign n9929 = x64 & n9928 ;
  assign n9930 = ~x46 & x47 ;
  assign n9931 = x46 & ~x47 ;
  assign n9932 = n9930 | n9931 ;
  assign n9933 = n9503 & ~n9932 ;
  assign n9934 = x65 & n9933 ;
  assign n9935 = n9929 | n9934 ;
  assign n9936 = n9503 & n9932 ;
  assign n9937 = x47 | n144 ;
  assign n9938 = ( x47 & n9936 ) | ( x47 & n9937 ) | ( n9936 & n9937 ) ;
  assign n9939 = ~x47 & n9938 ;
  assign n9940 = ( ~x47 & n9935 ) | ( ~x47 & n9939 ) | ( n9935 & n9939 ) ;
  assign n9941 = x47 & ~x64 ;
  assign n9942 = ( x47 & ~n9503 ) | ( x47 & n9941 ) | ( ~n9503 & n9941 ) ;
  assign n9943 = n9938 & n9942 ;
  assign n9944 = ( n9935 & n9942 ) | ( n9935 & n9943 ) | ( n9942 & n9943 ) ;
  assign n9945 = n144 & n9936 ;
  assign n9946 = n9942 & ~n9945 ;
  assign n9947 = ~n9935 & n9946 ;
  assign n9948 = ( n9940 & n9944 ) | ( n9940 & n9947 ) | ( n9944 & n9947 ) ;
  assign n9949 = n9938 | n9942 ;
  assign n9950 = n9935 | n9949 ;
  assign n9951 = ~n9942 & n9945 ;
  assign n9952 = ( n9935 & ~n9942 ) | ( n9935 & n9951 ) | ( ~n9942 & n9951 ) ;
  assign n9953 = ( n9940 & n9950 ) | ( n9940 & ~n9952 ) | ( n9950 & ~n9952 ) ;
  assign n9954 = ~n9948 & n9953 ;
  assign n9955 = n241 & n8727 ;
  assign n9956 = x68 & n8724 ;
  assign n9957 = x67 & n8719 ;
  assign n9958 = x66 & ~n8718 ;
  assign n9959 = n9149 & n9958 ;
  assign n9960 = n9957 | n9959 ;
  assign n9961 = n9956 | n9960 ;
  assign n9962 = n9955 | n9961 ;
  assign n9963 = x44 | n9956 ;
  assign n9964 = n9960 | n9963 ;
  assign n9965 = n9955 | n9964 ;
  assign n9966 = ~x44 & n9964 ;
  assign n9967 = ( ~x44 & n9955 ) | ( ~x44 & n9966 ) | ( n9955 & n9966 ) ;
  assign n9968 = ( ~n9962 & n9965 ) | ( ~n9962 & n9967 ) | ( n9965 & n9967 ) ;
  assign n9969 = n9954 | n9968 ;
  assign n9970 = n9954 & n9968 ;
  assign n9971 = n9969 & ~n9970 ;
  assign n9972 = ( n9163 & n9504 ) | ( n9163 & n9520 ) | ( n9504 & n9520 ) ;
  assign n9973 = n9971 | n9972 ;
  assign n9974 = n9971 & n9972 ;
  assign n9975 = n9973 & ~n9974 ;
  assign n9976 = x70 & n7561 ;
  assign n9977 = x69 & ~n7560 ;
  assign n9978 = n7953 & n9977 ;
  assign n9979 = n9976 | n9978 ;
  assign n9980 = x71 & n7566 ;
  assign n9981 = n7569 | n9980 ;
  assign n9982 = n9979 | n9981 ;
  assign n9983 = x41 & ~n9982 ;
  assign n9984 = x41 & ~n9980 ;
  assign n9985 = ~n9979 & n9984 ;
  assign n9986 = ( ~n438 & n9983 ) | ( ~n438 & n9985 ) | ( n9983 & n9985 ) ;
  assign n9987 = ~x41 & n9982 ;
  assign n9988 = ~x41 & n9980 ;
  assign n9989 = ( ~x41 & n9979 ) | ( ~x41 & n9988 ) | ( n9979 & n9988 ) ;
  assign n9990 = ( n438 & n9987 ) | ( n438 & n9989 ) | ( n9987 & n9989 ) ;
  assign n9991 = n9986 | n9990 ;
  assign n9992 = n9975 & n9991 ;
  assign n9993 = n9975 & ~n9992 ;
  assign n9994 = ~n9975 & n9991 ;
  assign n9995 = n9993 | n9994 ;
  assign n9996 = n9540 | n9545 ;
  assign n9997 = ( n9540 & n9543 ) | ( n9540 & n9996 ) | ( n9543 & n9996 ) ;
  assign n9998 = n9995 | n9997 ;
  assign n9999 = n9995 & n9997 ;
  assign n10000 = n9998 & ~n9999 ;
  assign n10001 = x74 & n6536 ;
  assign n10002 = x73 & n6531 ;
  assign n10003 = x72 & ~n6530 ;
  assign n10004 = n6871 & n10003 ;
  assign n10005 = n10002 | n10004 ;
  assign n10006 = n10001 | n10005 ;
  assign n10007 = n6539 | n10001 ;
  assign n10008 = n10005 | n10007 ;
  assign n10009 = ( n710 & n10006 ) | ( n710 & n10008 ) | ( n10006 & n10008 ) ;
  assign n10010 = x38 & n10008 ;
  assign n10011 = x38 & n10001 ;
  assign n10012 = ( x38 & n10005 ) | ( x38 & n10011 ) | ( n10005 & n10011 ) ;
  assign n10013 = ( n710 & n10010 ) | ( n710 & n10012 ) | ( n10010 & n10012 ) ;
  assign n10014 = x38 & ~n10012 ;
  assign n10015 = x38 & ~n10008 ;
  assign n10016 = ( ~n710 & n10014 ) | ( ~n710 & n10015 ) | ( n10014 & n10015 ) ;
  assign n10017 = ( n10009 & ~n10013 ) | ( n10009 & n10016 ) | ( ~n10013 & n10016 ) ;
  assign n10018 = n10000 & n10017 ;
  assign n10019 = n10000 | n10017 ;
  assign n10020 = ~n10018 & n10019 ;
  assign n10021 = n9924 & n10020 ;
  assign n10022 = n9924 & ~n10021 ;
  assign n10023 = x77 & n5554 ;
  assign n10024 = x76 & n5549 ;
  assign n10025 = x75 & ~n5548 ;
  assign n10026 = n5893 & n10025 ;
  assign n10027 = n10024 | n10026 ;
  assign n10028 = n10023 | n10027 ;
  assign n10029 = n5557 | n10023 ;
  assign n10030 = n10027 | n10029 ;
  assign n10031 = ( n1059 & n10028 ) | ( n1059 & n10030 ) | ( n10028 & n10030 ) ;
  assign n10032 = x35 & n10030 ;
  assign n10033 = x35 & n10023 ;
  assign n10034 = ( x35 & n10027 ) | ( x35 & n10033 ) | ( n10027 & n10033 ) ;
  assign n10035 = ( n1059 & n10032 ) | ( n1059 & n10034 ) | ( n10032 & n10034 ) ;
  assign n10036 = x35 & ~n10034 ;
  assign n10037 = x35 & ~n10030 ;
  assign n10038 = ( ~n1059 & n10036 ) | ( ~n1059 & n10037 ) | ( n10036 & n10037 ) ;
  assign n10039 = ( n10031 & ~n10035 ) | ( n10031 & n10038 ) | ( ~n10035 & n10038 ) ;
  assign n10040 = ~n10019 & n10020 ;
  assign n10041 = ( ~n9924 & n10020 ) | ( ~n9924 & n10040 ) | ( n10020 & n10040 ) ;
  assign n10042 = n10039 & n10041 ;
  assign n10043 = ( n10022 & n10039 ) | ( n10022 & n10042 ) | ( n10039 & n10042 ) ;
  assign n10044 = n10039 | n10041 ;
  assign n10045 = n10022 | n10044 ;
  assign n10046 = ~n10043 & n10045 ;
  assign n10047 = n9590 | n9594 ;
  assign n10048 = ( n9590 & n9593 ) | ( n9590 & n10047 ) | ( n9593 & n10047 ) ;
  assign n10049 = n10046 & n10048 ;
  assign n10050 = n10046 | n10048 ;
  assign n10051 = ~n10049 & n10050 ;
  assign n10052 = x80 & n4631 ;
  assign n10053 = x79 & n4626 ;
  assign n10054 = x78 & ~n4625 ;
  assign n10055 = n4943 & n10054 ;
  assign n10056 = n10053 | n10055 ;
  assign n10057 = n10052 | n10056 ;
  assign n10058 = n4634 | n10052 ;
  assign n10059 = n10056 | n10058 ;
  assign n10060 = ( n1499 & n10057 ) | ( n1499 & n10059 ) | ( n10057 & n10059 ) ;
  assign n10061 = x32 & n10059 ;
  assign n10062 = x32 & n10052 ;
  assign n10063 = ( x32 & n10056 ) | ( x32 & n10062 ) | ( n10056 & n10062 ) ;
  assign n10064 = ( n1499 & n10061 ) | ( n1499 & n10063 ) | ( n10061 & n10063 ) ;
  assign n10065 = x32 & ~n10063 ;
  assign n10066 = x32 & ~n10059 ;
  assign n10067 = ( ~n1499 & n10065 ) | ( ~n1499 & n10066 ) | ( n10065 & n10066 ) ;
  assign n10068 = ( n10060 & ~n10064 ) | ( n10060 & n10067 ) | ( ~n10064 & n10067 ) ;
  assign n10069 = n10051 & n10068 ;
  assign n10070 = n10051 & ~n10069 ;
  assign n10071 = ~n10051 & n10068 ;
  assign n10072 = n10070 | n10071 ;
  assign n10073 = n9594 & n9615 ;
  assign n10074 = ~n9593 & n10073 ;
  assign n10075 = ( n9596 & n9615 ) | ( n9596 & n10074 ) | ( n9615 & n10074 ) ;
  assign n10076 = n9598 & ~n10075 ;
  assign n10077 = ~n9594 & n9615 ;
  assign n10078 = ( n9593 & n9615 ) | ( n9593 & n10077 ) | ( n9615 & n10077 ) ;
  assign n10079 = ~n9596 & n10078 ;
  assign n10080 = n9617 & ~n10079 ;
  assign n10081 = ~n10076 & n10080 ;
  assign n10082 = ( n9617 & n10075 ) | ( n9617 & ~n10081 ) | ( n10075 & ~n10081 ) ;
  assign n10083 = n10072 | n10082 ;
  assign n10084 = n10072 & n10082 ;
  assign n10085 = n10083 & ~n10084 ;
  assign n10086 = x83 & n3816 ;
  assign n10087 = x82 & n3811 ;
  assign n10088 = x81 & ~n3810 ;
  assign n10089 = n4067 & n10088 ;
  assign n10090 = n10087 | n10089 ;
  assign n10091 = n10086 | n10090 ;
  assign n10092 = n3819 | n10086 ;
  assign n10093 = n10090 | n10092 ;
  assign n10094 = ( n2009 & n10091 ) | ( n2009 & n10093 ) | ( n10091 & n10093 ) ;
  assign n10095 = x29 & n10093 ;
  assign n10096 = x29 & n10086 ;
  assign n10097 = ( x29 & n10090 ) | ( x29 & n10096 ) | ( n10090 & n10096 ) ;
  assign n10098 = ( n2009 & n10095 ) | ( n2009 & n10097 ) | ( n10095 & n10097 ) ;
  assign n10099 = x29 & ~n10097 ;
  assign n10100 = x29 & ~n10093 ;
  assign n10101 = ( ~n2009 & n10099 ) | ( ~n2009 & n10100 ) | ( n10099 & n10100 ) ;
  assign n10102 = ( n10094 & ~n10098 ) | ( n10094 & n10101 ) | ( ~n10098 & n10101 ) ;
  assign n10103 = n10085 & n10102 ;
  assign n10104 = n10085 & ~n10103 ;
  assign n10105 = ~n10085 & n10102 ;
  assign n10106 = n10104 | n10105 ;
  assign n10107 = n9639 | n9645 ;
  assign n10108 = n10106 | n10107 ;
  assign n10109 = n10106 & n10107 ;
  assign n10110 = n10108 & ~n10109 ;
  assign n10111 = x86 & n3085 ;
  assign n10112 = x85 & n3080 ;
  assign n10113 = x84 & ~n3079 ;
  assign n10114 = n3309 & n10113 ;
  assign n10115 = n10112 | n10114 ;
  assign n10116 = n10111 | n10115 ;
  assign n10117 = n3088 | n10111 ;
  assign n10118 = n10115 | n10117 ;
  assign n10119 = ( n2606 & n10116 ) | ( n2606 & n10118 ) | ( n10116 & n10118 ) ;
  assign n10120 = x26 & n10118 ;
  assign n10121 = x26 & n10111 ;
  assign n10122 = ( x26 & n10115 ) | ( x26 & n10121 ) | ( n10115 & n10121 ) ;
  assign n10123 = ( n2606 & n10120 ) | ( n2606 & n10122 ) | ( n10120 & n10122 ) ;
  assign n10124 = x26 & ~n10122 ;
  assign n10125 = x26 & ~n10118 ;
  assign n10126 = ( ~n2606 & n10124 ) | ( ~n2606 & n10125 ) | ( n10124 & n10125 ) ;
  assign n10127 = ( n10119 & ~n10123 ) | ( n10119 & n10126 ) | ( ~n10123 & n10126 ) ;
  assign n10128 = n10110 & n10127 ;
  assign n10129 = n10110 & ~n10128 ;
  assign n10130 = ~n10110 & n10127 ;
  assign n10131 = n10129 | n10130 ;
  assign n10132 = n9666 | n9668 ;
  assign n10133 = n9667 | n10132 ;
  assign n10134 = ( n9666 & n9670 ) | ( n9666 & n10133 ) | ( n9670 & n10133 ) ;
  assign n10135 = n10131 | n10134 ;
  assign n10136 = n10131 & n10134 ;
  assign n10137 = n10135 & ~n10136 ;
  assign n10138 = x89 & n2429 ;
  assign n10139 = x88 & n2424 ;
  assign n10140 = x87 & ~n2423 ;
  assign n10141 = n2631 & n10140 ;
  assign n10142 = n10139 | n10141 ;
  assign n10143 = n10138 | n10142 ;
  assign n10144 = n2432 | n10138 ;
  assign n10145 = n10142 | n10144 ;
  assign n10146 = ( n3282 & n10143 ) | ( n3282 & n10145 ) | ( n10143 & n10145 ) ;
  assign n10147 = x23 & n10145 ;
  assign n10148 = x23 & n10138 ;
  assign n10149 = ( x23 & n10142 ) | ( x23 & n10148 ) | ( n10142 & n10148 ) ;
  assign n10150 = ( n3282 & n10147 ) | ( n3282 & n10149 ) | ( n10147 & n10149 ) ;
  assign n10151 = x23 & ~n10149 ;
  assign n10152 = x23 & ~n10145 ;
  assign n10153 = ( ~n3282 & n10151 ) | ( ~n3282 & n10152 ) | ( n10151 & n10152 ) ;
  assign n10154 = ( n10146 & ~n10150 ) | ( n10146 & n10153 ) | ( ~n10150 & n10153 ) ;
  assign n10155 = n10137 & n10154 ;
  assign n10156 = n10137 & ~n10155 ;
  assign n10157 = ~n10137 & n10154 ;
  assign n10158 = n10156 | n10157 ;
  assign n10159 = n9698 | n9701 ;
  assign n10160 = n10158 & n10159 ;
  assign n10161 = n10158 | n10159 ;
  assign n10162 = ~n10160 & n10161 ;
  assign n10163 = x92 & n1859 ;
  assign n10164 = x91 & n1854 ;
  assign n10165 = x90 & ~n1853 ;
  assign n10166 = n2037 & n10165 ;
  assign n10167 = n10164 | n10166 ;
  assign n10168 = n10163 | n10167 ;
  assign n10169 = n1862 | n10163 ;
  assign n10170 = n10167 | n10169 ;
  assign n10171 = ( n4040 & n10168 ) | ( n4040 & n10170 ) | ( n10168 & n10170 ) ;
  assign n10172 = x20 & n10170 ;
  assign n10173 = x20 & n10163 ;
  assign n10174 = ( x20 & n10167 ) | ( x20 & n10173 ) | ( n10167 & n10173 ) ;
  assign n10175 = ( n4040 & n10172 ) | ( n4040 & n10174 ) | ( n10172 & n10174 ) ;
  assign n10176 = x20 & ~n10174 ;
  assign n10177 = x20 & ~n10170 ;
  assign n10178 = ( ~n4040 & n10176 ) | ( ~n4040 & n10177 ) | ( n10176 & n10177 ) ;
  assign n10179 = ( n10171 & ~n10175 ) | ( n10171 & n10178 ) | ( ~n10175 & n10178 ) ;
  assign n10180 = n10162 & n10179 ;
  assign n10181 = n10162 & ~n10180 ;
  assign n10182 = ~n10162 & n10179 ;
  assign n10183 = ( n9322 & n9703 ) | ( n9322 & n9720 ) | ( n9703 & n9720 ) ;
  assign n10184 = n9703 | n9720 ;
  assign n10185 = ( n9328 & n10183 ) | ( n9328 & n10184 ) | ( n10183 & n10184 ) ;
  assign n10186 = ~n10182 & n10185 ;
  assign n10187 = ~n10181 & n10186 ;
  assign n10188 = n9922 & n10187 ;
  assign n10189 = n10182 & ~n10185 ;
  assign n10190 = ( n10181 & ~n10185 ) | ( n10181 & n10189 ) | ( ~n10185 & n10189 ) ;
  assign n10191 = ( n9922 & n10188 ) | ( n9922 & n10190 ) | ( n10188 & n10190 ) ;
  assign n10192 = n9922 | n10187 ;
  assign n10193 = n10190 | n10192 ;
  assign n10194 = ~n10191 & n10193 ;
  assign n10195 = n9905 & n10194 ;
  assign n10196 = n9905 | n10194 ;
  assign n10197 = ~n10195 & n10196 ;
  assign n10198 = x98 & n962 ;
  assign n10199 = x97 & n957 ;
  assign n10200 = x96 & ~n956 ;
  assign n10201 = n1105 & n10200 ;
  assign n10202 = n10199 | n10201 ;
  assign n10203 = n10198 | n10202 ;
  assign n10204 = n965 | n10198 ;
  assign n10205 = n10202 | n10204 ;
  assign n10206 = ( ~n5850 & n10203 ) | ( ~n5850 & n10205 ) | ( n10203 & n10205 ) ;
  assign n10207 = n10203 & n10205 ;
  assign n10208 = ( n5834 & n10206 ) | ( n5834 & n10207 ) | ( n10206 & n10207 ) ;
  assign n10209 = x14 & n10205 ;
  assign n10210 = x14 & n10198 ;
  assign n10211 = ( x14 & n10202 ) | ( x14 & n10210 ) | ( n10202 & n10210 ) ;
  assign n10212 = ( ~n5850 & n10209 ) | ( ~n5850 & n10211 ) | ( n10209 & n10211 ) ;
  assign n10213 = n10209 & n10211 ;
  assign n10214 = ( n5834 & n10212 ) | ( n5834 & n10213 ) | ( n10212 & n10213 ) ;
  assign n10215 = x14 & ~n10211 ;
  assign n10216 = x14 & ~n10205 ;
  assign n10217 = ( n5850 & n10215 ) | ( n5850 & n10216 ) | ( n10215 & n10216 ) ;
  assign n10218 = n10215 | n10216 ;
  assign n10219 = ( ~n5834 & n10217 ) | ( ~n5834 & n10218 ) | ( n10217 & n10218 ) ;
  assign n10220 = ( n10208 & ~n10214 ) | ( n10208 & n10219 ) | ( ~n10214 & n10219 ) ;
  assign n10221 = n10197 & n10220 ;
  assign n10222 = n10197 & ~n10221 ;
  assign n10223 = ( n9375 & n9754 ) | ( n9375 & n9771 ) | ( n9754 & n9771 ) ;
  assign n10224 = n9754 | n9771 ;
  assign n10225 = ( n9379 & n10223 ) | ( n9379 & n10224 ) | ( n10223 & n10224 ) ;
  assign n10226 = ~n10197 & n10220 ;
  assign n10227 = n10225 & n10226 ;
  assign n10228 = ( n10222 & n10225 ) | ( n10222 & n10227 ) | ( n10225 & n10227 ) ;
  assign n10229 = n10225 | n10226 ;
  assign n10230 = n10222 | n10229 ;
  assign n10231 = ~n10228 & n10230 ;
  assign n10232 = x101 & n636 ;
  assign n10233 = x100 & n631 ;
  assign n10234 = x99 & ~n630 ;
  assign n10235 = n764 & n10234 ;
  assign n10236 = n10233 | n10235 ;
  assign n10237 = n10232 | n10236 ;
  assign n10238 = n639 | n10232 ;
  assign n10239 = n10236 | n10238 ;
  assign n10240 = ( n6844 & n10237 ) | ( n6844 & n10239 ) | ( n10237 & n10239 ) ;
  assign n10241 = x11 & n10239 ;
  assign n10242 = x11 & n10232 ;
  assign n10243 = ( x11 & n10236 ) | ( x11 & n10242 ) | ( n10236 & n10242 ) ;
  assign n10244 = ( n6844 & n10241 ) | ( n6844 & n10243 ) | ( n10241 & n10243 ) ;
  assign n10245 = x11 & ~n10243 ;
  assign n10246 = x11 & ~n10239 ;
  assign n10247 = ( ~n6844 & n10245 ) | ( ~n6844 & n10246 ) | ( n10245 & n10246 ) ;
  assign n10248 = ( n10240 & ~n10244 ) | ( n10240 & n10247 ) | ( ~n10244 & n10247 ) ;
  assign n10249 = n10231 & n10248 ;
  assign n10250 = n10231 & ~n10249 ;
  assign n10251 = ~n10231 & n10248 ;
  assign n10252 = n10250 | n10251 ;
  assign n10253 = n9797 | n9799 ;
  assign n10254 = n9405 | n9797 ;
  assign n10255 = ( n9800 & n10253 ) | ( n9800 & n10254 ) | ( n10253 & n10254 ) ;
  assign n10256 = n10252 | n10255 ;
  assign n10257 = n10252 & n10255 ;
  assign n10258 = n10256 & ~n10257 ;
  assign n10259 = x104 & n389 ;
  assign n10260 = x103 & n384 ;
  assign n10261 = x102 & ~n383 ;
  assign n10262 = n463 & n10261 ;
  assign n10263 = n10260 | n10262 ;
  assign n10264 = n10259 | n10263 ;
  assign n10265 = n392 | n10259 ;
  assign n10266 = n10263 | n10265 ;
  assign n10267 = ( n7911 & n10264 ) | ( n7911 & n10266 ) | ( n10264 & n10266 ) ;
  assign n10268 = x8 & n10266 ;
  assign n10269 = x8 & n10259 ;
  assign n10270 = ( x8 & n10263 ) | ( x8 & n10269 ) | ( n10263 & n10269 ) ;
  assign n10271 = ( n7911 & n10268 ) | ( n7911 & n10270 ) | ( n10268 & n10270 ) ;
  assign n10272 = x8 & ~n10270 ;
  assign n10273 = x8 & ~n10266 ;
  assign n10274 = ( ~n7911 & n10272 ) | ( ~n7911 & n10273 ) | ( n10272 & n10273 ) ;
  assign n10275 = ( n10267 & ~n10271 ) | ( n10267 & n10274 ) | ( ~n10271 & n10274 ) ;
  assign n10276 = n10258 & n10275 ;
  assign n10277 = n10258 | n10275 ;
  assign n10278 = ~n10276 & n10277 ;
  assign n10279 = n9904 & n10278 ;
  assign n10280 = n9904 & ~n10279 ;
  assign n10281 = x107 & n212 ;
  assign n10282 = x106 & n207 ;
  assign n10283 = x105 & ~n206 ;
  assign n10284 = n267 & n10283 ;
  assign n10285 = n10282 | n10284 ;
  assign n10286 = n10281 | n10285 ;
  assign n10287 = n215 | n10281 ;
  assign n10288 = n10285 | n10287 ;
  assign n10289 = ( n9084 & n10286 ) | ( n9084 & n10288 ) | ( n10286 & n10288 ) ;
  assign n10290 = x5 & n10288 ;
  assign n10291 = x5 & n10281 ;
  assign n10292 = ( x5 & n10285 ) | ( x5 & n10291 ) | ( n10285 & n10291 ) ;
  assign n10293 = ( n9084 & n10290 ) | ( n9084 & n10292 ) | ( n10290 & n10292 ) ;
  assign n10294 = x5 & ~n10292 ;
  assign n10295 = x5 & ~n10288 ;
  assign n10296 = ( ~n9084 & n10294 ) | ( ~n9084 & n10295 ) | ( n10294 & n10295 ) ;
  assign n10297 = ( n10289 & ~n10293 ) | ( n10289 & n10296 ) | ( ~n10293 & n10296 ) ;
  assign n10298 = ~n10277 & n10278 ;
  assign n10299 = ( ~n9904 & n10278 ) | ( ~n9904 & n10298 ) | ( n10278 & n10298 ) ;
  assign n10300 = n10297 & n10299 ;
  assign n10301 = ( n10280 & n10297 ) | ( n10280 & n10300 ) | ( n10297 & n10300 ) ;
  assign n10302 = n10297 | n10299 ;
  assign n10303 = n10280 | n10302 ;
  assign n10304 = ~n10301 & n10303 ;
  assign n10305 = n9848 | n9852 ;
  assign n10306 = ( n9848 & n9851 ) | ( n9848 & n10305 ) | ( n9851 & n10305 ) ;
  assign n10307 = n10304 | n10306 ;
  assign n10308 = n10304 & n10306 ;
  assign n10309 = n10307 & ~n10308 ;
  assign n10310 = x109 | x110 ;
  assign n10311 = x109 & x110 ;
  assign n10312 = n10310 & ~n10311 ;
  assign n10313 = n9857 & n10312 ;
  assign n10314 = ( n9862 & n10312 ) | ( n9862 & n10313 ) | ( n10312 & n10313 ) ;
  assign n10315 = ( n9863 & n10312 ) | ( n9863 & n10313 ) | ( n10312 & n10313 ) ;
  assign n10316 = ( n8261 & n10314 ) | ( n8261 & n10315 ) | ( n10314 & n10315 ) ;
  assign n10317 = ( n8262 & n10314 ) | ( n8262 & n10315 ) | ( n10314 & n10315 ) ;
  assign n10318 = ( n6159 & n10316 ) | ( n6159 & n10317 ) | ( n10316 & n10317 ) ;
  assign n10319 = ( n6157 & n10316 ) | ( n6157 & n10317 ) | ( n10316 & n10317 ) ;
  assign n10320 = ( n5823 & n10318 ) | ( n5823 & n10319 ) | ( n10318 & n10319 ) ;
  assign n10321 = n9857 | n9862 ;
  assign n10322 = n9857 | n9863 ;
  assign n10323 = ( n8262 & n10321 ) | ( n8262 & n10322 ) | ( n10321 & n10322 ) ;
  assign n10324 = n10312 | n10323 ;
  assign n10325 = ( n8261 & n10321 ) | ( n8261 & n10322 ) | ( n10321 & n10322 ) ;
  assign n10326 = n10312 | n10325 ;
  assign n10327 = ( n6159 & n10324 ) | ( n6159 & n10326 ) | ( n10324 & n10326 ) ;
  assign n10328 = ( n6157 & n10324 ) | ( n6157 & n10326 ) | ( n10324 & n10326 ) ;
  assign n10329 = ( n5823 & n10327 ) | ( n5823 & n10328 ) | ( n10327 & n10328 ) ;
  assign n10330 = ~n10320 & n10329 ;
  assign n10331 = x109 & n133 ;
  assign n10332 = x108 & ~n162 ;
  assign n10333 = ( n137 & n10331 ) | ( n137 & n10332 ) | ( n10331 & n10332 ) ;
  assign n10334 = x0 & x110 ;
  assign n10335 = ( ~n137 & n10331 ) | ( ~n137 & n10334 ) | ( n10331 & n10334 ) ;
  assign n10336 = n10333 | n10335 ;
  assign n10337 = n141 | n10336 ;
  assign n10338 = ( n10330 & n10336 ) | ( n10330 & n10337 ) | ( n10336 & n10337 ) ;
  assign n10339 = x2 & n10336 ;
  assign n10340 = ( x2 & n523 ) | ( x2 & n10336 ) | ( n523 & n10336 ) ;
  assign n10341 = ( n10330 & n10339 ) | ( n10330 & n10340 ) | ( n10339 & n10340 ) ;
  assign n10342 = x2 & ~n10340 ;
  assign n10343 = x2 & ~n10336 ;
  assign n10344 = ( ~n10330 & n10342 ) | ( ~n10330 & n10343 ) | ( n10342 & n10343 ) ;
  assign n10345 = ( n10338 & ~n10341 ) | ( n10338 & n10344 ) | ( ~n10341 & n10344 ) ;
  assign n10346 = n10309 & n10345 ;
  assign n10347 = n10309 & ~n10346 ;
  assign n10348 = ~n10309 & n10345 ;
  assign n10349 = n10347 | n10348 ;
  assign n10350 = n9895 | n9899 ;
  assign n10351 = ( n9895 & n9896 ) | ( n9895 & n10350 ) | ( n9896 & n10350 ) ;
  assign n10352 = n10349 & n10351 ;
  assign n10353 = n10349 | n10351 ;
  assign n10354 = ~n10352 & n10353 ;
  assign n10355 = n10191 | n10195 ;
  assign n10356 = n10128 | n10134 ;
  assign n10357 = ( n10128 & n10131 ) | ( n10128 & n10356 ) | ( n10131 & n10356 ) ;
  assign n10358 = n10069 | n10084 ;
  assign n10359 = x75 & n6536 ;
  assign n10360 = x74 & n6531 ;
  assign n10361 = x73 & ~n6530 ;
  assign n10362 = n6871 & n10361 ;
  assign n10363 = n10360 | n10362 ;
  assign n10364 = n10359 | n10363 ;
  assign n10365 = n6539 | n10359 ;
  assign n10366 = n10363 | n10365 ;
  assign n10367 = ( n746 & n10364 ) | ( n746 & n10366 ) | ( n10364 & n10366 ) ;
  assign n10368 = x38 & n10366 ;
  assign n10369 = x38 & n10359 ;
  assign n10370 = ( x38 & n10363 ) | ( x38 & n10369 ) | ( n10363 & n10369 ) ;
  assign n10371 = ( n746 & n10368 ) | ( n746 & n10370 ) | ( n10368 & n10370 ) ;
  assign n10372 = x38 & ~n10370 ;
  assign n10373 = x38 & ~n10366 ;
  assign n10374 = ( ~n746 & n10372 ) | ( ~n746 & n10373 ) | ( n10372 & n10373 ) ;
  assign n10375 = ( n10367 & ~n10371 ) | ( n10367 & n10374 ) | ( ~n10371 & n10374 ) ;
  assign n10376 = n9992 | n9999 ;
  assign n10377 = x66 & n9933 ;
  assign n10378 = x65 & n9928 ;
  assign n10379 = ~n9503 & n9932 ;
  assign n10380 = x64 & ~n9927 ;
  assign n10381 = n10379 & n10380 ;
  assign n10382 = n10378 | n10381 ;
  assign n10383 = n10377 | n10382 ;
  assign n10384 = n159 & n9936 ;
  assign n10385 = n10383 | n10384 ;
  assign n10386 = x47 | n9936 ;
  assign n10387 = ( x47 & n159 ) | ( x47 & n10386 ) | ( n159 & n10386 ) ;
  assign n10388 = n10383 | n10387 ;
  assign n10389 = ~x47 & n10387 ;
  assign n10390 = ( ~x47 & n10383 ) | ( ~x47 & n10389 ) | ( n10383 & n10389 ) ;
  assign n10391 = ( ~n10385 & n10388 ) | ( ~n10385 & n10390 ) | ( n10388 & n10390 ) ;
  assign n10392 = n9948 | n10391 ;
  assign n10393 = n9948 & n10391 ;
  assign n10394 = n10392 & ~n10393 ;
  assign n10395 = n293 & n8727 ;
  assign n10396 = x69 & n8724 ;
  assign n10397 = x68 & n8719 ;
  assign n10398 = x67 & ~n8718 ;
  assign n10399 = n9149 & n10398 ;
  assign n10400 = n10397 | n10399 ;
  assign n10401 = n10396 | n10400 ;
  assign n10402 = n10395 | n10401 ;
  assign n10403 = x44 | n10396 ;
  assign n10404 = n10400 | n10403 ;
  assign n10405 = n10395 | n10404 ;
  assign n10406 = ~x44 & n10404 ;
  assign n10407 = ( ~x44 & n10395 ) | ( ~x44 & n10406 ) | ( n10395 & n10406 ) ;
  assign n10408 = ( ~n10402 & n10405 ) | ( ~n10402 & n10407 ) | ( n10405 & n10407 ) ;
  assign n10409 = n10394 & n10408 ;
  assign n10410 = n10394 & ~n10409 ;
  assign n10411 = ~n10394 & n10408 ;
  assign n10412 = n10410 | n10411 ;
  assign n10413 = n9970 | n9972 ;
  assign n10414 = ( n9970 & n9971 ) | ( n9970 & n10413 ) | ( n9971 & n10413 ) ;
  assign n10415 = n10412 & n10414 ;
  assign n10416 = n10412 | n10414 ;
  assign n10417 = ~n10415 & n10416 ;
  assign n10418 = x72 & n7566 ;
  assign n10419 = x71 & n7561 ;
  assign n10420 = x70 & ~n7560 ;
  assign n10421 = n7953 & n10420 ;
  assign n10422 = n10419 | n10421 ;
  assign n10423 = n10418 | n10422 ;
  assign n10424 = ( n513 & n7569 ) | ( n513 & n10423 ) | ( n7569 & n10423 ) ;
  assign n10425 = ( x41 & n7569 ) | ( x41 & ~n10418 ) | ( n7569 & ~n10418 ) ;
  assign n10426 = x41 & n7569 ;
  assign n10427 = ( ~n10422 & n10425 ) | ( ~n10422 & n10426 ) | ( n10425 & n10426 ) ;
  assign n10428 = ( x41 & n513 ) | ( x41 & n10427 ) | ( n513 & n10427 ) ;
  assign n10429 = ~n10424 & n10428 ;
  assign n10430 = n10423 | n10427 ;
  assign n10431 = x41 | n10423 ;
  assign n10432 = ( n513 & n10430 ) | ( n513 & n10431 ) | ( n10430 & n10431 ) ;
  assign n10433 = ( ~x41 & n10429 ) | ( ~x41 & n10432 ) | ( n10429 & n10432 ) ;
  assign n10434 = n10417 & n10433 ;
  assign n10435 = n10417 & ~n10434 ;
  assign n10436 = ~n10417 & n10433 ;
  assign n10437 = n10435 | n10436 ;
  assign n10438 = ~n10376 & n10437 ;
  assign n10439 = n10375 & n10438 ;
  assign n10440 = n10376 & ~n10437 ;
  assign n10441 = ( n10375 & n10439 ) | ( n10375 & n10440 ) | ( n10439 & n10440 ) ;
  assign n10442 = n10375 | n10438 ;
  assign n10443 = n10440 | n10442 ;
  assign n10444 = ~n10441 & n10443 ;
  assign n10445 = n10018 | n10019 ;
  assign n10446 = ( n9924 & n10018 ) | ( n9924 & n10445 ) | ( n10018 & n10445 ) ;
  assign n10447 = n10444 & n10446 ;
  assign n10448 = n10444 | n10446 ;
  assign n10449 = ~n10447 & n10448 ;
  assign n10450 = x78 & n5554 ;
  assign n10451 = x77 & n5549 ;
  assign n10452 = x76 & ~n5548 ;
  assign n10453 = n5893 & n10452 ;
  assign n10454 = n10451 | n10453 ;
  assign n10455 = n10450 | n10454 ;
  assign n10456 = n5557 | n10450 ;
  assign n10457 = n10454 | n10456 ;
  assign n10458 = ( n1192 & n10455 ) | ( n1192 & n10457 ) | ( n10455 & n10457 ) ;
  assign n10459 = x35 & n10457 ;
  assign n10460 = x35 & n10450 ;
  assign n10461 = ( x35 & n10454 ) | ( x35 & n10460 ) | ( n10454 & n10460 ) ;
  assign n10462 = ( n1192 & n10459 ) | ( n1192 & n10461 ) | ( n10459 & n10461 ) ;
  assign n10463 = x35 & ~n10461 ;
  assign n10464 = x35 & ~n10457 ;
  assign n10465 = ( ~n1192 & n10463 ) | ( ~n1192 & n10464 ) | ( n10463 & n10464 ) ;
  assign n10466 = ( n10458 & ~n10462 ) | ( n10458 & n10465 ) | ( ~n10462 & n10465 ) ;
  assign n10467 = n10449 & n10466 ;
  assign n10468 = n10449 & ~n10467 ;
  assign n10469 = ~n10449 & n10466 ;
  assign n10470 = n10468 | n10469 ;
  assign n10471 = n10043 | n10046 ;
  assign n10472 = ( n10043 & n10048 ) | ( n10043 & n10471 ) | ( n10048 & n10471 ) ;
  assign n10473 = n10470 & n10472 ;
  assign n10474 = n10470 | n10472 ;
  assign n10475 = ~n10473 & n10474 ;
  assign n10476 = x81 & n4631 ;
  assign n10477 = x80 & n4626 ;
  assign n10478 = x79 & ~n4625 ;
  assign n10479 = n4943 & n10478 ;
  assign n10480 = n10477 | n10479 ;
  assign n10481 = n10476 | n10480 ;
  assign n10482 = n4634 | n10476 ;
  assign n10483 = n10480 | n10482 ;
  assign n10484 = ( n1651 & n10481 ) | ( n1651 & n10483 ) | ( n10481 & n10483 ) ;
  assign n10485 = x32 & n10483 ;
  assign n10486 = x32 & n10476 ;
  assign n10487 = ( x32 & n10480 ) | ( x32 & n10486 ) | ( n10480 & n10486 ) ;
  assign n10488 = ( n1651 & n10485 ) | ( n1651 & n10487 ) | ( n10485 & n10487 ) ;
  assign n10489 = x32 & ~n10487 ;
  assign n10490 = x32 & ~n10483 ;
  assign n10491 = ( ~n1651 & n10489 ) | ( ~n1651 & n10490 ) | ( n10489 & n10490 ) ;
  assign n10492 = ( n10484 & ~n10488 ) | ( n10484 & n10491 ) | ( ~n10488 & n10491 ) ;
  assign n10493 = n10475 & n10492 ;
  assign n10494 = n10475 & ~n10493 ;
  assign n10495 = ~n10475 & n10492 ;
  assign n10496 = n10494 | n10495 ;
  assign n10497 = ~n10358 & n10496 ;
  assign n10498 = n10358 & ~n10496 ;
  assign n10499 = n10497 | n10498 ;
  assign n10500 = x84 & n3816 ;
  assign n10501 = x83 & n3811 ;
  assign n10502 = x82 & ~n3810 ;
  assign n10503 = n4067 & n10502 ;
  assign n10504 = n10501 | n10503 ;
  assign n10505 = n10500 | n10504 ;
  assign n10506 = n3819 | n10500 ;
  assign n10507 = n10504 | n10506 ;
  assign n10508 = ( n2194 & n10505 ) | ( n2194 & n10507 ) | ( n10505 & n10507 ) ;
  assign n10509 = x29 & n10507 ;
  assign n10510 = x29 & n10500 ;
  assign n10511 = ( x29 & n10504 ) | ( x29 & n10510 ) | ( n10504 & n10510 ) ;
  assign n10512 = ( n2194 & n10509 ) | ( n2194 & n10511 ) | ( n10509 & n10511 ) ;
  assign n10513 = x29 & ~n10511 ;
  assign n10514 = x29 & ~n10507 ;
  assign n10515 = ( ~n2194 & n10513 ) | ( ~n2194 & n10514 ) | ( n10513 & n10514 ) ;
  assign n10516 = ( n10508 & ~n10512 ) | ( n10508 & n10515 ) | ( ~n10512 & n10515 ) ;
  assign n10517 = n10499 & n10516 ;
  assign n10518 = n10499 | n10516 ;
  assign n10519 = ~n10517 & n10518 ;
  assign n10520 = n10103 | n10107 ;
  assign n10521 = ( n10103 & n10106 ) | ( n10103 & n10520 ) | ( n10106 & n10520 ) ;
  assign n10522 = n10519 | n10521 ;
  assign n10523 = n10519 & n10521 ;
  assign n10524 = n10522 & ~n10523 ;
  assign n10525 = x87 & n3085 ;
  assign n10526 = x86 & n3080 ;
  assign n10527 = x85 & ~n3079 ;
  assign n10528 = n3309 & n10527 ;
  assign n10529 = n10526 | n10528 ;
  assign n10530 = n10525 | n10529 ;
  assign n10531 = n3088 | n10525 ;
  assign n10532 = n10529 | n10531 ;
  assign n10533 = ( n2816 & n10530 ) | ( n2816 & n10532 ) | ( n10530 & n10532 ) ;
  assign n10534 = x26 & n10532 ;
  assign n10535 = x26 & n10525 ;
  assign n10536 = ( x26 & n10529 ) | ( x26 & n10535 ) | ( n10529 & n10535 ) ;
  assign n10537 = ( n2816 & n10534 ) | ( n2816 & n10536 ) | ( n10534 & n10536 ) ;
  assign n10538 = x26 & ~n10536 ;
  assign n10539 = x26 & ~n10532 ;
  assign n10540 = ( ~n2816 & n10538 ) | ( ~n2816 & n10539 ) | ( n10538 & n10539 ) ;
  assign n10541 = ( n10533 & ~n10537 ) | ( n10533 & n10540 ) | ( ~n10537 & n10540 ) ;
  assign n10542 = n10524 & n10541 ;
  assign n10543 = n10524 | n10541 ;
  assign n10544 = ~n10542 & n10543 ;
  assign n10545 = n10357 & n10544 ;
  assign n10546 = n10357 & ~n10545 ;
  assign n10547 = x90 & n2429 ;
  assign n10548 = x89 & n2424 ;
  assign n10549 = x88 & ~n2423 ;
  assign n10550 = n2631 & n10549 ;
  assign n10551 = n10548 | n10550 ;
  assign n10552 = n10547 | n10551 ;
  assign n10553 = n2432 | n10547 ;
  assign n10554 = n10551 | n10553 ;
  assign n10555 = ( n3519 & n10552 ) | ( n3519 & n10554 ) | ( n10552 & n10554 ) ;
  assign n10556 = x23 & n10554 ;
  assign n10557 = x23 & n10547 ;
  assign n10558 = ( x23 & n10551 ) | ( x23 & n10557 ) | ( n10551 & n10557 ) ;
  assign n10559 = ( n3519 & n10556 ) | ( n3519 & n10558 ) | ( n10556 & n10558 ) ;
  assign n10560 = x23 & ~n10558 ;
  assign n10561 = x23 & ~n10554 ;
  assign n10562 = ( ~n3519 & n10560 ) | ( ~n3519 & n10561 ) | ( n10560 & n10561 ) ;
  assign n10563 = ( n10555 & ~n10559 ) | ( n10555 & n10562 ) | ( ~n10559 & n10562 ) ;
  assign n10564 = ~n10543 & n10544 ;
  assign n10565 = ( ~n10357 & n10544 ) | ( ~n10357 & n10564 ) | ( n10544 & n10564 ) ;
  assign n10566 = n10563 & n10565 ;
  assign n10567 = ( n10546 & n10563 ) | ( n10546 & n10566 ) | ( n10563 & n10566 ) ;
  assign n10568 = n10563 | n10565 ;
  assign n10569 = n10546 | n10568 ;
  assign n10570 = ~n10567 & n10569 ;
  assign n10571 = n10155 | n10159 ;
  assign n10572 = ( n10155 & n10158 ) | ( n10155 & n10571 ) | ( n10158 & n10571 ) ;
  assign n10573 = n10570 & n10572 ;
  assign n10574 = n10570 | n10572 ;
  assign n10575 = ~n10573 & n10574 ;
  assign n10576 = x93 & n1859 ;
  assign n10577 = x92 & n1854 ;
  assign n10578 = x91 & ~n1853 ;
  assign n10579 = n2037 & n10578 ;
  assign n10580 = n10577 | n10579 ;
  assign n10581 = n10576 | n10580 ;
  assign n10582 = n1862 | n10576 ;
  assign n10583 = n10580 | n10582 ;
  assign n10584 = ( n4305 & n10581 ) | ( n4305 & n10583 ) | ( n10581 & n10583 ) ;
  assign n10585 = x20 & n10583 ;
  assign n10586 = x20 & n10576 ;
  assign n10587 = ( x20 & n10580 ) | ( x20 & n10586 ) | ( n10580 & n10586 ) ;
  assign n10588 = ( n4305 & n10585 ) | ( n4305 & n10587 ) | ( n10585 & n10587 ) ;
  assign n10589 = x20 & ~n10587 ;
  assign n10590 = x20 & ~n10583 ;
  assign n10591 = ( ~n4305 & n10589 ) | ( ~n4305 & n10590 ) | ( n10589 & n10590 ) ;
  assign n10592 = ( n10584 & ~n10588 ) | ( n10584 & n10591 ) | ( ~n10588 & n10591 ) ;
  assign n10593 = n10575 | n10592 ;
  assign n10594 = n10575 & n10592 ;
  assign n10595 = n10593 & ~n10594 ;
  assign n10596 = n10182 & n10185 ;
  assign n10597 = ( n10181 & n10185 ) | ( n10181 & n10596 ) | ( n10185 & n10596 ) ;
  assign n10598 = n10180 | n10597 ;
  assign n10599 = n10595 & n10598 ;
  assign n10600 = n10595 | n10598 ;
  assign n10601 = ~n10599 & n10600 ;
  assign n10602 = x96 & n1383 ;
  assign n10603 = x95 & n1378 ;
  assign n10604 = x94 & ~n1377 ;
  assign n10605 = n1542 & n10604 ;
  assign n10606 = n10603 | n10605 ;
  assign n10607 = n10602 | n10606 ;
  assign n10608 = n1386 | n10602 ;
  assign n10609 = n10606 | n10608 ;
  assign n10610 = ( n5202 & n10607 ) | ( n5202 & n10609 ) | ( n10607 & n10609 ) ;
  assign n10611 = x17 & n10609 ;
  assign n10612 = x17 & n10602 ;
  assign n10613 = ( x17 & n10606 ) | ( x17 & n10612 ) | ( n10606 & n10612 ) ;
  assign n10614 = ( n5202 & n10611 ) | ( n5202 & n10613 ) | ( n10611 & n10613 ) ;
  assign n10615 = x17 & ~n10613 ;
  assign n10616 = x17 & ~n10609 ;
  assign n10617 = ( ~n5202 & n10615 ) | ( ~n5202 & n10616 ) | ( n10615 & n10616 ) ;
  assign n10618 = ( n10610 & ~n10614 ) | ( n10610 & n10617 ) | ( ~n10614 & n10617 ) ;
  assign n10619 = n10601 | n10618 ;
  assign n10620 = n10601 & n10618 ;
  assign n10621 = n10619 & ~n10620 ;
  assign n10622 = n10355 & n10621 ;
  assign n10623 = n10355 | n10621 ;
  assign n10624 = ~n10622 & n10623 ;
  assign n10625 = x99 & n962 ;
  assign n10626 = x98 & n957 ;
  assign n10627 = x97 & ~n956 ;
  assign n10628 = n1105 & n10627 ;
  assign n10629 = n10626 | n10628 ;
  assign n10630 = n10625 | n10629 ;
  assign n10631 = n965 | n10625 ;
  assign n10632 = n10629 | n10631 ;
  assign n10633 = ( n6164 & n10630 ) | ( n6164 & n10632 ) | ( n10630 & n10632 ) ;
  assign n10634 = x14 & n10632 ;
  assign n10635 = x14 & n10625 ;
  assign n10636 = ( x14 & n10629 ) | ( x14 & n10635 ) | ( n10629 & n10635 ) ;
  assign n10637 = ( n6164 & n10634 ) | ( n6164 & n10636 ) | ( n10634 & n10636 ) ;
  assign n10638 = x14 & ~n10636 ;
  assign n10639 = x14 & ~n10632 ;
  assign n10640 = ( ~n6164 & n10638 ) | ( ~n6164 & n10639 ) | ( n10638 & n10639 ) ;
  assign n10641 = ( n10633 & ~n10637 ) | ( n10633 & n10640 ) | ( ~n10637 & n10640 ) ;
  assign n10642 = n10624 & n10641 ;
  assign n10643 = n10624 & ~n10642 ;
  assign n10644 = ~n10624 & n10641 ;
  assign n10645 = n10643 | n10644 ;
  assign n10646 = n10221 | n10228 ;
  assign n10647 = n10645 | n10646 ;
  assign n10648 = n10645 & n10646 ;
  assign n10649 = n10647 & ~n10648 ;
  assign n10650 = x102 & n636 ;
  assign n10651 = x101 & n631 ;
  assign n10652 = x100 & ~n630 ;
  assign n10653 = n764 & n10652 ;
  assign n10654 = n10651 | n10653 ;
  assign n10655 = n10650 | n10654 ;
  assign n10656 = n639 | n10650 ;
  assign n10657 = n10654 | n10656 ;
  assign n10658 = ( n7178 & n10655 ) | ( n7178 & n10657 ) | ( n10655 & n10657 ) ;
  assign n10659 = x11 & n10657 ;
  assign n10660 = x11 & n10650 ;
  assign n10661 = ( x11 & n10654 ) | ( x11 & n10660 ) | ( n10654 & n10660 ) ;
  assign n10662 = ( n7178 & n10659 ) | ( n7178 & n10661 ) | ( n10659 & n10661 ) ;
  assign n10663 = x11 & ~n10661 ;
  assign n10664 = x11 & ~n10657 ;
  assign n10665 = ( ~n7178 & n10663 ) | ( ~n7178 & n10664 ) | ( n10663 & n10664 ) ;
  assign n10666 = ( n10658 & ~n10662 ) | ( n10658 & n10665 ) | ( ~n10662 & n10665 ) ;
  assign n10667 = n10649 & n10666 ;
  assign n10668 = n10649 & ~n10667 ;
  assign n10669 = ~n10649 & n10666 ;
  assign n10670 = n10668 | n10669 ;
  assign n10671 = n10249 | n10257 ;
  assign n10672 = n10670 | n10671 ;
  assign n10673 = n10670 & n10671 ;
  assign n10674 = n10672 & ~n10673 ;
  assign n10675 = x105 & n389 ;
  assign n10676 = x104 & n384 ;
  assign n10677 = x103 & ~n383 ;
  assign n10678 = n463 & n10677 ;
  assign n10679 = n10676 | n10678 ;
  assign n10680 = n10675 | n10679 ;
  assign n10681 = n392 | n10675 ;
  assign n10682 = n10679 | n10681 ;
  assign n10683 = ( n8273 & n10680 ) | ( n8273 & n10682 ) | ( n10680 & n10682 ) ;
  assign n10684 = x8 & n10682 ;
  assign n10685 = x8 & n10675 ;
  assign n10686 = ( x8 & n10679 ) | ( x8 & n10685 ) | ( n10679 & n10685 ) ;
  assign n10687 = ( n8273 & n10684 ) | ( n8273 & n10686 ) | ( n10684 & n10686 ) ;
  assign n10688 = x8 & ~n10686 ;
  assign n10689 = x8 & ~n10682 ;
  assign n10690 = ( ~n8273 & n10688 ) | ( ~n8273 & n10689 ) | ( n10688 & n10689 ) ;
  assign n10691 = ( n10683 & ~n10687 ) | ( n10683 & n10690 ) | ( ~n10687 & n10690 ) ;
  assign n10692 = n10674 & n10691 ;
  assign n10693 = n10674 | n10691 ;
  assign n10694 = ~n10692 & n10693 ;
  assign n10695 = n10276 | n10277 ;
  assign n10696 = ( n9904 & n10276 ) | ( n9904 & n10695 ) | ( n10276 & n10695 ) ;
  assign n10697 = n10694 & n10696 ;
  assign n10698 = ~n10694 & n10696 ;
  assign n10699 = ( n10694 & ~n10697 ) | ( n10694 & n10698 ) | ( ~n10697 & n10698 ) ;
  assign n10700 = x108 & n212 ;
  assign n10701 = x107 & n207 ;
  assign n10702 = x106 & ~n206 ;
  assign n10703 = n267 & n10702 ;
  assign n10704 = n10701 | n10703 ;
  assign n10705 = n10700 | n10704 ;
  assign n10706 = n215 | n10700 ;
  assign n10707 = n10704 | n10706 ;
  assign n10708 = ( n9479 & n10705 ) | ( n9479 & n10707 ) | ( n10705 & n10707 ) ;
  assign n10709 = x5 & n10707 ;
  assign n10710 = x5 & n10700 ;
  assign n10711 = ( x5 & n10704 ) | ( x5 & n10710 ) | ( n10704 & n10710 ) ;
  assign n10712 = ( n9479 & n10709 ) | ( n9479 & n10711 ) | ( n10709 & n10711 ) ;
  assign n10713 = x5 & ~n10711 ;
  assign n10714 = x5 & ~n10707 ;
  assign n10715 = ( ~n9479 & n10713 ) | ( ~n9479 & n10714 ) | ( n10713 & n10714 ) ;
  assign n10716 = ( n10708 & ~n10712 ) | ( n10708 & n10715 ) | ( ~n10712 & n10715 ) ;
  assign n10717 = n10699 | n10716 ;
  assign n10718 = n10699 & n10716 ;
  assign n10719 = n10717 & ~n10718 ;
  assign n10720 = n10301 | n10304 ;
  assign n10721 = ( n10301 & n10306 ) | ( n10301 & n10720 ) | ( n10306 & n10720 ) ;
  assign n10722 = n10719 & n10721 ;
  assign n10723 = n10719 | n10721 ;
  assign n10724 = ~n10722 & n10723 ;
  assign n10725 = x110 | x111 ;
  assign n10726 = x110 & x111 ;
  assign n10727 = n10725 & ~n10726 ;
  assign n10728 = n9857 | n10311 ;
  assign n10729 = ( n10311 & n10312 ) | ( n10311 & n10728 ) | ( n10312 & n10728 ) ;
  assign n10730 = n10727 & n10729 ;
  assign n10731 = n10311 | n10312 ;
  assign n10732 = n10727 & n10731 ;
  assign n10733 = ( n9862 & n10730 ) | ( n9862 & n10732 ) | ( n10730 & n10732 ) ;
  assign n10734 = ( n9863 & n10730 ) | ( n9863 & n10732 ) | ( n10730 & n10732 ) ;
  assign n10735 = ( n8261 & n10733 ) | ( n8261 & n10734 ) | ( n10733 & n10734 ) ;
  assign n10736 = ( n8262 & n10733 ) | ( n8262 & n10734 ) | ( n10733 & n10734 ) ;
  assign n10737 = ( n6159 & n10735 ) | ( n6159 & n10736 ) | ( n10735 & n10736 ) ;
  assign n10738 = ( n6157 & n10735 ) | ( n6157 & n10736 ) | ( n10735 & n10736 ) ;
  assign n10739 = ( n5823 & n10737 ) | ( n5823 & n10738 ) | ( n10737 & n10738 ) ;
  assign n10740 = ( n9862 & n10729 ) | ( n9862 & n10731 ) | ( n10729 & n10731 ) ;
  assign n10741 = ( n9863 & n10729 ) | ( n9863 & n10731 ) | ( n10729 & n10731 ) ;
  assign n10742 = ( n8262 & n10740 ) | ( n8262 & n10741 ) | ( n10740 & n10741 ) ;
  assign n10743 = n10727 | n10742 ;
  assign n10744 = ( n8261 & n10740 ) | ( n8261 & n10741 ) | ( n10740 & n10741 ) ;
  assign n10745 = n10727 | n10744 ;
  assign n10746 = ( n6159 & n10743 ) | ( n6159 & n10745 ) | ( n10743 & n10745 ) ;
  assign n10747 = ( n6157 & n10743 ) | ( n6157 & n10745 ) | ( n10743 & n10745 ) ;
  assign n10748 = ( n5823 & n10746 ) | ( n5823 & n10747 ) | ( n10746 & n10747 ) ;
  assign n10749 = ~n10739 & n10748 ;
  assign n10750 = x110 & n133 ;
  assign n10751 = x109 & ~n162 ;
  assign n10752 = ( n137 & n10750 ) | ( n137 & n10751 ) | ( n10750 & n10751 ) ;
  assign n10753 = x0 & x111 ;
  assign n10754 = ( ~n137 & n10750 ) | ( ~n137 & n10753 ) | ( n10750 & n10753 ) ;
  assign n10755 = n10752 | n10754 ;
  assign n10756 = n141 | n10755 ;
  assign n10757 = ( n10749 & n10755 ) | ( n10749 & n10756 ) | ( n10755 & n10756 ) ;
  assign n10758 = x2 & n10755 ;
  assign n10759 = ( x2 & n523 ) | ( x2 & n10755 ) | ( n523 & n10755 ) ;
  assign n10760 = ( n10749 & n10758 ) | ( n10749 & n10759 ) | ( n10758 & n10759 ) ;
  assign n10761 = x2 & ~n10759 ;
  assign n10762 = x2 & ~n10755 ;
  assign n10763 = ( ~n10749 & n10761 ) | ( ~n10749 & n10762 ) | ( n10761 & n10762 ) ;
  assign n10764 = ( n10757 & ~n10760 ) | ( n10757 & n10763 ) | ( ~n10760 & n10763 ) ;
  assign n10765 = n10724 & n10764 ;
  assign n10766 = n10724 & ~n10765 ;
  assign n10767 = ~n10724 & n10764 ;
  assign n10768 = n10766 | n10767 ;
  assign n10769 = n10346 | n10351 ;
  assign n10770 = ( n10346 & n10349 ) | ( n10346 & n10769 ) | ( n10349 & n10769 ) ;
  assign n10771 = n10768 & n10770 ;
  assign n10772 = n10768 | n10770 ;
  assign n10773 = ~n10771 & n10772 ;
  assign n10774 = n10765 | n10771 ;
  assign n10775 = n10467 | n10473 ;
  assign n10776 = n10441 | n10447 ;
  assign n10777 = x47 & ~x48 ;
  assign n10778 = ~x47 & x48 ;
  assign n10779 = n10777 | n10778 ;
  assign n10780 = x64 & n10779 ;
  assign n10781 = ~n9948 & n10780 ;
  assign n10782 = ( ~n10391 & n10780 ) | ( ~n10391 & n10781 ) | ( n10780 & n10781 ) ;
  assign n10783 = n9948 & ~n10780 ;
  assign n10784 = n10391 & n10783 ;
  assign n10785 = n10782 | n10784 ;
  assign n10786 = x67 & n9933 ;
  assign n10787 = x66 & n9928 ;
  assign n10788 = x65 & ~n9927 ;
  assign n10789 = n10379 & n10788 ;
  assign n10790 = n10787 | n10789 ;
  assign n10791 = n10786 | n10790 ;
  assign n10792 = n186 & n9936 ;
  assign n10793 = n10791 | n10792 ;
  assign n10794 = x47 & ~n10793 ;
  assign n10795 = ~x47 & n10793 ;
  assign n10796 = n10794 | n10795 ;
  assign n10797 = n10785 & n10796 ;
  assign n10798 = n10785 | n10796 ;
  assign n10799 = ~n10797 & n10798 ;
  assign n10800 = x69 & n8719 ;
  assign n10801 = x68 & ~n8718 ;
  assign n10802 = n9149 & n10801 ;
  assign n10803 = n10800 | n10802 ;
  assign n10804 = x70 & n8724 ;
  assign n10805 = n8727 | n10804 ;
  assign n10806 = n10803 | n10805 ;
  assign n10807 = x44 & ~n10806 ;
  assign n10808 = x44 & ~n10804 ;
  assign n10809 = ~n10803 & n10808 ;
  assign n10810 = ( ~n340 & n10807 ) | ( ~n340 & n10809 ) | ( n10807 & n10809 ) ;
  assign n10811 = ~x44 & n10806 ;
  assign n10812 = ~x44 & n10804 ;
  assign n10813 = ( ~x44 & n10803 ) | ( ~x44 & n10812 ) | ( n10803 & n10812 ) ;
  assign n10814 = ( n340 & n10811 ) | ( n340 & n10813 ) | ( n10811 & n10813 ) ;
  assign n10815 = n10810 | n10814 ;
  assign n10816 = n10799 & n10815 ;
  assign n10817 = n10799 & ~n10816 ;
  assign n10818 = ~n10799 & n10815 ;
  assign n10819 = n10817 | n10818 ;
  assign n10820 = n10409 | n10414 ;
  assign n10821 = ( n10409 & n10412 ) | ( n10409 & n10820 ) | ( n10412 & n10820 ) ;
  assign n10822 = n10819 | n10821 ;
  assign n10823 = n10819 & n10821 ;
  assign n10824 = n10822 & ~n10823 ;
  assign n10825 = x73 & n7566 ;
  assign n10826 = x72 & n7561 ;
  assign n10827 = x71 & ~n7560 ;
  assign n10828 = n7953 & n10827 ;
  assign n10829 = n10826 | n10828 ;
  assign n10830 = n10825 | n10829 ;
  assign n10831 = ( ~n610 & n7569 ) | ( ~n610 & n10830 ) | ( n7569 & n10830 ) ;
  assign n10832 = n7569 & n10825 ;
  assign n10833 = ( n7569 & n10829 ) | ( n7569 & n10832 ) | ( n10829 & n10832 ) ;
  assign n10834 = ( n598 & n10831 ) | ( n598 & n10833 ) | ( n10831 & n10833 ) ;
  assign n10835 = ( x41 & ~n10830 ) | ( x41 & n10834 ) | ( ~n10830 & n10834 ) ;
  assign n10836 = ~n10834 & n10835 ;
  assign n10837 = x41 | n10825 ;
  assign n10838 = n10829 | n10837 ;
  assign n10839 = n10834 | n10838 ;
  assign n10840 = ( ~x41 & n10836 ) | ( ~x41 & n10839 ) | ( n10836 & n10839 ) ;
  assign n10841 = n10824 | n10840 ;
  assign n10842 = n10824 & n10840 ;
  assign n10843 = n10841 & ~n10842 ;
  assign n10844 = n10376 & n10437 ;
  assign n10845 = n10434 | n10844 ;
  assign n10846 = n10843 & n10845 ;
  assign n10847 = n10843 | n10845 ;
  assign n10848 = ~n10846 & n10847 ;
  assign n10849 = x76 & n6536 ;
  assign n10850 = x75 & n6531 ;
  assign n10851 = x74 & ~n6530 ;
  assign n10852 = n6871 & n10851 ;
  assign n10853 = n10850 | n10852 ;
  assign n10854 = n10849 | n10853 ;
  assign n10855 = n6539 | n10849 ;
  assign n10856 = n10853 | n10855 ;
  assign n10857 = ( n923 & n10854 ) | ( n923 & n10856 ) | ( n10854 & n10856 ) ;
  assign n10858 = x38 & n10856 ;
  assign n10859 = x38 & n10849 ;
  assign n10860 = ( x38 & n10853 ) | ( x38 & n10859 ) | ( n10853 & n10859 ) ;
  assign n10861 = ( n923 & n10858 ) | ( n923 & n10860 ) | ( n10858 & n10860 ) ;
  assign n10862 = x38 & ~n10860 ;
  assign n10863 = x38 & ~n10856 ;
  assign n10864 = ( ~n923 & n10862 ) | ( ~n923 & n10863 ) | ( n10862 & n10863 ) ;
  assign n10865 = ( n10857 & ~n10861 ) | ( n10857 & n10864 ) | ( ~n10861 & n10864 ) ;
  assign n10866 = n10848 & n10865 ;
  assign n10867 = n10848 & ~n10866 ;
  assign n10868 = ~n10848 & n10865 ;
  assign n10869 = n10867 | n10868 ;
  assign n10870 = n10776 & n10869 ;
  assign n10871 = n10776 | n10869 ;
  assign n10872 = ~n10870 & n10871 ;
  assign n10873 = x79 & n5554 ;
  assign n10874 = x78 & n5549 ;
  assign n10875 = x77 & ~n5548 ;
  assign n10876 = n5893 & n10875 ;
  assign n10877 = n10874 | n10876 ;
  assign n10878 = n10873 | n10877 ;
  assign n10879 = n5557 | n10873 ;
  assign n10880 = n10877 | n10879 ;
  assign n10881 = ( n1332 & n10878 ) | ( n1332 & n10880 ) | ( n10878 & n10880 ) ;
  assign n10882 = x35 & n10880 ;
  assign n10883 = x35 & n10873 ;
  assign n10884 = ( x35 & n10877 ) | ( x35 & n10883 ) | ( n10877 & n10883 ) ;
  assign n10885 = ( n1332 & n10882 ) | ( n1332 & n10884 ) | ( n10882 & n10884 ) ;
  assign n10886 = x35 & ~n10884 ;
  assign n10887 = x35 & ~n10880 ;
  assign n10888 = ( ~n1332 & n10886 ) | ( ~n1332 & n10887 ) | ( n10886 & n10887 ) ;
  assign n10889 = ( n10881 & ~n10885 ) | ( n10881 & n10888 ) | ( ~n10885 & n10888 ) ;
  assign n10890 = n10872 & n10889 ;
  assign n10891 = n10872 | n10889 ;
  assign n10892 = ~n10890 & n10891 ;
  assign n10893 = n10775 & n10892 ;
  assign n10894 = n10775 | n10892 ;
  assign n10895 = ~n10893 & n10894 ;
  assign n10896 = x82 & n4631 ;
  assign n10897 = x81 & n4626 ;
  assign n10898 = x80 & ~n4625 ;
  assign n10899 = n4943 & n10898 ;
  assign n10900 = n10897 | n10899 ;
  assign n10901 = n10896 | n10900 ;
  assign n10902 = n4634 | n10896 ;
  assign n10903 = n10900 | n10902 ;
  assign n10904 = ( n1811 & n10901 ) | ( n1811 & n10903 ) | ( n10901 & n10903 ) ;
  assign n10905 = x32 & n10903 ;
  assign n10906 = x32 & n10896 ;
  assign n10907 = ( x32 & n10900 ) | ( x32 & n10906 ) | ( n10900 & n10906 ) ;
  assign n10908 = ( n1811 & n10905 ) | ( n1811 & n10907 ) | ( n10905 & n10907 ) ;
  assign n10909 = x32 & ~n10907 ;
  assign n10910 = x32 & ~n10903 ;
  assign n10911 = ( ~n1811 & n10909 ) | ( ~n1811 & n10910 ) | ( n10909 & n10910 ) ;
  assign n10912 = ( n10904 & ~n10908 ) | ( n10904 & n10911 ) | ( ~n10908 & n10911 ) ;
  assign n10913 = n10895 & n10912 ;
  assign n10914 = n10895 & ~n10913 ;
  assign n10915 = ~n10895 & n10912 ;
  assign n10916 = n10914 | n10915 ;
  assign n10917 = n10493 | n10495 ;
  assign n10918 = n10494 | n10917 ;
  assign n10919 = ( n10358 & n10493 ) | ( n10358 & n10918 ) | ( n10493 & n10918 ) ;
  assign n10920 = n10916 | n10919 ;
  assign n10921 = n10916 & n10919 ;
  assign n10922 = n10920 & ~n10921 ;
  assign n10923 = x85 & n3816 ;
  assign n10924 = x84 & n3811 ;
  assign n10925 = x83 & ~n3810 ;
  assign n10926 = n4067 & n10925 ;
  assign n10927 = n10924 | n10926 ;
  assign n10928 = n10923 | n10927 ;
  assign n10929 = n3819 | n10923 ;
  assign n10930 = n10927 | n10929 ;
  assign n10931 = ( n2381 & n10928 ) | ( n2381 & n10930 ) | ( n10928 & n10930 ) ;
  assign n10932 = x29 & n10930 ;
  assign n10933 = x29 & n10923 ;
  assign n10934 = ( x29 & n10927 ) | ( x29 & n10933 ) | ( n10927 & n10933 ) ;
  assign n10935 = ( n2381 & n10932 ) | ( n2381 & n10934 ) | ( n10932 & n10934 ) ;
  assign n10936 = x29 & ~n10934 ;
  assign n10937 = x29 & ~n10930 ;
  assign n10938 = ( ~n2381 & n10936 ) | ( ~n2381 & n10937 ) | ( n10936 & n10937 ) ;
  assign n10939 = ( n10931 & ~n10935 ) | ( n10931 & n10938 ) | ( ~n10935 & n10938 ) ;
  assign n10940 = n10922 & n10939 ;
  assign n10941 = n10922 & ~n10940 ;
  assign n10942 = ~n10922 & n10939 ;
  assign n10943 = n10941 | n10942 ;
  assign n10944 = n10517 | n10523 ;
  assign n10945 = n10943 | n10944 ;
  assign n10946 = n10943 & n10944 ;
  assign n10947 = n10945 & ~n10946 ;
  assign n10948 = x88 & n3085 ;
  assign n10949 = x87 & n3080 ;
  assign n10950 = x86 & ~n3079 ;
  assign n10951 = n3309 & n10950 ;
  assign n10952 = n10949 | n10951 ;
  assign n10953 = n10948 | n10952 ;
  assign n10954 = n3088 | n10948 ;
  assign n10955 = n10952 | n10954 ;
  assign n10956 = ( ~n3039 & n10953 ) | ( ~n3039 & n10955 ) | ( n10953 & n10955 ) ;
  assign n10957 = n10953 & n10955 ;
  assign n10958 = ( n3023 & n10956 ) | ( n3023 & n10957 ) | ( n10956 & n10957 ) ;
  assign n10959 = x26 & n10955 ;
  assign n10960 = x26 & n10948 ;
  assign n10961 = ( x26 & n10952 ) | ( x26 & n10960 ) | ( n10952 & n10960 ) ;
  assign n10962 = ( ~n3039 & n10959 ) | ( ~n3039 & n10961 ) | ( n10959 & n10961 ) ;
  assign n10963 = n10959 & n10961 ;
  assign n10964 = ( n3023 & n10962 ) | ( n3023 & n10963 ) | ( n10962 & n10963 ) ;
  assign n10965 = x26 & ~n10961 ;
  assign n10966 = x26 & ~n10955 ;
  assign n10967 = ( n3039 & n10965 ) | ( n3039 & n10966 ) | ( n10965 & n10966 ) ;
  assign n10968 = n10965 | n10966 ;
  assign n10969 = ( ~n3023 & n10967 ) | ( ~n3023 & n10968 ) | ( n10967 & n10968 ) ;
  assign n10970 = ( n10958 & ~n10964 ) | ( n10958 & n10969 ) | ( ~n10964 & n10969 ) ;
  assign n10971 = n10947 | n10970 ;
  assign n10972 = n10947 & n10970 ;
  assign n10973 = n10971 & ~n10972 ;
  assign n10974 = n10542 | n10543 ;
  assign n10975 = ( n10357 & n10542 ) | ( n10357 & n10974 ) | ( n10542 & n10974 ) ;
  assign n10976 = n10973 & n10975 ;
  assign n10977 = n10973 | n10975 ;
  assign n10978 = ~n10976 & n10977 ;
  assign n10979 = x91 & n2429 ;
  assign n10980 = x90 & n2424 ;
  assign n10981 = x89 & ~n2423 ;
  assign n10982 = n2631 & n10981 ;
  assign n10983 = n10980 | n10982 ;
  assign n10984 = n10979 | n10983 ;
  assign n10985 = n2432 | n10979 ;
  assign n10986 = n10983 | n10985 ;
  assign n10987 = ( n3768 & n10984 ) | ( n3768 & n10986 ) | ( n10984 & n10986 ) ;
  assign n10988 = x23 & n10986 ;
  assign n10989 = x23 & n10979 ;
  assign n10990 = ( x23 & n10983 ) | ( x23 & n10989 ) | ( n10983 & n10989 ) ;
  assign n10991 = ( n3768 & n10988 ) | ( n3768 & n10990 ) | ( n10988 & n10990 ) ;
  assign n10992 = x23 & ~n10990 ;
  assign n10993 = x23 & ~n10986 ;
  assign n10994 = ( ~n3768 & n10992 ) | ( ~n3768 & n10993 ) | ( n10992 & n10993 ) ;
  assign n10995 = ( n10987 & ~n10991 ) | ( n10987 & n10994 ) | ( ~n10991 & n10994 ) ;
  assign n10996 = n10978 & n10995 ;
  assign n10997 = n10978 & ~n10996 ;
  assign n10998 = ~n10978 & n10995 ;
  assign n10999 = n10997 | n10998 ;
  assign n11000 = n10567 | n10570 ;
  assign n11001 = ( n10567 & n10572 ) | ( n10567 & n11000 ) | ( n10572 & n11000 ) ;
  assign n11002 = ~n10999 & n11001 ;
  assign n11003 = n10999 & ~n11001 ;
  assign n11004 = n11002 | n11003 ;
  assign n11005 = x94 & n1859 ;
  assign n11006 = x93 & n1854 ;
  assign n11007 = x92 & ~n1853 ;
  assign n11008 = n2037 & n11007 ;
  assign n11009 = n11006 | n11008 ;
  assign n11010 = n11005 | n11009 ;
  assign n11011 = n1862 | n11005 ;
  assign n11012 = n11009 | n11011 ;
  assign n11013 = ( n4583 & n11010 ) | ( n4583 & n11012 ) | ( n11010 & n11012 ) ;
  assign n11014 = x20 & n11012 ;
  assign n11015 = x20 & n11005 ;
  assign n11016 = ( x20 & n11009 ) | ( x20 & n11015 ) | ( n11009 & n11015 ) ;
  assign n11017 = ( n4583 & n11014 ) | ( n4583 & n11016 ) | ( n11014 & n11016 ) ;
  assign n11018 = x20 & ~n11016 ;
  assign n11019 = x20 & ~n11012 ;
  assign n11020 = ( ~n4583 & n11018 ) | ( ~n4583 & n11019 ) | ( n11018 & n11019 ) ;
  assign n11021 = ( n11013 & ~n11017 ) | ( n11013 & n11020 ) | ( ~n11017 & n11020 ) ;
  assign n11022 = n11004 & n11021 ;
  assign n11023 = n11004 | n11021 ;
  assign n11024 = ~n11022 & n11023 ;
  assign n11025 = n10594 | n10595 ;
  assign n11026 = ( n10594 & n10598 ) | ( n10594 & n11025 ) | ( n10598 & n11025 ) ;
  assign n11027 = n11024 & n11026 ;
  assign n11028 = n11024 | n11026 ;
  assign n11029 = ~n11027 & n11028 ;
  assign n11030 = x97 & n1383 ;
  assign n11031 = x96 & n1378 ;
  assign n11032 = x95 & ~n1377 ;
  assign n11033 = n1542 & n11032 ;
  assign n11034 = n11031 | n11033 ;
  assign n11035 = n11030 | n11034 ;
  assign n11036 = n1386 | n11030 ;
  assign n11037 = n11034 | n11036 ;
  assign n11038 = ( n5505 & n11035 ) | ( n5505 & n11037 ) | ( n11035 & n11037 ) ;
  assign n11039 = x17 & n11037 ;
  assign n11040 = x17 & n11030 ;
  assign n11041 = ( x17 & n11034 ) | ( x17 & n11040 ) | ( n11034 & n11040 ) ;
  assign n11042 = ( n5505 & n11039 ) | ( n5505 & n11041 ) | ( n11039 & n11041 ) ;
  assign n11043 = x17 & ~n11041 ;
  assign n11044 = x17 & ~n11037 ;
  assign n11045 = ( ~n5505 & n11043 ) | ( ~n5505 & n11044 ) | ( n11043 & n11044 ) ;
  assign n11046 = ( n11038 & ~n11042 ) | ( n11038 & n11045 ) | ( ~n11042 & n11045 ) ;
  assign n11047 = n11029 & n11046 ;
  assign n11048 = n11029 & ~n11047 ;
  assign n11049 = ~n11029 & n11046 ;
  assign n11050 = n11048 | n11049 ;
  assign n11051 = n10620 | n10622 ;
  assign n11052 = ~n11050 & n11051 ;
  assign n11053 = n11050 & ~n11051 ;
  assign n11054 = n11052 | n11053 ;
  assign n11055 = x100 & n962 ;
  assign n11056 = x99 & n957 ;
  assign n11057 = x98 & ~n956 ;
  assign n11058 = n1105 & n11057 ;
  assign n11059 = n11056 | n11058 ;
  assign n11060 = n11055 | n11059 ;
  assign n11061 = n965 | n11055 ;
  assign n11062 = n11059 | n11061 ;
  assign n11063 = ( n6483 & n11060 ) | ( n6483 & n11062 ) | ( n11060 & n11062 ) ;
  assign n11064 = x14 & n11062 ;
  assign n11065 = x14 & n11055 ;
  assign n11066 = ( x14 & n11059 ) | ( x14 & n11065 ) | ( n11059 & n11065 ) ;
  assign n11067 = ( n6483 & n11064 ) | ( n6483 & n11066 ) | ( n11064 & n11066 ) ;
  assign n11068 = x14 & ~n11066 ;
  assign n11069 = x14 & ~n11062 ;
  assign n11070 = ( ~n6483 & n11068 ) | ( ~n6483 & n11069 ) | ( n11068 & n11069 ) ;
  assign n11071 = ( n11063 & ~n11067 ) | ( n11063 & n11070 ) | ( ~n11067 & n11070 ) ;
  assign n11072 = n11054 & n11071 ;
  assign n11073 = n11054 | n11071 ;
  assign n11074 = ~n11072 & n11073 ;
  assign n11075 = n10642 & n11074 ;
  assign n11076 = ( n10648 & n11074 ) | ( n10648 & n11075 ) | ( n11074 & n11075 ) ;
  assign n11077 = n10642 | n11074 ;
  assign n11078 = n10648 | n11077 ;
  assign n11079 = ~n11076 & n11078 ;
  assign n11080 = x103 & n636 ;
  assign n11081 = x102 & n631 ;
  assign n11082 = x101 & ~n630 ;
  assign n11083 = n764 & n11082 ;
  assign n11084 = n11081 | n11083 ;
  assign n11085 = n11080 | n11084 ;
  assign n11086 = n639 | n11080 ;
  assign n11087 = n11084 | n11086 ;
  assign n11088 = ( n7529 & n11085 ) | ( n7529 & n11087 ) | ( n11085 & n11087 ) ;
  assign n11089 = x11 & n11087 ;
  assign n11090 = x11 & n11080 ;
  assign n11091 = ( x11 & n11084 ) | ( x11 & n11090 ) | ( n11084 & n11090 ) ;
  assign n11092 = ( n7529 & n11089 ) | ( n7529 & n11091 ) | ( n11089 & n11091 ) ;
  assign n11093 = x11 & ~n11091 ;
  assign n11094 = x11 & ~n11087 ;
  assign n11095 = ( ~n7529 & n11093 ) | ( ~n7529 & n11094 ) | ( n11093 & n11094 ) ;
  assign n11096 = ( n11088 & ~n11092 ) | ( n11088 & n11095 ) | ( ~n11092 & n11095 ) ;
  assign n11097 = n11079 & n11096 ;
  assign n11098 = n11079 & ~n11097 ;
  assign n11099 = ~n11079 & n11096 ;
  assign n11100 = n11098 | n11099 ;
  assign n11101 = n10667 | n10671 ;
  assign n11102 = ( n10667 & n10670 ) | ( n10667 & n11101 ) | ( n10670 & n11101 ) ;
  assign n11103 = n11100 | n11102 ;
  assign n11104 = n11100 & n11102 ;
  assign n11105 = n11103 & ~n11104 ;
  assign n11106 = x106 & n389 ;
  assign n11107 = x105 & n384 ;
  assign n11108 = x104 & ~n383 ;
  assign n11109 = n463 & n11108 ;
  assign n11110 = n11107 | n11109 ;
  assign n11111 = n11106 | n11110 ;
  assign n11112 = n392 | n11106 ;
  assign n11113 = n11110 | n11112 ;
  assign n11114 = ( n8656 & n11111 ) | ( n8656 & n11113 ) | ( n11111 & n11113 ) ;
  assign n11115 = x8 & n11113 ;
  assign n11116 = x8 & n11106 ;
  assign n11117 = ( x8 & n11110 ) | ( x8 & n11116 ) | ( n11110 & n11116 ) ;
  assign n11118 = ( n8656 & n11115 ) | ( n8656 & n11117 ) | ( n11115 & n11117 ) ;
  assign n11119 = x8 & ~n11117 ;
  assign n11120 = x8 & ~n11113 ;
  assign n11121 = ( ~n8656 & n11119 ) | ( ~n8656 & n11120 ) | ( n11119 & n11120 ) ;
  assign n11122 = ( n11114 & ~n11118 ) | ( n11114 & n11121 ) | ( ~n11118 & n11121 ) ;
  assign n11123 = n11105 & n11122 ;
  assign n11124 = n11105 & ~n11123 ;
  assign n11125 = ~n11105 & n11122 ;
  assign n11126 = n10692 | n10696 ;
  assign n11127 = ( n10692 & n10694 ) | ( n10692 & n11126 ) | ( n10694 & n11126 ) ;
  assign n11128 = ~n11125 & n11127 ;
  assign n11129 = ~n11124 & n11128 ;
  assign n11130 = n11125 & ~n11127 ;
  assign n11131 = ( n11124 & ~n11127 ) | ( n11124 & n11130 ) | ( ~n11127 & n11130 ) ;
  assign n11132 = n11129 | n11131 ;
  assign n11133 = x109 & n212 ;
  assign n11134 = x108 & n207 ;
  assign n11135 = x107 & ~n206 ;
  assign n11136 = n267 & n11135 ;
  assign n11137 = n11134 | n11136 ;
  assign n11138 = n11133 | n11137 ;
  assign n11139 = n215 | n11133 ;
  assign n11140 = n11137 | n11139 ;
  assign n11141 = ( n9878 & n11138 ) | ( n9878 & n11140 ) | ( n11138 & n11140 ) ;
  assign n11142 = x5 & n11140 ;
  assign n11143 = x5 & n11133 ;
  assign n11144 = ( x5 & n11137 ) | ( x5 & n11143 ) | ( n11137 & n11143 ) ;
  assign n11145 = ( n9878 & n11142 ) | ( n9878 & n11144 ) | ( n11142 & n11144 ) ;
  assign n11146 = x5 & ~n11144 ;
  assign n11147 = x5 & ~n11140 ;
  assign n11148 = ( ~n9878 & n11146 ) | ( ~n9878 & n11147 ) | ( n11146 & n11147 ) ;
  assign n11149 = ( n11141 & ~n11145 ) | ( n11141 & n11148 ) | ( ~n11145 & n11148 ) ;
  assign n11150 = n11132 & n11149 ;
  assign n11151 = n11132 | n11149 ;
  assign n11152 = ~n11150 & n11151 ;
  assign n11153 = n10718 | n10722 ;
  assign n11154 = n11152 & n11153 ;
  assign n11155 = n11152 | n11153 ;
  assign n11156 = ~n11154 & n11155 ;
  assign n11157 = x111 | x112 ;
  assign n11158 = x111 & x112 ;
  assign n11159 = n11157 & ~n11158 ;
  assign n11160 = n10726 & n11159 ;
  assign n11161 = ( n10735 & n11159 ) | ( n10735 & n11160 ) | ( n11159 & n11160 ) ;
  assign n11162 = ( n10736 & n11159 ) | ( n10736 & n11160 ) | ( n11159 & n11160 ) ;
  assign n11163 = ( n6159 & n11161 ) | ( n6159 & n11162 ) | ( n11161 & n11162 ) ;
  assign n11164 = ( n6157 & n11161 ) | ( n6157 & n11162 ) | ( n11161 & n11162 ) ;
  assign n11165 = ( n5823 & n11163 ) | ( n5823 & n11164 ) | ( n11163 & n11164 ) ;
  assign n11166 = n10726 | n11159 ;
  assign n11167 = n10735 | n11166 ;
  assign n11168 = n10736 | n11166 ;
  assign n11169 = ( n6159 & n11167 ) | ( n6159 & n11168 ) | ( n11167 & n11168 ) ;
  assign n11170 = ( n6157 & n11167 ) | ( n6157 & n11168 ) | ( n11167 & n11168 ) ;
  assign n11171 = ( n5823 & n11169 ) | ( n5823 & n11170 ) | ( n11169 & n11170 ) ;
  assign n11172 = ~n11165 & n11171 ;
  assign n11173 = x111 & n133 ;
  assign n11174 = x110 & ~n162 ;
  assign n11175 = ( n137 & n11173 ) | ( n137 & n11174 ) | ( n11173 & n11174 ) ;
  assign n11176 = x0 & x112 ;
  assign n11177 = ( ~n137 & n11173 ) | ( ~n137 & n11176 ) | ( n11173 & n11176 ) ;
  assign n11178 = n11175 | n11177 ;
  assign n11179 = n141 | n11178 ;
  assign n11180 = ( n11172 & n11178 ) | ( n11172 & n11179 ) | ( n11178 & n11179 ) ;
  assign n11181 = x2 & n11178 ;
  assign n11182 = ( x2 & n523 ) | ( x2 & n11178 ) | ( n523 & n11178 ) ;
  assign n11183 = ( n11172 & n11181 ) | ( n11172 & n11182 ) | ( n11181 & n11182 ) ;
  assign n11184 = x2 & ~n11182 ;
  assign n11185 = x2 & ~n11178 ;
  assign n11186 = ( ~n11172 & n11184 ) | ( ~n11172 & n11185 ) | ( n11184 & n11185 ) ;
  assign n11187 = ( n11180 & ~n11183 ) | ( n11180 & n11186 ) | ( ~n11183 & n11186 ) ;
  assign n11188 = n11156 | n11187 ;
  assign n11189 = n11156 & n11187 ;
  assign n11190 = n11188 & ~n11189 ;
  assign n11191 = n10774 | n11190 ;
  assign n11192 = n10774 & n11190 ;
  assign n11193 = n11191 & ~n11192 ;
  assign n11194 = ( n10978 & n10995 ) | ( n10978 & n11001 ) | ( n10995 & n11001 ) ;
  assign n11195 = n10842 | n10843 ;
  assign n11196 = ( n10842 & n10845 ) | ( n10842 & n11195 ) | ( n10845 & n11195 ) ;
  assign n11197 = ~x48 & x49 ;
  assign n11198 = x48 & ~x49 ;
  assign n11199 = n11197 | n11198 ;
  assign n11200 = ~n10779 & n11199 ;
  assign n11201 = x64 & n11200 ;
  assign n11202 = ~x49 & x50 ;
  assign n11203 = x49 & ~x50 ;
  assign n11204 = n11202 | n11203 ;
  assign n11205 = n10779 & ~n11204 ;
  assign n11206 = x65 & n11205 ;
  assign n11207 = n11201 | n11206 ;
  assign n11208 = n10779 & n11204 ;
  assign n11209 = x50 | n144 ;
  assign n11210 = ( x50 & n11208 ) | ( x50 & n11209 ) | ( n11208 & n11209 ) ;
  assign n11211 = ~x50 & n11210 ;
  assign n11212 = ( ~x50 & n11207 ) | ( ~x50 & n11211 ) | ( n11207 & n11211 ) ;
  assign n11213 = x50 & ~x64 ;
  assign n11214 = ( x50 & ~n10779 ) | ( x50 & n11213 ) | ( ~n10779 & n11213 ) ;
  assign n11215 = n11210 & n11214 ;
  assign n11216 = ( n11207 & n11214 ) | ( n11207 & n11215 ) | ( n11214 & n11215 ) ;
  assign n11217 = n144 & n11208 ;
  assign n11218 = n11214 & ~n11217 ;
  assign n11219 = ~n11207 & n11218 ;
  assign n11220 = ( n11212 & n11216 ) | ( n11212 & n11219 ) | ( n11216 & n11219 ) ;
  assign n11221 = n11210 | n11214 ;
  assign n11222 = n11207 | n11221 ;
  assign n11223 = ~n11214 & n11217 ;
  assign n11224 = ( n11207 & ~n11214 ) | ( n11207 & n11223 ) | ( ~n11214 & n11223 ) ;
  assign n11225 = ( n11212 & n11222 ) | ( n11212 & ~n11224 ) | ( n11222 & ~n11224 ) ;
  assign n11226 = ~n11220 & n11225 ;
  assign n11227 = n241 & n9936 ;
  assign n11228 = x68 & n9933 ;
  assign n11229 = x67 & n9928 ;
  assign n11230 = x66 & ~n9927 ;
  assign n11231 = n10379 & n11230 ;
  assign n11232 = n11229 | n11231 ;
  assign n11233 = n11228 | n11232 ;
  assign n11234 = n11227 | n11233 ;
  assign n11235 = x47 | n11228 ;
  assign n11236 = n11232 | n11235 ;
  assign n11237 = n11227 | n11236 ;
  assign n11238 = ~x47 & n11236 ;
  assign n11239 = ( ~x47 & n11227 ) | ( ~x47 & n11238 ) | ( n11227 & n11238 ) ;
  assign n11240 = ( ~n11234 & n11237 ) | ( ~n11234 & n11239 ) | ( n11237 & n11239 ) ;
  assign n11241 = n11226 | n11240 ;
  assign n11242 = n11226 & n11240 ;
  assign n11243 = n11241 & ~n11242 ;
  assign n11244 = ( n10393 & n10780 ) | ( n10393 & n10796 ) | ( n10780 & n10796 ) ;
  assign n11245 = n11243 | n11244 ;
  assign n11246 = n11243 & n11244 ;
  assign n11247 = n11245 & ~n11246 ;
  assign n11248 = x70 & n8719 ;
  assign n11249 = x69 & ~n8718 ;
  assign n11250 = n9149 & n11249 ;
  assign n11251 = n11248 | n11250 ;
  assign n11252 = x71 & n8724 ;
  assign n11253 = n8727 | n11252 ;
  assign n11254 = n11251 | n11253 ;
  assign n11255 = x44 & ~n11254 ;
  assign n11256 = x44 & ~n11252 ;
  assign n11257 = ~n11251 & n11256 ;
  assign n11258 = ( ~n438 & n11255 ) | ( ~n438 & n11257 ) | ( n11255 & n11257 ) ;
  assign n11259 = ~x44 & n11254 ;
  assign n11260 = ~x44 & n11252 ;
  assign n11261 = ( ~x44 & n11251 ) | ( ~x44 & n11260 ) | ( n11251 & n11260 ) ;
  assign n11262 = ( n438 & n11259 ) | ( n438 & n11261 ) | ( n11259 & n11261 ) ;
  assign n11263 = n11258 | n11262 ;
  assign n11264 = n11247 & n11263 ;
  assign n11265 = n11247 & ~n11264 ;
  assign n11266 = ~n11247 & n11263 ;
  assign n11267 = n11265 | n11266 ;
  assign n11268 = n10816 | n10821 ;
  assign n11269 = ( n10816 & n10819 ) | ( n10816 & n11268 ) | ( n10819 & n11268 ) ;
  assign n11270 = n11267 | n11269 ;
  assign n11271 = n11267 & n11269 ;
  assign n11272 = n11270 & ~n11271 ;
  assign n11273 = x74 & n7566 ;
  assign n11274 = x73 & n7561 ;
  assign n11275 = x72 & ~n7560 ;
  assign n11276 = n7953 & n11275 ;
  assign n11277 = n11274 | n11276 ;
  assign n11278 = n11273 | n11277 ;
  assign n11279 = n7569 | n11273 ;
  assign n11280 = n11277 | n11279 ;
  assign n11281 = ( n710 & n11278 ) | ( n710 & n11280 ) | ( n11278 & n11280 ) ;
  assign n11282 = x41 & n11280 ;
  assign n11283 = x41 & n11273 ;
  assign n11284 = ( x41 & n11277 ) | ( x41 & n11283 ) | ( n11277 & n11283 ) ;
  assign n11285 = ( n710 & n11282 ) | ( n710 & n11284 ) | ( n11282 & n11284 ) ;
  assign n11286 = x41 & ~n11284 ;
  assign n11287 = x41 & ~n11280 ;
  assign n11288 = ( ~n710 & n11286 ) | ( ~n710 & n11287 ) | ( n11286 & n11287 ) ;
  assign n11289 = ( n11281 & ~n11285 ) | ( n11281 & n11288 ) | ( ~n11285 & n11288 ) ;
  assign n11290 = n11272 & n11289 ;
  assign n11291 = n11272 | n11289 ;
  assign n11292 = ~n11290 & n11291 ;
  assign n11293 = n11196 & n11292 ;
  assign n11294 = n11196 & ~n11293 ;
  assign n11295 = x77 & n6536 ;
  assign n11296 = x76 & n6531 ;
  assign n11297 = x75 & ~n6530 ;
  assign n11298 = n6871 & n11297 ;
  assign n11299 = n11296 | n11298 ;
  assign n11300 = n11295 | n11299 ;
  assign n11301 = n6539 | n11295 ;
  assign n11302 = n11299 | n11301 ;
  assign n11303 = ( n1059 & n11300 ) | ( n1059 & n11302 ) | ( n11300 & n11302 ) ;
  assign n11304 = x38 & n11302 ;
  assign n11305 = x38 & n11295 ;
  assign n11306 = ( x38 & n11299 ) | ( x38 & n11305 ) | ( n11299 & n11305 ) ;
  assign n11307 = ( n1059 & n11304 ) | ( n1059 & n11306 ) | ( n11304 & n11306 ) ;
  assign n11308 = x38 & ~n11306 ;
  assign n11309 = x38 & ~n11302 ;
  assign n11310 = ( ~n1059 & n11308 ) | ( ~n1059 & n11309 ) | ( n11308 & n11309 ) ;
  assign n11311 = ( n11303 & ~n11307 ) | ( n11303 & n11310 ) | ( ~n11307 & n11310 ) ;
  assign n11312 = ~n11291 & n11292 ;
  assign n11313 = ( ~n11196 & n11292 ) | ( ~n11196 & n11312 ) | ( n11292 & n11312 ) ;
  assign n11314 = n11311 & n11313 ;
  assign n11315 = ( n11294 & n11311 ) | ( n11294 & n11314 ) | ( n11311 & n11314 ) ;
  assign n11316 = n11311 | n11313 ;
  assign n11317 = n11294 | n11316 ;
  assign n11318 = ~n11315 & n11317 ;
  assign n11319 = n10776 | n10866 ;
  assign n11320 = ( n10866 & n10869 ) | ( n10866 & n11319 ) | ( n10869 & n11319 ) ;
  assign n11321 = n11318 & n11320 ;
  assign n11322 = n11318 | n11320 ;
  assign n11323 = ~n11321 & n11322 ;
  assign n11324 = x80 & n5554 ;
  assign n11325 = x79 & n5549 ;
  assign n11326 = x78 & ~n5548 ;
  assign n11327 = n5893 & n11326 ;
  assign n11328 = n11325 | n11327 ;
  assign n11329 = n11324 | n11328 ;
  assign n11330 = n5557 | n11324 ;
  assign n11331 = n11328 | n11330 ;
  assign n11332 = ( n1499 & n11329 ) | ( n1499 & n11331 ) | ( n11329 & n11331 ) ;
  assign n11333 = x35 & n11331 ;
  assign n11334 = x35 & n11324 ;
  assign n11335 = ( x35 & n11328 ) | ( x35 & n11334 ) | ( n11328 & n11334 ) ;
  assign n11336 = ( n1499 & n11333 ) | ( n1499 & n11335 ) | ( n11333 & n11335 ) ;
  assign n11337 = x35 & ~n11335 ;
  assign n11338 = x35 & ~n11331 ;
  assign n11339 = ( ~n1499 & n11337 ) | ( ~n1499 & n11338 ) | ( n11337 & n11338 ) ;
  assign n11340 = ( n11332 & ~n11336 ) | ( n11332 & n11339 ) | ( ~n11336 & n11339 ) ;
  assign n11341 = n11323 & n11340 ;
  assign n11342 = n11323 & ~n11341 ;
  assign n11343 = ~n11323 & n11340 ;
  assign n11344 = n11342 | n11343 ;
  assign n11345 = n10890 | n10893 ;
  assign n11346 = n11344 | n11345 ;
  assign n11347 = n11344 & n11345 ;
  assign n11348 = n11346 & ~n11347 ;
  assign n11349 = x83 & n4631 ;
  assign n11350 = x82 & n4626 ;
  assign n11351 = x81 & ~n4625 ;
  assign n11352 = n4943 & n11351 ;
  assign n11353 = n11350 | n11352 ;
  assign n11354 = n11349 | n11353 ;
  assign n11355 = n4634 | n11349 ;
  assign n11356 = n11353 | n11355 ;
  assign n11357 = ( n2009 & n11354 ) | ( n2009 & n11356 ) | ( n11354 & n11356 ) ;
  assign n11358 = x32 & n11356 ;
  assign n11359 = x32 & n11349 ;
  assign n11360 = ( x32 & n11353 ) | ( x32 & n11359 ) | ( n11353 & n11359 ) ;
  assign n11361 = ( n2009 & n11358 ) | ( n2009 & n11360 ) | ( n11358 & n11360 ) ;
  assign n11362 = x32 & ~n11360 ;
  assign n11363 = x32 & ~n11356 ;
  assign n11364 = ( ~n2009 & n11362 ) | ( ~n2009 & n11363 ) | ( n11362 & n11363 ) ;
  assign n11365 = ( n11357 & ~n11361 ) | ( n11357 & n11364 ) | ( ~n11361 & n11364 ) ;
  assign n11366 = n11348 & n11365 ;
  assign n11367 = n11348 & ~n11366 ;
  assign n11368 = ~n11348 & n11365 ;
  assign n11369 = n11367 | n11368 ;
  assign n11370 = n10913 | n10921 ;
  assign n11371 = n11369 | n11370 ;
  assign n11372 = n11369 & n11370 ;
  assign n11373 = n11371 & ~n11372 ;
  assign n11374 = x86 & n3816 ;
  assign n11375 = x85 & n3811 ;
  assign n11376 = x84 & ~n3810 ;
  assign n11377 = n4067 & n11376 ;
  assign n11378 = n11375 | n11377 ;
  assign n11379 = n11374 | n11378 ;
  assign n11380 = n3819 | n11374 ;
  assign n11381 = n11378 | n11380 ;
  assign n11382 = ( n2606 & n11379 ) | ( n2606 & n11381 ) | ( n11379 & n11381 ) ;
  assign n11383 = x29 & n11381 ;
  assign n11384 = x29 & n11374 ;
  assign n11385 = ( x29 & n11378 ) | ( x29 & n11384 ) | ( n11378 & n11384 ) ;
  assign n11386 = ( n2606 & n11383 ) | ( n2606 & n11385 ) | ( n11383 & n11385 ) ;
  assign n11387 = x29 & ~n11385 ;
  assign n11388 = x29 & ~n11381 ;
  assign n11389 = ( ~n2606 & n11387 ) | ( ~n2606 & n11388 ) | ( n11387 & n11388 ) ;
  assign n11390 = ( n11382 & ~n11386 ) | ( n11382 & n11389 ) | ( ~n11386 & n11389 ) ;
  assign n11391 = n11373 & n11390 ;
  assign n11392 = n11373 & ~n11391 ;
  assign n11393 = ~n11373 & n11390 ;
  assign n11394 = n11392 | n11393 ;
  assign n11395 = n10940 | n10946 ;
  assign n11396 = n11394 | n11395 ;
  assign n11397 = n11394 & n11395 ;
  assign n11398 = n11396 & ~n11397 ;
  assign n11399 = x89 & n3085 ;
  assign n11400 = x88 & n3080 ;
  assign n11401 = x87 & ~n3079 ;
  assign n11402 = n3309 & n11401 ;
  assign n11403 = n11400 | n11402 ;
  assign n11404 = n11399 | n11403 ;
  assign n11405 = n3088 | n11399 ;
  assign n11406 = n11403 | n11405 ;
  assign n11407 = ( n3282 & n11404 ) | ( n3282 & n11406 ) | ( n11404 & n11406 ) ;
  assign n11408 = x26 & n11406 ;
  assign n11409 = x26 & n11399 ;
  assign n11410 = ( x26 & n11403 ) | ( x26 & n11409 ) | ( n11403 & n11409 ) ;
  assign n11411 = ( n3282 & n11408 ) | ( n3282 & n11410 ) | ( n11408 & n11410 ) ;
  assign n11412 = x26 & ~n11410 ;
  assign n11413 = x26 & ~n11406 ;
  assign n11414 = ( ~n3282 & n11412 ) | ( ~n3282 & n11413 ) | ( n11412 & n11413 ) ;
  assign n11415 = ( n11407 & ~n11411 ) | ( n11407 & n11414 ) | ( ~n11411 & n11414 ) ;
  assign n11416 = n11398 & n11415 ;
  assign n11417 = n11398 & ~n11416 ;
  assign n11418 = ~n11398 & n11415 ;
  assign n11419 = n11417 | n11418 ;
  assign n11420 = n10972 | n10976 ;
  assign n11421 = n11419 & n11420 ;
  assign n11422 = n11419 | n11420 ;
  assign n11423 = ~n11421 & n11422 ;
  assign n11424 = x92 & n2429 ;
  assign n11425 = x91 & n2424 ;
  assign n11426 = x90 & ~n2423 ;
  assign n11427 = n2631 & n11426 ;
  assign n11428 = n11425 | n11427 ;
  assign n11429 = n11424 | n11428 ;
  assign n11430 = n2432 | n11424 ;
  assign n11431 = n11428 | n11430 ;
  assign n11432 = ( n4040 & n11429 ) | ( n4040 & n11431 ) | ( n11429 & n11431 ) ;
  assign n11433 = x23 & n11431 ;
  assign n11434 = x23 & n11424 ;
  assign n11435 = ( x23 & n11428 ) | ( x23 & n11434 ) | ( n11428 & n11434 ) ;
  assign n11436 = ( n4040 & n11433 ) | ( n4040 & n11435 ) | ( n11433 & n11435 ) ;
  assign n11437 = x23 & ~n11435 ;
  assign n11438 = x23 & ~n11431 ;
  assign n11439 = ( ~n4040 & n11437 ) | ( ~n4040 & n11438 ) | ( n11437 & n11438 ) ;
  assign n11440 = ( n11432 & ~n11436 ) | ( n11432 & n11439 ) | ( ~n11436 & n11439 ) ;
  assign n11441 = n11423 & n11440 ;
  assign n11442 = n11423 & ~n11441 ;
  assign n11443 = ~n11423 & n11440 ;
  assign n11444 = n11194 & n11443 ;
  assign n11445 = ( n11194 & n11442 ) | ( n11194 & n11444 ) | ( n11442 & n11444 ) ;
  assign n11446 = n11194 & ~n11445 ;
  assign n11447 = n11442 | n11443 ;
  assign n11448 = ~n11445 & n11447 ;
  assign n11449 = n11446 | n11448 ;
  assign n11450 = x95 & n1859 ;
  assign n11451 = x94 & n1854 ;
  assign n11452 = x93 & ~n1853 ;
  assign n11453 = n2037 & n11452 ;
  assign n11454 = n11451 | n11453 ;
  assign n11455 = n11450 | n11454 ;
  assign n11456 = n1862 | n11450 ;
  assign n11457 = n11454 | n11456 ;
  assign n11458 = ( n4897 & n11455 ) | ( n4897 & n11457 ) | ( n11455 & n11457 ) ;
  assign n11459 = x20 & n11457 ;
  assign n11460 = x20 & n11450 ;
  assign n11461 = ( x20 & n11454 ) | ( x20 & n11460 ) | ( n11454 & n11460 ) ;
  assign n11462 = ( n4897 & n11459 ) | ( n4897 & n11461 ) | ( n11459 & n11461 ) ;
  assign n11463 = x20 & ~n11461 ;
  assign n11464 = x20 & ~n11457 ;
  assign n11465 = ( ~n4897 & n11463 ) | ( ~n4897 & n11464 ) | ( n11463 & n11464 ) ;
  assign n11466 = ( n11458 & ~n11462 ) | ( n11458 & n11465 ) | ( ~n11462 & n11465 ) ;
  assign n11467 = n11449 & n11466 ;
  assign n11468 = n11449 & ~n11467 ;
  assign n11470 = n11022 | n11024 ;
  assign n11471 = ( n11022 & n11026 ) | ( n11022 & n11470 ) | ( n11026 & n11470 ) ;
  assign n11469 = ~n11449 & n11466 ;
  assign n11472 = n11469 & n11471 ;
  assign n11473 = ( n11468 & n11471 ) | ( n11468 & n11472 ) | ( n11471 & n11472 ) ;
  assign n11474 = n11469 | n11471 ;
  assign n11475 = n11468 | n11474 ;
  assign n11476 = ~n11473 & n11475 ;
  assign n11477 = x98 & n1383 ;
  assign n11478 = x97 & n1378 ;
  assign n11479 = x96 & ~n1377 ;
  assign n11480 = n1542 & n11479 ;
  assign n11481 = n11478 | n11480 ;
  assign n11482 = n11477 | n11481 ;
  assign n11483 = n1386 | n11477 ;
  assign n11484 = n11481 | n11483 ;
  assign n11485 = ( ~n5850 & n11482 ) | ( ~n5850 & n11484 ) | ( n11482 & n11484 ) ;
  assign n11486 = n11482 & n11484 ;
  assign n11487 = ( n5834 & n11485 ) | ( n5834 & n11486 ) | ( n11485 & n11486 ) ;
  assign n11488 = x17 & n11484 ;
  assign n11489 = x17 & n11477 ;
  assign n11490 = ( x17 & n11481 ) | ( x17 & n11489 ) | ( n11481 & n11489 ) ;
  assign n11491 = ( ~n5850 & n11488 ) | ( ~n5850 & n11490 ) | ( n11488 & n11490 ) ;
  assign n11492 = n11488 & n11490 ;
  assign n11493 = ( n5834 & n11491 ) | ( n5834 & n11492 ) | ( n11491 & n11492 ) ;
  assign n11494 = x17 & ~n11490 ;
  assign n11495 = x17 & ~n11484 ;
  assign n11496 = ( n5850 & n11494 ) | ( n5850 & n11495 ) | ( n11494 & n11495 ) ;
  assign n11497 = n11494 | n11495 ;
  assign n11498 = ( ~n5834 & n11496 ) | ( ~n5834 & n11497 ) | ( n11496 & n11497 ) ;
  assign n11499 = ( n11487 & ~n11493 ) | ( n11487 & n11498 ) | ( ~n11493 & n11498 ) ;
  assign n11500 = n11476 & n11499 ;
  assign n11501 = n11476 & ~n11500 ;
  assign n11502 = ( n10620 & n11029 ) | ( n10620 & n11046 ) | ( n11029 & n11046 ) ;
  assign n11503 = n11029 | n11046 ;
  assign n11504 = ( n10622 & n11502 ) | ( n10622 & n11503 ) | ( n11502 & n11503 ) ;
  assign n11505 = ~n11476 & n11499 ;
  assign n11506 = n11504 & n11505 ;
  assign n11507 = ( n11501 & n11504 ) | ( n11501 & n11506 ) | ( n11504 & n11506 ) ;
  assign n11508 = n11504 | n11505 ;
  assign n11509 = n11501 | n11508 ;
  assign n11510 = ~n11507 & n11509 ;
  assign n11511 = x101 & n962 ;
  assign n11512 = x100 & n957 ;
  assign n11513 = x99 & ~n956 ;
  assign n11514 = n1105 & n11513 ;
  assign n11515 = n11512 | n11514 ;
  assign n11516 = n11511 | n11515 ;
  assign n11517 = n965 | n11511 ;
  assign n11518 = n11515 | n11517 ;
  assign n11519 = ( n6844 & n11516 ) | ( n6844 & n11518 ) | ( n11516 & n11518 ) ;
  assign n11520 = x14 & n11518 ;
  assign n11521 = x14 & n11511 ;
  assign n11522 = ( x14 & n11515 ) | ( x14 & n11521 ) | ( n11515 & n11521 ) ;
  assign n11523 = ( n6844 & n11520 ) | ( n6844 & n11522 ) | ( n11520 & n11522 ) ;
  assign n11524 = x14 & ~n11522 ;
  assign n11525 = x14 & ~n11518 ;
  assign n11526 = ( ~n6844 & n11524 ) | ( ~n6844 & n11525 ) | ( n11524 & n11525 ) ;
  assign n11527 = ( n11519 & ~n11523 ) | ( n11519 & n11526 ) | ( ~n11523 & n11526 ) ;
  assign n11528 = n11510 & n11527 ;
  assign n11529 = n11510 & ~n11528 ;
  assign n11530 = ~n11510 & n11527 ;
  assign n11531 = n11529 | n11530 ;
  assign n11532 = n11072 | n11074 ;
  assign n11533 = n10648 | n11072 ;
  assign n11534 = ( n11075 & n11532 ) | ( n11075 & n11533 ) | ( n11532 & n11533 ) ;
  assign n11535 = n11531 | n11534 ;
  assign n11536 = n11531 & n11534 ;
  assign n11537 = n11535 & ~n11536 ;
  assign n11538 = x104 & n636 ;
  assign n11539 = x103 & n631 ;
  assign n11540 = x102 & ~n630 ;
  assign n11541 = n764 & n11540 ;
  assign n11542 = n11539 | n11541 ;
  assign n11543 = n11538 | n11542 ;
  assign n11544 = n639 | n11538 ;
  assign n11545 = n11542 | n11544 ;
  assign n11546 = ( n7911 & n11543 ) | ( n7911 & n11545 ) | ( n11543 & n11545 ) ;
  assign n11547 = x11 & n11545 ;
  assign n11548 = x11 & n11538 ;
  assign n11549 = ( x11 & n11542 ) | ( x11 & n11548 ) | ( n11542 & n11548 ) ;
  assign n11550 = ( n7911 & n11547 ) | ( n7911 & n11549 ) | ( n11547 & n11549 ) ;
  assign n11551 = x11 & ~n11549 ;
  assign n11552 = x11 & ~n11545 ;
  assign n11553 = ( ~n7911 & n11551 ) | ( ~n7911 & n11552 ) | ( n11551 & n11552 ) ;
  assign n11554 = ( n11546 & ~n11550 ) | ( n11546 & n11553 ) | ( ~n11550 & n11553 ) ;
  assign n11555 = n11537 & n11554 ;
  assign n11556 = n11537 & ~n11555 ;
  assign n11557 = ~n11537 & n11554 ;
  assign n11558 = n11556 | n11557 ;
  assign n11559 = n11097 | n11102 ;
  assign n11560 = ( n11097 & n11100 ) | ( n11097 & n11559 ) | ( n11100 & n11559 ) ;
  assign n11561 = n11558 | n11560 ;
  assign n11562 = n11558 & n11560 ;
  assign n11563 = n11561 & ~n11562 ;
  assign n11564 = x107 & n389 ;
  assign n11565 = x106 & n384 ;
  assign n11566 = x105 & ~n383 ;
  assign n11567 = n463 & n11566 ;
  assign n11568 = n11565 | n11567 ;
  assign n11569 = n11564 | n11568 ;
  assign n11570 = n392 | n11564 ;
  assign n11571 = n11568 | n11570 ;
  assign n11572 = ( n9084 & n11569 ) | ( n9084 & n11571 ) | ( n11569 & n11571 ) ;
  assign n11573 = x8 & n11571 ;
  assign n11574 = x8 & n11564 ;
  assign n11575 = ( x8 & n11568 ) | ( x8 & n11574 ) | ( n11568 & n11574 ) ;
  assign n11576 = ( n9084 & n11573 ) | ( n9084 & n11575 ) | ( n11573 & n11575 ) ;
  assign n11577 = x8 & ~n11575 ;
  assign n11578 = x8 & ~n11571 ;
  assign n11579 = ( ~n9084 & n11577 ) | ( ~n9084 & n11578 ) | ( n11577 & n11578 ) ;
  assign n11580 = ( n11572 & ~n11576 ) | ( n11572 & n11579 ) | ( ~n11576 & n11579 ) ;
  assign n11581 = n11563 & n11580 ;
  assign n11582 = n11563 & ~n11581 ;
  assign n11583 = ( n11105 & n11122 ) | ( n11105 & n11127 ) | ( n11122 & n11127 ) ;
  assign n11584 = ~n11563 & n11580 ;
  assign n11585 = n11583 & n11584 ;
  assign n11586 = ( n11582 & n11583 ) | ( n11582 & n11585 ) | ( n11583 & n11585 ) ;
  assign n11587 = n11583 | n11584 ;
  assign n11588 = n11582 | n11587 ;
  assign n11589 = ~n11586 & n11588 ;
  assign n11590 = x110 & n212 ;
  assign n11591 = x109 & n207 ;
  assign n11592 = x108 & ~n206 ;
  assign n11593 = n267 & n11592 ;
  assign n11594 = n11591 | n11593 ;
  assign n11595 = n11590 | n11594 ;
  assign n11596 = n215 | n11590 ;
  assign n11597 = n11594 | n11596 ;
  assign n11598 = ( n10330 & n11595 ) | ( n10330 & n11597 ) | ( n11595 & n11597 ) ;
  assign n11599 = x5 & n11597 ;
  assign n11600 = x5 & n11590 ;
  assign n11601 = ( x5 & n11594 ) | ( x5 & n11600 ) | ( n11594 & n11600 ) ;
  assign n11602 = ( n10330 & n11599 ) | ( n10330 & n11601 ) | ( n11599 & n11601 ) ;
  assign n11603 = x5 & ~n11601 ;
  assign n11604 = x5 & ~n11597 ;
  assign n11605 = ( ~n10330 & n11603 ) | ( ~n10330 & n11604 ) | ( n11603 & n11604 ) ;
  assign n11606 = ( n11598 & ~n11602 ) | ( n11598 & n11605 ) | ( ~n11602 & n11605 ) ;
  assign n11607 = n11589 & n11606 ;
  assign n11608 = n11589 & ~n11607 ;
  assign n11609 = ~n11589 & n11606 ;
  assign n11610 = n11608 | n11609 ;
  assign n11611 = n11150 | n11154 ;
  assign n11612 = n11610 | n11611 ;
  assign n11613 = n11610 & n11611 ;
  assign n11614 = n11612 & ~n11613 ;
  assign n11615 = x112 | x113 ;
  assign n11616 = x112 & x113 ;
  assign n11617 = n11615 & ~n11616 ;
  assign n11618 = n11158 | n11159 ;
  assign n11619 = ( n10726 & n11158 ) | ( n10726 & n11618 ) | ( n11158 & n11618 ) ;
  assign n11620 = n11158 | n11618 ;
  assign n11621 = ( n10735 & n11619 ) | ( n10735 & n11620 ) | ( n11619 & n11620 ) ;
  assign n11622 = ( n10736 & n11619 ) | ( n10736 & n11620 ) | ( n11619 & n11620 ) ;
  assign n11623 = ( n6159 & n11621 ) | ( n6159 & n11622 ) | ( n11621 & n11622 ) ;
  assign n11624 = ( n6157 & n11621 ) | ( n6157 & n11622 ) | ( n11621 & n11622 ) ;
  assign n11625 = ( n5823 & n11623 ) | ( n5823 & n11624 ) | ( n11623 & n11624 ) ;
  assign n11626 = n11617 | n11625 ;
  assign n11627 = x112 & n133 ;
  assign n11628 = x111 & ~n162 ;
  assign n11629 = ( n137 & n11627 ) | ( n137 & n11628 ) | ( n11627 & n11628 ) ;
  assign n11630 = x0 & x113 ;
  assign n11631 = ( ~n137 & n11627 ) | ( ~n137 & n11630 ) | ( n11627 & n11630 ) ;
  assign n11632 = n11629 | n11631 ;
  assign n11633 = n141 | n11632 ;
  assign n11634 = n11617 & n11618 ;
  assign n11635 = n11158 & n11617 ;
  assign n11636 = ( n10726 & n11634 ) | ( n10726 & n11635 ) | ( n11634 & n11635 ) ;
  assign n11637 = n11634 | n11635 ;
  assign n11638 = ( n10735 & n11636 ) | ( n10735 & n11637 ) | ( n11636 & n11637 ) ;
  assign n11639 = ( n10736 & n11636 ) | ( n10736 & n11637 ) | ( n11636 & n11637 ) ;
  assign n11640 = ( n6159 & n11638 ) | ( n6159 & n11639 ) | ( n11638 & n11639 ) ;
  assign n11641 = ( n6157 & n11638 ) | ( n6157 & n11639 ) | ( n11638 & n11639 ) ;
  assign n11642 = ( n5823 & n11640 ) | ( n5823 & n11641 ) | ( n11640 & n11641 ) ;
  assign n11643 = ( n11632 & n11633 ) | ( n11632 & ~n11642 ) | ( n11633 & ~n11642 ) ;
  assign n11644 = n11632 & n11633 ;
  assign n11645 = ( n11626 & n11643 ) | ( n11626 & n11644 ) | ( n11643 & n11644 ) ;
  assign n11646 = x2 & n11645 ;
  assign n11647 = x2 & ~n11645 ;
  assign n11648 = ( n11645 & ~n11646 ) | ( n11645 & n11647 ) | ( ~n11646 & n11647 ) ;
  assign n11649 = n11614 | n11648 ;
  assign n11650 = n11614 & n11648 ;
  assign n11651 = n11649 & ~n11650 ;
  assign n11652 = n11189 | n11190 ;
  assign n11653 = ( n10774 & n11189 ) | ( n10774 & n11652 ) | ( n11189 & n11652 ) ;
  assign n11654 = n11651 & n11653 ;
  assign n11655 = n11651 | n11653 ;
  assign n11656 = ~n11654 & n11655 ;
  assign n11657 = n11391 | n11397 ;
  assign n11658 = n11341 | n11347 ;
  assign n11659 = x75 & n7566 ;
  assign n11660 = x74 & n7561 ;
  assign n11661 = x73 & ~n7560 ;
  assign n11662 = n7953 & n11661 ;
  assign n11663 = n11660 | n11662 ;
  assign n11664 = n11659 | n11663 ;
  assign n11665 = n7569 | n11659 ;
  assign n11666 = n11663 | n11665 ;
  assign n11667 = ( n746 & n11664 ) | ( n746 & n11666 ) | ( n11664 & n11666 ) ;
  assign n11668 = x41 & n11666 ;
  assign n11669 = x41 & n11659 ;
  assign n11670 = ( x41 & n11663 ) | ( x41 & n11669 ) | ( n11663 & n11669 ) ;
  assign n11671 = ( n746 & n11668 ) | ( n746 & n11670 ) | ( n11668 & n11670 ) ;
  assign n11672 = x41 & ~n11670 ;
  assign n11673 = x41 & ~n11666 ;
  assign n11674 = ( ~n746 & n11672 ) | ( ~n746 & n11673 ) | ( n11672 & n11673 ) ;
  assign n11675 = ( n11667 & ~n11671 ) | ( n11667 & n11674 ) | ( ~n11671 & n11674 ) ;
  assign n11676 = n11264 | n11271 ;
  assign n11677 = x66 & n11205 ;
  assign n11678 = x65 & n11200 ;
  assign n11679 = ~n10779 & n11204 ;
  assign n11680 = x64 & ~n11199 ;
  assign n11681 = n11679 & n11680 ;
  assign n11682 = n11678 | n11681 ;
  assign n11683 = n11677 | n11682 ;
  assign n11684 = n159 & n11208 ;
  assign n11685 = n11683 | n11684 ;
  assign n11686 = x50 | n11208 ;
  assign n11687 = ( x50 & n159 ) | ( x50 & n11686 ) | ( n159 & n11686 ) ;
  assign n11688 = n11683 | n11687 ;
  assign n11689 = ~x50 & n11687 ;
  assign n11690 = ( ~x50 & n11683 ) | ( ~x50 & n11689 ) | ( n11683 & n11689 ) ;
  assign n11691 = ( ~n11685 & n11688 ) | ( ~n11685 & n11690 ) | ( n11688 & n11690 ) ;
  assign n11692 = n11220 | n11691 ;
  assign n11693 = n11220 & n11691 ;
  assign n11694 = n11692 & ~n11693 ;
  assign n11695 = n293 & n9936 ;
  assign n11696 = x69 & n9933 ;
  assign n11697 = x68 & n9928 ;
  assign n11698 = x67 & ~n9927 ;
  assign n11699 = n10379 & n11698 ;
  assign n11700 = n11697 | n11699 ;
  assign n11701 = n11696 | n11700 ;
  assign n11702 = n11695 | n11701 ;
  assign n11703 = x47 | n11696 ;
  assign n11704 = n11700 | n11703 ;
  assign n11705 = n11695 | n11704 ;
  assign n11706 = ~x47 & n11704 ;
  assign n11707 = ( ~x47 & n11695 ) | ( ~x47 & n11706 ) | ( n11695 & n11706 ) ;
  assign n11708 = ( ~n11702 & n11705 ) | ( ~n11702 & n11707 ) | ( n11705 & n11707 ) ;
  assign n11709 = n11694 & n11708 ;
  assign n11710 = n11694 & ~n11709 ;
  assign n11711 = ~n11694 & n11708 ;
  assign n11712 = n11710 | n11711 ;
  assign n11713 = n11242 | n11244 ;
  assign n11714 = ( n11242 & n11243 ) | ( n11242 & n11713 ) | ( n11243 & n11713 ) ;
  assign n11715 = n11712 & n11714 ;
  assign n11716 = n11712 | n11714 ;
  assign n11717 = ~n11715 & n11716 ;
  assign n11718 = x72 & n8724 ;
  assign n11719 = x71 & n8719 ;
  assign n11720 = x70 & ~n8718 ;
  assign n11721 = n9149 & n11720 ;
  assign n11722 = n11719 | n11721 ;
  assign n11723 = n11718 | n11722 ;
  assign n11724 = ( n513 & n8727 ) | ( n513 & n11723 ) | ( n8727 & n11723 ) ;
  assign n11725 = ( x44 & n8727 ) | ( x44 & ~n11718 ) | ( n8727 & ~n11718 ) ;
  assign n11726 = x44 & n8727 ;
  assign n11727 = ( ~n11722 & n11725 ) | ( ~n11722 & n11726 ) | ( n11725 & n11726 ) ;
  assign n11728 = ( x44 & n513 ) | ( x44 & n11727 ) | ( n513 & n11727 ) ;
  assign n11729 = ~n11724 & n11728 ;
  assign n11730 = n11723 | n11727 ;
  assign n11731 = x44 | n11723 ;
  assign n11732 = ( n513 & n11730 ) | ( n513 & n11731 ) | ( n11730 & n11731 ) ;
  assign n11733 = ( ~x44 & n11729 ) | ( ~x44 & n11732 ) | ( n11729 & n11732 ) ;
  assign n11734 = n11717 & n11733 ;
  assign n11735 = n11717 & ~n11734 ;
  assign n11736 = ~n11717 & n11733 ;
  assign n11737 = n11735 | n11736 ;
  assign n11738 = ~n11676 & n11737 ;
  assign n11739 = n11675 & n11738 ;
  assign n11740 = n11676 & ~n11737 ;
  assign n11741 = ( n11675 & n11739 ) | ( n11675 & n11740 ) | ( n11739 & n11740 ) ;
  assign n11742 = n11675 | n11738 ;
  assign n11743 = n11740 | n11742 ;
  assign n11744 = ~n11741 & n11743 ;
  assign n11745 = n11290 | n11291 ;
  assign n11746 = ( n11196 & n11290 ) | ( n11196 & n11745 ) | ( n11290 & n11745 ) ;
  assign n11747 = n11744 & n11746 ;
  assign n11748 = n11744 | n11746 ;
  assign n11749 = ~n11747 & n11748 ;
  assign n11750 = x78 & n6536 ;
  assign n11751 = x77 & n6531 ;
  assign n11752 = x76 & ~n6530 ;
  assign n11753 = n6871 & n11752 ;
  assign n11754 = n11751 | n11753 ;
  assign n11755 = n11750 | n11754 ;
  assign n11756 = n6539 | n11750 ;
  assign n11757 = n11754 | n11756 ;
  assign n11758 = ( n1192 & n11755 ) | ( n1192 & n11757 ) | ( n11755 & n11757 ) ;
  assign n11759 = x38 & n11757 ;
  assign n11760 = x38 & n11750 ;
  assign n11761 = ( x38 & n11754 ) | ( x38 & n11760 ) | ( n11754 & n11760 ) ;
  assign n11762 = ( n1192 & n11759 ) | ( n1192 & n11761 ) | ( n11759 & n11761 ) ;
  assign n11763 = x38 & ~n11761 ;
  assign n11764 = x38 & ~n11757 ;
  assign n11765 = ( ~n1192 & n11763 ) | ( ~n1192 & n11764 ) | ( n11763 & n11764 ) ;
  assign n11766 = ( n11758 & ~n11762 ) | ( n11758 & n11765 ) | ( ~n11762 & n11765 ) ;
  assign n11767 = n11749 & n11766 ;
  assign n11768 = n11749 & ~n11767 ;
  assign n11769 = ~n11749 & n11766 ;
  assign n11770 = n11768 | n11769 ;
  assign n11771 = n11315 | n11318 ;
  assign n11772 = ( n11315 & n11320 ) | ( n11315 & n11771 ) | ( n11320 & n11771 ) ;
  assign n11773 = n11770 & n11772 ;
  assign n11774 = n11770 | n11772 ;
  assign n11775 = ~n11773 & n11774 ;
  assign n11776 = x81 & n5554 ;
  assign n11777 = x80 & n5549 ;
  assign n11778 = x79 & ~n5548 ;
  assign n11779 = n5893 & n11778 ;
  assign n11780 = n11777 | n11779 ;
  assign n11781 = n11776 | n11780 ;
  assign n11782 = n5557 | n11776 ;
  assign n11783 = n11780 | n11782 ;
  assign n11784 = ( n1651 & n11781 ) | ( n1651 & n11783 ) | ( n11781 & n11783 ) ;
  assign n11785 = x35 & n11783 ;
  assign n11786 = x35 & n11776 ;
  assign n11787 = ( x35 & n11780 ) | ( x35 & n11786 ) | ( n11780 & n11786 ) ;
  assign n11788 = ( n1651 & n11785 ) | ( n1651 & n11787 ) | ( n11785 & n11787 ) ;
  assign n11789 = x35 & ~n11787 ;
  assign n11790 = x35 & ~n11783 ;
  assign n11791 = ( ~n1651 & n11789 ) | ( ~n1651 & n11790 ) | ( n11789 & n11790 ) ;
  assign n11792 = ( n11784 & ~n11788 ) | ( n11784 & n11791 ) | ( ~n11788 & n11791 ) ;
  assign n11793 = n11775 & n11792 ;
  assign n11794 = n11775 & ~n11793 ;
  assign n11795 = ~n11775 & n11792 ;
  assign n11796 = n11794 | n11795 ;
  assign n11797 = n11658 & n11796 ;
  assign n11798 = n11658 & ~n11797 ;
  assign n11799 = ~n11658 & n11796 ;
  assign n11800 = n11798 | n11799 ;
  assign n11801 = x84 & n4631 ;
  assign n11802 = x83 & n4626 ;
  assign n11803 = x82 & ~n4625 ;
  assign n11804 = n4943 & n11803 ;
  assign n11805 = n11802 | n11804 ;
  assign n11806 = n11801 | n11805 ;
  assign n11807 = n4634 | n11801 ;
  assign n11808 = n11805 | n11807 ;
  assign n11809 = ( n2194 & n11806 ) | ( n2194 & n11808 ) | ( n11806 & n11808 ) ;
  assign n11810 = x32 & n11808 ;
  assign n11811 = x32 & n11801 ;
  assign n11812 = ( x32 & n11805 ) | ( x32 & n11811 ) | ( n11805 & n11811 ) ;
  assign n11813 = ( n2194 & n11810 ) | ( n2194 & n11812 ) | ( n11810 & n11812 ) ;
  assign n11814 = x32 & ~n11812 ;
  assign n11815 = x32 & ~n11808 ;
  assign n11816 = ( ~n2194 & n11814 ) | ( ~n2194 & n11815 ) | ( n11814 & n11815 ) ;
  assign n11817 = ( n11809 & ~n11813 ) | ( n11809 & n11816 ) | ( ~n11813 & n11816 ) ;
  assign n11818 = n11796 & n11817 ;
  assign n11819 = ~n11658 & n11818 ;
  assign n11820 = ( n11798 & n11817 ) | ( n11798 & n11819 ) | ( n11817 & n11819 ) ;
  assign n11821 = n11800 & ~n11820 ;
  assign n11822 = ~n11796 & n11817 ;
  assign n11823 = ( n11658 & n11817 ) | ( n11658 & n11822 ) | ( n11817 & n11822 ) ;
  assign n11824 = ~n11798 & n11823 ;
  assign n11825 = n11821 | n11824 ;
  assign n11826 = n11366 | n11372 ;
  assign n11827 = n11825 | n11826 ;
  assign n11828 = n11825 & n11826 ;
  assign n11829 = n11827 & ~n11828 ;
  assign n11830 = x87 & n3816 ;
  assign n11831 = x86 & n3811 ;
  assign n11832 = x85 & ~n3810 ;
  assign n11833 = n4067 & n11832 ;
  assign n11834 = n11831 | n11833 ;
  assign n11835 = n11830 | n11834 ;
  assign n11836 = n3819 | n11830 ;
  assign n11837 = n11834 | n11836 ;
  assign n11838 = ( n2816 & n11835 ) | ( n2816 & n11837 ) | ( n11835 & n11837 ) ;
  assign n11839 = x29 & n11837 ;
  assign n11840 = x29 & n11830 ;
  assign n11841 = ( x29 & n11834 ) | ( x29 & n11840 ) | ( n11834 & n11840 ) ;
  assign n11842 = ( n2816 & n11839 ) | ( n2816 & n11841 ) | ( n11839 & n11841 ) ;
  assign n11843 = x29 & ~n11841 ;
  assign n11844 = x29 & ~n11837 ;
  assign n11845 = ( ~n2816 & n11843 ) | ( ~n2816 & n11844 ) | ( n11843 & n11844 ) ;
  assign n11846 = ( n11838 & ~n11842 ) | ( n11838 & n11845 ) | ( ~n11842 & n11845 ) ;
  assign n11847 = n11829 & n11846 ;
  assign n11848 = n11829 | n11846 ;
  assign n11849 = ~n11847 & n11848 ;
  assign n11850 = n11391 & n11846 ;
  assign n11851 = ( n11391 & n11829 ) | ( n11391 & n11850 ) | ( n11829 & n11850 ) ;
  assign n11852 = ~n11847 & n11851 ;
  assign n11853 = ( n11397 & n11849 ) | ( n11397 & n11852 ) | ( n11849 & n11852 ) ;
  assign n11854 = n11657 & ~n11853 ;
  assign n11855 = x90 & n3085 ;
  assign n11856 = x89 & n3080 ;
  assign n11857 = x88 & ~n3079 ;
  assign n11858 = n3309 & n11857 ;
  assign n11859 = n11856 | n11858 ;
  assign n11860 = n11855 | n11859 ;
  assign n11861 = n3088 | n11855 ;
  assign n11862 = n11859 | n11861 ;
  assign n11863 = ( n3519 & n11860 ) | ( n3519 & n11862 ) | ( n11860 & n11862 ) ;
  assign n11864 = x26 & n11862 ;
  assign n11865 = x26 & n11855 ;
  assign n11866 = ( x26 & n11859 ) | ( x26 & n11865 ) | ( n11859 & n11865 ) ;
  assign n11867 = ( n3519 & n11864 ) | ( n3519 & n11866 ) | ( n11864 & n11866 ) ;
  assign n11868 = x26 & ~n11866 ;
  assign n11869 = x26 & ~n11862 ;
  assign n11870 = ( ~n3519 & n11868 ) | ( ~n3519 & n11869 ) | ( n11868 & n11869 ) ;
  assign n11871 = ( n11863 & ~n11867 ) | ( n11863 & n11870 ) | ( ~n11867 & n11870 ) ;
  assign n11872 = ( n11397 & n11848 ) | ( n11397 & n11851 ) | ( n11848 & n11851 ) ;
  assign n11873 = n11849 & n11871 ;
  assign n11874 = ~n11872 & n11873 ;
  assign n11875 = ( n11854 & n11871 ) | ( n11854 & n11874 ) | ( n11871 & n11874 ) ;
  assign n11876 = n11849 | n11871 ;
  assign n11877 = ( n11871 & ~n11872 ) | ( n11871 & n11876 ) | ( ~n11872 & n11876 ) ;
  assign n11878 = n11854 | n11877 ;
  assign n11879 = ~n11875 & n11878 ;
  assign n11880 = n11416 | n11420 ;
  assign n11881 = ( n11416 & n11419 ) | ( n11416 & n11880 ) | ( n11419 & n11880 ) ;
  assign n11882 = n11879 & n11881 ;
  assign n11883 = n11879 | n11881 ;
  assign n11884 = ~n11882 & n11883 ;
  assign n11885 = x93 & n2429 ;
  assign n11886 = x92 & n2424 ;
  assign n11887 = x91 & ~n2423 ;
  assign n11888 = n2631 & n11887 ;
  assign n11889 = n11886 | n11888 ;
  assign n11890 = n11885 | n11889 ;
  assign n11891 = n2432 | n11885 ;
  assign n11892 = n11889 | n11891 ;
  assign n11893 = ( n4305 & n11890 ) | ( n4305 & n11892 ) | ( n11890 & n11892 ) ;
  assign n11894 = x23 & n11892 ;
  assign n11895 = x23 & n11885 ;
  assign n11896 = ( x23 & n11889 ) | ( x23 & n11895 ) | ( n11889 & n11895 ) ;
  assign n11897 = ( n4305 & n11894 ) | ( n4305 & n11896 ) | ( n11894 & n11896 ) ;
  assign n11898 = x23 & ~n11896 ;
  assign n11899 = x23 & ~n11892 ;
  assign n11900 = ( ~n4305 & n11898 ) | ( ~n4305 & n11899 ) | ( n11898 & n11899 ) ;
  assign n11901 = ( n11893 & ~n11897 ) | ( n11893 & n11900 ) | ( ~n11897 & n11900 ) ;
  assign n11902 = n11884 | n11901 ;
  assign n11903 = n11884 & n11901 ;
  assign n11904 = n11902 & ~n11903 ;
  assign n11905 = n11441 & n11904 ;
  assign n11906 = ( n11445 & n11904 ) | ( n11445 & n11905 ) | ( n11904 & n11905 ) ;
  assign n11907 = n11441 | n11904 ;
  assign n11908 = n11445 | n11907 ;
  assign n11909 = ~n11906 & n11908 ;
  assign n11910 = x96 & n1859 ;
  assign n11911 = x95 & n1854 ;
  assign n11912 = x94 & ~n1853 ;
  assign n11913 = n2037 & n11912 ;
  assign n11914 = n11911 | n11913 ;
  assign n11915 = n11910 | n11914 ;
  assign n11916 = n1862 | n11910 ;
  assign n11917 = n11914 | n11916 ;
  assign n11918 = ( n5202 & n11915 ) | ( n5202 & n11917 ) | ( n11915 & n11917 ) ;
  assign n11919 = x20 & n11917 ;
  assign n11920 = x20 & n11910 ;
  assign n11921 = ( x20 & n11914 ) | ( x20 & n11920 ) | ( n11914 & n11920 ) ;
  assign n11922 = ( n5202 & n11919 ) | ( n5202 & n11921 ) | ( n11919 & n11921 ) ;
  assign n11923 = x20 & ~n11921 ;
  assign n11924 = x20 & ~n11917 ;
  assign n11925 = ( ~n5202 & n11923 ) | ( ~n5202 & n11924 ) | ( n11923 & n11924 ) ;
  assign n11926 = ( n11918 & ~n11922 ) | ( n11918 & n11925 ) | ( ~n11922 & n11925 ) ;
  assign n11927 = n11909 | n11926 ;
  assign n11928 = n11909 & n11926 ;
  assign n11929 = n11927 & ~n11928 ;
  assign n11930 = n11467 & n11929 ;
  assign n11931 = ( n11473 & n11929 ) | ( n11473 & n11930 ) | ( n11929 & n11930 ) ;
  assign n11932 = n11467 | n11929 ;
  assign n11933 = n11473 | n11932 ;
  assign n11934 = ~n11931 & n11933 ;
  assign n11935 = x99 & n1383 ;
  assign n11936 = x98 & n1378 ;
  assign n11937 = x97 & ~n1377 ;
  assign n11938 = n1542 & n11937 ;
  assign n11939 = n11936 | n11938 ;
  assign n11940 = n11935 | n11939 ;
  assign n11941 = n1386 | n11935 ;
  assign n11942 = n11939 | n11941 ;
  assign n11943 = ( n6164 & n11940 ) | ( n6164 & n11942 ) | ( n11940 & n11942 ) ;
  assign n11944 = x17 & n11942 ;
  assign n11945 = x17 & n11935 ;
  assign n11946 = ( x17 & n11939 ) | ( x17 & n11945 ) | ( n11939 & n11945 ) ;
  assign n11947 = ( n6164 & n11944 ) | ( n6164 & n11946 ) | ( n11944 & n11946 ) ;
  assign n11948 = x17 & ~n11946 ;
  assign n11949 = x17 & ~n11942 ;
  assign n11950 = ( ~n6164 & n11948 ) | ( ~n6164 & n11949 ) | ( n11948 & n11949 ) ;
  assign n11951 = ( n11943 & ~n11947 ) | ( n11943 & n11950 ) | ( ~n11947 & n11950 ) ;
  assign n11952 = n11934 & n11951 ;
  assign n11953 = n11934 & ~n11952 ;
  assign n11954 = ~n11934 & n11951 ;
  assign n11955 = n11953 | n11954 ;
  assign n11956 = n11500 | n11507 ;
  assign n11957 = n11955 | n11956 ;
  assign n11958 = n11955 & n11956 ;
  assign n11959 = n11957 & ~n11958 ;
  assign n11960 = x102 & n962 ;
  assign n11961 = x101 & n957 ;
  assign n11962 = x100 & ~n956 ;
  assign n11963 = n1105 & n11962 ;
  assign n11964 = n11961 | n11963 ;
  assign n11965 = n11960 | n11964 ;
  assign n11966 = n965 | n11960 ;
  assign n11967 = n11964 | n11966 ;
  assign n11968 = ( n7178 & n11965 ) | ( n7178 & n11967 ) | ( n11965 & n11967 ) ;
  assign n11969 = x14 & n11967 ;
  assign n11970 = x14 & n11960 ;
  assign n11971 = ( x14 & n11964 ) | ( x14 & n11970 ) | ( n11964 & n11970 ) ;
  assign n11972 = ( n7178 & n11969 ) | ( n7178 & n11971 ) | ( n11969 & n11971 ) ;
  assign n11973 = x14 & ~n11971 ;
  assign n11974 = x14 & ~n11967 ;
  assign n11975 = ( ~n7178 & n11973 ) | ( ~n7178 & n11974 ) | ( n11973 & n11974 ) ;
  assign n11976 = ( n11968 & ~n11972 ) | ( n11968 & n11975 ) | ( ~n11972 & n11975 ) ;
  assign n11977 = n11959 & n11976 ;
  assign n11978 = n11959 & ~n11977 ;
  assign n11979 = ~n11959 & n11976 ;
  assign n11980 = n11978 | n11979 ;
  assign n11981 = n11528 | n11536 ;
  assign n11982 = n11980 | n11981 ;
  assign n11983 = n11980 & n11981 ;
  assign n11984 = n11982 & ~n11983 ;
  assign n11985 = x105 & n636 ;
  assign n11986 = x104 & n631 ;
  assign n11987 = x103 & ~n630 ;
  assign n11988 = n764 & n11987 ;
  assign n11989 = n11986 | n11988 ;
  assign n11990 = n11985 | n11989 ;
  assign n11991 = n639 | n11985 ;
  assign n11992 = n11989 | n11991 ;
  assign n11993 = ( n8273 & n11990 ) | ( n8273 & n11992 ) | ( n11990 & n11992 ) ;
  assign n11994 = x11 & n11992 ;
  assign n11995 = x11 & n11985 ;
  assign n11996 = ( x11 & n11989 ) | ( x11 & n11995 ) | ( n11989 & n11995 ) ;
  assign n11997 = ( n8273 & n11994 ) | ( n8273 & n11996 ) | ( n11994 & n11996 ) ;
  assign n11998 = x11 & ~n11996 ;
  assign n11999 = x11 & ~n11992 ;
  assign n12000 = ( ~n8273 & n11998 ) | ( ~n8273 & n11999 ) | ( n11998 & n11999 ) ;
  assign n12001 = ( n11993 & ~n11997 ) | ( n11993 & n12000 ) | ( ~n11997 & n12000 ) ;
  assign n12002 = n11984 & n12001 ;
  assign n12003 = n11984 & ~n12002 ;
  assign n12004 = ~n11984 & n12001 ;
  assign n12005 = n12003 | n12004 ;
  assign n12006 = n11555 | n11562 ;
  assign n12007 = n12005 | n12006 ;
  assign n12008 = n12005 & n12006 ;
  assign n12009 = n12007 & ~n12008 ;
  assign n12010 = x108 & n389 ;
  assign n12011 = x107 & n384 ;
  assign n12012 = x106 & ~n383 ;
  assign n12013 = n463 & n12012 ;
  assign n12014 = n12011 | n12013 ;
  assign n12015 = n12010 | n12014 ;
  assign n12016 = n392 | n12010 ;
  assign n12017 = n12014 | n12016 ;
  assign n12018 = ( n9479 & n12015 ) | ( n9479 & n12017 ) | ( n12015 & n12017 ) ;
  assign n12019 = x8 & n12017 ;
  assign n12020 = x8 & n12010 ;
  assign n12021 = ( x8 & n12014 ) | ( x8 & n12020 ) | ( n12014 & n12020 ) ;
  assign n12022 = ( n9479 & n12019 ) | ( n9479 & n12021 ) | ( n12019 & n12021 ) ;
  assign n12023 = x8 & ~n12021 ;
  assign n12024 = x8 & ~n12017 ;
  assign n12025 = ( ~n9479 & n12023 ) | ( ~n9479 & n12024 ) | ( n12023 & n12024 ) ;
  assign n12026 = ( n12018 & ~n12022 ) | ( n12018 & n12025 ) | ( ~n12022 & n12025 ) ;
  assign n12027 = n12009 | n12026 ;
  assign n12028 = n12009 & n12026 ;
  assign n12029 = n12027 & ~n12028 ;
  assign n12030 = n11581 | n11586 ;
  assign n12031 = n12028 | n12030 ;
  assign n12032 = ( n12028 & n12029 ) | ( n12028 & n12031 ) | ( n12029 & n12031 ) ;
  assign n12033 = n12027 & ~n12032 ;
  assign n12034 = ~n12029 & n12030 ;
  assign n12035 = n12033 | n12034 ;
  assign n12036 = x111 & n212 ;
  assign n12037 = x110 & n207 ;
  assign n12038 = x109 & ~n206 ;
  assign n12039 = n267 & n12038 ;
  assign n12040 = n12037 | n12039 ;
  assign n12041 = n12036 | n12040 ;
  assign n12042 = n215 | n12036 ;
  assign n12043 = n12040 | n12042 ;
  assign n12044 = ( n10749 & n12041 ) | ( n10749 & n12043 ) | ( n12041 & n12043 ) ;
  assign n12045 = x5 & n12043 ;
  assign n12046 = x5 & n12036 ;
  assign n12047 = ( x5 & n12040 ) | ( x5 & n12046 ) | ( n12040 & n12046 ) ;
  assign n12048 = ( n10749 & n12045 ) | ( n10749 & n12047 ) | ( n12045 & n12047 ) ;
  assign n12049 = x5 & ~n12047 ;
  assign n12050 = x5 & ~n12043 ;
  assign n12051 = ( ~n10749 & n12049 ) | ( ~n10749 & n12050 ) | ( n12049 & n12050 ) ;
  assign n12052 = ( n12044 & ~n12048 ) | ( n12044 & n12051 ) | ( ~n12048 & n12051 ) ;
  assign n12053 = n12030 & n12052 ;
  assign n12054 = ~n12029 & n12053 ;
  assign n12055 = ( n12033 & n12052 ) | ( n12033 & n12054 ) | ( n12052 & n12054 ) ;
  assign n12056 = n12035 & ~n12055 ;
  assign n12057 = ~n12030 & n12052 ;
  assign n12058 = ( n12029 & n12052 ) | ( n12029 & n12057 ) | ( n12052 & n12057 ) ;
  assign n12059 = ~n12033 & n12058 ;
  assign n12060 = n12056 | n12059 ;
  assign n12061 = n11607 | n11613 ;
  assign n12062 = n12060 | n12061 ;
  assign n12063 = n12060 & n12061 ;
  assign n12064 = n12062 & ~n12063 ;
  assign n12065 = x113 | x114 ;
  assign n12066 = x113 & x114 ;
  assign n12067 = n12065 & ~n12066 ;
  assign n12068 = n11616 | n11617 ;
  assign n12069 = ( n11616 & n11618 ) | ( n11616 & n12068 ) | ( n11618 & n12068 ) ;
  assign n12070 = n11158 | n11616 ;
  assign n12071 = ( n11616 & n11617 ) | ( n11616 & n12070 ) | ( n11617 & n12070 ) ;
  assign n12072 = ( n10726 & n12069 ) | ( n10726 & n12071 ) | ( n12069 & n12071 ) ;
  assign n12073 = n12069 | n12071 ;
  assign n12074 = ( n10735 & n12072 ) | ( n10735 & n12073 ) | ( n12072 & n12073 ) ;
  assign n12075 = ( n10736 & n12072 ) | ( n10736 & n12073 ) | ( n12072 & n12073 ) ;
  assign n12076 = ( n6159 & n12074 ) | ( n6159 & n12075 ) | ( n12074 & n12075 ) ;
  assign n12077 = ( n6157 & n12074 ) | ( n6157 & n12075 ) | ( n12074 & n12075 ) ;
  assign n12078 = ( n5823 & n12076 ) | ( n5823 & n12077 ) | ( n12076 & n12077 ) ;
  assign n12079 = n12067 | n12078 ;
  assign n12080 = x113 & n133 ;
  assign n12081 = x112 & ~n162 ;
  assign n12082 = ( n137 & n12080 ) | ( n137 & n12081 ) | ( n12080 & n12081 ) ;
  assign n12083 = x0 & x114 ;
  assign n12084 = ( ~n137 & n12080 ) | ( ~n137 & n12083 ) | ( n12080 & n12083 ) ;
  assign n12085 = n12082 | n12084 ;
  assign n12086 = n141 | n12085 ;
  assign n12087 = n12067 & n12069 ;
  assign n12088 = n12067 & n12071 ;
  assign n12089 = ( n10726 & n12087 ) | ( n10726 & n12088 ) | ( n12087 & n12088 ) ;
  assign n12090 = n12087 | n12088 ;
  assign n12091 = ( n10735 & n12089 ) | ( n10735 & n12090 ) | ( n12089 & n12090 ) ;
  assign n12092 = ( n10736 & n12089 ) | ( n10736 & n12090 ) | ( n12089 & n12090 ) ;
  assign n12093 = ( n6159 & n12091 ) | ( n6159 & n12092 ) | ( n12091 & n12092 ) ;
  assign n12094 = ( n6157 & n12091 ) | ( n6157 & n12092 ) | ( n12091 & n12092 ) ;
  assign n12095 = ( n5823 & n12093 ) | ( n5823 & n12094 ) | ( n12093 & n12094 ) ;
  assign n12096 = ( n12085 & n12086 ) | ( n12085 & ~n12095 ) | ( n12086 & ~n12095 ) ;
  assign n12097 = n12085 & n12086 ;
  assign n12098 = ( n12079 & n12096 ) | ( n12079 & n12097 ) | ( n12096 & n12097 ) ;
  assign n12099 = x2 & n12098 ;
  assign n12100 = x2 & ~n12098 ;
  assign n12101 = ( n12098 & ~n12099 ) | ( n12098 & n12100 ) | ( ~n12099 & n12100 ) ;
  assign n12102 = n12064 & n12101 ;
  assign n12103 = n12064 & ~n12102 ;
  assign n12104 = ~n12064 & n12101 ;
  assign n12105 = n12103 | n12104 ;
  assign n12106 = n11650 | n11654 ;
  assign n12107 = n12105 | n12106 ;
  assign n12108 = n12104 & n12106 ;
  assign n12109 = ( n12103 & n12106 ) | ( n12103 & n12108 ) | ( n12106 & n12108 ) ;
  assign n12110 = n12107 & ~n12109 ;
  assign n12111 = n11767 | n11773 ;
  assign n12112 = n11741 | n11747 ;
  assign n12113 = x50 & ~x51 ;
  assign n12114 = ~x50 & x51 ;
  assign n12115 = n12113 | n12114 ;
  assign n12116 = x64 & n12115 ;
  assign n12117 = ~n11220 & n12116 ;
  assign n12118 = ( ~n11691 & n12116 ) | ( ~n11691 & n12117 ) | ( n12116 & n12117 ) ;
  assign n12119 = n11220 & ~n12116 ;
  assign n12120 = n11691 & n12119 ;
  assign n12121 = n12118 | n12120 ;
  assign n12122 = x67 & n11205 ;
  assign n12123 = x66 & n11200 ;
  assign n12124 = x65 & ~n11199 ;
  assign n12125 = n11679 & n12124 ;
  assign n12126 = n12123 | n12125 ;
  assign n12127 = n12122 | n12126 ;
  assign n12128 = n186 & n11208 ;
  assign n12129 = n12127 | n12128 ;
  assign n12130 = x50 & ~n12129 ;
  assign n12131 = ~x50 & n12129 ;
  assign n12132 = n12130 | n12131 ;
  assign n12133 = n12121 & n12132 ;
  assign n12134 = n12121 | n12132 ;
  assign n12135 = ~n12133 & n12134 ;
  assign n12136 = x69 & n9928 ;
  assign n12137 = x68 & ~n9927 ;
  assign n12138 = n10379 & n12137 ;
  assign n12139 = n12136 | n12138 ;
  assign n12140 = x70 & n9933 ;
  assign n12141 = n9936 | n12140 ;
  assign n12142 = n12139 | n12141 ;
  assign n12143 = x47 & ~n12142 ;
  assign n12144 = x47 & ~n12140 ;
  assign n12145 = ~n12139 & n12144 ;
  assign n12146 = ( ~n340 & n12143 ) | ( ~n340 & n12145 ) | ( n12143 & n12145 ) ;
  assign n12147 = ~x47 & n12142 ;
  assign n12148 = ~x47 & n12140 ;
  assign n12149 = ( ~x47 & n12139 ) | ( ~x47 & n12148 ) | ( n12139 & n12148 ) ;
  assign n12150 = ( n340 & n12147 ) | ( n340 & n12149 ) | ( n12147 & n12149 ) ;
  assign n12151 = n12146 | n12150 ;
  assign n12152 = n12135 & n12151 ;
  assign n12153 = n12135 & ~n12152 ;
  assign n12154 = ~n12135 & n12151 ;
  assign n12155 = n12153 | n12154 ;
  assign n12156 = n11709 | n11714 ;
  assign n12157 = ( n11709 & n11712 ) | ( n11709 & n12156 ) | ( n11712 & n12156 ) ;
  assign n12158 = n12155 | n12157 ;
  assign n12159 = n12155 & n12157 ;
  assign n12160 = n12158 & ~n12159 ;
  assign n12161 = x73 & n8724 ;
  assign n12162 = x72 & n8719 ;
  assign n12163 = x71 & ~n8718 ;
  assign n12164 = n9149 & n12163 ;
  assign n12165 = n12162 | n12164 ;
  assign n12166 = n12161 | n12165 ;
  assign n12167 = ( ~n610 & n8727 ) | ( ~n610 & n12166 ) | ( n8727 & n12166 ) ;
  assign n12168 = n8727 & n12161 ;
  assign n12169 = ( n8727 & n12165 ) | ( n8727 & n12168 ) | ( n12165 & n12168 ) ;
  assign n12170 = ( n598 & n12167 ) | ( n598 & n12169 ) | ( n12167 & n12169 ) ;
  assign n12171 = ( x44 & ~n12166 ) | ( x44 & n12170 ) | ( ~n12166 & n12170 ) ;
  assign n12172 = ~n12170 & n12171 ;
  assign n12173 = x44 | n12161 ;
  assign n12174 = n12165 | n12173 ;
  assign n12175 = n12170 | n12174 ;
  assign n12176 = ( ~x44 & n12172 ) | ( ~x44 & n12175 ) | ( n12172 & n12175 ) ;
  assign n12177 = n12160 | n12176 ;
  assign n12178 = n12160 & n12176 ;
  assign n12179 = n12177 & ~n12178 ;
  assign n12180 = n11676 & n11737 ;
  assign n12181 = n11734 | n12180 ;
  assign n12182 = n12179 & n12181 ;
  assign n12183 = n12179 | n12181 ;
  assign n12184 = ~n12182 & n12183 ;
  assign n12185 = x76 & n7566 ;
  assign n12186 = x75 & n7561 ;
  assign n12187 = x74 & ~n7560 ;
  assign n12188 = n7953 & n12187 ;
  assign n12189 = n12186 | n12188 ;
  assign n12190 = n12185 | n12189 ;
  assign n12191 = n7569 | n12185 ;
  assign n12192 = n12189 | n12191 ;
  assign n12193 = ( n923 & n12190 ) | ( n923 & n12192 ) | ( n12190 & n12192 ) ;
  assign n12194 = x41 & n12192 ;
  assign n12195 = x41 & n12185 ;
  assign n12196 = ( x41 & n12189 ) | ( x41 & n12195 ) | ( n12189 & n12195 ) ;
  assign n12197 = ( n923 & n12194 ) | ( n923 & n12196 ) | ( n12194 & n12196 ) ;
  assign n12198 = x41 & ~n12196 ;
  assign n12199 = x41 & ~n12192 ;
  assign n12200 = ( ~n923 & n12198 ) | ( ~n923 & n12199 ) | ( n12198 & n12199 ) ;
  assign n12201 = ( n12193 & ~n12197 ) | ( n12193 & n12200 ) | ( ~n12197 & n12200 ) ;
  assign n12202 = n12184 & n12201 ;
  assign n12203 = n12184 & ~n12202 ;
  assign n12204 = ~n12184 & n12201 ;
  assign n12205 = n12203 | n12204 ;
  assign n12206 = n12112 & n12205 ;
  assign n12207 = n12112 | n12205 ;
  assign n12208 = ~n12206 & n12207 ;
  assign n12209 = x79 & n6536 ;
  assign n12210 = x78 & n6531 ;
  assign n12211 = x77 & ~n6530 ;
  assign n12212 = n6871 & n12211 ;
  assign n12213 = n12210 | n12212 ;
  assign n12214 = n12209 | n12213 ;
  assign n12215 = n6539 | n12209 ;
  assign n12216 = n12213 | n12215 ;
  assign n12217 = ( n1332 & n12214 ) | ( n1332 & n12216 ) | ( n12214 & n12216 ) ;
  assign n12218 = x38 & n12216 ;
  assign n12219 = x38 & n12209 ;
  assign n12220 = ( x38 & n12213 ) | ( x38 & n12219 ) | ( n12213 & n12219 ) ;
  assign n12221 = ( n1332 & n12218 ) | ( n1332 & n12220 ) | ( n12218 & n12220 ) ;
  assign n12222 = x38 & ~n12220 ;
  assign n12223 = x38 & ~n12216 ;
  assign n12224 = ( ~n1332 & n12222 ) | ( ~n1332 & n12223 ) | ( n12222 & n12223 ) ;
  assign n12225 = ( n12217 & ~n12221 ) | ( n12217 & n12224 ) | ( ~n12221 & n12224 ) ;
  assign n12226 = n12208 & n12225 ;
  assign n12227 = n12208 | n12225 ;
  assign n12228 = ~n12226 & n12227 ;
  assign n12229 = n12111 & n12228 ;
  assign n12230 = n12111 | n12228 ;
  assign n12231 = ~n12229 & n12230 ;
  assign n12232 = x82 & n5554 ;
  assign n12233 = x81 & n5549 ;
  assign n12234 = x80 & ~n5548 ;
  assign n12235 = n5893 & n12234 ;
  assign n12236 = n12233 | n12235 ;
  assign n12237 = n12232 | n12236 ;
  assign n12238 = n5557 | n12232 ;
  assign n12239 = n12236 | n12238 ;
  assign n12240 = ( n1811 & n12237 ) | ( n1811 & n12239 ) | ( n12237 & n12239 ) ;
  assign n12241 = x35 & n12239 ;
  assign n12242 = x35 & n12232 ;
  assign n12243 = ( x35 & n12236 ) | ( x35 & n12242 ) | ( n12236 & n12242 ) ;
  assign n12244 = ( n1811 & n12241 ) | ( n1811 & n12243 ) | ( n12241 & n12243 ) ;
  assign n12245 = x35 & ~n12243 ;
  assign n12246 = x35 & ~n12239 ;
  assign n12247 = ( ~n1811 & n12245 ) | ( ~n1811 & n12246 ) | ( n12245 & n12246 ) ;
  assign n12248 = ( n12240 & ~n12244 ) | ( n12240 & n12247 ) | ( ~n12244 & n12247 ) ;
  assign n12249 = n12231 & n12248 ;
  assign n12250 = n12231 | n12248 ;
  assign n12251 = ~n12249 & n12250 ;
  assign n12252 = n11793 | n11795 ;
  assign n12253 = n11794 | n12252 ;
  assign n12254 = ( n11658 & n11793 ) | ( n11658 & n12253 ) | ( n11793 & n12253 ) ;
  assign n12255 = n12251 & n12254 ;
  assign n12256 = n12251 | n12254 ;
  assign n12257 = ~n12255 & n12256 ;
  assign n12258 = x85 & n4631 ;
  assign n12259 = x84 & n4626 ;
  assign n12260 = x83 & ~n4625 ;
  assign n12261 = n4943 & n12260 ;
  assign n12262 = n12259 | n12261 ;
  assign n12263 = n12258 | n12262 ;
  assign n12264 = n4634 | n12258 ;
  assign n12265 = n12262 | n12264 ;
  assign n12266 = ( n2381 & n12263 ) | ( n2381 & n12265 ) | ( n12263 & n12265 ) ;
  assign n12267 = x32 & n12265 ;
  assign n12268 = x32 & n12258 ;
  assign n12269 = ( x32 & n12262 ) | ( x32 & n12268 ) | ( n12262 & n12268 ) ;
  assign n12270 = ( n2381 & n12267 ) | ( n2381 & n12269 ) | ( n12267 & n12269 ) ;
  assign n12271 = x32 & ~n12269 ;
  assign n12272 = x32 & ~n12265 ;
  assign n12273 = ( ~n2381 & n12271 ) | ( ~n2381 & n12272 ) | ( n12271 & n12272 ) ;
  assign n12274 = ( n12266 & ~n12270 ) | ( n12266 & n12273 ) | ( ~n12270 & n12273 ) ;
  assign n12275 = n12257 & n12274 ;
  assign n12276 = n12257 & ~n12275 ;
  assign n12277 = ~n12257 & n12274 ;
  assign n12278 = n12276 | n12277 ;
  assign n12279 = n11820 | n11828 ;
  assign n12280 = n12278 | n12279 ;
  assign n12281 = n12278 & n12279 ;
  assign n12282 = n12280 & ~n12281 ;
  assign n12283 = x88 & n3816 ;
  assign n12284 = x87 & n3811 ;
  assign n12285 = x86 & ~n3810 ;
  assign n12286 = n4067 & n12285 ;
  assign n12287 = n12284 | n12286 ;
  assign n12288 = n12283 | n12287 ;
  assign n12289 = n3819 | n12283 ;
  assign n12290 = n12287 | n12289 ;
  assign n12291 = ( ~n3039 & n12288 ) | ( ~n3039 & n12290 ) | ( n12288 & n12290 ) ;
  assign n12292 = n12288 & n12290 ;
  assign n12293 = ( n3023 & n12291 ) | ( n3023 & n12292 ) | ( n12291 & n12292 ) ;
  assign n12294 = x29 & n12290 ;
  assign n12295 = x29 & n12283 ;
  assign n12296 = ( x29 & n12287 ) | ( x29 & n12295 ) | ( n12287 & n12295 ) ;
  assign n12297 = ( ~n3039 & n12294 ) | ( ~n3039 & n12296 ) | ( n12294 & n12296 ) ;
  assign n12298 = n12294 & n12296 ;
  assign n12299 = ( n3023 & n12297 ) | ( n3023 & n12298 ) | ( n12297 & n12298 ) ;
  assign n12300 = x29 & ~n12296 ;
  assign n12301 = x29 & ~n12290 ;
  assign n12302 = ( n3039 & n12300 ) | ( n3039 & n12301 ) | ( n12300 & n12301 ) ;
  assign n12303 = n12300 | n12301 ;
  assign n12304 = ( ~n3023 & n12302 ) | ( ~n3023 & n12303 ) | ( n12302 & n12303 ) ;
  assign n12305 = ( n12293 & ~n12299 ) | ( n12293 & n12304 ) | ( ~n12299 & n12304 ) ;
  assign n12306 = n12282 | n12305 ;
  assign n12307 = n12282 & n12305 ;
  assign n12308 = n12306 & ~n12307 ;
  assign n12309 = n11847 | n11851 ;
  assign n12310 = n11847 | n11848 ;
  assign n12311 = ( n11397 & n12309 ) | ( n11397 & n12310 ) | ( n12309 & n12310 ) ;
  assign n12312 = n12308 & n12311 ;
  assign n12313 = n12308 | n12311 ;
  assign n12314 = ~n12312 & n12313 ;
  assign n12315 = x91 & n3085 ;
  assign n12316 = x90 & n3080 ;
  assign n12317 = x89 & ~n3079 ;
  assign n12318 = n3309 & n12317 ;
  assign n12319 = n12316 | n12318 ;
  assign n12320 = n12315 | n12319 ;
  assign n12321 = n3088 | n12315 ;
  assign n12322 = n12319 | n12321 ;
  assign n12323 = ( n3768 & n12320 ) | ( n3768 & n12322 ) | ( n12320 & n12322 ) ;
  assign n12324 = x26 & n12322 ;
  assign n12325 = x26 & n12315 ;
  assign n12326 = ( x26 & n12319 ) | ( x26 & n12325 ) | ( n12319 & n12325 ) ;
  assign n12327 = ( n3768 & n12324 ) | ( n3768 & n12326 ) | ( n12324 & n12326 ) ;
  assign n12328 = x26 & ~n12326 ;
  assign n12329 = x26 & ~n12322 ;
  assign n12330 = ( ~n3768 & n12328 ) | ( ~n3768 & n12329 ) | ( n12328 & n12329 ) ;
  assign n12331 = ( n12323 & ~n12327 ) | ( n12323 & n12330 ) | ( ~n12327 & n12330 ) ;
  assign n12332 = n12314 & n12331 ;
  assign n12333 = n12314 & ~n12332 ;
  assign n12334 = ~n12314 & n12331 ;
  assign n12335 = n12333 | n12334 ;
  assign n12336 = n11875 | n11879 ;
  assign n12337 = ( n11875 & n11881 ) | ( n11875 & n12336 ) | ( n11881 & n12336 ) ;
  assign n12338 = ~n12335 & n12337 ;
  assign n12339 = n12335 & ~n12337 ;
  assign n12340 = n12338 | n12339 ;
  assign n12341 = x94 & n2429 ;
  assign n12342 = x93 & n2424 ;
  assign n12343 = x92 & ~n2423 ;
  assign n12344 = n2631 & n12343 ;
  assign n12345 = n12342 | n12344 ;
  assign n12346 = n12341 | n12345 ;
  assign n12347 = n2432 | n12341 ;
  assign n12348 = n12345 | n12347 ;
  assign n12349 = ( n4583 & n12346 ) | ( n4583 & n12348 ) | ( n12346 & n12348 ) ;
  assign n12350 = x23 & n12348 ;
  assign n12351 = x23 & n12341 ;
  assign n12352 = ( x23 & n12345 ) | ( x23 & n12351 ) | ( n12345 & n12351 ) ;
  assign n12353 = ( n4583 & n12350 ) | ( n4583 & n12352 ) | ( n12350 & n12352 ) ;
  assign n12354 = x23 & ~n12352 ;
  assign n12355 = x23 & ~n12348 ;
  assign n12356 = ( ~n4583 & n12354 ) | ( ~n4583 & n12355 ) | ( n12354 & n12355 ) ;
  assign n12357 = ( n12349 & ~n12353 ) | ( n12349 & n12356 ) | ( ~n12353 & n12356 ) ;
  assign n12358 = n12340 & n12357 ;
  assign n12359 = n12340 | n12357 ;
  assign n12360 = ~n12358 & n12359 ;
  assign n12361 = n11445 | n11903 ;
  assign n12362 = n11903 | n11904 ;
  assign n12363 = ( n11905 & n12361 ) | ( n11905 & n12362 ) | ( n12361 & n12362 ) ;
  assign n12364 = n12360 & n12363 ;
  assign n12365 = n12360 | n12363 ;
  assign n12366 = ~n12364 & n12365 ;
  assign n12367 = x97 & n1859 ;
  assign n12368 = x96 & n1854 ;
  assign n12369 = x95 & ~n1853 ;
  assign n12370 = n2037 & n12369 ;
  assign n12371 = n12368 | n12370 ;
  assign n12372 = n12367 | n12371 ;
  assign n12373 = n1862 | n12367 ;
  assign n12374 = n12371 | n12373 ;
  assign n12375 = ( n5505 & n12372 ) | ( n5505 & n12374 ) | ( n12372 & n12374 ) ;
  assign n12376 = x20 & n12374 ;
  assign n12377 = x20 & n12367 ;
  assign n12378 = ( x20 & n12371 ) | ( x20 & n12377 ) | ( n12371 & n12377 ) ;
  assign n12379 = ( n5505 & n12376 ) | ( n5505 & n12378 ) | ( n12376 & n12378 ) ;
  assign n12380 = x20 & ~n12378 ;
  assign n12381 = x20 & ~n12374 ;
  assign n12382 = ( ~n5505 & n12380 ) | ( ~n5505 & n12381 ) | ( n12380 & n12381 ) ;
  assign n12383 = ( n12375 & ~n12379 ) | ( n12375 & n12382 ) | ( ~n12379 & n12382 ) ;
  assign n12384 = n12366 & n12383 ;
  assign n12385 = n12366 & ~n12384 ;
  assign n12386 = ~n12366 & n12383 ;
  assign n12387 = n12385 | n12386 ;
  assign n12388 = n11928 | n11929 ;
  assign n12389 = n11473 | n11928 ;
  assign n12390 = ( n11930 & n12388 ) | ( n11930 & n12389 ) | ( n12388 & n12389 ) ;
  assign n12391 = ~n12387 & n12390 ;
  assign n12392 = n12387 & ~n12390 ;
  assign n12393 = n12391 | n12392 ;
  assign n12394 = x100 & n1383 ;
  assign n12395 = x99 & n1378 ;
  assign n12396 = x98 & ~n1377 ;
  assign n12397 = n1542 & n12396 ;
  assign n12398 = n12395 | n12397 ;
  assign n12399 = n12394 | n12398 ;
  assign n12400 = n1386 | n12394 ;
  assign n12401 = n12398 | n12400 ;
  assign n12402 = ( n6483 & n12399 ) | ( n6483 & n12401 ) | ( n12399 & n12401 ) ;
  assign n12403 = x17 & n12401 ;
  assign n12404 = x17 & n12394 ;
  assign n12405 = ( x17 & n12398 ) | ( x17 & n12404 ) | ( n12398 & n12404 ) ;
  assign n12406 = ( n6483 & n12403 ) | ( n6483 & n12405 ) | ( n12403 & n12405 ) ;
  assign n12407 = x17 & ~n12405 ;
  assign n12408 = x17 & ~n12401 ;
  assign n12409 = ( ~n6483 & n12407 ) | ( ~n6483 & n12408 ) | ( n12407 & n12408 ) ;
  assign n12410 = ( n12402 & ~n12406 ) | ( n12402 & n12409 ) | ( ~n12406 & n12409 ) ;
  assign n12411 = n12393 & n12410 ;
  assign n12412 = n12393 | n12410 ;
  assign n12413 = ~n12411 & n12412 ;
  assign n12414 = n11952 | n11956 ;
  assign n12415 = ( n11952 & n11955 ) | ( n11952 & n12414 ) | ( n11955 & n12414 ) ;
  assign n12416 = n12413 | n12415 ;
  assign n12417 = n12413 & n12415 ;
  assign n12418 = n12416 & ~n12417 ;
  assign n12419 = x103 & n962 ;
  assign n12420 = x102 & n957 ;
  assign n12421 = x101 & ~n956 ;
  assign n12422 = n1105 & n12421 ;
  assign n12423 = n12420 | n12422 ;
  assign n12424 = n12419 | n12423 ;
  assign n12425 = n965 | n12419 ;
  assign n12426 = n12423 | n12425 ;
  assign n12427 = ( n7529 & n12424 ) | ( n7529 & n12426 ) | ( n12424 & n12426 ) ;
  assign n12428 = x14 & n12426 ;
  assign n12429 = x14 & n12419 ;
  assign n12430 = ( x14 & n12423 ) | ( x14 & n12429 ) | ( n12423 & n12429 ) ;
  assign n12431 = ( n7529 & n12428 ) | ( n7529 & n12430 ) | ( n12428 & n12430 ) ;
  assign n12432 = x14 & ~n12430 ;
  assign n12433 = x14 & ~n12426 ;
  assign n12434 = ( ~n7529 & n12432 ) | ( ~n7529 & n12433 ) | ( n12432 & n12433 ) ;
  assign n12435 = ( n12427 & ~n12431 ) | ( n12427 & n12434 ) | ( ~n12431 & n12434 ) ;
  assign n12436 = n12418 & n12435 ;
  assign n12437 = n12418 & ~n12436 ;
  assign n12438 = ~n12418 & n12435 ;
  assign n12439 = n12437 | n12438 ;
  assign n12440 = n11977 | n11981 ;
  assign n12441 = ( n11977 & n11980 ) | ( n11977 & n12440 ) | ( n11980 & n12440 ) ;
  assign n12442 = n12439 | n12441 ;
  assign n12443 = n12439 & n12441 ;
  assign n12444 = n12442 & ~n12443 ;
  assign n12445 = x106 & n636 ;
  assign n12446 = x105 & n631 ;
  assign n12447 = x104 & ~n630 ;
  assign n12448 = n764 & n12447 ;
  assign n12449 = n12446 | n12448 ;
  assign n12450 = n12445 | n12449 ;
  assign n12451 = n639 | n12445 ;
  assign n12452 = n12449 | n12451 ;
  assign n12453 = ( n8656 & n12450 ) | ( n8656 & n12452 ) | ( n12450 & n12452 ) ;
  assign n12454 = x11 & n12452 ;
  assign n12455 = x11 & n12445 ;
  assign n12456 = ( x11 & n12449 ) | ( x11 & n12455 ) | ( n12449 & n12455 ) ;
  assign n12457 = ( n8656 & n12454 ) | ( n8656 & n12456 ) | ( n12454 & n12456 ) ;
  assign n12458 = x11 & ~n12456 ;
  assign n12459 = x11 & ~n12452 ;
  assign n12460 = ( ~n8656 & n12458 ) | ( ~n8656 & n12459 ) | ( n12458 & n12459 ) ;
  assign n12461 = ( n12453 & ~n12457 ) | ( n12453 & n12460 ) | ( ~n12457 & n12460 ) ;
  assign n12462 = n12444 | n12461 ;
  assign n12463 = n12444 & n12461 ;
  assign n12464 = n12462 & ~n12463 ;
  assign n12465 = n12002 | n12006 ;
  assign n12466 = ( n12002 & n12005 ) | ( n12002 & n12465 ) | ( n12005 & n12465 ) ;
  assign n12467 = n12464 & n12466 ;
  assign n12468 = n12464 | n12466 ;
  assign n12469 = ~n12467 & n12468 ;
  assign n12470 = x109 & n389 ;
  assign n12471 = x108 & n384 ;
  assign n12472 = x107 & ~n383 ;
  assign n12473 = n463 & n12472 ;
  assign n12474 = n12471 | n12473 ;
  assign n12475 = n12470 | n12474 ;
  assign n12476 = n392 | n12470 ;
  assign n12477 = n12474 | n12476 ;
  assign n12478 = ( n9878 & n12475 ) | ( n9878 & n12477 ) | ( n12475 & n12477 ) ;
  assign n12479 = x8 & n12477 ;
  assign n12480 = x8 & n12470 ;
  assign n12481 = ( x8 & n12474 ) | ( x8 & n12480 ) | ( n12474 & n12480 ) ;
  assign n12482 = ( n9878 & n12479 ) | ( n9878 & n12481 ) | ( n12479 & n12481 ) ;
  assign n12483 = x8 & ~n12481 ;
  assign n12484 = x8 & ~n12477 ;
  assign n12485 = ( ~n9878 & n12483 ) | ( ~n9878 & n12484 ) | ( n12483 & n12484 ) ;
  assign n12486 = ( n12478 & ~n12482 ) | ( n12478 & n12485 ) | ( ~n12482 & n12485 ) ;
  assign n12487 = n12469 & n12486 ;
  assign n12488 = n12469 & ~n12487 ;
  assign n12489 = ~n12469 & n12486 ;
  assign n12490 = n12488 | n12489 ;
  assign n12491 = n12032 & ~n12490 ;
  assign n12492 = ~n12032 & n12490 ;
  assign n12493 = n12491 | n12492 ;
  assign n12494 = x112 & n212 ;
  assign n12495 = x111 & n207 ;
  assign n12496 = x110 & ~n206 ;
  assign n12497 = n267 & n12496 ;
  assign n12498 = n12495 | n12497 ;
  assign n12499 = n12494 | n12498 ;
  assign n12500 = n215 | n12494 ;
  assign n12501 = n12498 | n12500 ;
  assign n12502 = ( n11172 & n12499 ) | ( n11172 & n12501 ) | ( n12499 & n12501 ) ;
  assign n12503 = x5 & n12501 ;
  assign n12504 = x5 & n12494 ;
  assign n12505 = ( x5 & n12498 ) | ( x5 & n12504 ) | ( n12498 & n12504 ) ;
  assign n12506 = ( n11172 & n12503 ) | ( n11172 & n12505 ) | ( n12503 & n12505 ) ;
  assign n12507 = x5 & ~n12505 ;
  assign n12508 = x5 & ~n12501 ;
  assign n12509 = ( ~n11172 & n12507 ) | ( ~n11172 & n12508 ) | ( n12507 & n12508 ) ;
  assign n12510 = ( n12502 & ~n12506 ) | ( n12502 & n12509 ) | ( ~n12506 & n12509 ) ;
  assign n12511 = n12493 | n12510 ;
  assign n12512 = n12493 & n12510 ;
  assign n12513 = n12511 & ~n12512 ;
  assign n12514 = n12055 | n12061 ;
  assign n12515 = ( n12055 & n12060 ) | ( n12055 & n12514 ) | ( n12060 & n12514 ) ;
  assign n12516 = n12513 & n12515 ;
  assign n12517 = n12513 | n12515 ;
  assign n12518 = ~n12516 & n12517 ;
  assign n12519 = x114 | x115 ;
  assign n12520 = x114 & x115 ;
  assign n12521 = n12519 & ~n12520 ;
  assign n12522 = n12066 | n12067 ;
  assign n12523 = ( n12066 & n12069 ) | ( n12066 & n12522 ) | ( n12069 & n12522 ) ;
  assign n12524 = ( n12066 & n12071 ) | ( n12066 & n12522 ) | ( n12071 & n12522 ) ;
  assign n12525 = ( n10726 & n12523 ) | ( n10726 & n12524 ) | ( n12523 & n12524 ) ;
  assign n12526 = n12523 | n12524 ;
  assign n12527 = ( n10735 & n12525 ) | ( n10735 & n12526 ) | ( n12525 & n12526 ) ;
  assign n12528 = ( n10736 & n12525 ) | ( n10736 & n12526 ) | ( n12525 & n12526 ) ;
  assign n12529 = ( n6159 & n12527 ) | ( n6159 & n12528 ) | ( n12527 & n12528 ) ;
  assign n12530 = ( n6157 & n12527 ) | ( n6157 & n12528 ) | ( n12527 & n12528 ) ;
  assign n12531 = ( n5823 & n12529 ) | ( n5823 & n12530 ) | ( n12529 & n12530 ) ;
  assign n12532 = n12521 | n12531 ;
  assign n12533 = x114 & n133 ;
  assign n12534 = x113 & ~n162 ;
  assign n12535 = ( n137 & n12533 ) | ( n137 & n12534 ) | ( n12533 & n12534 ) ;
  assign n12536 = x0 & x115 ;
  assign n12537 = ( ~n137 & n12533 ) | ( ~n137 & n12536 ) | ( n12533 & n12536 ) ;
  assign n12538 = n12535 | n12537 ;
  assign n12539 = n141 | n12538 ;
  assign n12540 = n12521 & n12524 ;
  assign n12541 = n12521 & n12522 ;
  assign n12542 = n12066 & n12521 ;
  assign n12543 = ( n12069 & n12541 ) | ( n12069 & n12542 ) | ( n12541 & n12542 ) ;
  assign n12544 = ( n10726 & n12540 ) | ( n10726 & n12543 ) | ( n12540 & n12543 ) ;
  assign n12545 = n12540 | n12543 ;
  assign n12546 = ( n10735 & n12544 ) | ( n10735 & n12545 ) | ( n12544 & n12545 ) ;
  assign n12547 = ( n10736 & n12544 ) | ( n10736 & n12545 ) | ( n12544 & n12545 ) ;
  assign n12548 = ( n6159 & n12546 ) | ( n6159 & n12547 ) | ( n12546 & n12547 ) ;
  assign n12549 = ( n6157 & n12546 ) | ( n6157 & n12547 ) | ( n12546 & n12547 ) ;
  assign n12550 = ( n5823 & n12548 ) | ( n5823 & n12549 ) | ( n12548 & n12549 ) ;
  assign n12551 = ( n12538 & n12539 ) | ( n12538 & ~n12550 ) | ( n12539 & ~n12550 ) ;
  assign n12552 = n12538 & n12539 ;
  assign n12553 = ( n12532 & n12551 ) | ( n12532 & n12552 ) | ( n12551 & n12552 ) ;
  assign n12554 = x2 & n12553 ;
  assign n12555 = x2 & ~n12553 ;
  assign n12556 = ( n12553 & ~n12554 ) | ( n12553 & n12555 ) | ( ~n12554 & n12555 ) ;
  assign n12557 = n12518 & n12556 ;
  assign n12558 = n12518 | n12556 ;
  assign n12559 = ~n12557 & n12558 ;
  assign n12560 = n12102 | n12109 ;
  assign n12561 = n12559 & n12560 ;
  assign n12562 = n12559 | n12560 ;
  assign n12563 = ~n12561 & n12562 ;
  assign n12564 = n12178 | n12179 ;
  assign n12565 = ( n12178 & n12181 ) | ( n12178 & n12564 ) | ( n12181 & n12564 ) ;
  assign n12566 = ~x51 & x52 ;
  assign n12567 = x51 & ~x52 ;
  assign n12568 = n12566 | n12567 ;
  assign n12569 = ~n12115 & n12568 ;
  assign n12570 = x64 & n12569 ;
  assign n12571 = ~x52 & x53 ;
  assign n12572 = x52 & ~x53 ;
  assign n12573 = n12571 | n12572 ;
  assign n12574 = n12115 & ~n12573 ;
  assign n12575 = x65 & n12574 ;
  assign n12576 = n12570 | n12575 ;
  assign n12577 = n12115 & n12573 ;
  assign n12578 = x53 | n144 ;
  assign n12579 = ( x53 & n12577 ) | ( x53 & n12578 ) | ( n12577 & n12578 ) ;
  assign n12580 = ~x53 & n12579 ;
  assign n12581 = ( ~x53 & n12576 ) | ( ~x53 & n12580 ) | ( n12576 & n12580 ) ;
  assign n12582 = x53 & ~x64 ;
  assign n12583 = ( x53 & ~n12115 ) | ( x53 & n12582 ) | ( ~n12115 & n12582 ) ;
  assign n12584 = n12579 & n12583 ;
  assign n12585 = ( n12576 & n12583 ) | ( n12576 & n12584 ) | ( n12583 & n12584 ) ;
  assign n12586 = n144 & n12577 ;
  assign n12587 = n12583 & ~n12586 ;
  assign n12588 = ~n12576 & n12587 ;
  assign n12589 = ( n12581 & n12585 ) | ( n12581 & n12588 ) | ( n12585 & n12588 ) ;
  assign n12590 = n12579 | n12583 ;
  assign n12591 = n12576 | n12590 ;
  assign n12592 = ~n12583 & n12586 ;
  assign n12593 = ( n12576 & ~n12583 ) | ( n12576 & n12592 ) | ( ~n12583 & n12592 ) ;
  assign n12594 = ( n12581 & n12591 ) | ( n12581 & ~n12593 ) | ( n12591 & ~n12593 ) ;
  assign n12595 = ~n12589 & n12594 ;
  assign n12596 = n241 & n11208 ;
  assign n12597 = x68 & n11205 ;
  assign n12598 = x67 & n11200 ;
  assign n12599 = x66 & ~n11199 ;
  assign n12600 = n11679 & n12599 ;
  assign n12601 = n12598 | n12600 ;
  assign n12602 = n12597 | n12601 ;
  assign n12603 = n12596 | n12602 ;
  assign n12604 = x50 | n12597 ;
  assign n12605 = n12601 | n12604 ;
  assign n12606 = n12596 | n12605 ;
  assign n12607 = ~x50 & n12605 ;
  assign n12608 = ( ~x50 & n12596 ) | ( ~x50 & n12607 ) | ( n12596 & n12607 ) ;
  assign n12609 = ( ~n12603 & n12606 ) | ( ~n12603 & n12608 ) | ( n12606 & n12608 ) ;
  assign n12610 = n12595 | n12609 ;
  assign n12611 = n12595 & n12609 ;
  assign n12612 = n12610 & ~n12611 ;
  assign n12613 = ( n11693 & n12116 ) | ( n11693 & n12132 ) | ( n12116 & n12132 ) ;
  assign n12614 = n12612 | n12613 ;
  assign n12615 = n12612 & n12613 ;
  assign n12616 = n12614 & ~n12615 ;
  assign n12617 = x70 & n9928 ;
  assign n12618 = x69 & ~n9927 ;
  assign n12619 = n10379 & n12618 ;
  assign n12620 = n12617 | n12619 ;
  assign n12621 = x71 & n9933 ;
  assign n12622 = n9936 | n12621 ;
  assign n12623 = n12620 | n12622 ;
  assign n12624 = x47 & ~n12623 ;
  assign n12625 = x47 & ~n12621 ;
  assign n12626 = ~n12620 & n12625 ;
  assign n12627 = ( ~n438 & n12624 ) | ( ~n438 & n12626 ) | ( n12624 & n12626 ) ;
  assign n12628 = ~x47 & n12623 ;
  assign n12629 = ~x47 & n12621 ;
  assign n12630 = ( ~x47 & n12620 ) | ( ~x47 & n12629 ) | ( n12620 & n12629 ) ;
  assign n12631 = ( n438 & n12628 ) | ( n438 & n12630 ) | ( n12628 & n12630 ) ;
  assign n12632 = n12627 | n12631 ;
  assign n12633 = n12616 & n12632 ;
  assign n12634 = n12616 & ~n12633 ;
  assign n12635 = ~n12616 & n12632 ;
  assign n12636 = n12634 | n12635 ;
  assign n12637 = n12152 | n12157 ;
  assign n12638 = ( n12152 & n12155 ) | ( n12152 & n12637 ) | ( n12155 & n12637 ) ;
  assign n12639 = n12636 | n12638 ;
  assign n12640 = n12636 & n12638 ;
  assign n12641 = n12639 & ~n12640 ;
  assign n12642 = x74 & n8724 ;
  assign n12643 = x73 & n8719 ;
  assign n12644 = x72 & ~n8718 ;
  assign n12645 = n9149 & n12644 ;
  assign n12646 = n12643 | n12645 ;
  assign n12647 = n12642 | n12646 ;
  assign n12648 = n8727 | n12642 ;
  assign n12649 = n12646 | n12648 ;
  assign n12650 = ( n710 & n12647 ) | ( n710 & n12649 ) | ( n12647 & n12649 ) ;
  assign n12651 = x44 & n12649 ;
  assign n12652 = x44 & n12642 ;
  assign n12653 = ( x44 & n12646 ) | ( x44 & n12652 ) | ( n12646 & n12652 ) ;
  assign n12654 = ( n710 & n12651 ) | ( n710 & n12653 ) | ( n12651 & n12653 ) ;
  assign n12655 = x44 & ~n12653 ;
  assign n12656 = x44 & ~n12649 ;
  assign n12657 = ( ~n710 & n12655 ) | ( ~n710 & n12656 ) | ( n12655 & n12656 ) ;
  assign n12658 = ( n12650 & ~n12654 ) | ( n12650 & n12657 ) | ( ~n12654 & n12657 ) ;
  assign n12659 = n12641 & n12658 ;
  assign n12660 = n12641 | n12658 ;
  assign n12661 = ~n12659 & n12660 ;
  assign n12662 = n12565 & n12661 ;
  assign n12663 = n12565 & ~n12662 ;
  assign n12664 = x77 & n7566 ;
  assign n12665 = x76 & n7561 ;
  assign n12666 = x75 & ~n7560 ;
  assign n12667 = n7953 & n12666 ;
  assign n12668 = n12665 | n12667 ;
  assign n12669 = n12664 | n12668 ;
  assign n12670 = n7569 | n12664 ;
  assign n12671 = n12668 | n12670 ;
  assign n12672 = ( n1059 & n12669 ) | ( n1059 & n12671 ) | ( n12669 & n12671 ) ;
  assign n12673 = x41 & n12671 ;
  assign n12674 = x41 & n12664 ;
  assign n12675 = ( x41 & n12668 ) | ( x41 & n12674 ) | ( n12668 & n12674 ) ;
  assign n12676 = ( n1059 & n12673 ) | ( n1059 & n12675 ) | ( n12673 & n12675 ) ;
  assign n12677 = x41 & ~n12675 ;
  assign n12678 = x41 & ~n12671 ;
  assign n12679 = ( ~n1059 & n12677 ) | ( ~n1059 & n12678 ) | ( n12677 & n12678 ) ;
  assign n12680 = ( n12672 & ~n12676 ) | ( n12672 & n12679 ) | ( ~n12676 & n12679 ) ;
  assign n12681 = ~n12660 & n12661 ;
  assign n12682 = ( ~n12565 & n12661 ) | ( ~n12565 & n12681 ) | ( n12661 & n12681 ) ;
  assign n12683 = n12680 & n12682 ;
  assign n12684 = ( n12663 & n12680 ) | ( n12663 & n12683 ) | ( n12680 & n12683 ) ;
  assign n12685 = n12680 | n12682 ;
  assign n12686 = n12663 | n12685 ;
  assign n12687 = ~n12684 & n12686 ;
  assign n12688 = n12112 | n12202 ;
  assign n12689 = ( n12202 & n12205 ) | ( n12202 & n12688 ) | ( n12205 & n12688 ) ;
  assign n12690 = n12687 & n12689 ;
  assign n12691 = n12687 | n12689 ;
  assign n12692 = ~n12690 & n12691 ;
  assign n12693 = x80 & n6536 ;
  assign n12694 = x79 & n6531 ;
  assign n12695 = x78 & ~n6530 ;
  assign n12696 = n6871 & n12695 ;
  assign n12697 = n12694 | n12696 ;
  assign n12698 = n12693 | n12697 ;
  assign n12699 = n6539 | n12693 ;
  assign n12700 = n12697 | n12699 ;
  assign n12701 = ( n1499 & n12698 ) | ( n1499 & n12700 ) | ( n12698 & n12700 ) ;
  assign n12702 = x38 & n12700 ;
  assign n12703 = x38 & n12693 ;
  assign n12704 = ( x38 & n12697 ) | ( x38 & n12703 ) | ( n12697 & n12703 ) ;
  assign n12705 = ( n1499 & n12702 ) | ( n1499 & n12704 ) | ( n12702 & n12704 ) ;
  assign n12706 = x38 & ~n12704 ;
  assign n12707 = x38 & ~n12700 ;
  assign n12708 = ( ~n1499 & n12706 ) | ( ~n1499 & n12707 ) | ( n12706 & n12707 ) ;
  assign n12709 = ( n12701 & ~n12705 ) | ( n12701 & n12708 ) | ( ~n12705 & n12708 ) ;
  assign n12710 = n12692 & n12709 ;
  assign n12711 = n12692 & ~n12710 ;
  assign n12712 = ~n12692 & n12709 ;
  assign n12713 = n12711 | n12712 ;
  assign n12714 = n12226 | n12229 ;
  assign n12715 = n12713 | n12714 ;
  assign n12716 = n12713 & n12714 ;
  assign n12717 = n12715 & ~n12716 ;
  assign n12718 = x83 & n5554 ;
  assign n12719 = x82 & n5549 ;
  assign n12720 = x81 & ~n5548 ;
  assign n12721 = n5893 & n12720 ;
  assign n12722 = n12719 | n12721 ;
  assign n12723 = n12718 | n12722 ;
  assign n12724 = n5557 | n12718 ;
  assign n12725 = n12722 | n12724 ;
  assign n12726 = ( n2009 & n12723 ) | ( n2009 & n12725 ) | ( n12723 & n12725 ) ;
  assign n12727 = x35 & n12725 ;
  assign n12728 = x35 & n12718 ;
  assign n12729 = ( x35 & n12722 ) | ( x35 & n12728 ) | ( n12722 & n12728 ) ;
  assign n12730 = ( n2009 & n12727 ) | ( n2009 & n12729 ) | ( n12727 & n12729 ) ;
  assign n12731 = x35 & ~n12729 ;
  assign n12732 = x35 & ~n12725 ;
  assign n12733 = ( ~n2009 & n12731 ) | ( ~n2009 & n12732 ) | ( n12731 & n12732 ) ;
  assign n12734 = ( n12726 & ~n12730 ) | ( n12726 & n12733 ) | ( ~n12730 & n12733 ) ;
  assign n12735 = n12717 & n12734 ;
  assign n12736 = n12717 | n12734 ;
  assign n12737 = ~n12735 & n12736 ;
  assign n12738 = n12249 | n12251 ;
  assign n12739 = ( n12249 & n12254 ) | ( n12249 & n12738 ) | ( n12254 & n12738 ) ;
  assign n12740 = n12737 & n12739 ;
  assign n12741 = n12739 & ~n12740 ;
  assign n12742 = ( n12737 & ~n12740 ) | ( n12737 & n12741 ) | ( ~n12740 & n12741 ) ;
  assign n12743 = x86 & n4631 ;
  assign n12744 = x85 & n4626 ;
  assign n12745 = x84 & ~n4625 ;
  assign n12746 = n4943 & n12745 ;
  assign n12747 = n12744 | n12746 ;
  assign n12748 = n12743 | n12747 ;
  assign n12749 = n4634 | n12743 ;
  assign n12750 = n12747 | n12749 ;
  assign n12751 = ( n2606 & n12748 ) | ( n2606 & n12750 ) | ( n12748 & n12750 ) ;
  assign n12752 = x32 & n12750 ;
  assign n12753 = x32 & n12743 ;
  assign n12754 = ( x32 & n12747 ) | ( x32 & n12753 ) | ( n12747 & n12753 ) ;
  assign n12755 = ( n2606 & n12752 ) | ( n2606 & n12754 ) | ( n12752 & n12754 ) ;
  assign n12756 = x32 & ~n12754 ;
  assign n12757 = x32 & ~n12750 ;
  assign n12758 = ( ~n2606 & n12756 ) | ( ~n2606 & n12757 ) | ( n12756 & n12757 ) ;
  assign n12759 = ( n12751 & ~n12755 ) | ( n12751 & n12758 ) | ( ~n12755 & n12758 ) ;
  assign n12760 = ~n12740 & n12759 ;
  assign n12761 = n12737 & n12759 ;
  assign n12762 = ( n12741 & n12760 ) | ( n12741 & n12761 ) | ( n12760 & n12761 ) ;
  assign n12763 = n12742 & ~n12762 ;
  assign n12764 = n12740 & n12759 ;
  assign n12765 = ~n12737 & n12759 ;
  assign n12766 = ( ~n12741 & n12764 ) | ( ~n12741 & n12765 ) | ( n12764 & n12765 ) ;
  assign n12767 = n12763 | n12766 ;
  assign n12768 = n12275 | n12277 ;
  assign n12769 = n12276 | n12768 ;
  assign n12770 = ( n12275 & n12279 ) | ( n12275 & n12769 ) | ( n12279 & n12769 ) ;
  assign n12771 = n12767 | n12770 ;
  assign n12772 = n12767 & n12770 ;
  assign n12773 = n12771 & ~n12772 ;
  assign n12774 = x89 & n3816 ;
  assign n12775 = x88 & n3811 ;
  assign n12776 = x87 & ~n3810 ;
  assign n12777 = n4067 & n12776 ;
  assign n12778 = n12775 | n12777 ;
  assign n12779 = n12774 | n12778 ;
  assign n12780 = n3819 | n12774 ;
  assign n12781 = n12778 | n12780 ;
  assign n12782 = ( n3282 & n12779 ) | ( n3282 & n12781 ) | ( n12779 & n12781 ) ;
  assign n12783 = x29 & n12781 ;
  assign n12784 = x29 & n12774 ;
  assign n12785 = ( x29 & n12778 ) | ( x29 & n12784 ) | ( n12778 & n12784 ) ;
  assign n12786 = ( n3282 & n12783 ) | ( n3282 & n12785 ) | ( n12783 & n12785 ) ;
  assign n12787 = x29 & ~n12785 ;
  assign n12788 = x29 & ~n12781 ;
  assign n12789 = ( ~n3282 & n12787 ) | ( ~n3282 & n12788 ) | ( n12787 & n12788 ) ;
  assign n12790 = ( n12782 & ~n12786 ) | ( n12782 & n12789 ) | ( ~n12786 & n12789 ) ;
  assign n12791 = n12773 & n12790 ;
  assign n12792 = n12773 & ~n12791 ;
  assign n12793 = ~n12773 & n12790 ;
  assign n12794 = n12792 | n12793 ;
  assign n12795 = n12307 | n12311 ;
  assign n12796 = ( n12307 & n12308 ) | ( n12307 & n12795 ) | ( n12308 & n12795 ) ;
  assign n12797 = ~n12794 & n12796 ;
  assign n12798 = n12794 & ~n12796 ;
  assign n12799 = n12797 | n12798 ;
  assign n12800 = x92 & n3085 ;
  assign n12801 = x91 & n3080 ;
  assign n12802 = x90 & ~n3079 ;
  assign n12803 = n3309 & n12802 ;
  assign n12804 = n12801 | n12803 ;
  assign n12805 = n12800 | n12804 ;
  assign n12806 = n3088 | n12800 ;
  assign n12807 = n12804 | n12806 ;
  assign n12808 = ( n4040 & n12805 ) | ( n4040 & n12807 ) | ( n12805 & n12807 ) ;
  assign n12809 = x26 & n12807 ;
  assign n12810 = x26 & n12800 ;
  assign n12811 = ( x26 & n12804 ) | ( x26 & n12810 ) | ( n12804 & n12810 ) ;
  assign n12812 = ( n4040 & n12809 ) | ( n4040 & n12811 ) | ( n12809 & n12811 ) ;
  assign n12813 = x26 & ~n12811 ;
  assign n12814 = x26 & ~n12807 ;
  assign n12815 = ( ~n4040 & n12813 ) | ( ~n4040 & n12814 ) | ( n12813 & n12814 ) ;
  assign n12816 = ( n12808 & ~n12812 ) | ( n12808 & n12815 ) | ( ~n12812 & n12815 ) ;
  assign n12817 = n12799 & n12816 ;
  assign n12818 = n12799 | n12816 ;
  assign n12819 = ~n12817 & n12818 ;
  assign n12820 = ( n11875 & n12314 ) | ( n11875 & n12331 ) | ( n12314 & n12331 ) ;
  assign n12821 = n12314 | n12331 ;
  assign n12822 = ( n11882 & n12820 ) | ( n11882 & n12821 ) | ( n12820 & n12821 ) ;
  assign n12823 = n12819 | n12822 ;
  assign n12824 = n12819 & n12822 ;
  assign n12825 = n12823 & ~n12824 ;
  assign n12826 = x95 & n2429 ;
  assign n12827 = x94 & n2424 ;
  assign n12828 = x93 & ~n2423 ;
  assign n12829 = n2631 & n12828 ;
  assign n12830 = n12827 | n12829 ;
  assign n12831 = n12826 | n12830 ;
  assign n12832 = n2432 | n12826 ;
  assign n12833 = n12830 | n12832 ;
  assign n12834 = ( n4897 & n12831 ) | ( n4897 & n12833 ) | ( n12831 & n12833 ) ;
  assign n12835 = x23 & n12833 ;
  assign n12836 = x23 & n12826 ;
  assign n12837 = ( x23 & n12830 ) | ( x23 & n12836 ) | ( n12830 & n12836 ) ;
  assign n12838 = ( n4897 & n12835 ) | ( n4897 & n12837 ) | ( n12835 & n12837 ) ;
  assign n12839 = x23 & ~n12837 ;
  assign n12840 = x23 & ~n12833 ;
  assign n12841 = ( ~n4897 & n12839 ) | ( ~n4897 & n12840 ) | ( n12839 & n12840 ) ;
  assign n12842 = ( n12834 & ~n12838 ) | ( n12834 & n12841 ) | ( ~n12838 & n12841 ) ;
  assign n12843 = n12825 & n12842 ;
  assign n12844 = n12825 & ~n12843 ;
  assign n12845 = ~n12825 & n12842 ;
  assign n12846 = n12844 | n12845 ;
  assign n12847 = n12358 | n12364 ;
  assign n12848 = n12846 | n12847 ;
  assign n12849 = n12846 & n12847 ;
  assign n12850 = n12848 & ~n12849 ;
  assign n12851 = x98 & n1859 ;
  assign n12852 = x97 & n1854 ;
  assign n12853 = x96 & ~n1853 ;
  assign n12854 = n2037 & n12853 ;
  assign n12855 = n12852 | n12854 ;
  assign n12856 = n12851 | n12855 ;
  assign n12857 = n1862 | n12851 ;
  assign n12858 = n12855 | n12857 ;
  assign n12859 = ( ~n5850 & n12856 ) | ( ~n5850 & n12858 ) | ( n12856 & n12858 ) ;
  assign n12860 = n12856 & n12858 ;
  assign n12861 = ( n5834 & n12859 ) | ( n5834 & n12860 ) | ( n12859 & n12860 ) ;
  assign n12862 = x20 & n12858 ;
  assign n12863 = x20 & n12851 ;
  assign n12864 = ( x20 & n12855 ) | ( x20 & n12863 ) | ( n12855 & n12863 ) ;
  assign n12865 = ( ~n5850 & n12862 ) | ( ~n5850 & n12864 ) | ( n12862 & n12864 ) ;
  assign n12866 = n12862 & n12864 ;
  assign n12867 = ( n5834 & n12865 ) | ( n5834 & n12866 ) | ( n12865 & n12866 ) ;
  assign n12868 = x20 & ~n12864 ;
  assign n12869 = x20 & ~n12858 ;
  assign n12870 = ( n5850 & n12868 ) | ( n5850 & n12869 ) | ( n12868 & n12869 ) ;
  assign n12871 = n12868 | n12869 ;
  assign n12872 = ( ~n5834 & n12870 ) | ( ~n5834 & n12871 ) | ( n12870 & n12871 ) ;
  assign n12873 = ( n12861 & ~n12867 ) | ( n12861 & n12872 ) | ( ~n12867 & n12872 ) ;
  assign n12874 = n12850 & n12873 ;
  assign n12875 = n12850 & ~n12874 ;
  assign n12876 = ~n12850 & n12873 ;
  assign n12877 = n12875 | n12876 ;
  assign n12878 = ( n12366 & n12383 ) | ( n12366 & n12390 ) | ( n12383 & n12390 ) ;
  assign n12879 = n12877 | n12878 ;
  assign n12880 = n12877 & n12878 ;
  assign n12881 = n12879 & ~n12880 ;
  assign n12882 = x101 & n1383 ;
  assign n12883 = x100 & n1378 ;
  assign n12884 = x99 & ~n1377 ;
  assign n12885 = n1542 & n12884 ;
  assign n12886 = n12883 | n12885 ;
  assign n12887 = n12882 | n12886 ;
  assign n12888 = n1386 | n12882 ;
  assign n12889 = n12886 | n12888 ;
  assign n12890 = ( n6844 & n12887 ) | ( n6844 & n12889 ) | ( n12887 & n12889 ) ;
  assign n12891 = x17 & n12889 ;
  assign n12892 = x17 & n12882 ;
  assign n12893 = ( x17 & n12886 ) | ( x17 & n12892 ) | ( n12886 & n12892 ) ;
  assign n12894 = ( n6844 & n12891 ) | ( n6844 & n12893 ) | ( n12891 & n12893 ) ;
  assign n12895 = x17 & ~n12893 ;
  assign n12896 = x17 & ~n12889 ;
  assign n12897 = ( ~n6844 & n12895 ) | ( ~n6844 & n12896 ) | ( n12895 & n12896 ) ;
  assign n12898 = ( n12890 & ~n12894 ) | ( n12890 & n12897 ) | ( ~n12894 & n12897 ) ;
  assign n12899 = n12881 & n12898 ;
  assign n12900 = n12881 & ~n12899 ;
  assign n12901 = ~n12881 & n12898 ;
  assign n12902 = n12900 | n12901 ;
  assign n12903 = n12411 | n12413 ;
  assign n12904 = ( n12411 & n12415 ) | ( n12411 & n12903 ) | ( n12415 & n12903 ) ;
  assign n12905 = n12902 | n12904 ;
  assign n12906 = n12902 & n12904 ;
  assign n12907 = n12905 & ~n12906 ;
  assign n12908 = x104 & n962 ;
  assign n12909 = x103 & n957 ;
  assign n12910 = x102 & ~n956 ;
  assign n12911 = n1105 & n12910 ;
  assign n12912 = n12909 | n12911 ;
  assign n12913 = n12908 | n12912 ;
  assign n12914 = n965 | n12908 ;
  assign n12915 = n12912 | n12914 ;
  assign n12916 = ( n7911 & n12913 ) | ( n7911 & n12915 ) | ( n12913 & n12915 ) ;
  assign n12917 = x14 & n12915 ;
  assign n12918 = x14 & n12908 ;
  assign n12919 = ( x14 & n12912 ) | ( x14 & n12918 ) | ( n12912 & n12918 ) ;
  assign n12920 = ( n7911 & n12917 ) | ( n7911 & n12919 ) | ( n12917 & n12919 ) ;
  assign n12921 = x14 & ~n12919 ;
  assign n12922 = x14 & ~n12915 ;
  assign n12923 = ( ~n7911 & n12921 ) | ( ~n7911 & n12922 ) | ( n12921 & n12922 ) ;
  assign n12924 = ( n12916 & ~n12920 ) | ( n12916 & n12923 ) | ( ~n12920 & n12923 ) ;
  assign n12925 = n12907 & n12924 ;
  assign n12926 = n12907 & ~n12925 ;
  assign n12927 = ~n12907 & n12924 ;
  assign n12928 = n12926 | n12927 ;
  assign n12929 = n12436 | n12443 ;
  assign n12930 = n12928 | n12929 ;
  assign n12931 = n12928 & n12929 ;
  assign n12932 = n12930 & ~n12931 ;
  assign n12933 = x107 & n636 ;
  assign n12934 = x106 & n631 ;
  assign n12935 = x105 & ~n630 ;
  assign n12936 = n764 & n12935 ;
  assign n12937 = n12934 | n12936 ;
  assign n12938 = n12933 | n12937 ;
  assign n12939 = n639 | n12933 ;
  assign n12940 = n12937 | n12939 ;
  assign n12941 = ( n9084 & n12938 ) | ( n9084 & n12940 ) | ( n12938 & n12940 ) ;
  assign n12942 = x11 & n12940 ;
  assign n12943 = x11 & n12933 ;
  assign n12944 = ( x11 & n12937 ) | ( x11 & n12943 ) | ( n12937 & n12943 ) ;
  assign n12945 = ( n9084 & n12942 ) | ( n9084 & n12944 ) | ( n12942 & n12944 ) ;
  assign n12946 = x11 & ~n12944 ;
  assign n12947 = x11 & ~n12940 ;
  assign n12948 = ( ~n9084 & n12946 ) | ( ~n9084 & n12947 ) | ( n12946 & n12947 ) ;
  assign n12949 = ( n12941 & ~n12945 ) | ( n12941 & n12948 ) | ( ~n12945 & n12948 ) ;
  assign n12950 = n12932 & n12949 ;
  assign n12951 = n12932 | n12949 ;
  assign n12952 = ~n12950 & n12951 ;
  assign n12953 = n12463 | n12464 ;
  assign n12954 = ( n12463 & n12466 ) | ( n12463 & n12953 ) | ( n12466 & n12953 ) ;
  assign n12955 = n12952 & n12954 ;
  assign n12956 = n12954 & ~n12955 ;
  assign n12957 = ( n12952 & ~n12955 ) | ( n12952 & n12956 ) | ( ~n12955 & n12956 ) ;
  assign n12958 = x110 & n389 ;
  assign n12959 = x109 & n384 ;
  assign n12960 = x108 & ~n383 ;
  assign n12961 = n463 & n12960 ;
  assign n12962 = n12959 | n12961 ;
  assign n12963 = n12958 | n12962 ;
  assign n12964 = n392 | n12958 ;
  assign n12965 = n12962 | n12964 ;
  assign n12966 = ( n10330 & n12963 ) | ( n10330 & n12965 ) | ( n12963 & n12965 ) ;
  assign n12967 = x8 & n12965 ;
  assign n12968 = x8 & n12958 ;
  assign n12969 = ( x8 & n12962 ) | ( x8 & n12968 ) | ( n12962 & n12968 ) ;
  assign n12970 = ( n10330 & n12967 ) | ( n10330 & n12969 ) | ( n12967 & n12969 ) ;
  assign n12971 = x8 & ~n12969 ;
  assign n12972 = x8 & ~n12965 ;
  assign n12973 = ( ~n10330 & n12971 ) | ( ~n10330 & n12972 ) | ( n12971 & n12972 ) ;
  assign n12974 = ( n12966 & ~n12970 ) | ( n12966 & n12973 ) | ( ~n12970 & n12973 ) ;
  assign n12975 = ~n12955 & n12974 ;
  assign n12976 = n12952 & n12974 ;
  assign n12977 = ( n12956 & n12975 ) | ( n12956 & n12976 ) | ( n12975 & n12976 ) ;
  assign n12978 = n12957 & ~n12977 ;
  assign n12979 = n12955 & n12974 ;
  assign n12980 = ~n12952 & n12974 ;
  assign n12981 = ( ~n12956 & n12979 ) | ( ~n12956 & n12980 ) | ( n12979 & n12980 ) ;
  assign n12982 = n12978 | n12981 ;
  assign n12983 = ( n12032 & n12469 ) | ( n12032 & n12486 ) | ( n12469 & n12486 ) ;
  assign n12984 = n12982 | n12983 ;
  assign n12985 = n12982 & n12983 ;
  assign n12986 = n12984 & ~n12985 ;
  assign n12987 = x113 & n212 ;
  assign n12988 = x112 & n207 ;
  assign n12989 = x111 & ~n206 ;
  assign n12990 = n267 & n12989 ;
  assign n12991 = n12988 | n12990 ;
  assign n12992 = n12987 | n12991 ;
  assign n12993 = n215 | n12987 ;
  assign n12994 = n12991 | n12993 ;
  assign n12995 = ( ~n11642 & n12992 ) | ( ~n11642 & n12994 ) | ( n12992 & n12994 ) ;
  assign n12996 = n12992 & n12994 ;
  assign n12997 = ( n11626 & n12995 ) | ( n11626 & n12996 ) | ( n12995 & n12996 ) ;
  assign n12998 = x5 & n12997 ;
  assign n12999 = x5 & ~n12997 ;
  assign n13000 = ( n12997 & ~n12998 ) | ( n12997 & n12999 ) | ( ~n12998 & n12999 ) ;
  assign n13001 = n12986 & n13000 ;
  assign n13002 = n12986 & ~n13001 ;
  assign n13003 = ~n12986 & n13000 ;
  assign n13004 = n13002 | n13003 ;
  assign n13005 = n12512 | n12516 ;
  assign n13006 = ~n13004 & n13005 ;
  assign n13007 = n13004 & ~n13005 ;
  assign n13008 = n13006 | n13007 ;
  assign n13009 = x115 | x116 ;
  assign n13010 = x115 & x116 ;
  assign n13011 = n13009 & ~n13010 ;
  assign n13012 = n12520 | n12543 ;
  assign n13013 = n12520 | n12521 ;
  assign n13014 = ( n12520 & n12524 ) | ( n12520 & n13013 ) | ( n12524 & n13013 ) ;
  assign n13015 = ( n10726 & n13012 ) | ( n10726 & n13014 ) | ( n13012 & n13014 ) ;
  assign n13016 = n13012 | n13014 ;
  assign n13017 = ( n10735 & n13015 ) | ( n10735 & n13016 ) | ( n13015 & n13016 ) ;
  assign n13018 = ( n10736 & n13015 ) | ( n10736 & n13016 ) | ( n13015 & n13016 ) ;
  assign n13019 = ( n6159 & n13017 ) | ( n6159 & n13018 ) | ( n13017 & n13018 ) ;
  assign n13020 = ( n6157 & n13017 ) | ( n6157 & n13018 ) | ( n13017 & n13018 ) ;
  assign n13021 = ( n5823 & n13019 ) | ( n5823 & n13020 ) | ( n13019 & n13020 ) ;
  assign n13022 = n13011 | n13021 ;
  assign n13023 = x115 & n133 ;
  assign n13024 = x114 & ~n162 ;
  assign n13025 = ( n137 & n13023 ) | ( n137 & n13024 ) | ( n13023 & n13024 ) ;
  assign n13026 = x0 & x116 ;
  assign n13027 = ( ~n137 & n13023 ) | ( ~n137 & n13026 ) | ( n13023 & n13026 ) ;
  assign n13028 = n13025 | n13027 ;
  assign n13029 = n141 | n13028 ;
  assign n13030 = n12520 & n13011 ;
  assign n13031 = ( n12543 & n13011 ) | ( n12543 & n13030 ) | ( n13011 & n13030 ) ;
  assign n13032 = n13011 & n13013 ;
  assign n13033 = ( n12524 & n13030 ) | ( n12524 & n13032 ) | ( n13030 & n13032 ) ;
  assign n13034 = ( n10726 & n13031 ) | ( n10726 & n13033 ) | ( n13031 & n13033 ) ;
  assign n13035 = n13031 | n13033 ;
  assign n13036 = ( n10735 & n13034 ) | ( n10735 & n13035 ) | ( n13034 & n13035 ) ;
  assign n13037 = ( n10736 & n13034 ) | ( n10736 & n13035 ) | ( n13034 & n13035 ) ;
  assign n13038 = ( n6159 & n13036 ) | ( n6159 & n13037 ) | ( n13036 & n13037 ) ;
  assign n13039 = ( n6157 & n13036 ) | ( n6157 & n13037 ) | ( n13036 & n13037 ) ;
  assign n13040 = ( n5823 & n13038 ) | ( n5823 & n13039 ) | ( n13038 & n13039 ) ;
  assign n13041 = ( n13028 & n13029 ) | ( n13028 & ~n13040 ) | ( n13029 & ~n13040 ) ;
  assign n13042 = n13028 & n13029 ;
  assign n13043 = ( n13022 & n13041 ) | ( n13022 & n13042 ) | ( n13041 & n13042 ) ;
  assign n13044 = x2 & n13043 ;
  assign n13045 = x2 & ~n13043 ;
  assign n13046 = ( n13043 & ~n13044 ) | ( n13043 & n13045 ) | ( ~n13044 & n13045 ) ;
  assign n13047 = n13008 & n13046 ;
  assign n13048 = n13008 | n13046 ;
  assign n13049 = ~n13047 & n13048 ;
  assign n13050 = n12557 | n12559 ;
  assign n13051 = ( n12557 & n12560 ) | ( n12557 & n13050 ) | ( n12560 & n13050 ) ;
  assign n13052 = n13049 & n13051 ;
  assign n13053 = n13049 | n13051 ;
  assign n13054 = ~n13052 & n13053 ;
  assign n13055 = n13047 | n13052 ;
  assign n13056 = n12735 | n12740 ;
  assign n13057 = n12710 | n12716 ;
  assign n13058 = x72 & n9933 ;
  assign n13059 = x71 & n9928 ;
  assign n13060 = x70 & ~n9927 ;
  assign n13061 = n10379 & n13060 ;
  assign n13062 = n13059 | n13061 ;
  assign n13063 = n13058 | n13062 ;
  assign n13064 = ( n513 & n9936 ) | ( n513 & n13063 ) | ( n9936 & n13063 ) ;
  assign n13065 = x47 & n9936 ;
  assign n13066 = ( x47 & n9936 ) | ( x47 & ~n13058 ) | ( n9936 & ~n13058 ) ;
  assign n13067 = ( ~n13062 & n13065 ) | ( ~n13062 & n13066 ) | ( n13065 & n13066 ) ;
  assign n13068 = ( x47 & n513 ) | ( x47 & n13067 ) | ( n513 & n13067 ) ;
  assign n13069 = ~n13064 & n13068 ;
  assign n13070 = n13063 | n13067 ;
  assign n13071 = x47 | n13063 ;
  assign n13072 = ( n513 & n13070 ) | ( n513 & n13071 ) | ( n13070 & n13071 ) ;
  assign n13073 = ( ~x47 & n13069 ) | ( ~x47 & n13072 ) | ( n13069 & n13072 ) ;
  assign n13074 = x66 & n12574 ;
  assign n13075 = x65 & n12569 ;
  assign n13076 = ~n12115 & n12573 ;
  assign n13077 = x64 & ~n12568 ;
  assign n13078 = n13076 & n13077 ;
  assign n13079 = n13075 | n13078 ;
  assign n13080 = n13074 | n13079 ;
  assign n13081 = n159 & n12577 ;
  assign n13082 = n13080 | n13081 ;
  assign n13083 = x53 | n12577 ;
  assign n13084 = ( x53 & n159 ) | ( x53 & n13083 ) | ( n159 & n13083 ) ;
  assign n13085 = n13080 | n13084 ;
  assign n13086 = ~x53 & n13084 ;
  assign n13087 = ( ~x53 & n13080 ) | ( ~x53 & n13086 ) | ( n13080 & n13086 ) ;
  assign n13088 = ( ~n13082 & n13085 ) | ( ~n13082 & n13087 ) | ( n13085 & n13087 ) ;
  assign n13089 = n12589 | n13088 ;
  assign n13090 = n12589 & n13088 ;
  assign n13091 = n13089 & ~n13090 ;
  assign n13092 = n293 & n11208 ;
  assign n13093 = x69 & n11205 ;
  assign n13094 = x68 & n11200 ;
  assign n13095 = x67 & ~n11199 ;
  assign n13096 = n11679 & n13095 ;
  assign n13097 = n13094 | n13096 ;
  assign n13098 = n13093 | n13097 ;
  assign n13099 = n13092 | n13098 ;
  assign n13100 = x50 | n13093 ;
  assign n13101 = n13097 | n13100 ;
  assign n13102 = n13092 | n13101 ;
  assign n13103 = ~x50 & n13101 ;
  assign n13104 = ( ~x50 & n13092 ) | ( ~x50 & n13103 ) | ( n13092 & n13103 ) ;
  assign n13105 = ( ~n13099 & n13102 ) | ( ~n13099 & n13104 ) | ( n13102 & n13104 ) ;
  assign n13106 = n13091 | n13105 ;
  assign n13107 = n13091 & n13105 ;
  assign n13108 = n13106 & ~n13107 ;
  assign n13109 = n12611 | n12613 ;
  assign n13110 = ( n12611 & n12612 ) | ( n12611 & n13109 ) | ( n12612 & n13109 ) ;
  assign n13111 = n13108 & n13110 ;
  assign n13112 = n13108 & ~n13111 ;
  assign n13113 = ~n13108 & n13110 ;
  assign n13114 = n13073 & n13113 ;
  assign n13115 = ( n13073 & n13112 ) | ( n13073 & n13114 ) | ( n13112 & n13114 ) ;
  assign n13116 = n13073 | n13113 ;
  assign n13117 = n13112 | n13116 ;
  assign n13118 = ~n13115 & n13117 ;
  assign n13119 = n12633 & n13118 ;
  assign n13120 = ( n12640 & n13118 ) | ( n12640 & n13119 ) | ( n13118 & n13119 ) ;
  assign n13121 = n12633 | n13118 ;
  assign n13122 = n12640 | n13121 ;
  assign n13123 = ~n13120 & n13122 ;
  assign n13124 = x75 & n8724 ;
  assign n13125 = x74 & n8719 ;
  assign n13126 = x73 & ~n8718 ;
  assign n13127 = n9149 & n13126 ;
  assign n13128 = n13125 | n13127 ;
  assign n13129 = n13124 | n13128 ;
  assign n13130 = n8727 | n13124 ;
  assign n13131 = n13128 | n13130 ;
  assign n13132 = ( n746 & n13129 ) | ( n746 & n13131 ) | ( n13129 & n13131 ) ;
  assign n13133 = x44 & n13131 ;
  assign n13134 = x44 & n13124 ;
  assign n13135 = ( x44 & n13128 ) | ( x44 & n13134 ) | ( n13128 & n13134 ) ;
  assign n13136 = ( n746 & n13133 ) | ( n746 & n13135 ) | ( n13133 & n13135 ) ;
  assign n13137 = x44 & ~n13135 ;
  assign n13138 = x44 & ~n13131 ;
  assign n13139 = ( ~n746 & n13137 ) | ( ~n746 & n13138 ) | ( n13137 & n13138 ) ;
  assign n13140 = ( n13132 & ~n13136 ) | ( n13132 & n13139 ) | ( ~n13136 & n13139 ) ;
  assign n13141 = n13123 | n13140 ;
  assign n13142 = n13123 & n13140 ;
  assign n13143 = n13141 & ~n13142 ;
  assign n13144 = n12659 | n12660 ;
  assign n13145 = ( n12565 & n12659 ) | ( n12565 & n13144 ) | ( n12659 & n13144 ) ;
  assign n13146 = n13143 & n13145 ;
  assign n13147 = n13143 | n13145 ;
  assign n13148 = ~n13146 & n13147 ;
  assign n13149 = x78 & n7566 ;
  assign n13150 = x77 & n7561 ;
  assign n13151 = x76 & ~n7560 ;
  assign n13152 = n7953 & n13151 ;
  assign n13153 = n13150 | n13152 ;
  assign n13154 = n13149 | n13153 ;
  assign n13155 = n7569 | n13149 ;
  assign n13156 = n13153 | n13155 ;
  assign n13157 = ( n1192 & n13154 ) | ( n1192 & n13156 ) | ( n13154 & n13156 ) ;
  assign n13158 = x41 & n13156 ;
  assign n13159 = x41 & n13149 ;
  assign n13160 = ( x41 & n13153 ) | ( x41 & n13159 ) | ( n13153 & n13159 ) ;
  assign n13161 = ( n1192 & n13158 ) | ( n1192 & n13160 ) | ( n13158 & n13160 ) ;
  assign n13162 = x41 & ~n13160 ;
  assign n13163 = x41 & ~n13156 ;
  assign n13164 = ( ~n1192 & n13162 ) | ( ~n1192 & n13163 ) | ( n13162 & n13163 ) ;
  assign n13165 = ( n13157 & ~n13161 ) | ( n13157 & n13164 ) | ( ~n13161 & n13164 ) ;
  assign n13166 = n13148 & n13165 ;
  assign n13167 = n13148 & ~n13166 ;
  assign n13168 = ~n13148 & n13165 ;
  assign n13169 = n13167 | n13168 ;
  assign n13170 = n12684 | n12687 ;
  assign n13171 = ( n12684 & n12689 ) | ( n12684 & n13170 ) | ( n12689 & n13170 ) ;
  assign n13172 = n13169 & n13171 ;
  assign n13173 = n13169 | n13171 ;
  assign n13174 = ~n13172 & n13173 ;
  assign n13175 = x81 & n6536 ;
  assign n13176 = x80 & n6531 ;
  assign n13177 = x79 & ~n6530 ;
  assign n13178 = n6871 & n13177 ;
  assign n13179 = n13176 | n13178 ;
  assign n13180 = n13175 | n13179 ;
  assign n13181 = n6539 | n13175 ;
  assign n13182 = n13179 | n13181 ;
  assign n13183 = ( n1651 & n13180 ) | ( n1651 & n13182 ) | ( n13180 & n13182 ) ;
  assign n13184 = x38 & n13182 ;
  assign n13185 = x38 & n13175 ;
  assign n13186 = ( x38 & n13179 ) | ( x38 & n13185 ) | ( n13179 & n13185 ) ;
  assign n13187 = ( n1651 & n13184 ) | ( n1651 & n13186 ) | ( n13184 & n13186 ) ;
  assign n13188 = x38 & ~n13186 ;
  assign n13189 = x38 & ~n13182 ;
  assign n13190 = ( ~n1651 & n13188 ) | ( ~n1651 & n13189 ) | ( n13188 & n13189 ) ;
  assign n13191 = ( n13183 & ~n13187 ) | ( n13183 & n13190 ) | ( ~n13187 & n13190 ) ;
  assign n13192 = n13174 & n13191 ;
  assign n13193 = n13174 & ~n13192 ;
  assign n13194 = ~n13174 & n13191 ;
  assign n13195 = n13193 | n13194 ;
  assign n13196 = n13057 & n13195 ;
  assign n13197 = n13057 & ~n13196 ;
  assign n13198 = ~n13057 & n13195 ;
  assign n13199 = n13197 | n13198 ;
  assign n13200 = x84 & n5554 ;
  assign n13201 = x83 & n5549 ;
  assign n13202 = x82 & ~n5548 ;
  assign n13203 = n5893 & n13202 ;
  assign n13204 = n13201 | n13203 ;
  assign n13205 = n13200 | n13204 ;
  assign n13206 = n5557 | n13200 ;
  assign n13207 = n13204 | n13206 ;
  assign n13208 = ( n2194 & n13205 ) | ( n2194 & n13207 ) | ( n13205 & n13207 ) ;
  assign n13209 = x35 & n13207 ;
  assign n13210 = x35 & n13200 ;
  assign n13211 = ( x35 & n13204 ) | ( x35 & n13210 ) | ( n13204 & n13210 ) ;
  assign n13212 = ( n2194 & n13209 ) | ( n2194 & n13211 ) | ( n13209 & n13211 ) ;
  assign n13213 = x35 & ~n13211 ;
  assign n13214 = x35 & ~n13207 ;
  assign n13215 = ( ~n2194 & n13213 ) | ( ~n2194 & n13214 ) | ( n13213 & n13214 ) ;
  assign n13216 = ( n13208 & ~n13212 ) | ( n13208 & n13215 ) | ( ~n13212 & n13215 ) ;
  assign n13217 = n13195 & n13216 ;
  assign n13218 = ~n13057 & n13217 ;
  assign n13219 = ( n13197 & n13216 ) | ( n13197 & n13218 ) | ( n13216 & n13218 ) ;
  assign n13220 = n13199 & ~n13219 ;
  assign n13221 = ~n13195 & n13216 ;
  assign n13222 = ( n13057 & n13216 ) | ( n13057 & n13221 ) | ( n13216 & n13221 ) ;
  assign n13223 = ~n13197 & n13222 ;
  assign n13224 = n13220 | n13223 ;
  assign n13225 = n13056 & n13224 ;
  assign n13226 = n13056 | n13224 ;
  assign n13227 = ~n13225 & n13226 ;
  assign n13228 = x87 & n4631 ;
  assign n13229 = x86 & n4626 ;
  assign n13230 = x85 & ~n4625 ;
  assign n13231 = n4943 & n13230 ;
  assign n13232 = n13229 | n13231 ;
  assign n13233 = n13228 | n13232 ;
  assign n13234 = n4634 | n13228 ;
  assign n13235 = n13232 | n13234 ;
  assign n13236 = ( n2816 & n13233 ) | ( n2816 & n13235 ) | ( n13233 & n13235 ) ;
  assign n13237 = x32 & n13235 ;
  assign n13238 = x32 & n13228 ;
  assign n13239 = ( x32 & n13232 ) | ( x32 & n13238 ) | ( n13232 & n13238 ) ;
  assign n13240 = ( n2816 & n13237 ) | ( n2816 & n13239 ) | ( n13237 & n13239 ) ;
  assign n13241 = x32 & ~n13239 ;
  assign n13242 = x32 & ~n13235 ;
  assign n13243 = ( ~n2816 & n13241 ) | ( ~n2816 & n13242 ) | ( n13241 & n13242 ) ;
  assign n13244 = ( n13236 & ~n13240 ) | ( n13236 & n13243 ) | ( ~n13240 & n13243 ) ;
  assign n13245 = n13227 & n13244 ;
  assign n13246 = n13227 & ~n13245 ;
  assign n13247 = ~n13227 & n13244 ;
  assign n13248 = n13246 | n13247 ;
  assign n13249 = n12762 | n12766 ;
  assign n13250 = n12763 | n13249 ;
  assign n13251 = ( n12762 & n12770 ) | ( n12762 & n13250 ) | ( n12770 & n13250 ) ;
  assign n13252 = n13248 & n13251 ;
  assign n13253 = n13248 & ~n13252 ;
  assign n13254 = x90 & n3816 ;
  assign n13255 = x89 & n3811 ;
  assign n13256 = x88 & ~n3810 ;
  assign n13257 = n4067 & n13256 ;
  assign n13258 = n13255 | n13257 ;
  assign n13259 = n13254 | n13258 ;
  assign n13260 = n3819 | n13254 ;
  assign n13261 = n13258 | n13260 ;
  assign n13262 = ( n3519 & n13259 ) | ( n3519 & n13261 ) | ( n13259 & n13261 ) ;
  assign n13263 = x29 & n13261 ;
  assign n13264 = x29 & n13254 ;
  assign n13265 = ( x29 & n13258 ) | ( x29 & n13264 ) | ( n13258 & n13264 ) ;
  assign n13266 = ( n3519 & n13263 ) | ( n3519 & n13265 ) | ( n13263 & n13265 ) ;
  assign n13267 = x29 & ~n13265 ;
  assign n13268 = x29 & ~n13261 ;
  assign n13269 = ( ~n3519 & n13267 ) | ( ~n3519 & n13268 ) | ( n13267 & n13268 ) ;
  assign n13270 = ( n13262 & ~n13266 ) | ( n13262 & n13269 ) | ( ~n13266 & n13269 ) ;
  assign n13271 = n13251 & n13270 ;
  assign n13272 = ~n13248 & n13271 ;
  assign n13273 = ( n13253 & n13270 ) | ( n13253 & n13272 ) | ( n13270 & n13272 ) ;
  assign n13274 = n13251 | n13270 ;
  assign n13275 = ( ~n13248 & n13270 ) | ( ~n13248 & n13274 ) | ( n13270 & n13274 ) ;
  assign n13276 = n13253 | n13275 ;
  assign n13277 = ~n13273 & n13276 ;
  assign n13278 = ( n12307 & n12773 ) | ( n12307 & n12790 ) | ( n12773 & n12790 ) ;
  assign n13279 = n12773 | n12790 ;
  assign n13280 = ( n12312 & n13278 ) | ( n12312 & n13279 ) | ( n13278 & n13279 ) ;
  assign n13281 = n13277 | n13280 ;
  assign n13282 = n13277 & n13280 ;
  assign n13283 = n13281 & ~n13282 ;
  assign n13284 = x93 & n3085 ;
  assign n13285 = x92 & n3080 ;
  assign n13286 = x91 & ~n3079 ;
  assign n13287 = n3309 & n13286 ;
  assign n13288 = n13285 | n13287 ;
  assign n13289 = n13284 | n13288 ;
  assign n13290 = n3088 | n13284 ;
  assign n13291 = n13288 | n13290 ;
  assign n13292 = ( n4305 & n13289 ) | ( n4305 & n13291 ) | ( n13289 & n13291 ) ;
  assign n13293 = x26 & n13291 ;
  assign n13294 = x26 & n13284 ;
  assign n13295 = ( x26 & n13288 ) | ( x26 & n13294 ) | ( n13288 & n13294 ) ;
  assign n13296 = ( n4305 & n13293 ) | ( n4305 & n13295 ) | ( n13293 & n13295 ) ;
  assign n13297 = x26 & ~n13295 ;
  assign n13298 = x26 & ~n13291 ;
  assign n13299 = ( ~n4305 & n13297 ) | ( ~n4305 & n13298 ) | ( n13297 & n13298 ) ;
  assign n13300 = ( n13292 & ~n13296 ) | ( n13292 & n13299 ) | ( ~n13296 & n13299 ) ;
  assign n13301 = n13283 | n13300 ;
  assign n13302 = n13283 & n13300 ;
  assign n13303 = n13301 & ~n13302 ;
  assign n13304 = n12817 | n12822 ;
  assign n13305 = ( n12817 & n12819 ) | ( n12817 & n13304 ) | ( n12819 & n13304 ) ;
  assign n13306 = n13303 & n13305 ;
  assign n13307 = n13303 | n13305 ;
  assign n13308 = ~n13306 & n13307 ;
  assign n13309 = x96 & n2429 ;
  assign n13310 = x95 & n2424 ;
  assign n13311 = x94 & ~n2423 ;
  assign n13312 = n2631 & n13311 ;
  assign n13313 = n13310 | n13312 ;
  assign n13314 = n13309 | n13313 ;
  assign n13315 = n2432 | n13309 ;
  assign n13316 = n13313 | n13315 ;
  assign n13317 = ( n5202 & n13314 ) | ( n5202 & n13316 ) | ( n13314 & n13316 ) ;
  assign n13318 = x23 & n13316 ;
  assign n13319 = x23 & n13309 ;
  assign n13320 = ( x23 & n13313 ) | ( x23 & n13319 ) | ( n13313 & n13319 ) ;
  assign n13321 = ( n5202 & n13318 ) | ( n5202 & n13320 ) | ( n13318 & n13320 ) ;
  assign n13322 = x23 & ~n13320 ;
  assign n13323 = x23 & ~n13316 ;
  assign n13324 = ( ~n5202 & n13322 ) | ( ~n5202 & n13323 ) | ( n13322 & n13323 ) ;
  assign n13325 = ( n13317 & ~n13321 ) | ( n13317 & n13324 ) | ( ~n13321 & n13324 ) ;
  assign n13326 = n13308 | n13325 ;
  assign n13327 = n13308 & n13325 ;
  assign n13328 = n13326 & ~n13327 ;
  assign n13329 = n12843 & n13328 ;
  assign n13330 = ( n12849 & n13328 ) | ( n12849 & n13329 ) | ( n13328 & n13329 ) ;
  assign n13331 = n12843 | n13328 ;
  assign n13332 = n12849 | n13331 ;
  assign n13333 = ~n13330 & n13332 ;
  assign n13334 = x99 & n1859 ;
  assign n13335 = x98 & n1854 ;
  assign n13336 = x97 & ~n1853 ;
  assign n13337 = n2037 & n13336 ;
  assign n13338 = n13335 | n13337 ;
  assign n13339 = n13334 | n13338 ;
  assign n13340 = n1862 | n13334 ;
  assign n13341 = n13338 | n13340 ;
  assign n13342 = ( n6164 & n13339 ) | ( n6164 & n13341 ) | ( n13339 & n13341 ) ;
  assign n13343 = x20 & n13341 ;
  assign n13344 = x20 & n13334 ;
  assign n13345 = ( x20 & n13338 ) | ( x20 & n13344 ) | ( n13338 & n13344 ) ;
  assign n13346 = ( n6164 & n13343 ) | ( n6164 & n13345 ) | ( n13343 & n13345 ) ;
  assign n13347 = x20 & ~n13345 ;
  assign n13348 = x20 & ~n13341 ;
  assign n13349 = ( ~n6164 & n13347 ) | ( ~n6164 & n13348 ) | ( n13347 & n13348 ) ;
  assign n13350 = ( n13342 & ~n13346 ) | ( n13342 & n13349 ) | ( ~n13346 & n13349 ) ;
  assign n13351 = n13333 & n13350 ;
  assign n13352 = n13333 & ~n13351 ;
  assign n13353 = ~n13333 & n13350 ;
  assign n13354 = n13352 | n13353 ;
  assign n13355 = n12874 | n12878 ;
  assign n13356 = ( n12874 & n12877 ) | ( n12874 & n13355 ) | ( n12877 & n13355 ) ;
  assign n13357 = n13354 | n13356 ;
  assign n13358 = n13354 & n13356 ;
  assign n13359 = n13357 & ~n13358 ;
  assign n13360 = x102 & n1383 ;
  assign n13361 = x101 & n1378 ;
  assign n13362 = x100 & ~n1377 ;
  assign n13363 = n1542 & n13362 ;
  assign n13364 = n13361 | n13363 ;
  assign n13365 = n13360 | n13364 ;
  assign n13366 = n1386 | n13360 ;
  assign n13367 = n13364 | n13366 ;
  assign n13368 = ( n7178 & n13365 ) | ( n7178 & n13367 ) | ( n13365 & n13367 ) ;
  assign n13369 = x17 & n13367 ;
  assign n13370 = x17 & n13360 ;
  assign n13371 = ( x17 & n13364 ) | ( x17 & n13370 ) | ( n13364 & n13370 ) ;
  assign n13372 = ( n7178 & n13369 ) | ( n7178 & n13371 ) | ( n13369 & n13371 ) ;
  assign n13373 = x17 & ~n13371 ;
  assign n13374 = x17 & ~n13367 ;
  assign n13375 = ( ~n7178 & n13373 ) | ( ~n7178 & n13374 ) | ( n13373 & n13374 ) ;
  assign n13376 = ( n13368 & ~n13372 ) | ( n13368 & n13375 ) | ( ~n13372 & n13375 ) ;
  assign n13377 = n13359 & n13376 ;
  assign n13378 = n13359 & ~n13377 ;
  assign n13379 = ~n13359 & n13376 ;
  assign n13380 = n13378 | n13379 ;
  assign n13381 = n12899 | n12904 ;
  assign n13382 = ( n12899 & n12902 ) | ( n12899 & n13381 ) | ( n12902 & n13381 ) ;
  assign n13383 = n13380 | n13382 ;
  assign n13384 = n13380 & n13382 ;
  assign n13385 = n13383 & ~n13384 ;
  assign n13386 = x105 & n962 ;
  assign n13387 = x104 & n957 ;
  assign n13388 = x103 & ~n956 ;
  assign n13389 = n1105 & n13388 ;
  assign n13390 = n13387 | n13389 ;
  assign n13391 = n13386 | n13390 ;
  assign n13392 = n965 | n13386 ;
  assign n13393 = n13390 | n13392 ;
  assign n13394 = ( n8273 & n13391 ) | ( n8273 & n13393 ) | ( n13391 & n13393 ) ;
  assign n13395 = x14 & n13393 ;
  assign n13396 = x14 & n13386 ;
  assign n13397 = ( x14 & n13390 ) | ( x14 & n13396 ) | ( n13390 & n13396 ) ;
  assign n13398 = ( n8273 & n13395 ) | ( n8273 & n13397 ) | ( n13395 & n13397 ) ;
  assign n13399 = x14 & ~n13397 ;
  assign n13400 = x14 & ~n13393 ;
  assign n13401 = ( ~n8273 & n13399 ) | ( ~n8273 & n13400 ) | ( n13399 & n13400 ) ;
  assign n13402 = ( n13394 & ~n13398 ) | ( n13394 & n13401 ) | ( ~n13398 & n13401 ) ;
  assign n13403 = n13385 & n13402 ;
  assign n13404 = n13385 & ~n13403 ;
  assign n13405 = ~n13385 & n13402 ;
  assign n13406 = n13404 | n13405 ;
  assign n13407 = n12925 | n12931 ;
  assign n13408 = n13406 | n13407 ;
  assign n13409 = n13406 & n13407 ;
  assign n13410 = n13408 & ~n13409 ;
  assign n13411 = x108 & n636 ;
  assign n13412 = x107 & n631 ;
  assign n13413 = x106 & ~n630 ;
  assign n13414 = n764 & n13413 ;
  assign n13415 = n13412 | n13414 ;
  assign n13416 = n13411 | n13415 ;
  assign n13417 = n639 | n13411 ;
  assign n13418 = n13415 | n13417 ;
  assign n13419 = ( n9479 & n13416 ) | ( n9479 & n13418 ) | ( n13416 & n13418 ) ;
  assign n13420 = x11 & n13418 ;
  assign n13421 = x11 & n13411 ;
  assign n13422 = ( x11 & n13415 ) | ( x11 & n13421 ) | ( n13415 & n13421 ) ;
  assign n13423 = ( n9479 & n13420 ) | ( n9479 & n13422 ) | ( n13420 & n13422 ) ;
  assign n13424 = x11 & ~n13422 ;
  assign n13425 = x11 & ~n13418 ;
  assign n13426 = ( ~n9479 & n13424 ) | ( ~n9479 & n13425 ) | ( n13424 & n13425 ) ;
  assign n13427 = ( n13419 & ~n13423 ) | ( n13419 & n13426 ) | ( ~n13423 & n13426 ) ;
  assign n13428 = n13410 & n13427 ;
  assign n13429 = n13410 | n13427 ;
  assign n13430 = ~n13428 & n13429 ;
  assign n13431 = n12950 | n12955 ;
  assign n13432 = n13430 & n13431 ;
  assign n13433 = n13431 & ~n13432 ;
  assign n13434 = ( n13430 & ~n13432 ) | ( n13430 & n13433 ) | ( ~n13432 & n13433 ) ;
  assign n13435 = x111 & n389 ;
  assign n13436 = x110 & n384 ;
  assign n13437 = x109 & ~n383 ;
  assign n13438 = n463 & n13437 ;
  assign n13439 = n13436 | n13438 ;
  assign n13440 = n13435 | n13439 ;
  assign n13441 = n392 | n13435 ;
  assign n13442 = n13439 | n13441 ;
  assign n13443 = ( n10749 & n13440 ) | ( n10749 & n13442 ) | ( n13440 & n13442 ) ;
  assign n13444 = x8 & n13442 ;
  assign n13445 = x8 & n13435 ;
  assign n13446 = ( x8 & n13439 ) | ( x8 & n13445 ) | ( n13439 & n13445 ) ;
  assign n13447 = ( n10749 & n13444 ) | ( n10749 & n13446 ) | ( n13444 & n13446 ) ;
  assign n13448 = x8 & ~n13446 ;
  assign n13449 = x8 & ~n13442 ;
  assign n13450 = ( ~n10749 & n13448 ) | ( ~n10749 & n13449 ) | ( n13448 & n13449 ) ;
  assign n13451 = ( n13443 & ~n13447 ) | ( n13443 & n13450 ) | ( ~n13447 & n13450 ) ;
  assign n13452 = ~n13432 & n13451 ;
  assign n13453 = n13430 & n13451 ;
  assign n13454 = ( n13433 & n13452 ) | ( n13433 & n13453 ) | ( n13452 & n13453 ) ;
  assign n13455 = n13434 & ~n13454 ;
  assign n13456 = n13432 & n13451 ;
  assign n13457 = ~n13430 & n13451 ;
  assign n13458 = ( ~n13433 & n13456 ) | ( ~n13433 & n13457 ) | ( n13456 & n13457 ) ;
  assign n13459 = n13455 | n13458 ;
  assign n13460 = n12977 | n12983 ;
  assign n13461 = ( n12977 & n12982 ) | ( n12977 & n13460 ) | ( n12982 & n13460 ) ;
  assign n13462 = n13459 | n13461 ;
  assign n13463 = n13459 & n13461 ;
  assign n13464 = n13462 & ~n13463 ;
  assign n13465 = x114 & n212 ;
  assign n13466 = x113 & n207 ;
  assign n13467 = x112 & ~n206 ;
  assign n13468 = n267 & n13467 ;
  assign n13469 = n13466 | n13468 ;
  assign n13470 = n13465 | n13469 ;
  assign n13471 = n215 | n13465 ;
  assign n13472 = n13469 | n13471 ;
  assign n13473 = ( ~n12095 & n13470 ) | ( ~n12095 & n13472 ) | ( n13470 & n13472 ) ;
  assign n13474 = n13470 & n13472 ;
  assign n13475 = ( n12079 & n13473 ) | ( n12079 & n13474 ) | ( n13473 & n13474 ) ;
  assign n13476 = x5 & n13475 ;
  assign n13477 = x5 & ~n13475 ;
  assign n13478 = ( n13475 & ~n13476 ) | ( n13475 & n13477 ) | ( ~n13476 & n13477 ) ;
  assign n13479 = n13464 & n13478 ;
  assign n13480 = n13464 | n13478 ;
  assign n13481 = ~n13479 & n13480 ;
  assign n13482 = ( n12512 & n12986 ) | ( n12512 & n13000 ) | ( n12986 & n13000 ) ;
  assign n13483 = n12986 | n13000 ;
  assign n13484 = ( n12516 & n13482 ) | ( n12516 & n13483 ) | ( n13482 & n13483 ) ;
  assign n13485 = n13481 & n13484 ;
  assign n13486 = ~n13481 & n13484 ;
  assign n13487 = ( n13481 & ~n13485 ) | ( n13481 & n13486 ) | ( ~n13485 & n13486 ) ;
  assign n13488 = x116 | x117 ;
  assign n13489 = x116 & x117 ;
  assign n13490 = n13488 & ~n13489 ;
  assign n13491 = n13010 | n13033 ;
  assign n13492 = n13010 | n13011 ;
  assign n13493 = n12520 | n13010 ;
  assign n13494 = ( n13010 & n13011 ) | ( n13010 & n13493 ) | ( n13011 & n13493 ) ;
  assign n13495 = ( n12543 & n13492 ) | ( n12543 & n13494 ) | ( n13492 & n13494 ) ;
  assign n13496 = ( n10726 & n13491 ) | ( n10726 & n13495 ) | ( n13491 & n13495 ) ;
  assign n13497 = n13491 | n13495 ;
  assign n13498 = ( n10735 & n13496 ) | ( n10735 & n13497 ) | ( n13496 & n13497 ) ;
  assign n13499 = ( n10736 & n13496 ) | ( n10736 & n13497 ) | ( n13496 & n13497 ) ;
  assign n13500 = ( n6159 & n13498 ) | ( n6159 & n13499 ) | ( n13498 & n13499 ) ;
  assign n13501 = ( n6157 & n13498 ) | ( n6157 & n13499 ) | ( n13498 & n13499 ) ;
  assign n13502 = ( n5823 & n13500 ) | ( n5823 & n13501 ) | ( n13500 & n13501 ) ;
  assign n13503 = n13490 | n13502 ;
  assign n13504 = x116 & n133 ;
  assign n13505 = x115 & ~n162 ;
  assign n13506 = ( n137 & n13504 ) | ( n137 & n13505 ) | ( n13504 & n13505 ) ;
  assign n13507 = x0 & x117 ;
  assign n13508 = ( ~n137 & n13504 ) | ( ~n137 & n13507 ) | ( n13504 & n13507 ) ;
  assign n13509 = n13506 | n13508 ;
  assign n13510 = n141 | n13509 ;
  assign n13511 = n13490 & n13494 ;
  assign n13512 = n13490 & n13492 ;
  assign n13513 = ( n12543 & n13511 ) | ( n12543 & n13512 ) | ( n13511 & n13512 ) ;
  assign n13514 = n13010 & n13490 ;
  assign n13515 = ( n13033 & n13490 ) | ( n13033 & n13514 ) | ( n13490 & n13514 ) ;
  assign n13516 = ( n10726 & n13513 ) | ( n10726 & n13515 ) | ( n13513 & n13515 ) ;
  assign n13517 = n13513 | n13515 ;
  assign n13518 = ( n10735 & n13516 ) | ( n10735 & n13517 ) | ( n13516 & n13517 ) ;
  assign n13519 = ( n10736 & n13516 ) | ( n10736 & n13517 ) | ( n13516 & n13517 ) ;
  assign n13520 = ( n6159 & n13518 ) | ( n6159 & n13519 ) | ( n13518 & n13519 ) ;
  assign n13521 = ( n6157 & n13518 ) | ( n6157 & n13519 ) | ( n13518 & n13519 ) ;
  assign n13522 = ( n5823 & n13520 ) | ( n5823 & n13521 ) | ( n13520 & n13521 ) ;
  assign n13523 = ( n13509 & n13510 ) | ( n13509 & ~n13522 ) | ( n13510 & ~n13522 ) ;
  assign n13524 = n13509 & n13510 ;
  assign n13525 = ( n13503 & n13523 ) | ( n13503 & n13524 ) | ( n13523 & n13524 ) ;
  assign n13526 = x2 & n13525 ;
  assign n13527 = x2 & ~n13525 ;
  assign n13528 = ( n13525 & ~n13526 ) | ( n13525 & n13527 ) | ( ~n13526 & n13527 ) ;
  assign n13529 = n13487 & ~n13528 ;
  assign n13530 = ~n13487 & n13528 ;
  assign n13531 = n13529 | n13530 ;
  assign n13532 = n13055 & n13531 ;
  assign n13533 = n13055 | n13531 ;
  assign n13534 = ~n13532 & n13533 ;
  assign n13535 = n13428 | n13432 ;
  assign n13536 = n13302 | n13306 ;
  assign n13537 = n13166 | n13172 ;
  assign n13538 = n13107 | n13111 ;
  assign n13539 = x53 & ~x54 ;
  assign n13540 = ~x53 & x54 ;
  assign n13541 = n13539 | n13540 ;
  assign n13542 = x64 & n13541 ;
  assign n13543 = ~n12589 & n13542 ;
  assign n13544 = ( ~n13088 & n13542 ) | ( ~n13088 & n13543 ) | ( n13542 & n13543 ) ;
  assign n13545 = n12589 & ~n13542 ;
  assign n13546 = n13088 & n13545 ;
  assign n13547 = n13544 | n13546 ;
  assign n13548 = x67 & n12574 ;
  assign n13549 = x66 & n12569 ;
  assign n13550 = x65 & ~n12568 ;
  assign n13551 = n13076 & n13550 ;
  assign n13552 = n13549 | n13551 ;
  assign n13553 = n13548 | n13552 ;
  assign n13554 = n186 & n12577 ;
  assign n13555 = n13553 | n13554 ;
  assign n13556 = x53 & ~n13555 ;
  assign n13557 = ~x53 & n13555 ;
  assign n13558 = n13556 | n13557 ;
  assign n13559 = n13547 & n13558 ;
  assign n13560 = n13547 | n13558 ;
  assign n13561 = ~n13559 & n13560 ;
  assign n13562 = x69 & n11200 ;
  assign n13563 = x68 & ~n11199 ;
  assign n13564 = n11679 & n13563 ;
  assign n13565 = n13562 | n13564 ;
  assign n13566 = x70 & n11205 ;
  assign n13567 = n11208 | n13566 ;
  assign n13568 = n13565 | n13567 ;
  assign n13569 = x50 & ~n13568 ;
  assign n13570 = x50 & ~n13566 ;
  assign n13571 = ~n13565 & n13570 ;
  assign n13572 = ( ~n340 & n13569 ) | ( ~n340 & n13571 ) | ( n13569 & n13571 ) ;
  assign n13573 = ~x50 & n13568 ;
  assign n13574 = ~x50 & n13566 ;
  assign n13575 = ( ~x50 & n13565 ) | ( ~x50 & n13574 ) | ( n13565 & n13574 ) ;
  assign n13576 = ( n340 & n13573 ) | ( n340 & n13575 ) | ( n13573 & n13575 ) ;
  assign n13577 = n13572 | n13576 ;
  assign n13578 = n13561 & n13577 ;
  assign n13579 = n13561 & ~n13578 ;
  assign n13580 = ~n13561 & n13577 ;
  assign n13581 = n13538 & n13580 ;
  assign n13582 = ( n13538 & n13579 ) | ( n13538 & n13581 ) | ( n13579 & n13581 ) ;
  assign n13583 = n13538 | n13580 ;
  assign n13584 = n13579 | n13583 ;
  assign n13585 = ~n13582 & n13584 ;
  assign n13586 = x73 & n9933 ;
  assign n13587 = x72 & n9928 ;
  assign n13588 = x71 & ~n9927 ;
  assign n13589 = n10379 & n13588 ;
  assign n13590 = n13587 | n13589 ;
  assign n13591 = n13586 | n13590 ;
  assign n13592 = ( ~n610 & n9936 ) | ( ~n610 & n13591 ) | ( n9936 & n13591 ) ;
  assign n13593 = n9936 & n13586 ;
  assign n13594 = ( n9936 & n13590 ) | ( n9936 & n13593 ) | ( n13590 & n13593 ) ;
  assign n13595 = ( n598 & n13592 ) | ( n598 & n13594 ) | ( n13592 & n13594 ) ;
  assign n13596 = ( x47 & ~n13591 ) | ( x47 & n13595 ) | ( ~n13591 & n13595 ) ;
  assign n13597 = ~n13595 & n13596 ;
  assign n13598 = x47 | n13586 ;
  assign n13599 = n13590 | n13598 ;
  assign n13600 = n13595 | n13599 ;
  assign n13601 = ( ~x47 & n13597 ) | ( ~x47 & n13600 ) | ( n13597 & n13600 ) ;
  assign n13602 = n13585 & n13601 ;
  assign n13603 = n13585 & ~n13602 ;
  assign n13604 = ~n13585 & n13601 ;
  assign n13605 = n13603 | n13604 ;
  assign n13606 = n13115 | n13120 ;
  assign n13607 = n13605 & n13606 ;
  assign n13608 = n13605 | n13606 ;
  assign n13609 = ~n13607 & n13608 ;
  assign n13610 = x76 & n8724 ;
  assign n13611 = x75 & n8719 ;
  assign n13612 = x74 & ~n8718 ;
  assign n13613 = n9149 & n13612 ;
  assign n13614 = n13611 | n13613 ;
  assign n13615 = n13610 | n13614 ;
  assign n13616 = n8727 | n13610 ;
  assign n13617 = n13614 | n13616 ;
  assign n13618 = ( n923 & n13615 ) | ( n923 & n13617 ) | ( n13615 & n13617 ) ;
  assign n13619 = x44 & n13617 ;
  assign n13620 = x44 & n13610 ;
  assign n13621 = ( x44 & n13614 ) | ( x44 & n13620 ) | ( n13614 & n13620 ) ;
  assign n13622 = ( n923 & n13619 ) | ( n923 & n13621 ) | ( n13619 & n13621 ) ;
  assign n13623 = x44 & ~n13621 ;
  assign n13624 = x44 & ~n13617 ;
  assign n13625 = ( ~n923 & n13623 ) | ( ~n923 & n13624 ) | ( n13623 & n13624 ) ;
  assign n13626 = ( n13618 & ~n13622 ) | ( n13618 & n13625 ) | ( ~n13622 & n13625 ) ;
  assign n13627 = n13609 & n13626 ;
  assign n13628 = n13609 & ~n13627 ;
  assign n13629 = n13142 | n13143 ;
  assign n13630 = ( n13142 & n13145 ) | ( n13142 & n13629 ) | ( n13145 & n13629 ) ;
  assign n13631 = ~n13609 & n13626 ;
  assign n13632 = n13630 & n13631 ;
  assign n13633 = ( n13628 & n13630 ) | ( n13628 & n13632 ) | ( n13630 & n13632 ) ;
  assign n13634 = n13630 | n13631 ;
  assign n13635 = n13628 | n13634 ;
  assign n13636 = ~n13633 & n13635 ;
  assign n13637 = x79 & n7566 ;
  assign n13638 = x78 & n7561 ;
  assign n13639 = x77 & ~n7560 ;
  assign n13640 = n7953 & n13639 ;
  assign n13641 = n13638 | n13640 ;
  assign n13642 = n13637 | n13641 ;
  assign n13643 = n7569 | n13637 ;
  assign n13644 = n13641 | n13643 ;
  assign n13645 = ( n1332 & n13642 ) | ( n1332 & n13644 ) | ( n13642 & n13644 ) ;
  assign n13646 = x41 & n13644 ;
  assign n13647 = x41 & n13637 ;
  assign n13648 = ( x41 & n13641 ) | ( x41 & n13647 ) | ( n13641 & n13647 ) ;
  assign n13649 = ( n1332 & n13646 ) | ( n1332 & n13648 ) | ( n13646 & n13648 ) ;
  assign n13650 = x41 & ~n13648 ;
  assign n13651 = x41 & ~n13644 ;
  assign n13652 = ( ~n1332 & n13650 ) | ( ~n1332 & n13651 ) | ( n13650 & n13651 ) ;
  assign n13653 = ( n13645 & ~n13649 ) | ( n13645 & n13652 ) | ( ~n13649 & n13652 ) ;
  assign n13654 = n13636 & n13653 ;
  assign n13655 = n13636 | n13653 ;
  assign n13656 = ~n13654 & n13655 ;
  assign n13657 = n13537 & n13656 ;
  assign n13658 = n13537 | n13656 ;
  assign n13659 = ~n13657 & n13658 ;
  assign n13660 = x82 & n6536 ;
  assign n13661 = x81 & n6531 ;
  assign n13662 = x80 & ~n6530 ;
  assign n13663 = n6871 & n13662 ;
  assign n13664 = n13661 | n13663 ;
  assign n13665 = n13660 | n13664 ;
  assign n13666 = n6539 | n13660 ;
  assign n13667 = n13664 | n13666 ;
  assign n13668 = ( n1811 & n13665 ) | ( n1811 & n13667 ) | ( n13665 & n13667 ) ;
  assign n13669 = x38 & n13667 ;
  assign n13670 = x38 & n13660 ;
  assign n13671 = ( x38 & n13664 ) | ( x38 & n13670 ) | ( n13664 & n13670 ) ;
  assign n13672 = ( n1811 & n13669 ) | ( n1811 & n13671 ) | ( n13669 & n13671 ) ;
  assign n13673 = x38 & ~n13671 ;
  assign n13674 = x38 & ~n13667 ;
  assign n13675 = ( ~n1811 & n13673 ) | ( ~n1811 & n13674 ) | ( n13673 & n13674 ) ;
  assign n13676 = ( n13668 & ~n13672 ) | ( n13668 & n13675 ) | ( ~n13672 & n13675 ) ;
  assign n13677 = n13659 & n13676 ;
  assign n13678 = n13659 & ~n13677 ;
  assign n13679 = ~n13659 & n13676 ;
  assign n13680 = n13678 | n13679 ;
  assign n13681 = n13192 | n13194 ;
  assign n13682 = n13193 | n13681 ;
  assign n13683 = ( n13057 & n13192 ) | ( n13057 & n13682 ) | ( n13192 & n13682 ) ;
  assign n13684 = n13680 & n13683 ;
  assign n13685 = n13680 | n13683 ;
  assign n13686 = ~n13684 & n13685 ;
  assign n13687 = x85 & n5554 ;
  assign n13688 = x84 & n5549 ;
  assign n13689 = x83 & ~n5548 ;
  assign n13690 = n5893 & n13689 ;
  assign n13691 = n13688 | n13690 ;
  assign n13692 = n13687 | n13691 ;
  assign n13693 = n5557 | n13687 ;
  assign n13694 = n13691 | n13693 ;
  assign n13695 = ( n2381 & n13692 ) | ( n2381 & n13694 ) | ( n13692 & n13694 ) ;
  assign n13696 = x35 & n13694 ;
  assign n13697 = x35 & n13687 ;
  assign n13698 = ( x35 & n13691 ) | ( x35 & n13697 ) | ( n13691 & n13697 ) ;
  assign n13699 = ( n2381 & n13696 ) | ( n2381 & n13698 ) | ( n13696 & n13698 ) ;
  assign n13700 = x35 & ~n13698 ;
  assign n13701 = x35 & ~n13694 ;
  assign n13702 = ( ~n2381 & n13700 ) | ( ~n2381 & n13701 ) | ( n13700 & n13701 ) ;
  assign n13703 = ( n13695 & ~n13699 ) | ( n13695 & n13702 ) | ( ~n13699 & n13702 ) ;
  assign n13704 = n13686 & n13703 ;
  assign n13705 = n13686 | n13703 ;
  assign n13706 = ~n13704 & n13705 ;
  assign n13707 = n13056 | n13219 ;
  assign n13708 = ( n13219 & n13224 ) | ( n13219 & n13707 ) | ( n13224 & n13707 ) ;
  assign n13709 = n13706 & n13708 ;
  assign n13710 = n13706 | n13708 ;
  assign n13711 = ~n13709 & n13710 ;
  assign n13712 = x88 & n4631 ;
  assign n13713 = x87 & n4626 ;
  assign n13714 = x86 & ~n4625 ;
  assign n13715 = n4943 & n13714 ;
  assign n13716 = n13713 | n13715 ;
  assign n13717 = n13712 | n13716 ;
  assign n13718 = n4634 | n13712 ;
  assign n13719 = n13716 | n13718 ;
  assign n13720 = ( ~n3039 & n13717 ) | ( ~n3039 & n13719 ) | ( n13717 & n13719 ) ;
  assign n13721 = n13717 & n13719 ;
  assign n13722 = ( n3023 & n13720 ) | ( n3023 & n13721 ) | ( n13720 & n13721 ) ;
  assign n13723 = x32 & n13719 ;
  assign n13724 = x32 & n13712 ;
  assign n13725 = ( x32 & n13716 ) | ( x32 & n13724 ) | ( n13716 & n13724 ) ;
  assign n13726 = ( ~n3039 & n13723 ) | ( ~n3039 & n13725 ) | ( n13723 & n13725 ) ;
  assign n13727 = n13723 & n13725 ;
  assign n13728 = ( n3023 & n13726 ) | ( n3023 & n13727 ) | ( n13726 & n13727 ) ;
  assign n13729 = x32 & ~n13725 ;
  assign n13730 = x32 & ~n13719 ;
  assign n13731 = ( n3039 & n13729 ) | ( n3039 & n13730 ) | ( n13729 & n13730 ) ;
  assign n13732 = n13729 | n13730 ;
  assign n13733 = ( ~n3023 & n13731 ) | ( ~n3023 & n13732 ) | ( n13731 & n13732 ) ;
  assign n13734 = ( n13722 & ~n13728 ) | ( n13722 & n13733 ) | ( ~n13728 & n13733 ) ;
  assign n13735 = n13711 & n13734 ;
  assign n13736 = n13711 | n13734 ;
  assign n13737 = ~n13735 & n13736 ;
  assign n13738 = n13245 & n13737 ;
  assign n13739 = ( n13252 & n13737 ) | ( n13252 & n13738 ) | ( n13737 & n13738 ) ;
  assign n13740 = n13245 | n13737 ;
  assign n13741 = n13252 | n13740 ;
  assign n13742 = ~n13739 & n13741 ;
  assign n13743 = x91 & n3816 ;
  assign n13744 = x90 & n3811 ;
  assign n13745 = x89 & ~n3810 ;
  assign n13746 = n4067 & n13745 ;
  assign n13747 = n13744 | n13746 ;
  assign n13748 = n13743 | n13747 ;
  assign n13749 = n3819 | n13743 ;
  assign n13750 = n13747 | n13749 ;
  assign n13751 = ( n3768 & n13748 ) | ( n3768 & n13750 ) | ( n13748 & n13750 ) ;
  assign n13752 = x29 & n13750 ;
  assign n13753 = x29 & n13743 ;
  assign n13754 = ( x29 & n13747 ) | ( x29 & n13753 ) | ( n13747 & n13753 ) ;
  assign n13755 = ( n3768 & n13752 ) | ( n3768 & n13754 ) | ( n13752 & n13754 ) ;
  assign n13756 = x29 & ~n13754 ;
  assign n13757 = x29 & ~n13750 ;
  assign n13758 = ( ~n3768 & n13756 ) | ( ~n3768 & n13757 ) | ( n13756 & n13757 ) ;
  assign n13759 = ( n13751 & ~n13755 ) | ( n13751 & n13758 ) | ( ~n13755 & n13758 ) ;
  assign n13760 = n13742 & n13759 ;
  assign n13761 = n13742 | n13759 ;
  assign n13762 = ~n13760 & n13761 ;
  assign n13763 = n13273 | n13762 ;
  assign n13764 = n13282 | n13763 ;
  assign n13765 = ( n13273 & n13282 ) | ( n13273 & n13762 ) | ( n13282 & n13762 ) ;
  assign n13766 = x94 & n3085 ;
  assign n13767 = x93 & n3080 ;
  assign n13768 = x92 & ~n3079 ;
  assign n13769 = n3309 & n13768 ;
  assign n13770 = n13767 | n13769 ;
  assign n13771 = n13766 | n13770 ;
  assign n13772 = n3088 | n13766 ;
  assign n13773 = n13770 | n13772 ;
  assign n13774 = ( n4583 & n13771 ) | ( n4583 & n13773 ) | ( n13771 & n13773 ) ;
  assign n13775 = x26 & n13773 ;
  assign n13776 = x26 & n13766 ;
  assign n13777 = ( x26 & n13770 ) | ( x26 & n13776 ) | ( n13770 & n13776 ) ;
  assign n13778 = ( n4583 & n13775 ) | ( n4583 & n13777 ) | ( n13775 & n13777 ) ;
  assign n13779 = x26 & ~n13777 ;
  assign n13780 = x26 & ~n13773 ;
  assign n13781 = ( ~n4583 & n13779 ) | ( ~n4583 & n13780 ) | ( n13779 & n13780 ) ;
  assign n13782 = ( n13774 & ~n13778 ) | ( n13774 & n13781 ) | ( ~n13778 & n13781 ) ;
  assign n13783 = ~n13765 & n13782 ;
  assign n13784 = n13764 & n13783 ;
  assign n13785 = n13765 & ~n13782 ;
  assign n13786 = ( n13764 & n13782 ) | ( n13764 & ~n13785 ) | ( n13782 & ~n13785 ) ;
  assign n13787 = ~n13784 & n13786 ;
  assign n13788 = n13536 & n13787 ;
  assign n13789 = n13536 | n13787 ;
  assign n13790 = ~n13788 & n13789 ;
  assign n13791 = x97 & n2429 ;
  assign n13792 = x96 & n2424 ;
  assign n13793 = x95 & ~n2423 ;
  assign n13794 = n2631 & n13793 ;
  assign n13795 = n13792 | n13794 ;
  assign n13796 = n13791 | n13795 ;
  assign n13797 = n2432 | n13791 ;
  assign n13798 = n13795 | n13797 ;
  assign n13799 = ( n5505 & n13796 ) | ( n5505 & n13798 ) | ( n13796 & n13798 ) ;
  assign n13800 = x23 & n13798 ;
  assign n13801 = x23 & n13791 ;
  assign n13802 = ( x23 & n13795 ) | ( x23 & n13801 ) | ( n13795 & n13801 ) ;
  assign n13803 = ( n5505 & n13800 ) | ( n5505 & n13802 ) | ( n13800 & n13802 ) ;
  assign n13804 = x23 & ~n13802 ;
  assign n13805 = x23 & ~n13798 ;
  assign n13806 = ( ~n5505 & n13804 ) | ( ~n5505 & n13805 ) | ( n13804 & n13805 ) ;
  assign n13807 = ( n13799 & ~n13803 ) | ( n13799 & n13806 ) | ( ~n13803 & n13806 ) ;
  assign n13808 = n13790 & n13807 ;
  assign n13809 = n13790 & ~n13808 ;
  assign n13810 = ~n13790 & n13807 ;
  assign n13811 = n13809 | n13810 ;
  assign n13812 = n13327 | n13330 ;
  assign n13813 = ~n13811 & n13812 ;
  assign n13814 = n13811 & ~n13812 ;
  assign n13815 = n13813 | n13814 ;
  assign n13816 = x100 & n1859 ;
  assign n13817 = x99 & n1854 ;
  assign n13818 = x98 & ~n1853 ;
  assign n13819 = n2037 & n13818 ;
  assign n13820 = n13817 | n13819 ;
  assign n13821 = n13816 | n13820 ;
  assign n13822 = n1862 | n13816 ;
  assign n13823 = n13820 | n13822 ;
  assign n13824 = ( n6483 & n13821 ) | ( n6483 & n13823 ) | ( n13821 & n13823 ) ;
  assign n13825 = x20 & n13823 ;
  assign n13826 = x20 & n13816 ;
  assign n13827 = ( x20 & n13820 ) | ( x20 & n13826 ) | ( n13820 & n13826 ) ;
  assign n13828 = ( n6483 & n13825 ) | ( n6483 & n13827 ) | ( n13825 & n13827 ) ;
  assign n13829 = x20 & ~n13827 ;
  assign n13830 = x20 & ~n13823 ;
  assign n13831 = ( ~n6483 & n13829 ) | ( ~n6483 & n13830 ) | ( n13829 & n13830 ) ;
  assign n13832 = ( n13824 & ~n13828 ) | ( n13824 & n13831 ) | ( ~n13828 & n13831 ) ;
  assign n13833 = n13815 & n13832 ;
  assign n13834 = n13815 | n13832 ;
  assign n13835 = ~n13833 & n13834 ;
  assign n13836 = n13351 | n13358 ;
  assign n13837 = n13835 | n13836 ;
  assign n13838 = n13835 & n13836 ;
  assign n13839 = n13837 & ~n13838 ;
  assign n13840 = x103 & n1383 ;
  assign n13841 = x102 & n1378 ;
  assign n13842 = x101 & ~n1377 ;
  assign n13843 = n1542 & n13842 ;
  assign n13844 = n13841 | n13843 ;
  assign n13845 = n13840 | n13844 ;
  assign n13846 = n1386 | n13840 ;
  assign n13847 = n13844 | n13846 ;
  assign n13848 = ( n7529 & n13845 ) | ( n7529 & n13847 ) | ( n13845 & n13847 ) ;
  assign n13849 = x17 & n13847 ;
  assign n13850 = x17 & n13840 ;
  assign n13851 = ( x17 & n13844 ) | ( x17 & n13850 ) | ( n13844 & n13850 ) ;
  assign n13852 = ( n7529 & n13849 ) | ( n7529 & n13851 ) | ( n13849 & n13851 ) ;
  assign n13853 = x17 & ~n13851 ;
  assign n13854 = x17 & ~n13847 ;
  assign n13855 = ( ~n7529 & n13853 ) | ( ~n7529 & n13854 ) | ( n13853 & n13854 ) ;
  assign n13856 = ( n13848 & ~n13852 ) | ( n13848 & n13855 ) | ( ~n13852 & n13855 ) ;
  assign n13857 = n13839 & n13856 ;
  assign n13858 = n13839 & ~n13857 ;
  assign n13859 = ~n13839 & n13856 ;
  assign n13860 = n13858 | n13859 ;
  assign n13861 = n13377 | n13384 ;
  assign n13862 = n13860 | n13861 ;
  assign n13863 = n13860 & n13861 ;
  assign n13864 = n13862 & ~n13863 ;
  assign n13865 = x106 & n962 ;
  assign n13866 = x105 & n957 ;
  assign n13867 = x104 & ~n956 ;
  assign n13868 = n1105 & n13867 ;
  assign n13869 = n13866 | n13868 ;
  assign n13870 = n13865 | n13869 ;
  assign n13871 = n965 | n13865 ;
  assign n13872 = n13869 | n13871 ;
  assign n13873 = ( n8656 & n13870 ) | ( n8656 & n13872 ) | ( n13870 & n13872 ) ;
  assign n13874 = x14 & n13872 ;
  assign n13875 = x14 & n13865 ;
  assign n13876 = ( x14 & n13869 ) | ( x14 & n13875 ) | ( n13869 & n13875 ) ;
  assign n13877 = ( n8656 & n13874 ) | ( n8656 & n13876 ) | ( n13874 & n13876 ) ;
  assign n13878 = x14 & ~n13876 ;
  assign n13879 = x14 & ~n13872 ;
  assign n13880 = ( ~n8656 & n13878 ) | ( ~n8656 & n13879 ) | ( n13878 & n13879 ) ;
  assign n13881 = ( n13873 & ~n13877 ) | ( n13873 & n13880 ) | ( ~n13877 & n13880 ) ;
  assign n13882 = n13864 | n13881 ;
  assign n13883 = n13864 & n13881 ;
  assign n13884 = n13882 & ~n13883 ;
  assign n13885 = n13403 & n13884 ;
  assign n13886 = ( n13409 & n13884 ) | ( n13409 & n13885 ) | ( n13884 & n13885 ) ;
  assign n13887 = n13403 | n13884 ;
  assign n13888 = n13409 | n13887 ;
  assign n13889 = ~n13886 & n13888 ;
  assign n13890 = x109 & n636 ;
  assign n13891 = x108 & n631 ;
  assign n13892 = x107 & ~n630 ;
  assign n13893 = n764 & n13892 ;
  assign n13894 = n13891 | n13893 ;
  assign n13895 = n13890 | n13894 ;
  assign n13896 = n639 | n13890 ;
  assign n13897 = n13894 | n13896 ;
  assign n13898 = ( n9878 & n13895 ) | ( n9878 & n13897 ) | ( n13895 & n13897 ) ;
  assign n13899 = x11 & n13897 ;
  assign n13900 = x11 & n13890 ;
  assign n13901 = ( x11 & n13894 ) | ( x11 & n13900 ) | ( n13894 & n13900 ) ;
  assign n13902 = ( n9878 & n13899 ) | ( n9878 & n13901 ) | ( n13899 & n13901 ) ;
  assign n13903 = x11 & ~n13901 ;
  assign n13904 = x11 & ~n13897 ;
  assign n13905 = ( ~n9878 & n13903 ) | ( ~n9878 & n13904 ) | ( n13903 & n13904 ) ;
  assign n13906 = ( n13898 & ~n13902 ) | ( n13898 & n13905 ) | ( ~n13902 & n13905 ) ;
  assign n13907 = n13889 & n13906 ;
  assign n13908 = n13889 & ~n13907 ;
  assign n13909 = ~n13889 & n13906 ;
  assign n13910 = n13908 | n13909 ;
  assign n13911 = n13535 & n13910 ;
  assign n13912 = n13535 & ~n13911 ;
  assign n13913 = n13910 & ~n13911 ;
  assign n13914 = n13912 | n13913 ;
  assign n13915 = x112 & n389 ;
  assign n13916 = x111 & n384 ;
  assign n13917 = x110 & ~n383 ;
  assign n13918 = n463 & n13917 ;
  assign n13919 = n13916 | n13918 ;
  assign n13920 = n13915 | n13919 ;
  assign n13921 = n392 | n13915 ;
  assign n13922 = n13919 | n13921 ;
  assign n13923 = ( n11172 & n13920 ) | ( n11172 & n13922 ) | ( n13920 & n13922 ) ;
  assign n13924 = x8 & n13922 ;
  assign n13925 = x8 & n13915 ;
  assign n13926 = ( x8 & n13919 ) | ( x8 & n13925 ) | ( n13919 & n13925 ) ;
  assign n13927 = ( n11172 & n13924 ) | ( n11172 & n13926 ) | ( n13924 & n13926 ) ;
  assign n13928 = x8 & ~n13926 ;
  assign n13929 = x8 & ~n13922 ;
  assign n13930 = ( ~n11172 & n13928 ) | ( ~n11172 & n13929 ) | ( n13928 & n13929 ) ;
  assign n13931 = ( n13923 & ~n13927 ) | ( n13923 & n13930 ) | ( ~n13927 & n13930 ) ;
  assign n13932 = n13914 & n13931 ;
  assign n13933 = n13914 & ~n13932 ;
  assign n13934 = n13454 | n13461 ;
  assign n13935 = ( n13454 & n13459 ) | ( n13454 & n13934 ) | ( n13459 & n13934 ) ;
  assign n13936 = ~n13914 & n13931 ;
  assign n13937 = n13935 & n13936 ;
  assign n13938 = ( n13933 & n13935 ) | ( n13933 & n13937 ) | ( n13935 & n13937 ) ;
  assign n13939 = n13935 | n13936 ;
  assign n13940 = n13933 | n13939 ;
  assign n13941 = ~n13938 & n13940 ;
  assign n13942 = x115 & n212 ;
  assign n13943 = x114 & n207 ;
  assign n13944 = x113 & ~n206 ;
  assign n13945 = n267 & n13944 ;
  assign n13946 = n13943 | n13945 ;
  assign n13947 = n13942 | n13946 ;
  assign n13948 = n215 | n13942 ;
  assign n13949 = n13946 | n13948 ;
  assign n13950 = ( ~n12550 & n13947 ) | ( ~n12550 & n13949 ) | ( n13947 & n13949 ) ;
  assign n13951 = n13947 & n13949 ;
  assign n13952 = ( n12532 & n13950 ) | ( n12532 & n13951 ) | ( n13950 & n13951 ) ;
  assign n13953 = x5 & n13952 ;
  assign n13954 = x5 & ~n13952 ;
  assign n13955 = ( n13952 & ~n13953 ) | ( n13952 & n13954 ) | ( ~n13953 & n13954 ) ;
  assign n13956 = n13941 | n13955 ;
  assign n13957 = n13941 & n13955 ;
  assign n13958 = n13956 & ~n13957 ;
  assign n13959 = n13479 | n13484 ;
  assign n13960 = ( n13479 & n13481 ) | ( n13479 & n13959 ) | ( n13481 & n13959 ) ;
  assign n13961 = n13958 & n13960 ;
  assign n13962 = n13958 | n13960 ;
  assign n13963 = ~n13961 & n13962 ;
  assign n13964 = x117 | x118 ;
  assign n13965 = x117 & x118 ;
  assign n13966 = n13964 & ~n13965 ;
  assign n13967 = n13489 | n13490 ;
  assign n13968 = n13010 | n13489 ;
  assign n13969 = ( n13489 & n13490 ) | ( n13489 & n13968 ) | ( n13490 & n13968 ) ;
  assign n13970 = ( n13033 & n13967 ) | ( n13033 & n13969 ) | ( n13967 & n13969 ) ;
  assign n13971 = n13489 | n13512 ;
  assign n13972 = n13489 | n13511 ;
  assign n13973 = ( n12543 & n13971 ) | ( n12543 & n13972 ) | ( n13971 & n13972 ) ;
  assign n13974 = ( n10726 & n13970 ) | ( n10726 & n13973 ) | ( n13970 & n13973 ) ;
  assign n13975 = n13970 | n13973 ;
  assign n13976 = ( n10735 & n13974 ) | ( n10735 & n13975 ) | ( n13974 & n13975 ) ;
  assign n13977 = ( n10736 & n13974 ) | ( n10736 & n13975 ) | ( n13974 & n13975 ) ;
  assign n13978 = ( n6159 & n13976 ) | ( n6159 & n13977 ) | ( n13976 & n13977 ) ;
  assign n13979 = ( n6157 & n13976 ) | ( n6157 & n13977 ) | ( n13976 & n13977 ) ;
  assign n13980 = ( n5823 & n13978 ) | ( n5823 & n13979 ) | ( n13978 & n13979 ) ;
  assign n13981 = n13966 | n13980 ;
  assign n13982 = x117 & n133 ;
  assign n13983 = x116 & ~n162 ;
  assign n13984 = ( n137 & n13982 ) | ( n137 & n13983 ) | ( n13982 & n13983 ) ;
  assign n13985 = x0 & x118 ;
  assign n13986 = ( ~n137 & n13982 ) | ( ~n137 & n13985 ) | ( n13982 & n13985 ) ;
  assign n13987 = n13984 | n13986 ;
  assign n13988 = n141 | n13987 ;
  assign n13989 = n13966 & n13969 ;
  assign n13990 = n13966 & n13967 ;
  assign n13991 = ( n13033 & n13989 ) | ( n13033 & n13990 ) | ( n13989 & n13990 ) ;
  assign n13992 = n13489 & n13966 ;
  assign n13993 = ( n13512 & n13966 ) | ( n13512 & n13992 ) | ( n13966 & n13992 ) ;
  assign n13994 = ( n13511 & n13966 ) | ( n13511 & n13992 ) | ( n13966 & n13992 ) ;
  assign n13995 = ( n12543 & n13993 ) | ( n12543 & n13994 ) | ( n13993 & n13994 ) ;
  assign n13996 = ( n10726 & n13991 ) | ( n10726 & n13995 ) | ( n13991 & n13995 ) ;
  assign n13997 = n13991 | n13995 ;
  assign n13998 = ( n10735 & n13996 ) | ( n10735 & n13997 ) | ( n13996 & n13997 ) ;
  assign n13999 = ( n10736 & n13996 ) | ( n10736 & n13997 ) | ( n13996 & n13997 ) ;
  assign n14000 = ( n6159 & n13998 ) | ( n6159 & n13999 ) | ( n13998 & n13999 ) ;
  assign n14001 = ( n6157 & n13998 ) | ( n6157 & n13999 ) | ( n13998 & n13999 ) ;
  assign n14002 = ( n5823 & n14000 ) | ( n5823 & n14001 ) | ( n14000 & n14001 ) ;
  assign n14003 = ( n13987 & n13988 ) | ( n13987 & ~n14002 ) | ( n13988 & ~n14002 ) ;
  assign n14004 = n13987 & n13988 ;
  assign n14005 = ( n13981 & n14003 ) | ( n13981 & n14004 ) | ( n14003 & n14004 ) ;
  assign n14006 = x2 & n14005 ;
  assign n14007 = x2 & ~n14005 ;
  assign n14008 = ( n14005 & ~n14006 ) | ( n14005 & n14007 ) | ( ~n14006 & n14007 ) ;
  assign n14009 = n13963 & n14008 ;
  assign n14010 = n13963 | n14008 ;
  assign n14011 = ~n14009 & n14010 ;
  assign n14012 = ( n13047 & n13487 ) | ( n13047 & n13528 ) | ( n13487 & n13528 ) ;
  assign n14013 = n13487 | n13528 ;
  assign n14014 = ( n13052 & n14012 ) | ( n13052 & n14013 ) | ( n14012 & n14013 ) ;
  assign n14015 = n14011 | n14014 ;
  assign n14016 = n14011 & n14014 ;
  assign n14017 = n14015 & ~n14016 ;
  assign n14018 = n13883 | n13886 ;
  assign n14019 = n13677 | n13684 ;
  assign n14020 = n13627 | n13633 ;
  assign n14021 = x70 & n11200 ;
  assign n14022 = x69 & ~n11199 ;
  assign n14023 = n11679 & n14022 ;
  assign n14024 = n14021 | n14023 ;
  assign n14025 = x71 & n11205 ;
  assign n14026 = n11208 | n14025 ;
  assign n14027 = n14024 | n14026 ;
  assign n14028 = x50 & ~n14027 ;
  assign n14029 = x50 & ~n14025 ;
  assign n14030 = ~n14024 & n14029 ;
  assign n14031 = ( ~n438 & n14028 ) | ( ~n438 & n14030 ) | ( n14028 & n14030 ) ;
  assign n14032 = ~x50 & n14027 ;
  assign n14033 = ~x50 & n14025 ;
  assign n14034 = ( ~x50 & n14024 ) | ( ~x50 & n14033 ) | ( n14024 & n14033 ) ;
  assign n14035 = ( n438 & n14032 ) | ( n438 & n14034 ) | ( n14032 & n14034 ) ;
  assign n14036 = n14031 | n14035 ;
  assign n14037 = ~x54 & x55 ;
  assign n14038 = x54 & ~x55 ;
  assign n14039 = n14037 | n14038 ;
  assign n14040 = ~n13541 & n14039 ;
  assign n14041 = x64 & n14040 ;
  assign n14042 = ~x55 & x56 ;
  assign n14043 = x55 & ~x56 ;
  assign n14044 = n14042 | n14043 ;
  assign n14045 = n13541 & ~n14044 ;
  assign n14046 = x65 & n14045 ;
  assign n14047 = n14041 | n14046 ;
  assign n14048 = n13541 & n14044 ;
  assign n14049 = x56 | n144 ;
  assign n14050 = ( x56 & n14048 ) | ( x56 & n14049 ) | ( n14048 & n14049 ) ;
  assign n14051 = ~x56 & n14050 ;
  assign n14052 = ( ~x56 & n14047 ) | ( ~x56 & n14051 ) | ( n14047 & n14051 ) ;
  assign n14053 = x56 & ~x64 ;
  assign n14054 = ( x56 & ~n13541 ) | ( x56 & n14053 ) | ( ~n13541 & n14053 ) ;
  assign n14055 = n14050 & n14054 ;
  assign n14056 = ( n14047 & n14054 ) | ( n14047 & n14055 ) | ( n14054 & n14055 ) ;
  assign n14057 = n144 & n14048 ;
  assign n14058 = n14054 & ~n14057 ;
  assign n14059 = ~n14047 & n14058 ;
  assign n14060 = ( n14052 & n14056 ) | ( n14052 & n14059 ) | ( n14056 & n14059 ) ;
  assign n14061 = n14050 | n14054 ;
  assign n14062 = n14047 | n14061 ;
  assign n14063 = ~n14054 & n14057 ;
  assign n14064 = ( n14047 & ~n14054 ) | ( n14047 & n14063 ) | ( ~n14054 & n14063 ) ;
  assign n14065 = ( n14052 & n14062 ) | ( n14052 & ~n14064 ) | ( n14062 & ~n14064 ) ;
  assign n14066 = ~n14060 & n14065 ;
  assign n14067 = n241 & n12577 ;
  assign n14068 = x68 & n12574 ;
  assign n14069 = x67 & n12569 ;
  assign n14070 = x66 & ~n12568 ;
  assign n14071 = n13076 & n14070 ;
  assign n14072 = n14069 | n14071 ;
  assign n14073 = n14068 | n14072 ;
  assign n14074 = n14067 | n14073 ;
  assign n14075 = x53 | n14068 ;
  assign n14076 = n14072 | n14075 ;
  assign n14077 = n14067 | n14076 ;
  assign n14078 = ~x53 & n14076 ;
  assign n14079 = ( ~x53 & n14067 ) | ( ~x53 & n14078 ) | ( n14067 & n14078 ) ;
  assign n14080 = ( ~n14074 & n14077 ) | ( ~n14074 & n14079 ) | ( n14077 & n14079 ) ;
  assign n14081 = n14066 | n14080 ;
  assign n14082 = n14066 & n14080 ;
  assign n14083 = n14081 & ~n14082 ;
  assign n14084 = ( n13090 & n13542 ) | ( n13090 & n13558 ) | ( n13542 & n13558 ) ;
  assign n14085 = n14083 | n14084 ;
  assign n14086 = n14083 & n14084 ;
  assign n14087 = n14085 & ~n14086 ;
  assign n14088 = n14036 | n14087 ;
  assign n14089 = n14036 & n14087 ;
  assign n14090 = n14088 & ~n14089 ;
  assign n14091 = n13578 | n13579 ;
  assign n14092 = n13538 | n13578 ;
  assign n14093 = ( n13581 & n14091 ) | ( n13581 & n14092 ) | ( n14091 & n14092 ) ;
  assign n14094 = n14090 & n14093 ;
  assign n14095 = n14090 | n14093 ;
  assign n14096 = ~n14094 & n14095 ;
  assign n14097 = x74 & n9933 ;
  assign n14098 = x73 & n9928 ;
  assign n14099 = x72 & ~n9927 ;
  assign n14100 = n10379 & n14099 ;
  assign n14101 = n14098 | n14100 ;
  assign n14102 = n14097 | n14101 ;
  assign n14103 = n9936 | n14097 ;
  assign n14104 = n14101 | n14103 ;
  assign n14105 = ( n710 & n14102 ) | ( n710 & n14104 ) | ( n14102 & n14104 ) ;
  assign n14106 = x47 & n14104 ;
  assign n14107 = x47 & n14097 ;
  assign n14108 = ( x47 & n14101 ) | ( x47 & n14107 ) | ( n14101 & n14107 ) ;
  assign n14109 = ( n710 & n14106 ) | ( n710 & n14108 ) | ( n14106 & n14108 ) ;
  assign n14110 = x47 & ~n14108 ;
  assign n14111 = x47 & ~n14104 ;
  assign n14112 = ( ~n710 & n14110 ) | ( ~n710 & n14111 ) | ( n14110 & n14111 ) ;
  assign n14113 = ( n14105 & ~n14109 ) | ( n14105 & n14112 ) | ( ~n14109 & n14112 ) ;
  assign n14114 = n14096 | n14113 ;
  assign n14115 = n14096 & n14113 ;
  assign n14116 = n14114 & ~n14115 ;
  assign n14117 = n13602 | n13606 ;
  assign n14118 = ( n13602 & n13605 ) | ( n13602 & n14117 ) | ( n13605 & n14117 ) ;
  assign n14119 = n14116 & n14118 ;
  assign n14120 = n14116 | n14118 ;
  assign n14121 = ~n14119 & n14120 ;
  assign n14122 = x77 & n8724 ;
  assign n14123 = x76 & n8719 ;
  assign n14124 = x75 & ~n8718 ;
  assign n14125 = n9149 & n14124 ;
  assign n14126 = n14123 | n14125 ;
  assign n14127 = n14122 | n14126 ;
  assign n14128 = n8727 | n14122 ;
  assign n14129 = n14126 | n14128 ;
  assign n14130 = ( n1059 & n14127 ) | ( n1059 & n14129 ) | ( n14127 & n14129 ) ;
  assign n14131 = x44 & n14129 ;
  assign n14132 = x44 & n14122 ;
  assign n14133 = ( x44 & n14126 ) | ( x44 & n14132 ) | ( n14126 & n14132 ) ;
  assign n14134 = ( n1059 & n14131 ) | ( n1059 & n14133 ) | ( n14131 & n14133 ) ;
  assign n14135 = x44 & ~n14133 ;
  assign n14136 = x44 & ~n14129 ;
  assign n14137 = ( ~n1059 & n14135 ) | ( ~n1059 & n14136 ) | ( n14135 & n14136 ) ;
  assign n14138 = ( n14130 & ~n14134 ) | ( n14130 & n14137 ) | ( ~n14134 & n14137 ) ;
  assign n14139 = n14121 | n14138 ;
  assign n14140 = n14121 & n14138 ;
  assign n14141 = n14139 & ~n14140 ;
  assign n14142 = n14020 & n14141 ;
  assign n14143 = n14020 | n14141 ;
  assign n14144 = ~n14142 & n14143 ;
  assign n14145 = x80 & n7566 ;
  assign n14146 = x79 & n7561 ;
  assign n14147 = x78 & ~n7560 ;
  assign n14148 = n7953 & n14147 ;
  assign n14149 = n14146 | n14148 ;
  assign n14150 = n14145 | n14149 ;
  assign n14151 = n7569 | n14145 ;
  assign n14152 = n14149 | n14151 ;
  assign n14153 = ( n1499 & n14150 ) | ( n1499 & n14152 ) | ( n14150 & n14152 ) ;
  assign n14154 = x41 & n14152 ;
  assign n14155 = x41 & n14145 ;
  assign n14156 = ( x41 & n14149 ) | ( x41 & n14155 ) | ( n14149 & n14155 ) ;
  assign n14157 = ( n1499 & n14154 ) | ( n1499 & n14156 ) | ( n14154 & n14156 ) ;
  assign n14158 = x41 & ~n14156 ;
  assign n14159 = x41 & ~n14152 ;
  assign n14160 = ( ~n1499 & n14158 ) | ( ~n1499 & n14159 ) | ( n14158 & n14159 ) ;
  assign n14161 = ( n14153 & ~n14157 ) | ( n14153 & n14160 ) | ( ~n14157 & n14160 ) ;
  assign n14162 = n14144 & n14161 ;
  assign n14163 = n14144 & ~n14162 ;
  assign n14164 = ~n14144 & n14161 ;
  assign n14165 = n14163 | n14164 ;
  assign n14166 = n13654 | n13656 ;
  assign n14167 = ( n13537 & n13654 ) | ( n13537 & n14166 ) | ( n13654 & n14166 ) ;
  assign n14168 = n14165 | n14167 ;
  assign n14169 = n14165 & n14167 ;
  assign n14170 = n14168 & ~n14169 ;
  assign n14171 = x83 & n6536 ;
  assign n14172 = x82 & n6531 ;
  assign n14173 = x81 & ~n6530 ;
  assign n14174 = n6871 & n14173 ;
  assign n14175 = n14172 | n14174 ;
  assign n14176 = n14171 | n14175 ;
  assign n14177 = n6539 | n14171 ;
  assign n14178 = n14175 | n14177 ;
  assign n14179 = ( n2009 & n14176 ) | ( n2009 & n14178 ) | ( n14176 & n14178 ) ;
  assign n14180 = x38 & n14178 ;
  assign n14181 = x38 & n14171 ;
  assign n14182 = ( x38 & n14175 ) | ( x38 & n14181 ) | ( n14175 & n14181 ) ;
  assign n14183 = ( n2009 & n14180 ) | ( n2009 & n14182 ) | ( n14180 & n14182 ) ;
  assign n14184 = x38 & ~n14182 ;
  assign n14185 = x38 & ~n14178 ;
  assign n14186 = ( ~n2009 & n14184 ) | ( ~n2009 & n14185 ) | ( n14184 & n14185 ) ;
  assign n14187 = ( n14179 & ~n14183 ) | ( n14179 & n14186 ) | ( ~n14183 & n14186 ) ;
  assign n14188 = n14170 & n14187 ;
  assign n14189 = n14170 | n14187 ;
  assign n14190 = ~n14188 & n14189 ;
  assign n14191 = n13677 & n14187 ;
  assign n14192 = ( n13677 & n14170 ) | ( n13677 & n14191 ) | ( n14170 & n14191 ) ;
  assign n14193 = ~n14188 & n14192 ;
  assign n14194 = ( n13684 & n14190 ) | ( n13684 & n14193 ) | ( n14190 & n14193 ) ;
  assign n14195 = n14019 & ~n14194 ;
  assign n14196 = x86 & n5554 ;
  assign n14197 = x85 & n5549 ;
  assign n14198 = x84 & ~n5548 ;
  assign n14199 = n5893 & n14198 ;
  assign n14200 = n14197 | n14199 ;
  assign n14201 = n14196 | n14200 ;
  assign n14202 = n5557 | n14196 ;
  assign n14203 = n14200 | n14202 ;
  assign n14204 = ( n2606 & n14201 ) | ( n2606 & n14203 ) | ( n14201 & n14203 ) ;
  assign n14205 = x35 & n14203 ;
  assign n14206 = x35 & n14196 ;
  assign n14207 = ( x35 & n14200 ) | ( x35 & n14206 ) | ( n14200 & n14206 ) ;
  assign n14208 = ( n2606 & n14205 ) | ( n2606 & n14207 ) | ( n14205 & n14207 ) ;
  assign n14209 = x35 & ~n14207 ;
  assign n14210 = x35 & ~n14203 ;
  assign n14211 = ( ~n2606 & n14209 ) | ( ~n2606 & n14210 ) | ( n14209 & n14210 ) ;
  assign n14212 = ( n14204 & ~n14208 ) | ( n14204 & n14211 ) | ( ~n14208 & n14211 ) ;
  assign n14213 = ( n13684 & n14189 ) | ( n13684 & n14192 ) | ( n14189 & n14192 ) ;
  assign n14214 = n14190 & n14212 ;
  assign n14215 = ~n14213 & n14214 ;
  assign n14216 = ( n14195 & n14212 ) | ( n14195 & n14215 ) | ( n14212 & n14215 ) ;
  assign n14217 = n14190 | n14212 ;
  assign n14218 = ( n14212 & ~n14213 ) | ( n14212 & n14217 ) | ( ~n14213 & n14217 ) ;
  assign n14219 = n14195 | n14218 ;
  assign n14220 = ~n14216 & n14219 ;
  assign n14221 = n13704 | n13706 ;
  assign n14222 = ( n13704 & n13708 ) | ( n13704 & n14221 ) | ( n13708 & n14221 ) ;
  assign n14223 = n14220 | n14222 ;
  assign n14224 = n14220 & n14222 ;
  assign n14225 = n14223 & ~n14224 ;
  assign n14226 = x89 & n4631 ;
  assign n14227 = x88 & n4626 ;
  assign n14228 = x87 & ~n4625 ;
  assign n14229 = n4943 & n14228 ;
  assign n14230 = n14227 | n14229 ;
  assign n14231 = n14226 | n14230 ;
  assign n14232 = n4634 | n14226 ;
  assign n14233 = n14230 | n14232 ;
  assign n14234 = ( n3282 & n14231 ) | ( n3282 & n14233 ) | ( n14231 & n14233 ) ;
  assign n14235 = x32 & n14233 ;
  assign n14236 = x32 & n14226 ;
  assign n14237 = ( x32 & n14230 ) | ( x32 & n14236 ) | ( n14230 & n14236 ) ;
  assign n14238 = ( n3282 & n14235 ) | ( n3282 & n14237 ) | ( n14235 & n14237 ) ;
  assign n14239 = x32 & ~n14237 ;
  assign n14240 = x32 & ~n14233 ;
  assign n14241 = ( ~n3282 & n14239 ) | ( ~n3282 & n14240 ) | ( n14239 & n14240 ) ;
  assign n14242 = ( n14234 & ~n14238 ) | ( n14234 & n14241 ) | ( ~n14238 & n14241 ) ;
  assign n14243 = n14225 & n14242 ;
  assign n14244 = n14225 & ~n14243 ;
  assign n14245 = ~n14225 & n14242 ;
  assign n14246 = n14244 | n14245 ;
  assign n14247 = n13735 | n13739 ;
  assign n14248 = n14246 | n14247 ;
  assign n14249 = n14246 & n14247 ;
  assign n14250 = n14248 & ~n14249 ;
  assign n14251 = x92 & n3816 ;
  assign n14252 = x91 & n3811 ;
  assign n14253 = x90 & ~n3810 ;
  assign n14254 = n4067 & n14253 ;
  assign n14255 = n14252 | n14254 ;
  assign n14256 = n14251 | n14255 ;
  assign n14257 = n3819 | n14251 ;
  assign n14258 = n14255 | n14257 ;
  assign n14259 = ( n4040 & n14256 ) | ( n4040 & n14258 ) | ( n14256 & n14258 ) ;
  assign n14260 = x29 & n14258 ;
  assign n14261 = x29 & n14251 ;
  assign n14262 = ( x29 & n14255 ) | ( x29 & n14261 ) | ( n14255 & n14261 ) ;
  assign n14263 = ( n4040 & n14260 ) | ( n4040 & n14262 ) | ( n14260 & n14262 ) ;
  assign n14264 = x29 & ~n14262 ;
  assign n14265 = x29 & ~n14258 ;
  assign n14266 = ( ~n4040 & n14264 ) | ( ~n4040 & n14265 ) | ( n14264 & n14265 ) ;
  assign n14267 = ( n14259 & ~n14263 ) | ( n14259 & n14266 ) | ( ~n14263 & n14266 ) ;
  assign n14268 = n14250 & n14267 ;
  assign n14269 = n14250 & ~n14268 ;
  assign n14270 = ~n14250 & n14267 ;
  assign n14271 = n14269 | n14270 ;
  assign n14272 = n13760 | n13765 ;
  assign n14273 = n14271 | n14272 ;
  assign n14274 = n14271 & n14272 ;
  assign n14275 = n14273 & ~n14274 ;
  assign n14276 = x95 & n3085 ;
  assign n14277 = x94 & n3080 ;
  assign n14278 = x93 & ~n3079 ;
  assign n14279 = n3309 & n14278 ;
  assign n14280 = n14277 | n14279 ;
  assign n14281 = n14276 | n14280 ;
  assign n14282 = n3088 | n14276 ;
  assign n14283 = n14280 | n14282 ;
  assign n14284 = ( n4897 & n14281 ) | ( n4897 & n14283 ) | ( n14281 & n14283 ) ;
  assign n14285 = x26 & n14283 ;
  assign n14286 = x26 & n14276 ;
  assign n14287 = ( x26 & n14280 ) | ( x26 & n14286 ) | ( n14280 & n14286 ) ;
  assign n14288 = ( n4897 & n14285 ) | ( n4897 & n14287 ) | ( n14285 & n14287 ) ;
  assign n14289 = x26 & ~n14287 ;
  assign n14290 = x26 & ~n14283 ;
  assign n14291 = ( ~n4897 & n14289 ) | ( ~n4897 & n14290 ) | ( n14289 & n14290 ) ;
  assign n14292 = ( n14284 & ~n14288 ) | ( n14284 & n14291 ) | ( ~n14288 & n14291 ) ;
  assign n14293 = n14275 & n14292 ;
  assign n14294 = n14275 & ~n14293 ;
  assign n14295 = n13784 | n13787 ;
  assign n14296 = ( n13536 & n13784 ) | ( n13536 & n14295 ) | ( n13784 & n14295 ) ;
  assign n14297 = ~n14275 & n14292 ;
  assign n14298 = n14296 & n14297 ;
  assign n14299 = ( n14294 & n14296 ) | ( n14294 & n14298 ) | ( n14296 & n14298 ) ;
  assign n14300 = n14296 | n14297 ;
  assign n14301 = n14294 | n14300 ;
  assign n14302 = ~n14299 & n14301 ;
  assign n14303 = x98 & n2429 ;
  assign n14304 = x97 & n2424 ;
  assign n14305 = x96 & ~n2423 ;
  assign n14306 = n2631 & n14305 ;
  assign n14307 = n14304 | n14306 ;
  assign n14308 = n14303 | n14307 ;
  assign n14309 = n2432 | n14303 ;
  assign n14310 = n14307 | n14309 ;
  assign n14311 = ( ~n5850 & n14308 ) | ( ~n5850 & n14310 ) | ( n14308 & n14310 ) ;
  assign n14312 = n14308 & n14310 ;
  assign n14313 = ( n5834 & n14311 ) | ( n5834 & n14312 ) | ( n14311 & n14312 ) ;
  assign n14314 = x23 & n14310 ;
  assign n14315 = x23 & n14303 ;
  assign n14316 = ( x23 & n14307 ) | ( x23 & n14315 ) | ( n14307 & n14315 ) ;
  assign n14317 = ( ~n5850 & n14314 ) | ( ~n5850 & n14316 ) | ( n14314 & n14316 ) ;
  assign n14318 = n14314 & n14316 ;
  assign n14319 = ( n5834 & n14317 ) | ( n5834 & n14318 ) | ( n14317 & n14318 ) ;
  assign n14320 = x23 & ~n14316 ;
  assign n14321 = x23 & ~n14310 ;
  assign n14322 = ( n5850 & n14320 ) | ( n5850 & n14321 ) | ( n14320 & n14321 ) ;
  assign n14323 = n14320 | n14321 ;
  assign n14324 = ( ~n5834 & n14322 ) | ( ~n5834 & n14323 ) | ( n14322 & n14323 ) ;
  assign n14325 = ( n14313 & ~n14319 ) | ( n14313 & n14324 ) | ( ~n14319 & n14324 ) ;
  assign n14326 = n14302 & n14325 ;
  assign n14327 = n14302 & ~n14326 ;
  assign n14328 = ( n13327 & n13790 ) | ( n13327 & n13807 ) | ( n13790 & n13807 ) ;
  assign n14329 = n13790 | n13807 ;
  assign n14330 = ( n13330 & n14328 ) | ( n13330 & n14329 ) | ( n14328 & n14329 ) ;
  assign n14331 = ~n14302 & n14325 ;
  assign n14332 = n14330 & n14331 ;
  assign n14333 = ( n14327 & n14330 ) | ( n14327 & n14332 ) | ( n14330 & n14332 ) ;
  assign n14334 = n14330 | n14331 ;
  assign n14335 = n14327 | n14334 ;
  assign n14336 = ~n14333 & n14335 ;
  assign n14337 = x101 & n1859 ;
  assign n14338 = x100 & n1854 ;
  assign n14339 = x99 & ~n1853 ;
  assign n14340 = n2037 & n14339 ;
  assign n14341 = n14338 | n14340 ;
  assign n14342 = n14337 | n14341 ;
  assign n14343 = n1862 | n14337 ;
  assign n14344 = n14341 | n14343 ;
  assign n14345 = ( n6844 & n14342 ) | ( n6844 & n14344 ) | ( n14342 & n14344 ) ;
  assign n14346 = x20 & n14344 ;
  assign n14347 = x20 & n14337 ;
  assign n14348 = ( x20 & n14341 ) | ( x20 & n14347 ) | ( n14341 & n14347 ) ;
  assign n14349 = ( n6844 & n14346 ) | ( n6844 & n14348 ) | ( n14346 & n14348 ) ;
  assign n14350 = x20 & ~n14348 ;
  assign n14351 = x20 & ~n14344 ;
  assign n14352 = ( ~n6844 & n14350 ) | ( ~n6844 & n14351 ) | ( n14350 & n14351 ) ;
  assign n14353 = ( n14345 & ~n14349 ) | ( n14345 & n14352 ) | ( ~n14349 & n14352 ) ;
  assign n14354 = n14336 & n14353 ;
  assign n14355 = n14336 & ~n14354 ;
  assign n14356 = ~n14336 & n14353 ;
  assign n14357 = n14355 | n14356 ;
  assign n14358 = n13833 | n13835 ;
  assign n14359 = ( n13833 & n13836 ) | ( n13833 & n14358 ) | ( n13836 & n14358 ) ;
  assign n14360 = n14357 | n14359 ;
  assign n14361 = n14357 & n14359 ;
  assign n14362 = n14360 & ~n14361 ;
  assign n14363 = x104 & n1383 ;
  assign n14364 = x103 & n1378 ;
  assign n14365 = x102 & ~n1377 ;
  assign n14366 = n1542 & n14365 ;
  assign n14367 = n14364 | n14366 ;
  assign n14368 = n14363 | n14367 ;
  assign n14369 = n1386 | n14363 ;
  assign n14370 = n14367 | n14369 ;
  assign n14371 = ( n7911 & n14368 ) | ( n7911 & n14370 ) | ( n14368 & n14370 ) ;
  assign n14372 = x17 & n14370 ;
  assign n14373 = x17 & n14363 ;
  assign n14374 = ( x17 & n14367 ) | ( x17 & n14373 ) | ( n14367 & n14373 ) ;
  assign n14375 = ( n7911 & n14372 ) | ( n7911 & n14374 ) | ( n14372 & n14374 ) ;
  assign n14376 = x17 & ~n14374 ;
  assign n14377 = x17 & ~n14370 ;
  assign n14378 = ( ~n7911 & n14376 ) | ( ~n7911 & n14377 ) | ( n14376 & n14377 ) ;
  assign n14379 = ( n14371 & ~n14375 ) | ( n14371 & n14378 ) | ( ~n14375 & n14378 ) ;
  assign n14380 = n14362 & n14379 ;
  assign n14381 = n14362 & ~n14380 ;
  assign n14382 = ~n14362 & n14379 ;
  assign n14383 = n14381 | n14382 ;
  assign n14384 = n13857 | n13863 ;
  assign n14385 = n14383 | n14384 ;
  assign n14386 = n14383 & n14384 ;
  assign n14387 = n14385 & ~n14386 ;
  assign n14388 = x107 & n962 ;
  assign n14389 = x106 & n957 ;
  assign n14390 = x105 & ~n956 ;
  assign n14391 = n1105 & n14390 ;
  assign n14392 = n14389 | n14391 ;
  assign n14393 = n14388 | n14392 ;
  assign n14394 = n965 | n14388 ;
  assign n14395 = n14392 | n14394 ;
  assign n14396 = ( n9084 & n14393 ) | ( n9084 & n14395 ) | ( n14393 & n14395 ) ;
  assign n14397 = x14 & n14395 ;
  assign n14398 = x14 & n14388 ;
  assign n14399 = ( x14 & n14392 ) | ( x14 & n14398 ) | ( n14392 & n14398 ) ;
  assign n14400 = ( n9084 & n14397 ) | ( n9084 & n14399 ) | ( n14397 & n14399 ) ;
  assign n14401 = x14 & ~n14399 ;
  assign n14402 = x14 & ~n14395 ;
  assign n14403 = ( ~n9084 & n14401 ) | ( ~n9084 & n14402 ) | ( n14401 & n14402 ) ;
  assign n14404 = ( n14396 & ~n14400 ) | ( n14396 & n14403 ) | ( ~n14400 & n14403 ) ;
  assign n14405 = n14387 & n14404 ;
  assign n14406 = n14387 | n14404 ;
  assign n14407 = ~n14405 & n14406 ;
  assign n14408 = n13883 & n14404 ;
  assign n14409 = ( n13883 & n14387 ) | ( n13883 & n14408 ) | ( n14387 & n14408 ) ;
  assign n14410 = ~n14405 & n14409 ;
  assign n14411 = ( n13886 & n14407 ) | ( n13886 & n14410 ) | ( n14407 & n14410 ) ;
  assign n14412 = n14018 & ~n14411 ;
  assign n14413 = x110 & n636 ;
  assign n14414 = x109 & n631 ;
  assign n14415 = x108 & ~n630 ;
  assign n14416 = n764 & n14415 ;
  assign n14417 = n14414 | n14416 ;
  assign n14418 = n14413 | n14417 ;
  assign n14419 = n639 | n14413 ;
  assign n14420 = n14417 | n14419 ;
  assign n14421 = ( n10330 & n14418 ) | ( n10330 & n14420 ) | ( n14418 & n14420 ) ;
  assign n14422 = x11 & n14420 ;
  assign n14423 = x11 & n14413 ;
  assign n14424 = ( x11 & n14417 ) | ( x11 & n14423 ) | ( n14417 & n14423 ) ;
  assign n14425 = ( n10330 & n14422 ) | ( n10330 & n14424 ) | ( n14422 & n14424 ) ;
  assign n14426 = x11 & ~n14424 ;
  assign n14427 = x11 & ~n14420 ;
  assign n14428 = ( ~n10330 & n14426 ) | ( ~n10330 & n14427 ) | ( n14426 & n14427 ) ;
  assign n14429 = ( n14421 & ~n14425 ) | ( n14421 & n14428 ) | ( ~n14425 & n14428 ) ;
  assign n14430 = ( n13886 & n14406 ) | ( n13886 & n14409 ) | ( n14406 & n14409 ) ;
  assign n14431 = n14407 & n14429 ;
  assign n14432 = ~n14430 & n14431 ;
  assign n14433 = ( n14412 & n14429 ) | ( n14412 & n14432 ) | ( n14429 & n14432 ) ;
  assign n14434 = n14407 | n14429 ;
  assign n14435 = ( n14429 & ~n14430 ) | ( n14429 & n14434 ) | ( ~n14430 & n14434 ) ;
  assign n14436 = n14412 | n14435 ;
  assign n14437 = ~n14433 & n14436 ;
  assign n14438 = n13907 & n14437 ;
  assign n14439 = ( n13911 & n14437 ) | ( n13911 & n14438 ) | ( n14437 & n14438 ) ;
  assign n14440 = n13907 | n14437 ;
  assign n14441 = n13911 | n14440 ;
  assign n14442 = ~n14439 & n14441 ;
  assign n14443 = x113 & n389 ;
  assign n14444 = x112 & n384 ;
  assign n14445 = x111 & ~n383 ;
  assign n14446 = n463 & n14445 ;
  assign n14447 = n14444 | n14446 ;
  assign n14448 = n14443 | n14447 ;
  assign n14449 = n392 | n14443 ;
  assign n14450 = n14447 | n14449 ;
  assign n14451 = ( ~n11642 & n14448 ) | ( ~n11642 & n14450 ) | ( n14448 & n14450 ) ;
  assign n14452 = n14448 & n14450 ;
  assign n14453 = ( n11626 & n14451 ) | ( n11626 & n14452 ) | ( n14451 & n14452 ) ;
  assign n14454 = x8 & n14453 ;
  assign n14455 = x8 & ~n14453 ;
  assign n14456 = ( n14453 & ~n14454 ) | ( n14453 & n14455 ) | ( ~n14454 & n14455 ) ;
  assign n14457 = n14442 | n14456 ;
  assign n14458 = n14442 & n14456 ;
  assign n14459 = n14457 & ~n14458 ;
  assign n14460 = n13932 & n14459 ;
  assign n14461 = ( n13938 & n14459 ) | ( n13938 & n14460 ) | ( n14459 & n14460 ) ;
  assign n14462 = n13932 | n14459 ;
  assign n14463 = n13938 | n14462 ;
  assign n14464 = ~n14461 & n14463 ;
  assign n14465 = x116 & n212 ;
  assign n14466 = x115 & n207 ;
  assign n14467 = x114 & ~n206 ;
  assign n14468 = n267 & n14467 ;
  assign n14469 = n14466 | n14468 ;
  assign n14470 = n14465 | n14469 ;
  assign n14471 = n215 | n14465 ;
  assign n14472 = n14469 | n14471 ;
  assign n14473 = ( ~n13040 & n14470 ) | ( ~n13040 & n14472 ) | ( n14470 & n14472 ) ;
  assign n14474 = n14470 & n14472 ;
  assign n14475 = ( n13022 & n14473 ) | ( n13022 & n14474 ) | ( n14473 & n14474 ) ;
  assign n14476 = x5 & n14475 ;
  assign n14477 = x5 & ~n14475 ;
  assign n14478 = ( n14475 & ~n14476 ) | ( n14475 & n14477 ) | ( ~n14476 & n14477 ) ;
  assign n14479 = n14464 & n14478 ;
  assign n14480 = n14464 & ~n14479 ;
  assign n14481 = ~n14464 & n14478 ;
  assign n14482 = n13957 | n13960 ;
  assign n14483 = ( n13957 & n13958 ) | ( n13957 & n14482 ) | ( n13958 & n14482 ) ;
  assign n14484 = ~n14481 & n14483 ;
  assign n14485 = ~n14480 & n14484 ;
  assign n14486 = n14481 & ~n14483 ;
  assign n14487 = ( n14480 & ~n14483 ) | ( n14480 & n14486 ) | ( ~n14483 & n14486 ) ;
  assign n14488 = n14485 | n14487 ;
  assign n14489 = x118 | x119 ;
  assign n14490 = x118 & x119 ;
  assign n14491 = n14489 & ~n14490 ;
  assign n14492 = n13965 & n14491 ;
  assign n14493 = ( n14002 & n14491 ) | ( n14002 & n14492 ) | ( n14491 & n14492 ) ;
  assign n14494 = n13965 | n14491 ;
  assign n14495 = n14002 | n14494 ;
  assign n14496 = ~n14493 & n14495 ;
  assign n14497 = x118 & n133 ;
  assign n14498 = x117 & ~n162 ;
  assign n14499 = ( n137 & n14497 ) | ( n137 & n14498 ) | ( n14497 & n14498 ) ;
  assign n14500 = x0 & x119 ;
  assign n14501 = ( ~n137 & n14497 ) | ( ~n137 & n14500 ) | ( n14497 & n14500 ) ;
  assign n14502 = n14499 | n14501 ;
  assign n14503 = n141 | n14502 ;
  assign n14504 = ( n14496 & n14502 ) | ( n14496 & n14503 ) | ( n14502 & n14503 ) ;
  assign n14505 = x2 & n14502 ;
  assign n14506 = ( x2 & n523 ) | ( x2 & n14502 ) | ( n523 & n14502 ) ;
  assign n14507 = ( n14496 & n14505 ) | ( n14496 & n14506 ) | ( n14505 & n14506 ) ;
  assign n14508 = x2 & ~n14506 ;
  assign n14509 = x2 & ~n14502 ;
  assign n14510 = ( ~n14496 & n14508 ) | ( ~n14496 & n14509 ) | ( n14508 & n14509 ) ;
  assign n14511 = ( n14504 & ~n14507 ) | ( n14504 & n14510 ) | ( ~n14507 & n14510 ) ;
  assign n14512 = n14488 & n14511 ;
  assign n14513 = n14488 | n14511 ;
  assign n14514 = ~n14512 & n14513 ;
  assign n14515 = n14009 | n14014 ;
  assign n14516 = ( n14009 & n14011 ) | ( n14009 & n14515 ) | ( n14011 & n14515 ) ;
  assign n14517 = n14514 & n14516 ;
  assign n14518 = n14514 | n14516 ;
  assign n14519 = ~n14517 & n14518 ;
  assign n14520 = x117 & n212 ;
  assign n14521 = x116 & n207 ;
  assign n14522 = x115 & ~n206 ;
  assign n14523 = n267 & n14522 ;
  assign n14524 = n14521 | n14523 ;
  assign n14525 = n14520 | n14524 ;
  assign n14526 = n215 | n14520 ;
  assign n14527 = n14524 | n14526 ;
  assign n14528 = ( ~n13522 & n14525 ) | ( ~n13522 & n14527 ) | ( n14525 & n14527 ) ;
  assign n14529 = n14525 & n14527 ;
  assign n14530 = ( n13503 & n14528 ) | ( n13503 & n14529 ) | ( n14528 & n14529 ) ;
  assign n14531 = x5 & n14530 ;
  assign n14532 = x5 & ~n14530 ;
  assign n14533 = ( n14530 & ~n14531 ) | ( n14530 & n14532 ) | ( ~n14531 & n14532 ) ;
  assign n14672 = n14162 | n14167 ;
  assign n14673 = ( n14162 & n14165 ) | ( n14162 & n14672 ) | ( n14165 & n14672 ) ;
  assign n14534 = x72 & n11205 ;
  assign n14535 = x71 & n11200 ;
  assign n14536 = x70 & ~n11199 ;
  assign n14537 = n11679 & n14536 ;
  assign n14538 = n14535 | n14537 ;
  assign n14539 = n14534 | n14538 ;
  assign n14540 = ( n513 & n11208 ) | ( n513 & n14539 ) | ( n11208 & n14539 ) ;
  assign n14541 = x50 & n11208 ;
  assign n14542 = ( x50 & n11208 ) | ( x50 & ~n14534 ) | ( n11208 & ~n14534 ) ;
  assign n14543 = ( ~n14538 & n14541 ) | ( ~n14538 & n14542 ) | ( n14541 & n14542 ) ;
  assign n14544 = ( x50 & n513 ) | ( x50 & n14543 ) | ( n513 & n14543 ) ;
  assign n14545 = ~n14540 & n14544 ;
  assign n14546 = n14539 | n14543 ;
  assign n14547 = x50 | n14539 ;
  assign n14548 = ( n513 & n14546 ) | ( n513 & n14547 ) | ( n14546 & n14547 ) ;
  assign n14549 = ( ~x50 & n14545 ) | ( ~x50 & n14548 ) | ( n14545 & n14548 ) ;
  assign n14550 = x66 & n14045 ;
  assign n14551 = x65 & n14040 ;
  assign n14552 = ~n13541 & n14044 ;
  assign n14553 = x64 & ~n14039 ;
  assign n14554 = n14552 & n14553 ;
  assign n14555 = n14551 | n14554 ;
  assign n14556 = n14550 | n14555 ;
  assign n14557 = n159 & n14048 ;
  assign n14558 = n14556 | n14557 ;
  assign n14559 = x56 | n14048 ;
  assign n14560 = ( x56 & n159 ) | ( x56 & n14559 ) | ( n159 & n14559 ) ;
  assign n14561 = n14556 | n14560 ;
  assign n14562 = ~x56 & n14560 ;
  assign n14563 = ( ~x56 & n14556 ) | ( ~x56 & n14562 ) | ( n14556 & n14562 ) ;
  assign n14564 = ( ~n14558 & n14561 ) | ( ~n14558 & n14563 ) | ( n14561 & n14563 ) ;
  assign n14565 = n14060 | n14564 ;
  assign n14566 = n14060 & n14564 ;
  assign n14567 = n14565 & ~n14566 ;
  assign n14568 = n293 & n12577 ;
  assign n14569 = x69 & n12574 ;
  assign n14570 = x68 & n12569 ;
  assign n14571 = x67 & ~n12568 ;
  assign n14572 = n13076 & n14571 ;
  assign n14573 = n14570 | n14572 ;
  assign n14574 = n14569 | n14573 ;
  assign n14575 = n14568 | n14574 ;
  assign n14576 = x53 | n14569 ;
  assign n14577 = n14573 | n14576 ;
  assign n14578 = n14568 | n14577 ;
  assign n14579 = ~x53 & n14577 ;
  assign n14580 = ( ~x53 & n14568 ) | ( ~x53 & n14579 ) | ( n14568 & n14579 ) ;
  assign n14581 = ( ~n14575 & n14578 ) | ( ~n14575 & n14580 ) | ( n14578 & n14580 ) ;
  assign n14582 = n14567 | n14581 ;
  assign n14583 = n14567 & n14581 ;
  assign n14584 = n14582 & ~n14583 ;
  assign n14585 = n14082 | n14084 ;
  assign n14586 = ( n14082 & n14083 ) | ( n14082 & n14585 ) | ( n14083 & n14585 ) ;
  assign n14587 = n14584 & n14586 ;
  assign n14588 = n14584 & ~n14587 ;
  assign n14589 = ~n14584 & n14586 ;
  assign n14590 = n14549 & n14589 ;
  assign n14591 = ( n14549 & n14588 ) | ( n14549 & n14590 ) | ( n14588 & n14590 ) ;
  assign n14592 = n14549 | n14589 ;
  assign n14593 = n14588 | n14592 ;
  assign n14594 = ~n14591 & n14593 ;
  assign n14595 = n14089 | n14090 ;
  assign n14596 = ( n14089 & n14093 ) | ( n14089 & n14595 ) | ( n14093 & n14595 ) ;
  assign n14597 = n14594 & n14596 ;
  assign n14598 = n14594 | n14596 ;
  assign n14599 = ~n14597 & n14598 ;
  assign n14600 = x75 & n9933 ;
  assign n14601 = x74 & n9928 ;
  assign n14602 = x73 & ~n9927 ;
  assign n14603 = n10379 & n14602 ;
  assign n14604 = n14601 | n14603 ;
  assign n14605 = n14600 | n14604 ;
  assign n14606 = n9936 | n14600 ;
  assign n14607 = n14604 | n14606 ;
  assign n14608 = ( n746 & n14605 ) | ( n746 & n14607 ) | ( n14605 & n14607 ) ;
  assign n14609 = x47 & n14607 ;
  assign n14610 = x47 & n14600 ;
  assign n14611 = ( x47 & n14604 ) | ( x47 & n14610 ) | ( n14604 & n14610 ) ;
  assign n14612 = ( n746 & n14609 ) | ( n746 & n14611 ) | ( n14609 & n14611 ) ;
  assign n14613 = x47 & ~n14611 ;
  assign n14614 = x47 & ~n14607 ;
  assign n14615 = ( ~n746 & n14613 ) | ( ~n746 & n14614 ) | ( n14613 & n14614 ) ;
  assign n14616 = ( n14608 & ~n14612 ) | ( n14608 & n14615 ) | ( ~n14612 & n14615 ) ;
  assign n14617 = n14599 | n14616 ;
  assign n14618 = n14599 & n14616 ;
  assign n14619 = n14617 & ~n14618 ;
  assign n14620 = n14115 | n14116 ;
  assign n14621 = ( n14115 & n14118 ) | ( n14115 & n14620 ) | ( n14118 & n14620 ) ;
  assign n14622 = n14619 & n14621 ;
  assign n14623 = n14619 | n14621 ;
  assign n14624 = ~n14622 & n14623 ;
  assign n14625 = x78 & n8724 ;
  assign n14626 = x77 & n8719 ;
  assign n14627 = x76 & ~n8718 ;
  assign n14628 = n9149 & n14627 ;
  assign n14629 = n14626 | n14628 ;
  assign n14630 = n14625 | n14629 ;
  assign n14631 = n8727 | n14625 ;
  assign n14632 = n14629 | n14631 ;
  assign n14633 = ( n1192 & n14630 ) | ( n1192 & n14632 ) | ( n14630 & n14632 ) ;
  assign n14634 = x44 & n14632 ;
  assign n14635 = x44 & n14625 ;
  assign n14636 = ( x44 & n14629 ) | ( x44 & n14635 ) | ( n14629 & n14635 ) ;
  assign n14637 = ( n1192 & n14634 ) | ( n1192 & n14636 ) | ( n14634 & n14636 ) ;
  assign n14638 = x44 & ~n14636 ;
  assign n14639 = x44 & ~n14632 ;
  assign n14640 = ( ~n1192 & n14638 ) | ( ~n1192 & n14639 ) | ( n14638 & n14639 ) ;
  assign n14641 = ( n14633 & ~n14637 ) | ( n14633 & n14640 ) | ( ~n14637 & n14640 ) ;
  assign n14642 = n14624 & n14641 ;
  assign n14643 = n14624 & ~n14642 ;
  assign n14644 = ~n14624 & n14641 ;
  assign n14645 = n14643 | n14644 ;
  assign n14646 = n14140 | n14141 ;
  assign n14647 = ( n14020 & n14140 ) | ( n14020 & n14646 ) | ( n14140 & n14646 ) ;
  assign n14648 = n14645 & n14647 ;
  assign n14649 = n14645 | n14647 ;
  assign n14650 = ~n14648 & n14649 ;
  assign n14651 = x81 & n7566 ;
  assign n14652 = x80 & n7561 ;
  assign n14653 = x79 & ~n7560 ;
  assign n14654 = n7953 & n14653 ;
  assign n14655 = n14652 | n14654 ;
  assign n14656 = n14651 | n14655 ;
  assign n14657 = n7569 | n14651 ;
  assign n14658 = n14655 | n14657 ;
  assign n14659 = ( n1651 & n14656 ) | ( n1651 & n14658 ) | ( n14656 & n14658 ) ;
  assign n14660 = x41 & n14658 ;
  assign n14661 = x41 & n14651 ;
  assign n14662 = ( x41 & n14655 ) | ( x41 & n14661 ) | ( n14655 & n14661 ) ;
  assign n14663 = ( n1651 & n14660 ) | ( n1651 & n14662 ) | ( n14660 & n14662 ) ;
  assign n14664 = x41 & ~n14662 ;
  assign n14665 = x41 & ~n14658 ;
  assign n14666 = ( ~n1651 & n14664 ) | ( ~n1651 & n14665 ) | ( n14664 & n14665 ) ;
  assign n14667 = ( n14659 & ~n14663 ) | ( n14659 & n14666 ) | ( ~n14663 & n14666 ) ;
  assign n14668 = n14650 & n14667 ;
  assign n14669 = n14650 & ~n14668 ;
  assign n14670 = ~n14650 & n14667 ;
  assign n14671 = n14669 | n14670 ;
  assign n14674 = n14671 & n14673 ;
  assign n14675 = n14673 & ~n14674 ;
  assign n14676 = n14671 & ~n14674 ;
  assign n14677 = n14675 | n14676 ;
  assign n14678 = x84 & n6536 ;
  assign n14679 = x83 & n6531 ;
  assign n14680 = x82 & ~n6530 ;
  assign n14681 = n6871 & n14680 ;
  assign n14682 = n14679 | n14681 ;
  assign n14683 = n14678 | n14682 ;
  assign n14684 = n6539 | n14678 ;
  assign n14685 = n14682 | n14684 ;
  assign n14686 = ( n2194 & n14683 ) | ( n2194 & n14685 ) | ( n14683 & n14685 ) ;
  assign n14687 = x38 & n14685 ;
  assign n14688 = x38 & n14678 ;
  assign n14689 = ( x38 & n14682 ) | ( x38 & n14688 ) | ( n14682 & n14688 ) ;
  assign n14690 = ( n2194 & n14687 ) | ( n2194 & n14689 ) | ( n14687 & n14689 ) ;
  assign n14691 = x38 & ~n14689 ;
  assign n14692 = x38 & ~n14685 ;
  assign n14693 = ( ~n2194 & n14691 ) | ( ~n2194 & n14692 ) | ( n14691 & n14692 ) ;
  assign n14694 = ( n14686 & ~n14690 ) | ( n14686 & n14693 ) | ( ~n14690 & n14693 ) ;
  assign n14695 = n14677 & n14694 ;
  assign n14696 = n14677 & ~n14695 ;
  assign n14697 = ~n14677 & n14694 ;
  assign n14698 = n14188 | n14192 ;
  assign n14699 = n14188 | n14189 ;
  assign n14700 = ( n13684 & n14698 ) | ( n13684 & n14699 ) | ( n14698 & n14699 ) ;
  assign n14701 = ~n14697 & n14700 ;
  assign n14702 = ~n14696 & n14701 ;
  assign n14703 = n14697 & ~n14700 ;
  assign n14704 = ( n14696 & ~n14700 ) | ( n14696 & n14703 ) | ( ~n14700 & n14703 ) ;
  assign n14705 = n14702 | n14704 ;
  assign n14706 = x87 & n5554 ;
  assign n14707 = x86 & n5549 ;
  assign n14708 = x85 & ~n5548 ;
  assign n14709 = n5893 & n14708 ;
  assign n14710 = n14707 | n14709 ;
  assign n14711 = n14706 | n14710 ;
  assign n14712 = n5557 | n14706 ;
  assign n14713 = n14710 | n14712 ;
  assign n14714 = ( n2816 & n14711 ) | ( n2816 & n14713 ) | ( n14711 & n14713 ) ;
  assign n14715 = x35 & n14713 ;
  assign n14716 = x35 & n14706 ;
  assign n14717 = ( x35 & n14710 ) | ( x35 & n14716 ) | ( n14710 & n14716 ) ;
  assign n14718 = ( n2816 & n14715 ) | ( n2816 & n14717 ) | ( n14715 & n14717 ) ;
  assign n14719 = x35 & ~n14717 ;
  assign n14720 = x35 & ~n14713 ;
  assign n14721 = ( ~n2816 & n14719 ) | ( ~n2816 & n14720 ) | ( n14719 & n14720 ) ;
  assign n14722 = ( n14714 & ~n14718 ) | ( n14714 & n14721 ) | ( ~n14718 & n14721 ) ;
  assign n14723 = n14705 & n14722 ;
  assign n14724 = n14705 | n14722 ;
  assign n14725 = ~n14723 & n14724 ;
  assign n14726 = n14216 | n14220 ;
  assign n14727 = ( n14216 & n14222 ) | ( n14216 & n14726 ) | ( n14222 & n14726 ) ;
  assign n14728 = n14725 | n14727 ;
  assign n14729 = n14725 & n14727 ;
  assign n14730 = n14728 & ~n14729 ;
  assign n14731 = x90 & n4631 ;
  assign n14732 = x89 & n4626 ;
  assign n14733 = x88 & ~n4625 ;
  assign n14734 = n4943 & n14733 ;
  assign n14735 = n14732 | n14734 ;
  assign n14736 = n14731 | n14735 ;
  assign n14737 = n4634 | n14731 ;
  assign n14738 = n14735 | n14737 ;
  assign n14739 = ( n3519 & n14736 ) | ( n3519 & n14738 ) | ( n14736 & n14738 ) ;
  assign n14740 = x32 & n14738 ;
  assign n14741 = x32 & n14731 ;
  assign n14742 = ( x32 & n14735 ) | ( x32 & n14741 ) | ( n14735 & n14741 ) ;
  assign n14743 = ( n3519 & n14740 ) | ( n3519 & n14742 ) | ( n14740 & n14742 ) ;
  assign n14744 = x32 & ~n14742 ;
  assign n14745 = x32 & ~n14738 ;
  assign n14746 = ( ~n3519 & n14744 ) | ( ~n3519 & n14745 ) | ( n14744 & n14745 ) ;
  assign n14747 = ( n14739 & ~n14743 ) | ( n14739 & n14746 ) | ( ~n14743 & n14746 ) ;
  assign n14748 = n14730 & n14747 ;
  assign n14749 = n14730 | n14747 ;
  assign n14750 = ~n14748 & n14749 ;
  assign n14751 = n14243 & n14750 ;
  assign n14752 = ( n14249 & n14750 ) | ( n14249 & n14751 ) | ( n14750 & n14751 ) ;
  assign n14753 = x93 & n3816 ;
  assign n14754 = x92 & n3811 ;
  assign n14755 = x91 & ~n3810 ;
  assign n14756 = n4067 & n14755 ;
  assign n14757 = n14754 | n14756 ;
  assign n14758 = n14753 | n14757 ;
  assign n14759 = n3819 | n14753 ;
  assign n14760 = n14757 | n14759 ;
  assign n14761 = ( n4305 & n14758 ) | ( n4305 & n14760 ) | ( n14758 & n14760 ) ;
  assign n14762 = x29 & n14760 ;
  assign n14763 = x29 & n14753 ;
  assign n14764 = ( x29 & n14757 ) | ( x29 & n14763 ) | ( n14757 & n14763 ) ;
  assign n14765 = ( n4305 & n14762 ) | ( n4305 & n14764 ) | ( n14762 & n14764 ) ;
  assign n14766 = x29 & ~n14764 ;
  assign n14767 = x29 & ~n14760 ;
  assign n14768 = ( ~n4305 & n14766 ) | ( ~n4305 & n14767 ) | ( n14766 & n14767 ) ;
  assign n14769 = ( n14761 & ~n14765 ) | ( n14761 & n14768 ) | ( ~n14765 & n14768 ) ;
  assign n14770 = n14243 | n14245 ;
  assign n14771 = n14244 | n14770 ;
  assign n14772 = n14750 | n14771 ;
  assign n14773 = n14243 | n14750 ;
  assign n14774 = ( n14247 & n14772 ) | ( n14247 & n14773 ) | ( n14772 & n14773 ) ;
  assign n14775 = n14769 & n14774 ;
  assign n14776 = ~n14752 & n14775 ;
  assign n14777 = n14769 | n14774 ;
  assign n14778 = ( ~n14752 & n14769 ) | ( ~n14752 & n14777 ) | ( n14769 & n14777 ) ;
  assign n14779 = ~n14776 & n14778 ;
  assign n14780 = n14268 | n14272 ;
  assign n14781 = ( n14268 & n14271 ) | ( n14268 & n14780 ) | ( n14271 & n14780 ) ;
  assign n14782 = n14779 & n14781 ;
  assign n14783 = n14779 | n14781 ;
  assign n14784 = ~n14782 & n14783 ;
  assign n14785 = x96 & n3085 ;
  assign n14786 = x95 & n3080 ;
  assign n14787 = x94 & ~n3079 ;
  assign n14788 = n3309 & n14787 ;
  assign n14789 = n14786 | n14788 ;
  assign n14790 = n14785 | n14789 ;
  assign n14791 = n3088 | n14785 ;
  assign n14792 = n14789 | n14791 ;
  assign n14793 = ( n5202 & n14790 ) | ( n5202 & n14792 ) | ( n14790 & n14792 ) ;
  assign n14794 = x26 & n14792 ;
  assign n14795 = x26 & n14785 ;
  assign n14796 = ( x26 & n14789 ) | ( x26 & n14795 ) | ( n14789 & n14795 ) ;
  assign n14797 = ( n5202 & n14794 ) | ( n5202 & n14796 ) | ( n14794 & n14796 ) ;
  assign n14798 = x26 & ~n14796 ;
  assign n14799 = x26 & ~n14792 ;
  assign n14800 = ( ~n5202 & n14798 ) | ( ~n5202 & n14799 ) | ( n14798 & n14799 ) ;
  assign n14801 = ( n14793 & ~n14797 ) | ( n14793 & n14800 ) | ( ~n14797 & n14800 ) ;
  assign n14802 = n14784 | n14801 ;
  assign n14803 = n14784 & n14801 ;
  assign n14804 = n14802 & ~n14803 ;
  assign n14805 = n14293 | n14299 ;
  assign n14806 = n14804 & n14805 ;
  assign n14807 = n14804 | n14805 ;
  assign n14808 = ~n14806 & n14807 ;
  assign n14809 = x99 & n2429 ;
  assign n14810 = x98 & n2424 ;
  assign n14811 = x97 & ~n2423 ;
  assign n14812 = n2631 & n14811 ;
  assign n14813 = n14810 | n14812 ;
  assign n14814 = n14809 | n14813 ;
  assign n14815 = n2432 | n14809 ;
  assign n14816 = n14813 | n14815 ;
  assign n14817 = ( n6164 & n14814 ) | ( n6164 & n14816 ) | ( n14814 & n14816 ) ;
  assign n14818 = x23 & n14816 ;
  assign n14819 = x23 & n14809 ;
  assign n14820 = ( x23 & n14813 ) | ( x23 & n14819 ) | ( n14813 & n14819 ) ;
  assign n14821 = ( n6164 & n14818 ) | ( n6164 & n14820 ) | ( n14818 & n14820 ) ;
  assign n14822 = x23 & ~n14820 ;
  assign n14823 = x23 & ~n14816 ;
  assign n14824 = ( ~n6164 & n14822 ) | ( ~n6164 & n14823 ) | ( n14822 & n14823 ) ;
  assign n14825 = ( n14817 & ~n14821 ) | ( n14817 & n14824 ) | ( ~n14821 & n14824 ) ;
  assign n14826 = n14808 & n14825 ;
  assign n14827 = n14808 & ~n14826 ;
  assign n14828 = ~n14808 & n14825 ;
  assign n14829 = n14827 | n14828 ;
  assign n14830 = n14326 | n14333 ;
  assign n14831 = n14829 | n14830 ;
  assign n14832 = n14829 & n14830 ;
  assign n14833 = n14831 & ~n14832 ;
  assign n14834 = x102 & n1859 ;
  assign n14835 = x101 & n1854 ;
  assign n14836 = x100 & ~n1853 ;
  assign n14837 = n2037 & n14836 ;
  assign n14838 = n14835 | n14837 ;
  assign n14839 = n14834 | n14838 ;
  assign n14840 = n1862 | n14834 ;
  assign n14841 = n14838 | n14840 ;
  assign n14842 = ( n7178 & n14839 ) | ( n7178 & n14841 ) | ( n14839 & n14841 ) ;
  assign n14843 = x20 & n14841 ;
  assign n14844 = x20 & n14834 ;
  assign n14845 = ( x20 & n14838 ) | ( x20 & n14844 ) | ( n14838 & n14844 ) ;
  assign n14846 = ( n7178 & n14843 ) | ( n7178 & n14845 ) | ( n14843 & n14845 ) ;
  assign n14847 = x20 & ~n14845 ;
  assign n14848 = x20 & ~n14841 ;
  assign n14849 = ( ~n7178 & n14847 ) | ( ~n7178 & n14848 ) | ( n14847 & n14848 ) ;
  assign n14850 = ( n14842 & ~n14846 ) | ( n14842 & n14849 ) | ( ~n14846 & n14849 ) ;
  assign n14851 = n14833 & n14850 ;
  assign n14852 = n14833 & ~n14851 ;
  assign n14853 = ~n14833 & n14850 ;
  assign n14854 = n14852 | n14853 ;
  assign n14855 = n14354 | n14361 ;
  assign n14856 = n14854 | n14855 ;
  assign n14857 = n14854 & n14855 ;
  assign n14858 = n14856 & ~n14857 ;
  assign n14859 = x105 & n1383 ;
  assign n14860 = x104 & n1378 ;
  assign n14861 = x103 & ~n1377 ;
  assign n14862 = n1542 & n14861 ;
  assign n14863 = n14860 | n14862 ;
  assign n14864 = n14859 | n14863 ;
  assign n14865 = n1386 | n14859 ;
  assign n14866 = n14863 | n14865 ;
  assign n14867 = ( n8273 & n14864 ) | ( n8273 & n14866 ) | ( n14864 & n14866 ) ;
  assign n14868 = x17 & n14866 ;
  assign n14869 = x17 & n14859 ;
  assign n14870 = ( x17 & n14863 ) | ( x17 & n14869 ) | ( n14863 & n14869 ) ;
  assign n14871 = ( n8273 & n14868 ) | ( n8273 & n14870 ) | ( n14868 & n14870 ) ;
  assign n14872 = x17 & ~n14870 ;
  assign n14873 = x17 & ~n14866 ;
  assign n14874 = ( ~n8273 & n14872 ) | ( ~n8273 & n14873 ) | ( n14872 & n14873 ) ;
  assign n14875 = ( n14867 & ~n14871 ) | ( n14867 & n14874 ) | ( ~n14871 & n14874 ) ;
  assign n14876 = n14858 & n14875 ;
  assign n14877 = n14858 & ~n14876 ;
  assign n14878 = ~n14858 & n14875 ;
  assign n14879 = n14877 | n14878 ;
  assign n14880 = n14380 | n14382 ;
  assign n14881 = n14381 | n14880 ;
  assign n14882 = ( n14380 & n14384 ) | ( n14380 & n14881 ) | ( n14384 & n14881 ) ;
  assign n14883 = n14879 | n14882 ;
  assign n14884 = n14879 & n14882 ;
  assign n14885 = n14883 & ~n14884 ;
  assign n14886 = x108 & n962 ;
  assign n14887 = x107 & n957 ;
  assign n14888 = x106 & ~n956 ;
  assign n14889 = n1105 & n14888 ;
  assign n14890 = n14887 | n14889 ;
  assign n14891 = n14886 | n14890 ;
  assign n14892 = n965 | n14886 ;
  assign n14893 = n14890 | n14892 ;
  assign n14894 = ( n9479 & n14891 ) | ( n9479 & n14893 ) | ( n14891 & n14893 ) ;
  assign n14895 = x14 & n14893 ;
  assign n14896 = x14 & n14886 ;
  assign n14897 = ( x14 & n14890 ) | ( x14 & n14896 ) | ( n14890 & n14896 ) ;
  assign n14898 = ( n9479 & n14895 ) | ( n9479 & n14897 ) | ( n14895 & n14897 ) ;
  assign n14899 = x14 & ~n14897 ;
  assign n14900 = x14 & ~n14893 ;
  assign n14901 = ( ~n9479 & n14899 ) | ( ~n9479 & n14900 ) | ( n14899 & n14900 ) ;
  assign n14902 = ( n14894 & ~n14898 ) | ( n14894 & n14901 ) | ( ~n14898 & n14901 ) ;
  assign n14903 = n14885 & n14902 ;
  assign n14904 = n14885 | n14902 ;
  assign n14905 = ~n14903 & n14904 ;
  assign n14906 = n14405 | n14409 ;
  assign n14907 = n14405 | n14406 ;
  assign n14908 = ( n13886 & n14906 ) | ( n13886 & n14907 ) | ( n14906 & n14907 ) ;
  assign n14909 = n14905 & n14908 ;
  assign n14910 = ~n14905 & n14908 ;
  assign n14911 = ( n14905 & ~n14909 ) | ( n14905 & n14910 ) | ( ~n14909 & n14910 ) ;
  assign n14912 = x111 & n636 ;
  assign n14913 = x110 & n631 ;
  assign n14914 = x109 & ~n630 ;
  assign n14915 = n764 & n14914 ;
  assign n14916 = n14913 | n14915 ;
  assign n14917 = n14912 | n14916 ;
  assign n14918 = n639 | n14912 ;
  assign n14919 = n14916 | n14918 ;
  assign n14920 = ( n10749 & n14917 ) | ( n10749 & n14919 ) | ( n14917 & n14919 ) ;
  assign n14921 = x11 & n14919 ;
  assign n14922 = x11 & n14912 ;
  assign n14923 = ( x11 & n14916 ) | ( x11 & n14922 ) | ( n14916 & n14922 ) ;
  assign n14924 = ( n10749 & n14921 ) | ( n10749 & n14923 ) | ( n14921 & n14923 ) ;
  assign n14925 = x11 & ~n14923 ;
  assign n14926 = x11 & ~n14919 ;
  assign n14927 = ( ~n10749 & n14925 ) | ( ~n10749 & n14926 ) | ( n14925 & n14926 ) ;
  assign n14928 = ( n14920 & ~n14924 ) | ( n14920 & n14927 ) | ( ~n14924 & n14927 ) ;
  assign n14929 = n14905 & n14928 ;
  assign n14930 = ~n14908 & n14928 ;
  assign n14931 = ( ~n14905 & n14928 ) | ( ~n14905 & n14930 ) | ( n14928 & n14930 ) ;
  assign n14932 = ( n14910 & n14929 ) | ( n14910 & n14931 ) | ( n14929 & n14931 ) ;
  assign n14933 = n14911 & ~n14932 ;
  assign n14934 = ~n14905 & n14928 ;
  assign n14935 = n14908 & n14928 ;
  assign n14936 = n14905 & n14935 ;
  assign n14937 = ( ~n14910 & n14934 ) | ( ~n14910 & n14936 ) | ( n14934 & n14936 ) ;
  assign n14938 = n14933 | n14937 ;
  assign n14939 = n13907 | n13911 ;
  assign n14940 = n14433 | n14437 ;
  assign n14941 = ( n14433 & n14939 ) | ( n14433 & n14940 ) | ( n14939 & n14940 ) ;
  assign n14942 = n14938 & n14941 ;
  assign n14943 = n14938 | n14941 ;
  assign n14944 = ~n14942 & n14943 ;
  assign n14945 = x114 & n389 ;
  assign n14946 = x113 & n384 ;
  assign n14947 = x112 & ~n383 ;
  assign n14948 = n463 & n14947 ;
  assign n14949 = n14946 | n14948 ;
  assign n14950 = n14945 | n14949 ;
  assign n14951 = n392 | n14945 ;
  assign n14952 = n14949 | n14951 ;
  assign n14953 = ( ~n12095 & n14950 ) | ( ~n12095 & n14952 ) | ( n14950 & n14952 ) ;
  assign n14954 = n14950 & n14952 ;
  assign n14955 = ( n12079 & n14953 ) | ( n12079 & n14954 ) | ( n14953 & n14954 ) ;
  assign n14956 = x8 & n14955 ;
  assign n14957 = x8 & ~n14955 ;
  assign n14958 = ( n14955 & ~n14956 ) | ( n14955 & n14957 ) | ( ~n14956 & n14957 ) ;
  assign n14959 = n14944 & n14958 ;
  assign n14960 = n14944 & ~n14959 ;
  assign n14961 = ~n14944 & n14958 ;
  assign n14962 = n14960 | n14961 ;
  assign n14963 = n13932 | n13938 ;
  assign n14964 = n14458 | n14459 ;
  assign n14965 = ( n14458 & n14963 ) | ( n14458 & n14964 ) | ( n14963 & n14964 ) ;
  assign n14966 = ~n14962 & n14965 ;
  assign n14967 = n14533 & n14966 ;
  assign n14968 = n14962 & ~n14965 ;
  assign n14969 = ( n14533 & n14967 ) | ( n14533 & n14968 ) | ( n14967 & n14968 ) ;
  assign n14970 = n14533 | n14966 ;
  assign n14971 = n14968 | n14970 ;
  assign n14972 = ~n14969 & n14971 ;
  assign n14973 = ( n14464 & n14478 ) | ( n14464 & n14483 ) | ( n14478 & n14483 ) ;
  assign n14974 = n14972 | n14973 ;
  assign n14975 = n14972 & n14973 ;
  assign n14976 = n14974 & ~n14975 ;
  assign n14977 = x119 | x120 ;
  assign n14978 = x119 & x120 ;
  assign n14979 = n14977 & ~n14978 ;
  assign n14980 = n14490 | n14491 ;
  assign n14981 = n14979 & n14980 ;
  assign n14982 = n14490 & n14979 ;
  assign n14983 = ( n13965 & n14981 ) | ( n13965 & n14982 ) | ( n14981 & n14982 ) ;
  assign n14984 = n14981 | n14982 ;
  assign n14985 = ( n14002 & n14983 ) | ( n14002 & n14984 ) | ( n14983 & n14984 ) ;
  assign n14986 = n14979 | n14980 ;
  assign n14987 = n13965 | n14490 ;
  assign n14988 = ( n14490 & n14491 ) | ( n14490 & n14987 ) | ( n14491 & n14987 ) ;
  assign n14989 = n14979 | n14988 ;
  assign n14990 = ( n14002 & n14986 ) | ( n14002 & n14989 ) | ( n14986 & n14989 ) ;
  assign n14991 = ~n14985 & n14990 ;
  assign n14992 = x119 & n133 ;
  assign n14993 = x118 & ~n162 ;
  assign n14994 = ( n137 & n14992 ) | ( n137 & n14993 ) | ( n14992 & n14993 ) ;
  assign n14995 = x0 & x120 ;
  assign n14996 = ( ~n137 & n14992 ) | ( ~n137 & n14995 ) | ( n14992 & n14995 ) ;
  assign n14997 = n14994 | n14996 ;
  assign n14998 = n141 | n14997 ;
  assign n14999 = ( n14991 & n14997 ) | ( n14991 & n14998 ) | ( n14997 & n14998 ) ;
  assign n15000 = x2 & n14997 ;
  assign n15001 = ( x2 & n523 ) | ( x2 & n14997 ) | ( n523 & n14997 ) ;
  assign n15002 = ( n14991 & n15000 ) | ( n14991 & n15001 ) | ( n15000 & n15001 ) ;
  assign n15003 = x2 & ~n15001 ;
  assign n15004 = x2 & ~n14997 ;
  assign n15005 = ( ~n14991 & n15003 ) | ( ~n14991 & n15004 ) | ( n15003 & n15004 ) ;
  assign n15006 = ( n14999 & ~n15002 ) | ( n14999 & n15005 ) | ( ~n15002 & n15005 ) ;
  assign n15007 = n14976 & n15006 ;
  assign n15008 = n14976 & ~n15007 ;
  assign n15009 = ~n14976 & n15006 ;
  assign n15010 = n15008 | n15009 ;
  assign n15011 = n14512 | n14516 ;
  assign n15012 = ( n14512 & n14514 ) | ( n14512 & n15011 ) | ( n14514 & n15011 ) ;
  assign n15013 = n15010 & n15012 ;
  assign n15014 = n15010 | n15012 ;
  assign n15015 = ~n15013 & n15014 ;
  assign n15016 = n14969 | n14973 ;
  assign n15017 = ( n14969 & n14972 ) | ( n14969 & n15016 ) | ( n14972 & n15016 ) ;
  assign n15018 = n14668 | n14674 ;
  assign n15019 = x82 & n7566 ;
  assign n15020 = x81 & n7561 ;
  assign n15021 = x80 & ~n7560 ;
  assign n15022 = n7953 & n15021 ;
  assign n15023 = n15020 | n15022 ;
  assign n15024 = n15019 | n15023 ;
  assign n15025 = n7569 | n15019 ;
  assign n15026 = n15023 | n15025 ;
  assign n15027 = ( n1811 & n15024 ) | ( n1811 & n15026 ) | ( n15024 & n15026 ) ;
  assign n15028 = x41 & n15026 ;
  assign n15029 = x41 & n15019 ;
  assign n15030 = ( x41 & n15023 ) | ( x41 & n15029 ) | ( n15023 & n15029 ) ;
  assign n15031 = ( n1811 & n15028 ) | ( n1811 & n15030 ) | ( n15028 & n15030 ) ;
  assign n15032 = x41 & ~n15030 ;
  assign n15033 = x41 & ~n15026 ;
  assign n15034 = ( ~n1811 & n15032 ) | ( ~n1811 & n15033 ) | ( n15032 & n15033 ) ;
  assign n15035 = ( n15027 & ~n15031 ) | ( n15027 & n15034 ) | ( ~n15031 & n15034 ) ;
  assign n15036 = n14583 | n14587 ;
  assign n15037 = x56 & ~x57 ;
  assign n15038 = ~x56 & x57 ;
  assign n15039 = n15037 | n15038 ;
  assign n15040 = x64 & n15039 ;
  assign n15041 = ~n14060 & n15040 ;
  assign n15042 = ( ~n14564 & n15040 ) | ( ~n14564 & n15041 ) | ( n15040 & n15041 ) ;
  assign n15043 = n14060 & ~n15040 ;
  assign n15044 = n14564 & n15043 ;
  assign n15045 = n15042 | n15044 ;
  assign n15046 = x67 & n14045 ;
  assign n15047 = x66 & n14040 ;
  assign n15048 = x65 & ~n14039 ;
  assign n15049 = n14552 & n15048 ;
  assign n15050 = n15047 | n15049 ;
  assign n15051 = n15046 | n15050 ;
  assign n15052 = n186 & n14048 ;
  assign n15053 = n15051 | n15052 ;
  assign n15054 = x56 & ~n15053 ;
  assign n15055 = ~x56 & n15053 ;
  assign n15056 = n15054 | n15055 ;
  assign n15057 = n15045 & n15056 ;
  assign n15058 = n15045 | n15056 ;
  assign n15059 = ~n15057 & n15058 ;
  assign n15060 = x69 & n12569 ;
  assign n15061 = x68 & ~n12568 ;
  assign n15062 = n13076 & n15061 ;
  assign n15063 = n15060 | n15062 ;
  assign n15064 = x70 & n12574 ;
  assign n15065 = n12577 | n15064 ;
  assign n15066 = n15063 | n15065 ;
  assign n15067 = x53 & ~n15066 ;
  assign n15068 = x53 & ~n15064 ;
  assign n15069 = ~n15063 & n15068 ;
  assign n15070 = ( ~n340 & n15067 ) | ( ~n340 & n15069 ) | ( n15067 & n15069 ) ;
  assign n15071 = ~x53 & n15066 ;
  assign n15072 = ~x53 & n15064 ;
  assign n15073 = ( ~x53 & n15063 ) | ( ~x53 & n15072 ) | ( n15063 & n15072 ) ;
  assign n15074 = ( n340 & n15071 ) | ( n340 & n15073 ) | ( n15071 & n15073 ) ;
  assign n15075 = n15070 | n15074 ;
  assign n15076 = ( n14583 & ~n15059 ) | ( n14583 & n15075 ) | ( ~n15059 & n15075 ) ;
  assign n15077 = n15059 & ~n15075 ;
  assign n15078 = ( n14587 & n15076 ) | ( n14587 & ~n15077 ) | ( n15076 & ~n15077 ) ;
  assign n15079 = ( ~n15036 & n15059 ) | ( ~n15036 & n15078 ) | ( n15059 & n15078 ) ;
  assign n15080 = x73 & n11205 ;
  assign n15081 = x72 & n11200 ;
  assign n15082 = x71 & ~n11199 ;
  assign n15083 = n11679 & n15082 ;
  assign n15084 = n15081 | n15083 ;
  assign n15085 = n15080 | n15084 ;
  assign n15086 = ( ~n610 & n11208 ) | ( ~n610 & n15085 ) | ( n11208 & n15085 ) ;
  assign n15087 = n11208 & n15080 ;
  assign n15088 = ( n11208 & n15084 ) | ( n11208 & n15087 ) | ( n15084 & n15087 ) ;
  assign n15089 = ( n598 & n15086 ) | ( n598 & n15088 ) | ( n15086 & n15088 ) ;
  assign n15090 = ( x50 & ~n15085 ) | ( x50 & n15089 ) | ( ~n15085 & n15089 ) ;
  assign n15091 = ~n15089 & n15090 ;
  assign n15092 = x50 | n15080 ;
  assign n15093 = n15084 | n15092 ;
  assign n15094 = n15089 | n15093 ;
  assign n15095 = ( ~x50 & n15091 ) | ( ~x50 & n15094 ) | ( n15091 & n15094 ) ;
  assign n15096 = n15078 & n15095 ;
  assign n15097 = ~n15075 & n15094 ;
  assign n15098 = x50 | n15075 ;
  assign n15099 = ( n15091 & n15097 ) | ( n15091 & ~n15098 ) | ( n15097 & ~n15098 ) ;
  assign n15100 = ( n15079 & n15096 ) | ( n15079 & n15099 ) | ( n15096 & n15099 ) ;
  assign n15101 = n15078 | n15095 ;
  assign n15102 = n15075 & ~n15094 ;
  assign n15103 = x50 & n15075 ;
  assign n15104 = ( ~n15091 & n15102 ) | ( ~n15091 & n15103 ) | ( n15102 & n15103 ) ;
  assign n15105 = ( n15079 & n15101 ) | ( n15079 & ~n15104 ) | ( n15101 & ~n15104 ) ;
  assign n15106 = ~n15100 & n15105 ;
  assign n15107 = n14591 | n14594 ;
  assign n15108 = ( n14591 & n14596 ) | ( n14591 & n15107 ) | ( n14596 & n15107 ) ;
  assign n15109 = n15106 & n15108 ;
  assign n15110 = n15106 | n15108 ;
  assign n15111 = ~n15109 & n15110 ;
  assign n15112 = x76 & n9933 ;
  assign n15113 = x75 & n9928 ;
  assign n15114 = x74 & ~n9927 ;
  assign n15115 = n10379 & n15114 ;
  assign n15116 = n15113 | n15115 ;
  assign n15117 = n15112 | n15116 ;
  assign n15118 = n9936 | n15112 ;
  assign n15119 = n15116 | n15118 ;
  assign n15120 = ( n923 & n15117 ) | ( n923 & n15119 ) | ( n15117 & n15119 ) ;
  assign n15121 = x47 & n15119 ;
  assign n15122 = x47 & n15112 ;
  assign n15123 = ( x47 & n15116 ) | ( x47 & n15122 ) | ( n15116 & n15122 ) ;
  assign n15124 = ( n923 & n15121 ) | ( n923 & n15123 ) | ( n15121 & n15123 ) ;
  assign n15125 = x47 & ~n15123 ;
  assign n15126 = x47 & ~n15119 ;
  assign n15127 = ( ~n923 & n15125 ) | ( ~n923 & n15126 ) | ( n15125 & n15126 ) ;
  assign n15128 = ( n15120 & ~n15124 ) | ( n15120 & n15127 ) | ( ~n15124 & n15127 ) ;
  assign n15129 = n15111 | n15128 ;
  assign n15130 = n15111 & n15128 ;
  assign n15131 = n15129 & ~n15130 ;
  assign n15132 = n14618 | n14619 ;
  assign n15133 = ( n14618 & n14621 ) | ( n14618 & n15132 ) | ( n14621 & n15132 ) ;
  assign n15134 = n15131 & n15133 ;
  assign n15135 = n15131 | n15133 ;
  assign n15136 = ~n15134 & n15135 ;
  assign n15137 = x79 & n8724 ;
  assign n15138 = x78 & n8719 ;
  assign n15139 = x77 & ~n8718 ;
  assign n15140 = n9149 & n15139 ;
  assign n15141 = n15138 | n15140 ;
  assign n15142 = n15137 | n15141 ;
  assign n15143 = n8727 | n15137 ;
  assign n15144 = n15141 | n15143 ;
  assign n15145 = ( n1332 & n15142 ) | ( n1332 & n15144 ) | ( n15142 & n15144 ) ;
  assign n15146 = x44 & n15144 ;
  assign n15147 = x44 & n15137 ;
  assign n15148 = ( x44 & n15141 ) | ( x44 & n15147 ) | ( n15141 & n15147 ) ;
  assign n15149 = ( n1332 & n15146 ) | ( n1332 & n15148 ) | ( n15146 & n15148 ) ;
  assign n15150 = x44 & ~n15148 ;
  assign n15151 = x44 & ~n15144 ;
  assign n15152 = ( ~n1332 & n15150 ) | ( ~n1332 & n15151 ) | ( n15150 & n15151 ) ;
  assign n15153 = ( n15145 & ~n15149 ) | ( n15145 & n15152 ) | ( ~n15149 & n15152 ) ;
  assign n15154 = n15136 & n15153 ;
  assign n15155 = n15136 | n15153 ;
  assign n15156 = ~n15154 & n15155 ;
  assign n15157 = n14642 & n15156 ;
  assign n15158 = ( n14648 & n15156 ) | ( n14648 & n15157 ) | ( n15156 & n15157 ) ;
  assign n15159 = n14642 | n15156 ;
  assign n15160 = n14648 | n15159 ;
  assign n15161 = ~n15158 & n15160 ;
  assign n15162 = n15035 & n15161 ;
  assign n15163 = ( ~n14668 & n15035 ) | ( ~n14668 & n15161 ) | ( n15035 & n15161 ) ;
  assign n15164 = ( ~n14674 & n15162 ) | ( ~n14674 & n15163 ) | ( n15162 & n15163 ) ;
  assign n15165 = ( n15018 & ~n15035 ) | ( n15018 & n15164 ) | ( ~n15035 & n15164 ) ;
  assign n15166 = x85 & n6536 ;
  assign n15167 = x84 & n6531 ;
  assign n15168 = x83 & ~n6530 ;
  assign n15169 = n6871 & n15168 ;
  assign n15170 = n15167 | n15169 ;
  assign n15171 = n15166 | n15170 ;
  assign n15172 = n6539 | n15166 ;
  assign n15173 = n15170 | n15172 ;
  assign n15174 = ( n2381 & n15171 ) | ( n2381 & n15173 ) | ( n15171 & n15173 ) ;
  assign n15175 = x38 & n15173 ;
  assign n15176 = x38 & n15166 ;
  assign n15177 = ( x38 & n15170 ) | ( x38 & n15176 ) | ( n15170 & n15176 ) ;
  assign n15178 = ( n2381 & n15175 ) | ( n2381 & n15177 ) | ( n15175 & n15177 ) ;
  assign n15179 = x38 & ~n15177 ;
  assign n15180 = x38 & ~n15173 ;
  assign n15181 = ( ~n2381 & n15179 ) | ( ~n2381 & n15180 ) | ( n15179 & n15180 ) ;
  assign n15182 = ( n15174 & ~n15178 ) | ( n15174 & n15181 ) | ( ~n15178 & n15181 ) ;
  assign n15183 = ~n15161 & n15182 ;
  assign n15184 = n15163 & n15182 ;
  assign n15185 = n15162 & n15182 ;
  assign n15186 = ( ~n14674 & n15184 ) | ( ~n14674 & n15185 ) | ( n15184 & n15185 ) ;
  assign n15187 = ( n15165 & n15183 ) | ( n15165 & n15186 ) | ( n15183 & n15186 ) ;
  assign n15188 = n15161 & ~n15182 ;
  assign n15189 = n15163 | n15182 ;
  assign n15190 = n15162 | n15182 ;
  assign n15191 = ( ~n14674 & n15189 ) | ( ~n14674 & n15190 ) | ( n15189 & n15190 ) ;
  assign n15192 = ( n15165 & ~n15188 ) | ( n15165 & n15191 ) | ( ~n15188 & n15191 ) ;
  assign n15193 = ~n15187 & n15192 ;
  assign n15194 = ( n14188 & n14677 ) | ( n14188 & n14694 ) | ( n14677 & n14694 ) ;
  assign n15195 = n14677 | n14694 ;
  assign n15196 = ( n14213 & n15194 ) | ( n14213 & n15195 ) | ( n15194 & n15195 ) ;
  assign n15197 = n15193 | n15196 ;
  assign n15198 = n15193 & n15196 ;
  assign n15199 = n15197 & ~n15198 ;
  assign n15200 = x88 & n5554 ;
  assign n15201 = x87 & n5549 ;
  assign n15202 = x86 & ~n5548 ;
  assign n15203 = n5893 & n15202 ;
  assign n15204 = n15201 | n15203 ;
  assign n15205 = n15200 | n15204 ;
  assign n15206 = n5557 | n15200 ;
  assign n15207 = n15204 | n15206 ;
  assign n15208 = ( ~n3039 & n15205 ) | ( ~n3039 & n15207 ) | ( n15205 & n15207 ) ;
  assign n15209 = n15205 & n15207 ;
  assign n15210 = ( n3023 & n15208 ) | ( n3023 & n15209 ) | ( n15208 & n15209 ) ;
  assign n15211 = x35 & n15207 ;
  assign n15212 = x35 & n15200 ;
  assign n15213 = ( x35 & n15204 ) | ( x35 & n15212 ) | ( n15204 & n15212 ) ;
  assign n15214 = ( ~n3039 & n15211 ) | ( ~n3039 & n15213 ) | ( n15211 & n15213 ) ;
  assign n15215 = n15211 & n15213 ;
  assign n15216 = ( n3023 & n15214 ) | ( n3023 & n15215 ) | ( n15214 & n15215 ) ;
  assign n15217 = x35 & ~n15213 ;
  assign n15218 = x35 & ~n15207 ;
  assign n15219 = ( n3039 & n15217 ) | ( n3039 & n15218 ) | ( n15217 & n15218 ) ;
  assign n15220 = n15217 | n15218 ;
  assign n15221 = ( ~n3023 & n15219 ) | ( ~n3023 & n15220 ) | ( n15219 & n15220 ) ;
  assign n15222 = ( n15210 & ~n15216 ) | ( n15210 & n15221 ) | ( ~n15216 & n15221 ) ;
  assign n15223 = n15199 & n15222 ;
  assign n15224 = n15199 & ~n15223 ;
  assign n15225 = ~n15199 & n15222 ;
  assign n15226 = n15224 | n15225 ;
  assign n15227 = n14723 & n15225 ;
  assign n15228 = ( n14723 & n15224 ) | ( n14723 & n15227 ) | ( n15224 & n15227 ) ;
  assign n15229 = ( n14729 & n15226 ) | ( n14729 & n15228 ) | ( n15226 & n15228 ) ;
  assign n15230 = n14723 | n15225 ;
  assign n15231 = n15224 | n15230 ;
  assign n15232 = n14729 | n15231 ;
  assign n15233 = ~n15229 & n15232 ;
  assign n15234 = x91 & n4631 ;
  assign n15235 = x90 & n4626 ;
  assign n15236 = x89 & ~n4625 ;
  assign n15237 = n4943 & n15236 ;
  assign n15238 = n15235 | n15237 ;
  assign n15239 = n15234 | n15238 ;
  assign n15240 = n4634 | n15234 ;
  assign n15241 = n15238 | n15240 ;
  assign n15242 = ( n3768 & n15239 ) | ( n3768 & n15241 ) | ( n15239 & n15241 ) ;
  assign n15243 = x32 & n15241 ;
  assign n15244 = x32 & n15234 ;
  assign n15245 = ( x32 & n15238 ) | ( x32 & n15244 ) | ( n15238 & n15244 ) ;
  assign n15246 = ( n3768 & n15243 ) | ( n3768 & n15245 ) | ( n15243 & n15245 ) ;
  assign n15247 = x32 & ~n15245 ;
  assign n15248 = x32 & ~n15241 ;
  assign n15249 = ( ~n3768 & n15247 ) | ( ~n3768 & n15248 ) | ( n15247 & n15248 ) ;
  assign n15250 = ( n15242 & ~n15246 ) | ( n15242 & n15249 ) | ( ~n15246 & n15249 ) ;
  assign n15251 = n15233 | n15250 ;
  assign n15252 = n15233 & n15250 ;
  assign n15253 = n15251 & ~n15252 ;
  assign n15254 = n14748 & n15253 ;
  assign n15255 = ( n14752 & n15253 ) | ( n14752 & n15254 ) | ( n15253 & n15254 ) ;
  assign n15256 = n14748 | n15253 ;
  assign n15257 = n14752 | n15256 ;
  assign n15258 = ~n15255 & n15257 ;
  assign n15259 = x94 & n3816 ;
  assign n15260 = x93 & n3811 ;
  assign n15261 = x92 & ~n3810 ;
  assign n15262 = n4067 & n15261 ;
  assign n15263 = n15260 | n15262 ;
  assign n15264 = n15259 | n15263 ;
  assign n15265 = n3819 | n15259 ;
  assign n15266 = n15263 | n15265 ;
  assign n15267 = ( n4583 & n15264 ) | ( n4583 & n15266 ) | ( n15264 & n15266 ) ;
  assign n15268 = x29 & n15266 ;
  assign n15269 = x29 & n15259 ;
  assign n15270 = ( x29 & n15263 ) | ( x29 & n15269 ) | ( n15263 & n15269 ) ;
  assign n15271 = ( n4583 & n15268 ) | ( n4583 & n15270 ) | ( n15268 & n15270 ) ;
  assign n15272 = x29 & ~n15270 ;
  assign n15273 = x29 & ~n15266 ;
  assign n15274 = ( ~n4583 & n15272 ) | ( ~n4583 & n15273 ) | ( n15272 & n15273 ) ;
  assign n15275 = ( n15267 & ~n15271 ) | ( n15267 & n15274 ) | ( ~n15271 & n15274 ) ;
  assign n15276 = n15258 & n15275 ;
  assign n15277 = n15258 | n15275 ;
  assign n15278 = ~n15276 & n15277 ;
  assign n15279 = n14776 | n14779 ;
  assign n15280 = ( n14776 & n14781 ) | ( n14776 & n15279 ) | ( n14781 & n15279 ) ;
  assign n15281 = n15278 & n15280 ;
  assign n15282 = n15278 | n15280 ;
  assign n15283 = ~n15281 & n15282 ;
  assign n15284 = x97 & n3085 ;
  assign n15285 = x96 & n3080 ;
  assign n15286 = x95 & ~n3079 ;
  assign n15287 = n3309 & n15286 ;
  assign n15288 = n15285 | n15287 ;
  assign n15289 = n15284 | n15288 ;
  assign n15290 = n3088 | n15284 ;
  assign n15291 = n15288 | n15290 ;
  assign n15292 = ( n5505 & n15289 ) | ( n5505 & n15291 ) | ( n15289 & n15291 ) ;
  assign n15293 = x26 & n15291 ;
  assign n15294 = x26 & n15284 ;
  assign n15295 = ( x26 & n15288 ) | ( x26 & n15294 ) | ( n15288 & n15294 ) ;
  assign n15296 = ( n5505 & n15293 ) | ( n5505 & n15295 ) | ( n15293 & n15295 ) ;
  assign n15297 = x26 & ~n15295 ;
  assign n15298 = x26 & ~n15291 ;
  assign n15299 = ( ~n5505 & n15297 ) | ( ~n5505 & n15298 ) | ( n15297 & n15298 ) ;
  assign n15300 = ( n15292 & ~n15296 ) | ( n15292 & n15299 ) | ( ~n15296 & n15299 ) ;
  assign n15301 = n15283 & n15300 ;
  assign n15302 = n15283 & ~n15301 ;
  assign n15303 = ~n15283 & n15300 ;
  assign n15304 = n15302 | n15303 ;
  assign n15305 = n14803 | n14804 ;
  assign n15306 = ( n14803 & n14805 ) | ( n14803 & n15305 ) | ( n14805 & n15305 ) ;
  assign n15307 = ~n15304 & n15306 ;
  assign n15308 = n15304 & ~n15306 ;
  assign n15309 = n15307 | n15308 ;
  assign n15310 = x100 & n2429 ;
  assign n15311 = x99 & n2424 ;
  assign n15312 = x98 & ~n2423 ;
  assign n15313 = n2631 & n15312 ;
  assign n15314 = n15311 | n15313 ;
  assign n15315 = n15310 | n15314 ;
  assign n15316 = n2432 | n15310 ;
  assign n15317 = n15314 | n15316 ;
  assign n15318 = ( n6483 & n15315 ) | ( n6483 & n15317 ) | ( n15315 & n15317 ) ;
  assign n15319 = x23 & n15317 ;
  assign n15320 = x23 & n15310 ;
  assign n15321 = ( x23 & n15314 ) | ( x23 & n15320 ) | ( n15314 & n15320 ) ;
  assign n15322 = ( n6483 & n15319 ) | ( n6483 & n15321 ) | ( n15319 & n15321 ) ;
  assign n15323 = x23 & ~n15321 ;
  assign n15324 = x23 & ~n15317 ;
  assign n15325 = ( ~n6483 & n15323 ) | ( ~n6483 & n15324 ) | ( n15323 & n15324 ) ;
  assign n15326 = ( n15318 & ~n15322 ) | ( n15318 & n15325 ) | ( ~n15322 & n15325 ) ;
  assign n15327 = n15309 & n15326 ;
  assign n15328 = n15309 | n15326 ;
  assign n15329 = ~n15327 & n15328 ;
  assign n15330 = n14826 | n14830 ;
  assign n15331 = ( n14826 & n14829 ) | ( n14826 & n15330 ) | ( n14829 & n15330 ) ;
  assign n15332 = n15329 | n15331 ;
  assign n15333 = n15329 & n15331 ;
  assign n15334 = n15332 & ~n15333 ;
  assign n15335 = x103 & n1859 ;
  assign n15336 = x102 & n1854 ;
  assign n15337 = x101 & ~n1853 ;
  assign n15338 = n2037 & n15337 ;
  assign n15339 = n15336 | n15338 ;
  assign n15340 = n15335 | n15339 ;
  assign n15341 = n1862 | n15335 ;
  assign n15342 = n15339 | n15341 ;
  assign n15343 = ( n7529 & n15340 ) | ( n7529 & n15342 ) | ( n15340 & n15342 ) ;
  assign n15344 = x20 & n15342 ;
  assign n15345 = x20 & n15335 ;
  assign n15346 = ( x20 & n15339 ) | ( x20 & n15345 ) | ( n15339 & n15345 ) ;
  assign n15347 = ( n7529 & n15344 ) | ( n7529 & n15346 ) | ( n15344 & n15346 ) ;
  assign n15348 = x20 & ~n15346 ;
  assign n15349 = x20 & ~n15342 ;
  assign n15350 = ( ~n7529 & n15348 ) | ( ~n7529 & n15349 ) | ( n15348 & n15349 ) ;
  assign n15351 = ( n15343 & ~n15347 ) | ( n15343 & n15350 ) | ( ~n15347 & n15350 ) ;
  assign n15352 = n15334 & n15351 ;
  assign n15353 = n15334 & ~n15352 ;
  assign n15354 = ~n15334 & n15351 ;
  assign n15355 = n15353 | n15354 ;
  assign n15356 = n14851 | n14855 ;
  assign n15357 = ( n14851 & n14854 ) | ( n14851 & n15356 ) | ( n14854 & n15356 ) ;
  assign n15358 = n15355 | n15357 ;
  assign n15359 = n15355 & n15357 ;
  assign n15360 = n15358 & ~n15359 ;
  assign n15361 = x106 & n1383 ;
  assign n15362 = x105 & n1378 ;
  assign n15363 = x104 & ~n1377 ;
  assign n15364 = n1542 & n15363 ;
  assign n15365 = n15362 | n15364 ;
  assign n15366 = n15361 | n15365 ;
  assign n15367 = n1386 | n15361 ;
  assign n15368 = n15365 | n15367 ;
  assign n15369 = ( n8656 & n15366 ) | ( n8656 & n15368 ) | ( n15366 & n15368 ) ;
  assign n15370 = x17 & n15368 ;
  assign n15371 = x17 & n15361 ;
  assign n15372 = ( x17 & n15365 ) | ( x17 & n15371 ) | ( n15365 & n15371 ) ;
  assign n15373 = ( n8656 & n15370 ) | ( n8656 & n15372 ) | ( n15370 & n15372 ) ;
  assign n15374 = x17 & ~n15372 ;
  assign n15375 = x17 & ~n15368 ;
  assign n15376 = ( ~n8656 & n15374 ) | ( ~n8656 & n15375 ) | ( n15374 & n15375 ) ;
  assign n15377 = ( n15369 & ~n15373 ) | ( n15369 & n15376 ) | ( ~n15373 & n15376 ) ;
  assign n15378 = n15360 | n15377 ;
  assign n15379 = n15360 & n15377 ;
  assign n15380 = n15378 & ~n15379 ;
  assign n15381 = n14876 | n14882 ;
  assign n15382 = ( n14876 & n14879 ) | ( n14876 & n15381 ) | ( n14879 & n15381 ) ;
  assign n15383 = n15380 & n15382 ;
  assign n15384 = n15380 | n15382 ;
  assign n15385 = ~n15383 & n15384 ;
  assign n15386 = x109 & n962 ;
  assign n15387 = x108 & n957 ;
  assign n15388 = x107 & ~n956 ;
  assign n15389 = n1105 & n15388 ;
  assign n15390 = n15387 | n15389 ;
  assign n15391 = n15386 | n15390 ;
  assign n15392 = n965 | n15386 ;
  assign n15393 = n15390 | n15392 ;
  assign n15394 = ( n9878 & n15391 ) | ( n9878 & n15393 ) | ( n15391 & n15393 ) ;
  assign n15395 = x14 & n15393 ;
  assign n15396 = x14 & n15386 ;
  assign n15397 = ( x14 & n15390 ) | ( x14 & n15396 ) | ( n15390 & n15396 ) ;
  assign n15398 = ( n9878 & n15395 ) | ( n9878 & n15397 ) | ( n15395 & n15397 ) ;
  assign n15399 = x14 & ~n15397 ;
  assign n15400 = x14 & ~n15393 ;
  assign n15401 = ( ~n9878 & n15399 ) | ( ~n9878 & n15400 ) | ( n15399 & n15400 ) ;
  assign n15402 = ( n15394 & ~n15398 ) | ( n15394 & n15401 ) | ( ~n15398 & n15401 ) ;
  assign n15403 = n15385 & n15402 ;
  assign n15404 = n15385 & ~n15403 ;
  assign n15405 = ~n15385 & n15402 ;
  assign n15406 = n15404 | n15405 ;
  assign n15407 = n14903 | n14908 ;
  assign n15408 = ( n14903 & n14905 ) | ( n14903 & n15407 ) | ( n14905 & n15407 ) ;
  assign n15409 = n15406 & n15408 ;
  assign n15410 = n15406 | n15408 ;
  assign n15411 = ~n15409 & n15410 ;
  assign n15412 = x112 & n636 ;
  assign n15413 = x111 & n631 ;
  assign n15414 = x110 & ~n630 ;
  assign n15415 = n764 & n15414 ;
  assign n15416 = n15413 | n15415 ;
  assign n15417 = n15412 | n15416 ;
  assign n15418 = n639 | n15412 ;
  assign n15419 = n15416 | n15418 ;
  assign n15420 = ( n11172 & n15417 ) | ( n11172 & n15419 ) | ( n15417 & n15419 ) ;
  assign n15421 = x11 & n15419 ;
  assign n15422 = x11 & n15412 ;
  assign n15423 = ( x11 & n15416 ) | ( x11 & n15422 ) | ( n15416 & n15422 ) ;
  assign n15424 = ( n11172 & n15421 ) | ( n11172 & n15423 ) | ( n15421 & n15423 ) ;
  assign n15425 = x11 & ~n15423 ;
  assign n15426 = x11 & ~n15419 ;
  assign n15427 = ( ~n11172 & n15425 ) | ( ~n11172 & n15426 ) | ( n15425 & n15426 ) ;
  assign n15428 = ( n15420 & ~n15424 ) | ( n15420 & n15427 ) | ( ~n15424 & n15427 ) ;
  assign n15429 = n15411 & n15428 ;
  assign n15430 = n15411 & ~n15429 ;
  assign n15431 = ~n15411 & n15428 ;
  assign n15432 = n15430 | n15431 ;
  assign n15433 = n14932 | n14938 ;
  assign n15434 = ( n14932 & n14941 ) | ( n14932 & n15433 ) | ( n14941 & n15433 ) ;
  assign n15435 = n15432 & n15434 ;
  assign n15436 = n15432 | n15434 ;
  assign n15437 = ~n15435 & n15436 ;
  assign n15438 = x115 & n389 ;
  assign n15439 = x114 & n384 ;
  assign n15440 = x113 & ~n383 ;
  assign n15441 = n463 & n15440 ;
  assign n15442 = n15439 | n15441 ;
  assign n15443 = n15438 | n15442 ;
  assign n15444 = n392 | n15438 ;
  assign n15445 = n15442 | n15444 ;
  assign n15446 = ( ~n12550 & n15443 ) | ( ~n12550 & n15445 ) | ( n15443 & n15445 ) ;
  assign n15447 = n15443 & n15445 ;
  assign n15448 = ( n12532 & n15446 ) | ( n12532 & n15447 ) | ( n15446 & n15447 ) ;
  assign n15449 = x8 & n15448 ;
  assign n15450 = x8 & ~n15448 ;
  assign n15451 = ( n15448 & ~n15449 ) | ( n15448 & n15450 ) | ( ~n15449 & n15450 ) ;
  assign n15452 = n15437 & n15451 ;
  assign n15453 = n15437 & ~n15452 ;
  assign n15454 = ~n15437 & n15451 ;
  assign n15455 = n15453 | n15454 ;
  assign n15456 = n14962 & n14965 ;
  assign n15457 = n14959 | n15456 ;
  assign n15458 = n15455 & n15457 ;
  assign n15459 = n15455 | n15457 ;
  assign n15460 = ~n15458 & n15459 ;
  assign n15461 = x118 & n212 ;
  assign n15462 = x117 & n207 ;
  assign n15463 = x116 & ~n206 ;
  assign n15464 = n267 & n15463 ;
  assign n15465 = n15462 | n15464 ;
  assign n15466 = n15461 | n15465 ;
  assign n15467 = n215 | n15461 ;
  assign n15468 = n15465 | n15467 ;
  assign n15469 = ( ~n14002 & n15466 ) | ( ~n14002 & n15468 ) | ( n15466 & n15468 ) ;
  assign n15470 = n15466 & n15468 ;
  assign n15471 = ( n13981 & n15469 ) | ( n13981 & n15470 ) | ( n15469 & n15470 ) ;
  assign n15472 = x5 & n15471 ;
  assign n15473 = x5 & ~n15471 ;
  assign n15474 = ( n15471 & ~n15472 ) | ( n15471 & n15473 ) | ( ~n15472 & n15473 ) ;
  assign n15475 = n15460 & n15474 ;
  assign n15476 = n15460 & ~n15475 ;
  assign n15477 = ~n15460 & n15474 ;
  assign n15478 = n15017 & n15477 ;
  assign n15479 = ( n15017 & n15476 ) | ( n15017 & n15478 ) | ( n15476 & n15478 ) ;
  assign n15480 = n15017 & ~n15479 ;
  assign n15481 = n15476 | n15477 ;
  assign n15482 = ~n15479 & n15481 ;
  assign n15483 = n15480 | n15482 ;
  assign n15484 = x120 | x121 ;
  assign n15485 = x120 & x121 ;
  assign n15486 = n15484 & ~n15485 ;
  assign n15487 = n14978 | n14979 ;
  assign n15488 = ( n14978 & n14980 ) | ( n14978 & n15487 ) | ( n14980 & n15487 ) ;
  assign n15489 = n15486 & n15488 ;
  assign n15490 = n14490 | n14978 ;
  assign n15491 = ( n14978 & n14979 ) | ( n14978 & n15490 ) | ( n14979 & n15490 ) ;
  assign n15492 = n15486 & n15491 ;
  assign n15493 = ( n13965 & n15489 ) | ( n13965 & n15492 ) | ( n15489 & n15492 ) ;
  assign n15494 = n15489 | n15492 ;
  assign n15495 = ( n14002 & n15493 ) | ( n14002 & n15494 ) | ( n15493 & n15494 ) ;
  assign n15496 = n15486 | n15491 ;
  assign n15497 = n15488 | n15496 ;
  assign n15498 = n13965 | n15486 ;
  assign n15499 = ( n15488 & n15496 ) | ( n15488 & n15498 ) | ( n15496 & n15498 ) ;
  assign n15500 = ( n14002 & n15497 ) | ( n14002 & n15499 ) | ( n15497 & n15499 ) ;
  assign n15501 = ~n15495 & n15500 ;
  assign n15502 = x120 & n133 ;
  assign n15503 = x119 & ~n162 ;
  assign n15504 = ( n137 & n15502 ) | ( n137 & n15503 ) | ( n15502 & n15503 ) ;
  assign n15505 = x0 & x121 ;
  assign n15506 = ( ~n137 & n15502 ) | ( ~n137 & n15505 ) | ( n15502 & n15505 ) ;
  assign n15507 = n15504 | n15506 ;
  assign n15508 = n141 | n15507 ;
  assign n15509 = ( n15501 & n15507 ) | ( n15501 & n15508 ) | ( n15507 & n15508 ) ;
  assign n15510 = x2 & n15507 ;
  assign n15511 = ( x2 & n523 ) | ( x2 & n15507 ) | ( n523 & n15507 ) ;
  assign n15512 = ( n15501 & n15510 ) | ( n15501 & n15511 ) | ( n15510 & n15511 ) ;
  assign n15513 = x2 & ~n15511 ;
  assign n15514 = x2 & ~n15507 ;
  assign n15515 = ( ~n15501 & n15513 ) | ( ~n15501 & n15514 ) | ( n15513 & n15514 ) ;
  assign n15516 = ( n15509 & ~n15512 ) | ( n15509 & n15515 ) | ( ~n15512 & n15515 ) ;
  assign n15517 = n15483 & n15516 ;
  assign n15518 = n15483 & ~n15517 ;
  assign n15519 = ~n15483 & n15516 ;
  assign n15520 = n15518 | n15519 ;
  assign n15521 = n15007 | n15012 ;
  assign n15522 = ( n15007 & n15010 ) | ( n15007 & n15521 ) | ( n15010 & n15521 ) ;
  assign n15523 = n15520 | n15522 ;
  assign n15524 = n15519 & n15522 ;
  assign n15525 = ( n15518 & n15522 ) | ( n15518 & n15524 ) | ( n15522 & n15524 ) ;
  assign n15526 = n15523 & ~n15525 ;
  assign n15527 = n15475 | n15479 ;
  assign n15925 = n15379 | n15380 ;
  assign n15926 = ( n15379 & n15382 ) | ( n15379 & n15925 ) | ( n15382 & n15925 ) ;
  assign n15528 = x70 & n12569 ;
  assign n15529 = x69 & ~n12568 ;
  assign n15530 = n13076 & n15529 ;
  assign n15531 = n15528 | n15530 ;
  assign n15532 = x71 & n12574 ;
  assign n15533 = n12577 | n15532 ;
  assign n15534 = n15531 | n15533 ;
  assign n15535 = x53 & ~n15534 ;
  assign n15536 = x53 & ~n15532 ;
  assign n15537 = ~n15531 & n15536 ;
  assign n15538 = ( ~n438 & n15535 ) | ( ~n438 & n15537 ) | ( n15535 & n15537 ) ;
  assign n15539 = ~x53 & n15534 ;
  assign n15540 = ~x53 & n15532 ;
  assign n15541 = ( ~x53 & n15531 ) | ( ~x53 & n15540 ) | ( n15531 & n15540 ) ;
  assign n15542 = ( n438 & n15539 ) | ( n438 & n15541 ) | ( n15539 & n15541 ) ;
  assign n15543 = n15538 | n15542 ;
  assign n15544 = ~x57 & x58 ;
  assign n15545 = x57 & ~x58 ;
  assign n15546 = n15544 | n15545 ;
  assign n15547 = ~n15039 & n15546 ;
  assign n15548 = x64 & n15547 ;
  assign n15549 = ~x58 & x59 ;
  assign n15550 = x58 & ~x59 ;
  assign n15551 = n15549 | n15550 ;
  assign n15552 = n15039 & ~n15551 ;
  assign n15553 = x65 & n15552 ;
  assign n15554 = n15548 | n15553 ;
  assign n15555 = n15039 & n15551 ;
  assign n15556 = x59 | n144 ;
  assign n15557 = ( x59 & n15555 ) | ( x59 & n15556 ) | ( n15555 & n15556 ) ;
  assign n15558 = ~x59 & n15557 ;
  assign n15559 = ( ~x59 & n15554 ) | ( ~x59 & n15558 ) | ( n15554 & n15558 ) ;
  assign n15560 = x59 & ~x64 ;
  assign n15561 = ( x59 & ~n15039 ) | ( x59 & n15560 ) | ( ~n15039 & n15560 ) ;
  assign n15562 = n15557 & n15561 ;
  assign n15563 = ( n15554 & n15561 ) | ( n15554 & n15562 ) | ( n15561 & n15562 ) ;
  assign n15564 = n144 & n15555 ;
  assign n15565 = n15561 & ~n15564 ;
  assign n15566 = ~n15554 & n15565 ;
  assign n15567 = ( n15559 & n15563 ) | ( n15559 & n15566 ) | ( n15563 & n15566 ) ;
  assign n15568 = n15557 | n15561 ;
  assign n15569 = n15554 | n15568 ;
  assign n15570 = ~n15561 & n15564 ;
  assign n15571 = ( n15554 & ~n15561 ) | ( n15554 & n15570 ) | ( ~n15561 & n15570 ) ;
  assign n15572 = ( n15559 & n15569 ) | ( n15559 & ~n15571 ) | ( n15569 & ~n15571 ) ;
  assign n15573 = ~n15567 & n15572 ;
  assign n15574 = n241 & n14048 ;
  assign n15575 = x68 & n14045 ;
  assign n15576 = x67 & n14040 ;
  assign n15577 = x66 & ~n14039 ;
  assign n15578 = n14552 & n15577 ;
  assign n15579 = n15576 | n15578 ;
  assign n15580 = n15575 | n15579 ;
  assign n15581 = n15574 | n15580 ;
  assign n15582 = x56 | n15575 ;
  assign n15583 = n15579 | n15582 ;
  assign n15584 = n15574 | n15583 ;
  assign n15585 = ~x56 & n15583 ;
  assign n15586 = ( ~x56 & n15574 ) | ( ~x56 & n15585 ) | ( n15574 & n15585 ) ;
  assign n15587 = ( ~n15581 & n15584 ) | ( ~n15581 & n15586 ) | ( n15584 & n15586 ) ;
  assign n15588 = n15573 | n15587 ;
  assign n15589 = n15573 & n15587 ;
  assign n15590 = n15588 & ~n15589 ;
  assign n15591 = ( n14566 & n15040 ) | ( n14566 & n15056 ) | ( n15040 & n15056 ) ;
  assign n15592 = n15590 | n15591 ;
  assign n15593 = n15590 & n15591 ;
  assign n15594 = n15592 & ~n15593 ;
  assign n15595 = n15543 | n15594 ;
  assign n15596 = n15543 & n15594 ;
  assign n15597 = n15595 & ~n15596 ;
  assign n15598 = ~n15059 & n15075 ;
  assign n15599 = n15036 & ~n15598 ;
  assign n15600 = n15059 & n15075 ;
  assign n15601 = n15059 & ~n15600 ;
  assign n15602 = ( n15036 & n15600 ) | ( n15036 & n15601 ) | ( n15600 & n15601 ) ;
  assign n15603 = n15036 | n15600 ;
  assign n15604 = ( ~n15599 & n15602 ) | ( ~n15599 & n15603 ) | ( n15602 & n15603 ) ;
  assign n15605 = n15597 & n15604 ;
  assign n15606 = n15597 | n15604 ;
  assign n15607 = ~n15605 & n15606 ;
  assign n15608 = x74 & n11205 ;
  assign n15609 = x73 & n11200 ;
  assign n15610 = x72 & ~n11199 ;
  assign n15611 = n11679 & n15610 ;
  assign n15612 = n15609 | n15611 ;
  assign n15613 = n15608 | n15612 ;
  assign n15614 = n11208 | n15608 ;
  assign n15615 = n15612 | n15614 ;
  assign n15616 = ( n710 & n15613 ) | ( n710 & n15615 ) | ( n15613 & n15615 ) ;
  assign n15617 = x50 & n15615 ;
  assign n15618 = x50 & n15608 ;
  assign n15619 = ( x50 & n15612 ) | ( x50 & n15618 ) | ( n15612 & n15618 ) ;
  assign n15620 = ( n710 & n15617 ) | ( n710 & n15619 ) | ( n15617 & n15619 ) ;
  assign n15621 = x50 & ~n15619 ;
  assign n15622 = x50 & ~n15615 ;
  assign n15623 = ( ~n710 & n15621 ) | ( ~n710 & n15622 ) | ( n15621 & n15622 ) ;
  assign n15624 = ( n15616 & ~n15620 ) | ( n15616 & n15623 ) | ( ~n15620 & n15623 ) ;
  assign n15625 = n15607 & n15624 ;
  assign n15626 = n15607 & ~n15625 ;
  assign n15627 = n15100 | n15106 ;
  assign n15628 = ( n15100 & n15108 ) | ( n15100 & n15627 ) | ( n15108 & n15627 ) ;
  assign n15629 = ~n15607 & n15624 ;
  assign n15630 = n15628 & n15629 ;
  assign n15631 = ( n15626 & n15628 ) | ( n15626 & n15630 ) | ( n15628 & n15630 ) ;
  assign n15632 = n15628 | n15629 ;
  assign n15633 = n15626 | n15632 ;
  assign n15634 = ~n15631 & n15633 ;
  assign n15635 = x77 & n9933 ;
  assign n15636 = x76 & n9928 ;
  assign n15637 = x75 & ~n9927 ;
  assign n15638 = n10379 & n15637 ;
  assign n15639 = n15636 | n15638 ;
  assign n15640 = n15635 | n15639 ;
  assign n15641 = n9936 | n15635 ;
  assign n15642 = n15639 | n15641 ;
  assign n15643 = ( n1059 & n15640 ) | ( n1059 & n15642 ) | ( n15640 & n15642 ) ;
  assign n15644 = x47 & n15642 ;
  assign n15645 = x47 & n15635 ;
  assign n15646 = ( x47 & n15639 ) | ( x47 & n15645 ) | ( n15639 & n15645 ) ;
  assign n15647 = ( n1059 & n15644 ) | ( n1059 & n15646 ) | ( n15644 & n15646 ) ;
  assign n15648 = x47 & ~n15646 ;
  assign n15649 = x47 & ~n15642 ;
  assign n15650 = ( ~n1059 & n15648 ) | ( ~n1059 & n15649 ) | ( n15648 & n15649 ) ;
  assign n15651 = ( n15643 & ~n15647 ) | ( n15643 & n15650 ) | ( ~n15647 & n15650 ) ;
  assign n15652 = n15634 & n15651 ;
  assign n15653 = n15634 | n15651 ;
  assign n15654 = ~n15652 & n15653 ;
  assign n15655 = n15130 | n15131 ;
  assign n15656 = ( n15130 & n15133 ) | ( n15130 & n15655 ) | ( n15133 & n15655 ) ;
  assign n15657 = n15654 & n15656 ;
  assign n15658 = n15656 & ~n15657 ;
  assign n15659 = ( n15654 & ~n15657 ) | ( n15654 & n15658 ) | ( ~n15657 & n15658 ) ;
  assign n15660 = x80 & n8724 ;
  assign n15661 = x79 & n8719 ;
  assign n15662 = x78 & ~n8718 ;
  assign n15663 = n9149 & n15662 ;
  assign n15664 = n15661 | n15663 ;
  assign n15665 = n15660 | n15664 ;
  assign n15666 = n8727 | n15660 ;
  assign n15667 = n15664 | n15666 ;
  assign n15668 = ( n1499 & n15665 ) | ( n1499 & n15667 ) | ( n15665 & n15667 ) ;
  assign n15669 = x44 & n15667 ;
  assign n15670 = x44 & n15660 ;
  assign n15671 = ( x44 & n15664 ) | ( x44 & n15670 ) | ( n15664 & n15670 ) ;
  assign n15672 = ( n1499 & n15669 ) | ( n1499 & n15671 ) | ( n15669 & n15671 ) ;
  assign n15673 = x44 & ~n15671 ;
  assign n15674 = x44 & ~n15667 ;
  assign n15675 = ( ~n1499 & n15673 ) | ( ~n1499 & n15674 ) | ( n15673 & n15674 ) ;
  assign n15676 = ( n15668 & ~n15672 ) | ( n15668 & n15675 ) | ( ~n15672 & n15675 ) ;
  assign n15677 = ~n15657 & n15676 ;
  assign n15678 = n15654 & n15676 ;
  assign n15679 = ( n15658 & n15677 ) | ( n15658 & n15678 ) | ( n15677 & n15678 ) ;
  assign n15680 = n15659 & ~n15679 ;
  assign n15681 = n15657 & n15676 ;
  assign n15682 = ~n15654 & n15676 ;
  assign n15683 = ( ~n15658 & n15681 ) | ( ~n15658 & n15682 ) | ( n15681 & n15682 ) ;
  assign n15684 = n15680 | n15683 ;
  assign n15685 = n15154 | n15158 ;
  assign n15686 = n15684 | n15685 ;
  assign n15687 = n15684 & n15685 ;
  assign n15688 = n15686 & ~n15687 ;
  assign n15689 = x83 & n7566 ;
  assign n15690 = x82 & n7561 ;
  assign n15691 = x81 & ~n7560 ;
  assign n15692 = n7953 & n15691 ;
  assign n15693 = n15690 | n15692 ;
  assign n15694 = n15689 | n15693 ;
  assign n15695 = n7569 | n15689 ;
  assign n15696 = n15693 | n15695 ;
  assign n15697 = ( n2009 & n15694 ) | ( n2009 & n15696 ) | ( n15694 & n15696 ) ;
  assign n15698 = x41 & n15696 ;
  assign n15699 = x41 & n15689 ;
  assign n15700 = ( x41 & n15693 ) | ( x41 & n15699 ) | ( n15693 & n15699 ) ;
  assign n15701 = ( n2009 & n15698 ) | ( n2009 & n15700 ) | ( n15698 & n15700 ) ;
  assign n15702 = x41 & ~n15700 ;
  assign n15703 = x41 & ~n15696 ;
  assign n15704 = ( ~n2009 & n15702 ) | ( ~n2009 & n15703 ) | ( n15702 & n15703 ) ;
  assign n15705 = ( n15697 & ~n15701 ) | ( n15697 & n15704 ) | ( ~n15701 & n15704 ) ;
  assign n15706 = n15688 & n15705 ;
  assign n15707 = n15688 | n15705 ;
  assign n15708 = ~n15706 & n15707 ;
  assign n15709 = n15161 & ~n15162 ;
  assign n15710 = n15035 & ~n15161 ;
  assign n15711 = n15162 | n15710 ;
  assign n15712 = n15709 | n15711 ;
  assign n15713 = ( n15018 & n15162 ) | ( n15018 & n15712 ) | ( n15162 & n15712 ) ;
  assign n15714 = n15708 & n15713 ;
  assign n15715 = n15713 & ~n15714 ;
  assign n15716 = ( n15708 & ~n15714 ) | ( n15708 & n15715 ) | ( ~n15714 & n15715 ) ;
  assign n15717 = x86 & n6536 ;
  assign n15718 = x85 & n6531 ;
  assign n15719 = x84 & ~n6530 ;
  assign n15720 = n6871 & n15719 ;
  assign n15721 = n15718 | n15720 ;
  assign n15722 = n15717 | n15721 ;
  assign n15723 = n6539 | n15717 ;
  assign n15724 = n15721 | n15723 ;
  assign n15725 = ( n2606 & n15722 ) | ( n2606 & n15724 ) | ( n15722 & n15724 ) ;
  assign n15726 = x38 & n15724 ;
  assign n15727 = x38 & n15717 ;
  assign n15728 = ( x38 & n15721 ) | ( x38 & n15727 ) | ( n15721 & n15727 ) ;
  assign n15729 = ( n2606 & n15726 ) | ( n2606 & n15728 ) | ( n15726 & n15728 ) ;
  assign n15730 = x38 & ~n15728 ;
  assign n15731 = x38 & ~n15724 ;
  assign n15732 = ( ~n2606 & n15730 ) | ( ~n2606 & n15731 ) | ( n15730 & n15731 ) ;
  assign n15733 = ( n15725 & ~n15729 ) | ( n15725 & n15732 ) | ( ~n15729 & n15732 ) ;
  assign n15734 = n15708 & n15733 ;
  assign n15735 = ~n15708 & n15733 ;
  assign n15736 = ( ~n15713 & n15733 ) | ( ~n15713 & n15735 ) | ( n15733 & n15735 ) ;
  assign n15737 = ( n15715 & n15734 ) | ( n15715 & n15736 ) | ( n15734 & n15736 ) ;
  assign n15738 = n15716 & ~n15737 ;
  assign n15739 = n15713 & n15734 ;
  assign n15740 = ( ~n15715 & n15735 ) | ( ~n15715 & n15739 ) | ( n15735 & n15739 ) ;
  assign n15741 = n15738 | n15740 ;
  assign n15742 = n15187 | n15198 ;
  assign n15743 = n15741 | n15742 ;
  assign n15744 = n15741 & n15742 ;
  assign n15745 = n15743 & ~n15744 ;
  assign n15746 = x89 & n5554 ;
  assign n15747 = x88 & n5549 ;
  assign n15748 = x87 & ~n5548 ;
  assign n15749 = n5893 & n15748 ;
  assign n15750 = n15747 | n15749 ;
  assign n15751 = n15746 | n15750 ;
  assign n15752 = n5557 | n15746 ;
  assign n15753 = n15750 | n15752 ;
  assign n15754 = ( n3282 & n15751 ) | ( n3282 & n15753 ) | ( n15751 & n15753 ) ;
  assign n15755 = x35 & n15753 ;
  assign n15756 = x35 & n15746 ;
  assign n15757 = ( x35 & n15750 ) | ( x35 & n15756 ) | ( n15750 & n15756 ) ;
  assign n15758 = ( n3282 & n15755 ) | ( n3282 & n15757 ) | ( n15755 & n15757 ) ;
  assign n15759 = x35 & ~n15757 ;
  assign n15760 = x35 & ~n15753 ;
  assign n15761 = ( ~n3282 & n15759 ) | ( ~n3282 & n15760 ) | ( n15759 & n15760 ) ;
  assign n15762 = ( n15754 & ~n15758 ) | ( n15754 & n15761 ) | ( ~n15758 & n15761 ) ;
  assign n15763 = n15745 & n15762 ;
  assign n15764 = n15745 & ~n15763 ;
  assign n15765 = ~n15745 & n15762 ;
  assign n15766 = n15764 | n15765 ;
  assign n15767 = n15223 | n15229 ;
  assign n15768 = n15766 | n15767 ;
  assign n15769 = n15766 & n15767 ;
  assign n15770 = n15768 & ~n15769 ;
  assign n15771 = x92 & n4631 ;
  assign n15772 = x91 & n4626 ;
  assign n15773 = x90 & ~n4625 ;
  assign n15774 = n4943 & n15773 ;
  assign n15775 = n15772 | n15774 ;
  assign n15776 = n15771 | n15775 ;
  assign n15777 = n4634 | n15771 ;
  assign n15778 = n15775 | n15777 ;
  assign n15779 = ( n4040 & n15776 ) | ( n4040 & n15778 ) | ( n15776 & n15778 ) ;
  assign n15780 = x32 & n15778 ;
  assign n15781 = x32 & n15771 ;
  assign n15782 = ( x32 & n15775 ) | ( x32 & n15781 ) | ( n15775 & n15781 ) ;
  assign n15783 = ( n4040 & n15780 ) | ( n4040 & n15782 ) | ( n15780 & n15782 ) ;
  assign n15784 = x32 & ~n15782 ;
  assign n15785 = x32 & ~n15778 ;
  assign n15786 = ( ~n4040 & n15784 ) | ( ~n4040 & n15785 ) | ( n15784 & n15785 ) ;
  assign n15787 = ( n15779 & ~n15783 ) | ( n15779 & n15786 ) | ( ~n15783 & n15786 ) ;
  assign n15788 = n15770 & n15787 ;
  assign n15789 = n15770 & ~n15788 ;
  assign n15790 = ~n15770 & n15787 ;
  assign n15791 = n15789 | n15790 ;
  assign n15792 = n15252 | n15254 ;
  assign n15793 = n15252 | n15253 ;
  assign n15794 = ( n14752 & n15792 ) | ( n14752 & n15793 ) | ( n15792 & n15793 ) ;
  assign n15795 = ~n15791 & n15794 ;
  assign n15796 = n15791 & ~n15794 ;
  assign n15797 = n15795 | n15796 ;
  assign n15798 = x95 & n3816 ;
  assign n15799 = x94 & n3811 ;
  assign n15800 = x93 & ~n3810 ;
  assign n15801 = n4067 & n15800 ;
  assign n15802 = n15799 | n15801 ;
  assign n15803 = n15798 | n15802 ;
  assign n15804 = n3819 | n15798 ;
  assign n15805 = n15802 | n15804 ;
  assign n15806 = ( n4897 & n15803 ) | ( n4897 & n15805 ) | ( n15803 & n15805 ) ;
  assign n15807 = x29 & n15805 ;
  assign n15808 = x29 & n15798 ;
  assign n15809 = ( x29 & n15802 ) | ( x29 & n15808 ) | ( n15802 & n15808 ) ;
  assign n15810 = ( n4897 & n15807 ) | ( n4897 & n15809 ) | ( n15807 & n15809 ) ;
  assign n15811 = x29 & ~n15809 ;
  assign n15812 = x29 & ~n15805 ;
  assign n15813 = ( ~n4897 & n15811 ) | ( ~n4897 & n15812 ) | ( n15811 & n15812 ) ;
  assign n15814 = ( n15806 & ~n15810 ) | ( n15806 & n15813 ) | ( ~n15810 & n15813 ) ;
  assign n15815 = n15797 & n15814 ;
  assign n15816 = n15797 | n15814 ;
  assign n15817 = ~n15815 & n15816 ;
  assign n15818 = n15276 | n15278 ;
  assign n15819 = ( n15276 & n15280 ) | ( n15276 & n15818 ) | ( n15280 & n15818 ) ;
  assign n15820 = n15817 | n15819 ;
  assign n15821 = n15817 & n15819 ;
  assign n15822 = n15820 & ~n15821 ;
  assign n15823 = x98 & n3085 ;
  assign n15824 = x97 & n3080 ;
  assign n15825 = x96 & ~n3079 ;
  assign n15826 = n3309 & n15825 ;
  assign n15827 = n15824 | n15826 ;
  assign n15828 = n15823 | n15827 ;
  assign n15829 = n3088 | n15823 ;
  assign n15830 = n15827 | n15829 ;
  assign n15831 = ( ~n5850 & n15828 ) | ( ~n5850 & n15830 ) | ( n15828 & n15830 ) ;
  assign n15832 = n15828 & n15830 ;
  assign n15833 = ( n5834 & n15831 ) | ( n5834 & n15832 ) | ( n15831 & n15832 ) ;
  assign n15834 = x26 & n15830 ;
  assign n15835 = x26 & n15823 ;
  assign n15836 = ( x26 & n15827 ) | ( x26 & n15835 ) | ( n15827 & n15835 ) ;
  assign n15837 = ( ~n5850 & n15834 ) | ( ~n5850 & n15836 ) | ( n15834 & n15836 ) ;
  assign n15838 = n15834 & n15836 ;
  assign n15839 = ( n5834 & n15837 ) | ( n5834 & n15838 ) | ( n15837 & n15838 ) ;
  assign n15840 = x26 & ~n15836 ;
  assign n15841 = x26 & ~n15830 ;
  assign n15842 = ( n5850 & n15840 ) | ( n5850 & n15841 ) | ( n15840 & n15841 ) ;
  assign n15843 = n15840 | n15841 ;
  assign n15844 = ( ~n5834 & n15842 ) | ( ~n5834 & n15843 ) | ( n15842 & n15843 ) ;
  assign n15845 = ( n15833 & ~n15839 ) | ( n15833 & n15844 ) | ( ~n15839 & n15844 ) ;
  assign n15846 = n15822 & n15845 ;
  assign n15847 = n15822 & ~n15846 ;
  assign n15848 = ~n15822 & n15845 ;
  assign n15849 = n15847 | n15848 ;
  assign n15850 = ( n15283 & n15300 ) | ( n15283 & n15306 ) | ( n15300 & n15306 ) ;
  assign n15851 = n15849 | n15850 ;
  assign n15852 = n15849 & n15850 ;
  assign n15853 = n15851 & ~n15852 ;
  assign n15854 = x101 & n2429 ;
  assign n15855 = x100 & n2424 ;
  assign n15856 = x99 & ~n2423 ;
  assign n15857 = n2631 & n15856 ;
  assign n15858 = n15855 | n15857 ;
  assign n15859 = n15854 | n15858 ;
  assign n15860 = n2432 | n15854 ;
  assign n15861 = n15858 | n15860 ;
  assign n15862 = ( n6844 & n15859 ) | ( n6844 & n15861 ) | ( n15859 & n15861 ) ;
  assign n15863 = x23 & n15861 ;
  assign n15864 = x23 & n15854 ;
  assign n15865 = ( x23 & n15858 ) | ( x23 & n15864 ) | ( n15858 & n15864 ) ;
  assign n15866 = ( n6844 & n15863 ) | ( n6844 & n15865 ) | ( n15863 & n15865 ) ;
  assign n15867 = x23 & ~n15865 ;
  assign n15868 = x23 & ~n15861 ;
  assign n15869 = ( ~n6844 & n15867 ) | ( ~n6844 & n15868 ) | ( n15867 & n15868 ) ;
  assign n15870 = ( n15862 & ~n15866 ) | ( n15862 & n15869 ) | ( ~n15866 & n15869 ) ;
  assign n15871 = n15853 & n15870 ;
  assign n15872 = n15853 & ~n15871 ;
  assign n15873 = ~n15853 & n15870 ;
  assign n15874 = n15872 | n15873 ;
  assign n15875 = n15327 | n15329 ;
  assign n15876 = ( n15327 & n15331 ) | ( n15327 & n15875 ) | ( n15331 & n15875 ) ;
  assign n15877 = n15874 | n15876 ;
  assign n15878 = n15874 & n15876 ;
  assign n15879 = n15877 & ~n15878 ;
  assign n15880 = x104 & n1859 ;
  assign n15881 = x103 & n1854 ;
  assign n15882 = x102 & ~n1853 ;
  assign n15883 = n2037 & n15882 ;
  assign n15884 = n15881 | n15883 ;
  assign n15885 = n15880 | n15884 ;
  assign n15886 = n1862 | n15880 ;
  assign n15887 = n15884 | n15886 ;
  assign n15888 = ( n7911 & n15885 ) | ( n7911 & n15887 ) | ( n15885 & n15887 ) ;
  assign n15889 = x20 & n15887 ;
  assign n15890 = x20 & n15880 ;
  assign n15891 = ( x20 & n15884 ) | ( x20 & n15890 ) | ( n15884 & n15890 ) ;
  assign n15892 = ( n7911 & n15889 ) | ( n7911 & n15891 ) | ( n15889 & n15891 ) ;
  assign n15893 = x20 & ~n15891 ;
  assign n15894 = x20 & ~n15887 ;
  assign n15895 = ( ~n7911 & n15893 ) | ( ~n7911 & n15894 ) | ( n15893 & n15894 ) ;
  assign n15896 = ( n15888 & ~n15892 ) | ( n15888 & n15895 ) | ( ~n15892 & n15895 ) ;
  assign n15897 = n15879 & n15896 ;
  assign n15898 = n15879 & ~n15897 ;
  assign n15899 = ~n15879 & n15896 ;
  assign n15900 = n15898 | n15899 ;
  assign n15901 = n15352 | n15359 ;
  assign n15902 = n15900 | n15901 ;
  assign n15903 = n15900 & n15901 ;
  assign n15904 = n15902 & ~n15903 ;
  assign n15905 = x107 & n1383 ;
  assign n15906 = x106 & n1378 ;
  assign n15907 = x105 & ~n1377 ;
  assign n15908 = n1542 & n15907 ;
  assign n15909 = n15906 | n15908 ;
  assign n15910 = n15905 | n15909 ;
  assign n15911 = n1386 | n15905 ;
  assign n15912 = n15909 | n15911 ;
  assign n15913 = ( n9084 & n15910 ) | ( n9084 & n15912 ) | ( n15910 & n15912 ) ;
  assign n15914 = x17 & n15912 ;
  assign n15915 = x17 & n15905 ;
  assign n15916 = ( x17 & n15909 ) | ( x17 & n15915 ) | ( n15909 & n15915 ) ;
  assign n15917 = ( n9084 & n15914 ) | ( n9084 & n15916 ) | ( n15914 & n15916 ) ;
  assign n15918 = x17 & ~n15916 ;
  assign n15919 = x17 & ~n15912 ;
  assign n15920 = ( ~n9084 & n15918 ) | ( ~n9084 & n15919 ) | ( n15918 & n15919 ) ;
  assign n15921 = ( n15913 & ~n15917 ) | ( n15913 & n15920 ) | ( ~n15917 & n15920 ) ;
  assign n15922 = n15904 & n15921 ;
  assign n15923 = n15904 | n15921 ;
  assign n15924 = ~n15922 & n15923 ;
  assign n15927 = n15924 & n15926 ;
  assign n15928 = n15926 & ~n15927 ;
  assign n15929 = x110 & n962 ;
  assign n15930 = x109 & n957 ;
  assign n15931 = x108 & ~n956 ;
  assign n15932 = n1105 & n15931 ;
  assign n15933 = n15930 | n15932 ;
  assign n15934 = n15929 | n15933 ;
  assign n15935 = n965 | n15929 ;
  assign n15936 = n15933 | n15935 ;
  assign n15937 = ( n10330 & n15934 ) | ( n10330 & n15936 ) | ( n15934 & n15936 ) ;
  assign n15938 = x14 & n15936 ;
  assign n15939 = x14 & n15929 ;
  assign n15940 = ( x14 & n15933 ) | ( x14 & n15939 ) | ( n15933 & n15939 ) ;
  assign n15941 = ( n10330 & n15938 ) | ( n10330 & n15940 ) | ( n15938 & n15940 ) ;
  assign n15942 = x14 & ~n15940 ;
  assign n15943 = x14 & ~n15936 ;
  assign n15944 = ( ~n10330 & n15942 ) | ( ~n10330 & n15943 ) | ( n15942 & n15943 ) ;
  assign n15945 = ( n15937 & ~n15941 ) | ( n15937 & n15944 ) | ( ~n15941 & n15944 ) ;
  assign n15946 = ~n15927 & n15945 ;
  assign n15947 = n15924 & n15945 ;
  assign n15948 = ( n15928 & n15946 ) | ( n15928 & n15947 ) | ( n15946 & n15947 ) ;
  assign n15949 = n15927 & ~n15945 ;
  assign n15950 = n15924 | n15945 ;
  assign n15951 = ( n15928 & ~n15949 ) | ( n15928 & n15950 ) | ( ~n15949 & n15950 ) ;
  assign n15952 = ~n15948 & n15951 ;
  assign n15953 = n15403 & n15952 ;
  assign n15954 = ( n15409 & n15952 ) | ( n15409 & n15953 ) | ( n15952 & n15953 ) ;
  assign n15955 = n15403 | n15952 ;
  assign n15956 = n15409 | n15955 ;
  assign n15957 = ~n15954 & n15956 ;
  assign n15958 = x113 & n636 ;
  assign n15959 = x112 & n631 ;
  assign n15960 = x111 & ~n630 ;
  assign n15961 = n764 & n15960 ;
  assign n15962 = n15959 | n15961 ;
  assign n15963 = n15958 | n15962 ;
  assign n15964 = n639 | n15958 ;
  assign n15965 = n15962 | n15964 ;
  assign n15966 = ( ~n11642 & n15963 ) | ( ~n11642 & n15965 ) | ( n15963 & n15965 ) ;
  assign n15967 = n15963 & n15965 ;
  assign n15968 = ( n11626 & n15966 ) | ( n11626 & n15967 ) | ( n15966 & n15967 ) ;
  assign n15969 = x11 & n15968 ;
  assign n15970 = x11 & ~n15968 ;
  assign n15971 = ( n15968 & ~n15969 ) | ( n15968 & n15970 ) | ( ~n15969 & n15970 ) ;
  assign n15972 = n15957 | n15971 ;
  assign n15973 = n15957 & n15971 ;
  assign n15974 = n15972 & ~n15973 ;
  assign n15975 = n15429 & n15974 ;
  assign n15976 = ( n15435 & n15974 ) | ( n15435 & n15975 ) | ( n15974 & n15975 ) ;
  assign n15977 = n15429 | n15974 ;
  assign n15978 = n15435 | n15977 ;
  assign n15979 = ~n15976 & n15978 ;
  assign n15980 = x116 & n389 ;
  assign n15981 = x115 & n384 ;
  assign n15982 = x114 & ~n383 ;
  assign n15983 = n463 & n15982 ;
  assign n15984 = n15981 | n15983 ;
  assign n15985 = n15980 | n15984 ;
  assign n15986 = n392 | n15980 ;
  assign n15987 = n15984 | n15986 ;
  assign n15988 = ( ~n13040 & n15985 ) | ( ~n13040 & n15987 ) | ( n15985 & n15987 ) ;
  assign n15989 = n15985 & n15987 ;
  assign n15990 = ( n13022 & n15988 ) | ( n13022 & n15989 ) | ( n15988 & n15989 ) ;
  assign n15991 = x8 & n15990 ;
  assign n15992 = x8 & ~n15990 ;
  assign n15993 = ( n15990 & ~n15991 ) | ( n15990 & n15992 ) | ( ~n15991 & n15992 ) ;
  assign n15994 = n15979 | n15993 ;
  assign n15995 = n15979 & n15993 ;
  assign n15996 = n15994 & ~n15995 ;
  assign n15997 = n15452 & n15996 ;
  assign n15998 = ( n15458 & n15996 ) | ( n15458 & n15997 ) | ( n15996 & n15997 ) ;
  assign n15999 = n15452 | n15996 ;
  assign n16000 = n15458 | n15999 ;
  assign n16001 = ~n15998 & n16000 ;
  assign n16002 = x119 & n212 ;
  assign n16003 = x118 & n207 ;
  assign n16004 = x117 & ~n206 ;
  assign n16005 = n267 & n16004 ;
  assign n16006 = n16003 | n16005 ;
  assign n16007 = n16002 | n16006 ;
  assign n16008 = n215 | n16002 ;
  assign n16009 = n16006 | n16008 ;
  assign n16010 = ( n14496 & n16007 ) | ( n14496 & n16009 ) | ( n16007 & n16009 ) ;
  assign n16011 = x5 & n16009 ;
  assign n16012 = x5 & n16002 ;
  assign n16013 = ( x5 & n16006 ) | ( x5 & n16012 ) | ( n16006 & n16012 ) ;
  assign n16014 = ( n14496 & n16011 ) | ( n14496 & n16013 ) | ( n16011 & n16013 ) ;
  assign n16015 = x5 & ~n16013 ;
  assign n16016 = x5 & ~n16009 ;
  assign n16017 = ( ~n14496 & n16015 ) | ( ~n14496 & n16016 ) | ( n16015 & n16016 ) ;
  assign n16018 = ( n16010 & ~n16014 ) | ( n16010 & n16017 ) | ( ~n16014 & n16017 ) ;
  assign n16019 = n16001 | n16018 ;
  assign n16020 = n16001 & n16018 ;
  assign n16021 = n16019 & ~n16020 ;
  assign n16022 = n15527 & n16021 ;
  assign n16023 = n15527 | n16021 ;
  assign n16024 = ~n16022 & n16023 ;
  assign n16025 = x121 | x122 ;
  assign n16026 = x121 & x122 ;
  assign n16027 = n16025 & ~n16026 ;
  assign n16028 = n15485 | n15486 ;
  assign n16029 = ( n15485 & n15491 ) | ( n15485 & n16028 ) | ( n15491 & n16028 ) ;
  assign n16030 = n16027 & n16029 ;
  assign n16031 = n16027 & n16028 ;
  assign n16032 = n15485 & n16027 ;
  assign n16033 = ( n15488 & n16031 ) | ( n15488 & n16032 ) | ( n16031 & n16032 ) ;
  assign n16034 = ( n13965 & n16030 ) | ( n13965 & n16033 ) | ( n16030 & n16033 ) ;
  assign n16035 = n16030 | n16033 ;
  assign n16036 = ( n14002 & n16034 ) | ( n14002 & n16035 ) | ( n16034 & n16035 ) ;
  assign n16037 = ( n15485 & n15488 ) | ( n15485 & n16028 ) | ( n15488 & n16028 ) ;
  assign n16038 = n16027 | n16029 ;
  assign n16039 = n16037 | n16038 ;
  assign n16040 = n13965 | n16027 ;
  assign n16041 = ( n16037 & n16038 ) | ( n16037 & n16040 ) | ( n16038 & n16040 ) ;
  assign n16042 = ( n14002 & n16039 ) | ( n14002 & n16041 ) | ( n16039 & n16041 ) ;
  assign n16043 = ~n16036 & n16042 ;
  assign n16044 = x121 & n133 ;
  assign n16045 = x120 & ~n162 ;
  assign n16046 = ( n137 & n16044 ) | ( n137 & n16045 ) | ( n16044 & n16045 ) ;
  assign n16047 = x0 & x122 ;
  assign n16048 = ( ~n137 & n16044 ) | ( ~n137 & n16047 ) | ( n16044 & n16047 ) ;
  assign n16049 = n16046 | n16048 ;
  assign n16050 = n141 | n16049 ;
  assign n16051 = ( n16043 & n16049 ) | ( n16043 & n16050 ) | ( n16049 & n16050 ) ;
  assign n16052 = x2 & n16049 ;
  assign n16053 = ( x2 & n523 ) | ( x2 & n16049 ) | ( n523 & n16049 ) ;
  assign n16054 = ( n16043 & n16052 ) | ( n16043 & n16053 ) | ( n16052 & n16053 ) ;
  assign n16055 = x2 & ~n16053 ;
  assign n16056 = x2 & ~n16049 ;
  assign n16057 = ( ~n16043 & n16055 ) | ( ~n16043 & n16056 ) | ( n16055 & n16056 ) ;
  assign n16058 = ( n16051 & ~n16054 ) | ( n16051 & n16057 ) | ( ~n16054 & n16057 ) ;
  assign n16059 = n16024 & n16058 ;
  assign n16060 = n16024 & ~n16059 ;
  assign n16061 = ~n16024 & n16058 ;
  assign n16062 = n16060 | n16061 ;
  assign n16063 = n15517 | n15525 ;
  assign n16064 = n16062 & n16063 ;
  assign n16065 = n16062 | n16063 ;
  assign n16066 = ~n16064 & n16065 ;
  assign n16067 = n16059 | n16064 ;
  assign n16068 = x122 | x123 ;
  assign n16069 = x122 & x123 ;
  assign n16070 = n16068 & ~n16069 ;
  assign n16071 = n16026 & n16070 ;
  assign n16072 = ( n16033 & n16070 ) | ( n16033 & n16071 ) | ( n16070 & n16071 ) ;
  assign n16073 = n16026 | n16027 ;
  assign n16074 = n16070 & n16073 ;
  assign n16075 = ( n16029 & n16071 ) | ( n16029 & n16074 ) | ( n16071 & n16074 ) ;
  assign n16076 = ( n13965 & n16072 ) | ( n13965 & n16075 ) | ( n16072 & n16075 ) ;
  assign n16077 = n16072 | n16075 ;
  assign n16078 = ( n14002 & n16076 ) | ( n14002 & n16077 ) | ( n16076 & n16077 ) ;
  assign n16079 = n16026 | n16033 ;
  assign n16080 = ( n16026 & n16029 ) | ( n16026 & n16073 ) | ( n16029 & n16073 ) ;
  assign n16081 = n16070 | n16080 ;
  assign n16082 = n16079 | n16081 ;
  assign n16083 = n13965 | n16070 ;
  assign n16084 = ( n16079 & n16081 ) | ( n16079 & n16083 ) | ( n16081 & n16083 ) ;
  assign n16085 = ( n14002 & n16082 ) | ( n14002 & n16084 ) | ( n16082 & n16084 ) ;
  assign n16086 = ~n16078 & n16085 ;
  assign n16087 = x122 & n133 ;
  assign n16088 = x121 & ~n162 ;
  assign n16089 = ( n137 & n16087 ) | ( n137 & n16088 ) | ( n16087 & n16088 ) ;
  assign n16090 = x0 & x123 ;
  assign n16091 = ( ~n137 & n16087 ) | ( ~n137 & n16090 ) | ( n16087 & n16090 ) ;
  assign n16092 = n16089 | n16091 ;
  assign n16093 = n141 | n16092 ;
  assign n16094 = ( n16086 & n16092 ) | ( n16086 & n16093 ) | ( n16092 & n16093 ) ;
  assign n16095 = x2 & n16092 ;
  assign n16096 = ( x2 & n523 ) | ( x2 & n16092 ) | ( n523 & n16092 ) ;
  assign n16097 = ( n16086 & n16095 ) | ( n16086 & n16096 ) | ( n16095 & n16096 ) ;
  assign n16098 = x2 & ~n16096 ;
  assign n16099 = x2 & ~n16092 ;
  assign n16100 = ( ~n16086 & n16098 ) | ( ~n16086 & n16099 ) | ( n16098 & n16099 ) ;
  assign n16101 = ( n16094 & ~n16097 ) | ( n16094 & n16100 ) | ( ~n16097 & n16100 ) ;
  assign n16102 = n15995 | n15998 ;
  assign n16103 = n15922 | n15927 ;
  assign n16104 = n15652 | n15657 ;
  assign n16105 = x72 & n12574 ;
  assign n16106 = x71 & n12569 ;
  assign n16107 = x70 & ~n12568 ;
  assign n16108 = n13076 & n16107 ;
  assign n16109 = n16106 | n16108 ;
  assign n16110 = n16105 | n16109 ;
  assign n16111 = ( n513 & n12577 ) | ( n513 & n16110 ) | ( n12577 & n16110 ) ;
  assign n16112 = x53 & n12577 ;
  assign n16113 = ( x53 & n12577 ) | ( x53 & ~n16105 ) | ( n12577 & ~n16105 ) ;
  assign n16114 = ( ~n16109 & n16112 ) | ( ~n16109 & n16113 ) | ( n16112 & n16113 ) ;
  assign n16115 = ( x53 & n513 ) | ( x53 & n16114 ) | ( n513 & n16114 ) ;
  assign n16116 = ~n16111 & n16115 ;
  assign n16117 = n16110 | n16114 ;
  assign n16118 = x53 | n16110 ;
  assign n16119 = ( n513 & n16117 ) | ( n513 & n16118 ) | ( n16117 & n16118 ) ;
  assign n16120 = ( ~x53 & n16116 ) | ( ~x53 & n16119 ) | ( n16116 & n16119 ) ;
  assign n16121 = x66 & n15552 ;
  assign n16122 = x65 & n15547 ;
  assign n16123 = ~n15039 & n15551 ;
  assign n16124 = x64 & ~n15546 ;
  assign n16125 = n16123 & n16124 ;
  assign n16126 = n16122 | n16125 ;
  assign n16127 = n16121 | n16126 ;
  assign n16128 = n159 & n15555 ;
  assign n16129 = n16127 | n16128 ;
  assign n16130 = x59 | n15555 ;
  assign n16131 = ( x59 & n159 ) | ( x59 & n16130 ) | ( n159 & n16130 ) ;
  assign n16132 = n16127 | n16131 ;
  assign n16133 = ~x59 & n16131 ;
  assign n16134 = ( ~x59 & n16127 ) | ( ~x59 & n16133 ) | ( n16127 & n16133 ) ;
  assign n16135 = ( ~n16129 & n16132 ) | ( ~n16129 & n16134 ) | ( n16132 & n16134 ) ;
  assign n16136 = n15567 | n16135 ;
  assign n16137 = n15567 & n16135 ;
  assign n16138 = n16136 & ~n16137 ;
  assign n16139 = n293 & n14048 ;
  assign n16140 = x69 & n14045 ;
  assign n16141 = x68 & n14040 ;
  assign n16142 = x67 & ~n14039 ;
  assign n16143 = n14552 & n16142 ;
  assign n16144 = n16141 | n16143 ;
  assign n16145 = n16140 | n16144 ;
  assign n16146 = n16139 | n16145 ;
  assign n16147 = x56 | n16140 ;
  assign n16148 = n16144 | n16147 ;
  assign n16149 = n16139 | n16148 ;
  assign n16150 = ~x56 & n16148 ;
  assign n16151 = ( ~x56 & n16139 ) | ( ~x56 & n16150 ) | ( n16139 & n16150 ) ;
  assign n16152 = ( ~n16146 & n16149 ) | ( ~n16146 & n16151 ) | ( n16149 & n16151 ) ;
  assign n16153 = n16138 | n16152 ;
  assign n16154 = n16138 & n16152 ;
  assign n16155 = n16153 & ~n16154 ;
  assign n16156 = n15589 | n15591 ;
  assign n16157 = ( n15589 & n15590 ) | ( n15589 & n16156 ) | ( n15590 & n16156 ) ;
  assign n16158 = n16155 & n16157 ;
  assign n16159 = n16155 & ~n16158 ;
  assign n16160 = ~n16155 & n16157 ;
  assign n16161 = n16120 & n16160 ;
  assign n16162 = ( n16120 & n16159 ) | ( n16120 & n16161 ) | ( n16159 & n16161 ) ;
  assign n16163 = n16120 | n16160 ;
  assign n16164 = n16159 | n16163 ;
  assign n16165 = ~n16162 & n16164 ;
  assign n16166 = n15596 | n15597 ;
  assign n16167 = ( n15596 & n15604 ) | ( n15596 & n16166 ) | ( n15604 & n16166 ) ;
  assign n16168 = n16165 & n16167 ;
  assign n16169 = n16165 | n16167 ;
  assign n16170 = ~n16168 & n16169 ;
  assign n16171 = x75 & n11205 ;
  assign n16172 = x74 & n11200 ;
  assign n16173 = x73 & ~n11199 ;
  assign n16174 = n11679 & n16173 ;
  assign n16175 = n16172 | n16174 ;
  assign n16176 = n16171 | n16175 ;
  assign n16177 = n11208 | n16171 ;
  assign n16178 = n16175 | n16177 ;
  assign n16179 = ( n746 & n16176 ) | ( n746 & n16178 ) | ( n16176 & n16178 ) ;
  assign n16180 = x50 & n16178 ;
  assign n16181 = x50 & n16171 ;
  assign n16182 = ( x50 & n16175 ) | ( x50 & n16181 ) | ( n16175 & n16181 ) ;
  assign n16183 = ( n746 & n16180 ) | ( n746 & n16182 ) | ( n16180 & n16182 ) ;
  assign n16184 = x50 & ~n16182 ;
  assign n16185 = x50 & ~n16178 ;
  assign n16186 = ( ~n746 & n16184 ) | ( ~n746 & n16185 ) | ( n16184 & n16185 ) ;
  assign n16187 = ( n16179 & ~n16183 ) | ( n16179 & n16186 ) | ( ~n16183 & n16186 ) ;
  assign n16188 = n16170 | n16187 ;
  assign n16189 = n16170 & n16187 ;
  assign n16190 = n16188 & ~n16189 ;
  assign n16191 = n15625 | n15631 ;
  assign n16192 = n16190 & n16191 ;
  assign n16193 = n16190 | n16191 ;
  assign n16194 = ~n16192 & n16193 ;
  assign n16195 = x78 & n9933 ;
  assign n16196 = x77 & n9928 ;
  assign n16197 = x76 & ~n9927 ;
  assign n16198 = n10379 & n16197 ;
  assign n16199 = n16196 | n16198 ;
  assign n16200 = n16195 | n16199 ;
  assign n16201 = n9936 | n16195 ;
  assign n16202 = n16199 | n16201 ;
  assign n16203 = ( n1192 & n16200 ) | ( n1192 & n16202 ) | ( n16200 & n16202 ) ;
  assign n16204 = x47 & n16202 ;
  assign n16205 = x47 & n16195 ;
  assign n16206 = ( x47 & n16199 ) | ( x47 & n16205 ) | ( n16199 & n16205 ) ;
  assign n16207 = ( n1192 & n16204 ) | ( n1192 & n16206 ) | ( n16204 & n16206 ) ;
  assign n16208 = x47 & ~n16206 ;
  assign n16209 = x47 & ~n16202 ;
  assign n16210 = ( ~n1192 & n16208 ) | ( ~n1192 & n16209 ) | ( n16208 & n16209 ) ;
  assign n16211 = ( n16203 & ~n16207 ) | ( n16203 & n16210 ) | ( ~n16207 & n16210 ) ;
  assign n16212 = n16194 & n16211 ;
  assign n16213 = n16194 & ~n16212 ;
  assign n16214 = ~n16194 & n16211 ;
  assign n16215 = n16213 | n16214 ;
  assign n16216 = n16104 & n16215 ;
  assign n16217 = n16104 | n16215 ;
  assign n16218 = ~n16216 & n16217 ;
  assign n16219 = x81 & n8724 ;
  assign n16220 = x80 & n8719 ;
  assign n16221 = x79 & ~n8718 ;
  assign n16222 = n9149 & n16221 ;
  assign n16223 = n16220 | n16222 ;
  assign n16224 = n16219 | n16223 ;
  assign n16225 = n8727 | n16219 ;
  assign n16226 = n16223 | n16225 ;
  assign n16227 = ( n1651 & n16224 ) | ( n1651 & n16226 ) | ( n16224 & n16226 ) ;
  assign n16228 = x44 & n16226 ;
  assign n16229 = x44 & n16219 ;
  assign n16230 = ( x44 & n16223 ) | ( x44 & n16229 ) | ( n16223 & n16229 ) ;
  assign n16231 = ( n1651 & n16228 ) | ( n1651 & n16230 ) | ( n16228 & n16230 ) ;
  assign n16232 = x44 & ~n16230 ;
  assign n16233 = x44 & ~n16226 ;
  assign n16234 = ( ~n1651 & n16232 ) | ( ~n1651 & n16233 ) | ( n16232 & n16233 ) ;
  assign n16235 = ( n16227 & ~n16231 ) | ( n16227 & n16234 ) | ( ~n16231 & n16234 ) ;
  assign n16236 = n16218 & n16235 ;
  assign n16237 = n16218 & ~n16236 ;
  assign n16238 = ~n16218 & n16235 ;
  assign n16239 = n16237 | n16238 ;
  assign n16240 = n15679 | n15683 ;
  assign n16241 = n15680 | n16240 ;
  assign n16242 = ( n15679 & n15685 ) | ( n15679 & n16241 ) | ( n15685 & n16241 ) ;
  assign n16243 = n16239 & n16242 ;
  assign n16244 = n16239 & ~n16243 ;
  assign n16245 = ~n16239 & n16242 ;
  assign n16246 = n16244 | n16245 ;
  assign n16247 = x84 & n7566 ;
  assign n16248 = x83 & n7561 ;
  assign n16249 = x82 & ~n7560 ;
  assign n16250 = n7953 & n16249 ;
  assign n16251 = n16248 | n16250 ;
  assign n16252 = n16247 | n16251 ;
  assign n16253 = n7569 | n16247 ;
  assign n16254 = n16251 | n16253 ;
  assign n16255 = ( n2194 & n16252 ) | ( n2194 & n16254 ) | ( n16252 & n16254 ) ;
  assign n16256 = x41 & n16254 ;
  assign n16257 = x41 & n16247 ;
  assign n16258 = ( x41 & n16251 ) | ( x41 & n16257 ) | ( n16251 & n16257 ) ;
  assign n16259 = ( n2194 & n16256 ) | ( n2194 & n16258 ) | ( n16256 & n16258 ) ;
  assign n16260 = x41 & ~n16258 ;
  assign n16261 = x41 & ~n16254 ;
  assign n16262 = ( ~n2194 & n16260 ) | ( ~n2194 & n16261 ) | ( n16260 & n16261 ) ;
  assign n16263 = ( n16255 & ~n16259 ) | ( n16255 & n16262 ) | ( ~n16259 & n16262 ) ;
  assign n16264 = n16242 & n16263 ;
  assign n16265 = ~n16239 & n16264 ;
  assign n16266 = ( n16244 & n16263 ) | ( n16244 & n16265 ) | ( n16263 & n16265 ) ;
  assign n16267 = n16246 & ~n16266 ;
  assign n16268 = ~n16242 & n16263 ;
  assign n16269 = ( n16239 & n16263 ) | ( n16239 & n16268 ) | ( n16263 & n16268 ) ;
  assign n16270 = ~n16244 & n16269 ;
  assign n16271 = n16267 | n16270 ;
  assign n16272 = n15706 | n15708 ;
  assign n16273 = ( n15706 & n15713 ) | ( n15706 & n16272 ) | ( n15713 & n16272 ) ;
  assign n16274 = ~n16271 & n16273 ;
  assign n16275 = n16271 & ~n16273 ;
  assign n16276 = n16274 | n16275 ;
  assign n16277 = x87 & n6536 ;
  assign n16278 = x86 & n6531 ;
  assign n16279 = x85 & ~n6530 ;
  assign n16280 = n6871 & n16279 ;
  assign n16281 = n16278 | n16280 ;
  assign n16282 = n16277 | n16281 ;
  assign n16283 = n6539 | n16277 ;
  assign n16284 = n16281 | n16283 ;
  assign n16285 = ( n2816 & n16282 ) | ( n2816 & n16284 ) | ( n16282 & n16284 ) ;
  assign n16286 = x38 & n16284 ;
  assign n16287 = x38 & n16277 ;
  assign n16288 = ( x38 & n16281 ) | ( x38 & n16287 ) | ( n16281 & n16287 ) ;
  assign n16289 = ( n2816 & n16286 ) | ( n2816 & n16288 ) | ( n16286 & n16288 ) ;
  assign n16290 = x38 & ~n16288 ;
  assign n16291 = x38 & ~n16284 ;
  assign n16292 = ( ~n2816 & n16290 ) | ( ~n2816 & n16291 ) | ( n16290 & n16291 ) ;
  assign n16293 = ( n16285 & ~n16289 ) | ( n16285 & n16292 ) | ( ~n16289 & n16292 ) ;
  assign n16294 = n16276 & n16293 ;
  assign n16295 = n16276 | n16293 ;
  assign n16296 = ~n16294 & n16295 ;
  assign n16297 = n15737 | n15742 ;
  assign n16298 = ( n15737 & n15741 ) | ( n15737 & n16297 ) | ( n15741 & n16297 ) ;
  assign n16299 = n16296 | n16298 ;
  assign n16300 = n16296 & n16298 ;
  assign n16301 = n16299 & ~n16300 ;
  assign n16302 = x90 & n5554 ;
  assign n16303 = x89 & n5549 ;
  assign n16304 = x88 & ~n5548 ;
  assign n16305 = n5893 & n16304 ;
  assign n16306 = n16303 | n16305 ;
  assign n16307 = n16302 | n16306 ;
  assign n16308 = n5557 | n16302 ;
  assign n16309 = n16306 | n16308 ;
  assign n16310 = ( n3519 & n16307 ) | ( n3519 & n16309 ) | ( n16307 & n16309 ) ;
  assign n16311 = x35 & n16309 ;
  assign n16312 = x35 & n16302 ;
  assign n16313 = ( x35 & n16306 ) | ( x35 & n16312 ) | ( n16306 & n16312 ) ;
  assign n16314 = ( n3519 & n16311 ) | ( n3519 & n16313 ) | ( n16311 & n16313 ) ;
  assign n16315 = x35 & ~n16313 ;
  assign n16316 = x35 & ~n16309 ;
  assign n16317 = ( ~n3519 & n16315 ) | ( ~n3519 & n16316 ) | ( n16315 & n16316 ) ;
  assign n16318 = ( n16310 & ~n16314 ) | ( n16310 & n16317 ) | ( ~n16314 & n16317 ) ;
  assign n16319 = n16301 & n16318 ;
  assign n16320 = n16301 & ~n16319 ;
  assign n16321 = ~n16301 & n16318 ;
  assign n16322 = n16320 | n16321 ;
  assign n16323 = n15763 | n15767 ;
  assign n16324 = ( n15763 & n15766 ) | ( n15763 & n16323 ) | ( n15766 & n16323 ) ;
  assign n16325 = n16322 | n16324 ;
  assign n16326 = n16322 & n16324 ;
  assign n16327 = n16325 & ~n16326 ;
  assign n16328 = x93 & n4631 ;
  assign n16329 = x92 & n4626 ;
  assign n16330 = x91 & ~n4625 ;
  assign n16331 = n4943 & n16330 ;
  assign n16332 = n16329 | n16331 ;
  assign n16333 = n16328 | n16332 ;
  assign n16334 = n4634 | n16328 ;
  assign n16335 = n16332 | n16334 ;
  assign n16336 = ( n4305 & n16333 ) | ( n4305 & n16335 ) | ( n16333 & n16335 ) ;
  assign n16337 = x32 & n16335 ;
  assign n16338 = x32 & n16328 ;
  assign n16339 = ( x32 & n16332 ) | ( x32 & n16338 ) | ( n16332 & n16338 ) ;
  assign n16340 = ( n4305 & n16337 ) | ( n4305 & n16339 ) | ( n16337 & n16339 ) ;
  assign n16341 = x32 & ~n16339 ;
  assign n16342 = x32 & ~n16335 ;
  assign n16343 = ( ~n4305 & n16341 ) | ( ~n4305 & n16342 ) | ( n16341 & n16342 ) ;
  assign n16344 = ( n16336 & ~n16340 ) | ( n16336 & n16343 ) | ( ~n16340 & n16343 ) ;
  assign n16345 = n16327 & n16344 ;
  assign n16346 = n16327 | n16344 ;
  assign n16347 = ~n16345 & n16346 ;
  assign n16348 = ( n15252 & n15770 ) | ( n15252 & n15787 ) | ( n15770 & n15787 ) ;
  assign n16349 = n15770 | n15787 ;
  assign n16350 = ( n15255 & n16348 ) | ( n15255 & n16349 ) | ( n16348 & n16349 ) ;
  assign n16351 = n16347 & n16350 ;
  assign n16352 = ~n16347 & n16350 ;
  assign n16353 = ( n16347 & ~n16351 ) | ( n16347 & n16352 ) | ( ~n16351 & n16352 ) ;
  assign n16354 = x96 & n3816 ;
  assign n16355 = x95 & n3811 ;
  assign n16356 = x94 & ~n3810 ;
  assign n16357 = n4067 & n16356 ;
  assign n16358 = n16355 | n16357 ;
  assign n16359 = n16354 | n16358 ;
  assign n16360 = n3819 | n16354 ;
  assign n16361 = n16358 | n16360 ;
  assign n16362 = ( n5202 & n16359 ) | ( n5202 & n16361 ) | ( n16359 & n16361 ) ;
  assign n16363 = x29 & n16361 ;
  assign n16364 = x29 & n16354 ;
  assign n16365 = ( x29 & n16358 ) | ( x29 & n16364 ) | ( n16358 & n16364 ) ;
  assign n16366 = ( n5202 & n16363 ) | ( n5202 & n16365 ) | ( n16363 & n16365 ) ;
  assign n16367 = x29 & ~n16365 ;
  assign n16368 = x29 & ~n16361 ;
  assign n16369 = ( ~n5202 & n16367 ) | ( ~n5202 & n16368 ) | ( n16367 & n16368 ) ;
  assign n16370 = ( n16362 & ~n16366 ) | ( n16362 & n16369 ) | ( ~n16366 & n16369 ) ;
  assign n16371 = n16353 | n16370 ;
  assign n16372 = n16353 & n16370 ;
  assign n16373 = n16371 & ~n16372 ;
  assign n16374 = n15815 & n16373 ;
  assign n16375 = ( n15821 & n16373 ) | ( n15821 & n16374 ) | ( n16373 & n16374 ) ;
  assign n16376 = n15815 | n16373 ;
  assign n16377 = n15821 | n16376 ;
  assign n16378 = ~n16375 & n16377 ;
  assign n16379 = x99 & n3085 ;
  assign n16380 = x98 & n3080 ;
  assign n16381 = x97 & ~n3079 ;
  assign n16382 = n3309 & n16381 ;
  assign n16383 = n16380 | n16382 ;
  assign n16384 = n16379 | n16383 ;
  assign n16385 = n3088 | n16379 ;
  assign n16386 = n16383 | n16385 ;
  assign n16387 = ( n6164 & n16384 ) | ( n6164 & n16386 ) | ( n16384 & n16386 ) ;
  assign n16388 = x26 & n16386 ;
  assign n16389 = x26 & n16379 ;
  assign n16390 = ( x26 & n16383 ) | ( x26 & n16389 ) | ( n16383 & n16389 ) ;
  assign n16391 = ( n6164 & n16388 ) | ( n6164 & n16390 ) | ( n16388 & n16390 ) ;
  assign n16392 = x26 & ~n16390 ;
  assign n16393 = x26 & ~n16386 ;
  assign n16394 = ( ~n6164 & n16392 ) | ( ~n6164 & n16393 ) | ( n16392 & n16393 ) ;
  assign n16395 = ( n16387 & ~n16391 ) | ( n16387 & n16394 ) | ( ~n16391 & n16394 ) ;
  assign n16396 = n16378 & n16395 ;
  assign n16397 = n16378 & ~n16396 ;
  assign n16398 = ~n16378 & n16395 ;
  assign n16399 = n16397 | n16398 ;
  assign n16400 = n15846 | n15852 ;
  assign n16401 = n16399 | n16400 ;
  assign n16402 = n16399 & n16400 ;
  assign n16403 = n16401 & ~n16402 ;
  assign n16404 = x102 & n2429 ;
  assign n16405 = x101 & n2424 ;
  assign n16406 = x100 & ~n2423 ;
  assign n16407 = n2631 & n16406 ;
  assign n16408 = n16405 | n16407 ;
  assign n16409 = n16404 | n16408 ;
  assign n16410 = n2432 | n16404 ;
  assign n16411 = n16408 | n16410 ;
  assign n16412 = ( n7178 & n16409 ) | ( n7178 & n16411 ) | ( n16409 & n16411 ) ;
  assign n16413 = x23 & n16411 ;
  assign n16414 = x23 & n16404 ;
  assign n16415 = ( x23 & n16408 ) | ( x23 & n16414 ) | ( n16408 & n16414 ) ;
  assign n16416 = ( n7178 & n16413 ) | ( n7178 & n16415 ) | ( n16413 & n16415 ) ;
  assign n16417 = x23 & ~n16415 ;
  assign n16418 = x23 & ~n16411 ;
  assign n16419 = ( ~n7178 & n16417 ) | ( ~n7178 & n16418 ) | ( n16417 & n16418 ) ;
  assign n16420 = ( n16412 & ~n16416 ) | ( n16412 & n16419 ) | ( ~n16416 & n16419 ) ;
  assign n16421 = n16403 & n16420 ;
  assign n16422 = n16403 & ~n16421 ;
  assign n16423 = ~n16403 & n16420 ;
  assign n16424 = n16422 | n16423 ;
  assign n16425 = n15871 | n15878 ;
  assign n16426 = n16424 | n16425 ;
  assign n16427 = n16424 & n16425 ;
  assign n16428 = n16426 & ~n16427 ;
  assign n16429 = x105 & n1859 ;
  assign n16430 = x104 & n1854 ;
  assign n16431 = x103 & ~n1853 ;
  assign n16432 = n2037 & n16431 ;
  assign n16433 = n16430 | n16432 ;
  assign n16434 = n16429 | n16433 ;
  assign n16435 = n1862 | n16429 ;
  assign n16436 = n16433 | n16435 ;
  assign n16437 = ( n8273 & n16434 ) | ( n8273 & n16436 ) | ( n16434 & n16436 ) ;
  assign n16438 = x20 & n16436 ;
  assign n16439 = x20 & n16429 ;
  assign n16440 = ( x20 & n16433 ) | ( x20 & n16439 ) | ( n16433 & n16439 ) ;
  assign n16441 = ( n8273 & n16438 ) | ( n8273 & n16440 ) | ( n16438 & n16440 ) ;
  assign n16442 = x20 & ~n16440 ;
  assign n16443 = x20 & ~n16436 ;
  assign n16444 = ( ~n8273 & n16442 ) | ( ~n8273 & n16443 ) | ( n16442 & n16443 ) ;
  assign n16445 = ( n16437 & ~n16441 ) | ( n16437 & n16444 ) | ( ~n16441 & n16444 ) ;
  assign n16446 = n16428 & n16445 ;
  assign n16447 = n16428 | n16445 ;
  assign n16448 = ~n16446 & n16447 ;
  assign n16449 = n15897 & n16448 ;
  assign n16450 = ( n15903 & n16448 ) | ( n15903 & n16449 ) | ( n16448 & n16449 ) ;
  assign n16451 = n15897 | n15899 ;
  assign n16452 = n15898 | n16451 ;
  assign n16453 = ( n15897 & n15901 ) | ( n15897 & n16452 ) | ( n15901 & n16452 ) ;
  assign n16454 = n16448 | n16453 ;
  assign n16455 = ~n16450 & n16454 ;
  assign n16456 = x108 & n1383 ;
  assign n16457 = x107 & n1378 ;
  assign n16458 = x106 & ~n1377 ;
  assign n16459 = n1542 & n16458 ;
  assign n16460 = n16457 | n16459 ;
  assign n16461 = n16456 | n16460 ;
  assign n16462 = n1386 | n16456 ;
  assign n16463 = n16460 | n16462 ;
  assign n16464 = ( n9479 & n16461 ) | ( n9479 & n16463 ) | ( n16461 & n16463 ) ;
  assign n16465 = x17 & n16463 ;
  assign n16466 = x17 & n16456 ;
  assign n16467 = ( x17 & n16460 ) | ( x17 & n16466 ) | ( n16460 & n16466 ) ;
  assign n16468 = ( n9479 & n16465 ) | ( n9479 & n16467 ) | ( n16465 & n16467 ) ;
  assign n16469 = x17 & ~n16467 ;
  assign n16470 = x17 & ~n16463 ;
  assign n16471 = ( ~n9479 & n16469 ) | ( ~n9479 & n16470 ) | ( n16469 & n16470 ) ;
  assign n16472 = ( n16464 & ~n16468 ) | ( n16464 & n16471 ) | ( ~n16468 & n16471 ) ;
  assign n16473 = n16455 & n16472 ;
  assign n16474 = n16455 & ~n16473 ;
  assign n16475 = ~n16455 & n16472 ;
  assign n16476 = n16474 | n16475 ;
  assign n16477 = n16103 & ~n16476 ;
  assign n16478 = ~n16103 & n16476 ;
  assign n16479 = n16477 | n16478 ;
  assign n16480 = x111 & n962 ;
  assign n16481 = x110 & n957 ;
  assign n16482 = x109 & ~n956 ;
  assign n16483 = n1105 & n16482 ;
  assign n16484 = n16481 | n16483 ;
  assign n16485 = n16480 | n16484 ;
  assign n16486 = n965 | n16480 ;
  assign n16487 = n16484 | n16486 ;
  assign n16488 = ( n10749 & n16485 ) | ( n10749 & n16487 ) | ( n16485 & n16487 ) ;
  assign n16489 = x14 & n16487 ;
  assign n16490 = x14 & n16480 ;
  assign n16491 = ( x14 & n16484 ) | ( x14 & n16490 ) | ( n16484 & n16490 ) ;
  assign n16492 = ( n10749 & n16489 ) | ( n10749 & n16491 ) | ( n16489 & n16491 ) ;
  assign n16493 = x14 & ~n16491 ;
  assign n16494 = x14 & ~n16487 ;
  assign n16495 = ( ~n10749 & n16493 ) | ( ~n10749 & n16494 ) | ( n16493 & n16494 ) ;
  assign n16496 = ( n16488 & ~n16492 ) | ( n16488 & n16495 ) | ( ~n16492 & n16495 ) ;
  assign n16497 = n16479 & n16496 ;
  assign n16498 = n16479 | n16496 ;
  assign n16499 = ~n16497 & n16498 ;
  assign n16500 = n15948 | n15954 ;
  assign n16501 = n16499 & n16500 ;
  assign n16502 = n16499 | n16500 ;
  assign n16503 = ~n16501 & n16502 ;
  assign n16504 = x114 & n636 ;
  assign n16505 = x113 & n631 ;
  assign n16506 = x112 & ~n630 ;
  assign n16507 = n764 & n16506 ;
  assign n16508 = n16505 | n16507 ;
  assign n16509 = n16504 | n16508 ;
  assign n16510 = n639 | n16504 ;
  assign n16511 = n16508 | n16510 ;
  assign n16512 = ( ~n12095 & n16509 ) | ( ~n12095 & n16511 ) | ( n16509 & n16511 ) ;
  assign n16513 = n16509 & n16511 ;
  assign n16514 = ( n12079 & n16512 ) | ( n12079 & n16513 ) | ( n16512 & n16513 ) ;
  assign n16515 = x11 & n16514 ;
  assign n16516 = x11 & ~n16514 ;
  assign n16517 = ( n16514 & ~n16515 ) | ( n16514 & n16516 ) | ( ~n16515 & n16516 ) ;
  assign n16518 = n16503 & n16517 ;
  assign n16519 = n16503 & ~n16518 ;
  assign n16520 = ~n16503 & n16517 ;
  assign n16521 = n16519 | n16520 ;
  assign n16522 = n15973 | n15976 ;
  assign n16523 = n16521 & n16522 ;
  assign n16524 = n16521 | n16522 ;
  assign n16525 = ~n16523 & n16524 ;
  assign n16526 = x117 & n389 ;
  assign n16527 = x116 & n384 ;
  assign n16528 = x115 & ~n383 ;
  assign n16529 = n463 & n16528 ;
  assign n16530 = n16527 | n16529 ;
  assign n16531 = n16526 | n16530 ;
  assign n16532 = n392 | n16526 ;
  assign n16533 = n16530 | n16532 ;
  assign n16534 = ( ~n13522 & n16531 ) | ( ~n13522 & n16533 ) | ( n16531 & n16533 ) ;
  assign n16535 = n16531 & n16533 ;
  assign n16536 = ( n13503 & n16534 ) | ( n13503 & n16535 ) | ( n16534 & n16535 ) ;
  assign n16537 = x8 & n16536 ;
  assign n16538 = x8 & ~n16536 ;
  assign n16539 = ( n16536 & ~n16537 ) | ( n16536 & n16538 ) | ( ~n16537 & n16538 ) ;
  assign n16540 = n16525 & n16539 ;
  assign n16541 = n16525 & ~n16540 ;
  assign n16542 = ~n16525 & n16539 ;
  assign n16543 = n16541 | n16542 ;
  assign n16544 = n16102 & n16543 ;
  assign n16545 = n16102 & ~n16544 ;
  assign n16546 = n16543 & ~n16544 ;
  assign n16547 = n16545 | n16546 ;
  assign n16548 = x120 & n212 ;
  assign n16549 = x119 & n207 ;
  assign n16550 = x118 & ~n206 ;
  assign n16551 = n267 & n16550 ;
  assign n16552 = n16549 | n16551 ;
  assign n16553 = n16548 | n16552 ;
  assign n16554 = n215 | n16548 ;
  assign n16555 = n16552 | n16554 ;
  assign n16556 = ( n14991 & n16553 ) | ( n14991 & n16555 ) | ( n16553 & n16555 ) ;
  assign n16557 = x5 & n16555 ;
  assign n16558 = x5 & n16548 ;
  assign n16559 = ( x5 & n16552 ) | ( x5 & n16558 ) | ( n16552 & n16558 ) ;
  assign n16560 = ( n14991 & n16557 ) | ( n14991 & n16559 ) | ( n16557 & n16559 ) ;
  assign n16561 = x5 & ~n16559 ;
  assign n16562 = x5 & ~n16555 ;
  assign n16563 = ( ~n14991 & n16561 ) | ( ~n14991 & n16562 ) | ( n16561 & n16562 ) ;
  assign n16564 = ( n16556 & ~n16560 ) | ( n16556 & n16563 ) | ( ~n16560 & n16563 ) ;
  assign n16565 = ( n16101 & n16547 ) | ( n16101 & ~n16564 ) | ( n16547 & ~n16564 ) ;
  assign n16566 = ( ~n16547 & n16564 ) | ( ~n16547 & n16565 ) | ( n16564 & n16565 ) ;
  assign n16567 = ( ~n16101 & n16565 ) | ( ~n16101 & n16566 ) | ( n16565 & n16566 ) ;
  assign n16568 = n16020 | n16021 ;
  assign n16569 = ( n15527 & n16020 ) | ( n15527 & n16568 ) | ( n16020 & n16568 ) ;
  assign n16570 = n16565 & n16569 ;
  assign n16571 = ~n16101 & n16569 ;
  assign n16572 = ( n16566 & n16570 ) | ( n16566 & n16571 ) | ( n16570 & n16571 ) ;
  assign n16573 = n16567 & ~n16572 ;
  assign n16574 = ~n16565 & n16569 ;
  assign n16575 = n16101 & n16569 ;
  assign n16576 = ( ~n16566 & n16574 ) | ( ~n16566 & n16575 ) | ( n16574 & n16575 ) ;
  assign n16577 = n16573 | n16576 ;
  assign n16578 = n16067 | n16577 ;
  assign n16579 = n16059 & n16576 ;
  assign n16580 = ( n16059 & n16573 ) | ( n16059 & n16579 ) | ( n16573 & n16579 ) ;
  assign n16581 = ( n16064 & n16577 ) | ( n16064 & n16580 ) | ( n16577 & n16580 ) ;
  assign n16582 = n16578 & ~n16581 ;
  assign n16583 = n16540 | n16544 ;
  assign n16584 = n16518 | n16523 ;
  assign n16585 = n16446 | n16450 ;
  assign n16586 = x82 & n8724 ;
  assign n16587 = x81 & n8719 ;
  assign n16588 = x80 & ~n8718 ;
  assign n16589 = n9149 & n16588 ;
  assign n16590 = n16587 | n16589 ;
  assign n16591 = n16586 | n16590 ;
  assign n16592 = n8727 | n16586 ;
  assign n16593 = n16590 | n16592 ;
  assign n16594 = ( n1811 & n16591 ) | ( n1811 & n16593 ) | ( n16591 & n16593 ) ;
  assign n16595 = x44 & n16593 ;
  assign n16596 = x44 & n16586 ;
  assign n16597 = ( x44 & n16590 ) | ( x44 & n16596 ) | ( n16590 & n16596 ) ;
  assign n16598 = ( n1811 & n16595 ) | ( n1811 & n16597 ) | ( n16595 & n16597 ) ;
  assign n16599 = x44 & ~n16597 ;
  assign n16600 = x44 & ~n16593 ;
  assign n16601 = ( ~n1811 & n16599 ) | ( ~n1811 & n16600 ) | ( n16599 & n16600 ) ;
  assign n16602 = ( n16594 & ~n16598 ) | ( n16594 & n16601 ) | ( ~n16598 & n16601 ) ;
  assign n16729 = n16236 | n16242 ;
  assign n16730 = ( n16236 & n16239 ) | ( n16236 & n16729 ) | ( n16239 & n16729 ) ;
  assign n16603 = n16154 | n16158 ;
  assign n16604 = x59 & ~x60 ;
  assign n16605 = ~x59 & x60 ;
  assign n16606 = n16604 | n16605 ;
  assign n16607 = x64 & n16606 ;
  assign n16608 = ~n15567 & n16607 ;
  assign n16609 = ( ~n16135 & n16607 ) | ( ~n16135 & n16608 ) | ( n16607 & n16608 ) ;
  assign n16610 = n15567 & ~n16607 ;
  assign n16611 = n16135 & n16610 ;
  assign n16612 = n16609 | n16611 ;
  assign n16613 = x67 & n15552 ;
  assign n16614 = x66 & n15547 ;
  assign n16615 = x65 & ~n15546 ;
  assign n16616 = n16123 & n16615 ;
  assign n16617 = n16614 | n16616 ;
  assign n16618 = n16613 | n16617 ;
  assign n16619 = n186 & n15555 ;
  assign n16620 = n16618 | n16619 ;
  assign n16621 = x59 & ~n16620 ;
  assign n16622 = ~x59 & n16620 ;
  assign n16623 = n16621 | n16622 ;
  assign n16624 = n16612 & n16623 ;
  assign n16625 = n16612 | n16623 ;
  assign n16626 = ~n16624 & n16625 ;
  assign n16627 = x69 & n14040 ;
  assign n16628 = x68 & ~n14039 ;
  assign n16629 = n14552 & n16628 ;
  assign n16630 = n16627 | n16629 ;
  assign n16631 = x70 & n14045 ;
  assign n16632 = n14048 | n16631 ;
  assign n16633 = n16630 | n16632 ;
  assign n16634 = x56 & ~n16633 ;
  assign n16635 = x56 & ~n16631 ;
  assign n16636 = ~n16630 & n16635 ;
  assign n16637 = ( ~n340 & n16634 ) | ( ~n340 & n16636 ) | ( n16634 & n16636 ) ;
  assign n16638 = ~x56 & n16633 ;
  assign n16639 = ~x56 & n16631 ;
  assign n16640 = ( ~x56 & n16630 ) | ( ~x56 & n16639 ) | ( n16630 & n16639 ) ;
  assign n16641 = ( n340 & n16638 ) | ( n340 & n16640 ) | ( n16638 & n16640 ) ;
  assign n16642 = n16637 | n16641 ;
  assign n16643 = ( n16154 & ~n16626 ) | ( n16154 & n16642 ) | ( ~n16626 & n16642 ) ;
  assign n16644 = n16626 & ~n16642 ;
  assign n16645 = ( n16158 & n16643 ) | ( n16158 & ~n16644 ) | ( n16643 & ~n16644 ) ;
  assign n16646 = ( ~n16603 & n16626 ) | ( ~n16603 & n16645 ) | ( n16626 & n16645 ) ;
  assign n16647 = x73 & n12574 ;
  assign n16648 = x72 & n12569 ;
  assign n16649 = x71 & ~n12568 ;
  assign n16650 = n13076 & n16649 ;
  assign n16651 = n16648 | n16650 ;
  assign n16652 = n16647 | n16651 ;
  assign n16653 = ( ~n610 & n12577 ) | ( ~n610 & n16652 ) | ( n12577 & n16652 ) ;
  assign n16654 = n12577 & n16647 ;
  assign n16655 = ( n12577 & n16651 ) | ( n12577 & n16654 ) | ( n16651 & n16654 ) ;
  assign n16656 = ( n598 & n16653 ) | ( n598 & n16655 ) | ( n16653 & n16655 ) ;
  assign n16657 = ( x53 & ~n16652 ) | ( x53 & n16656 ) | ( ~n16652 & n16656 ) ;
  assign n16658 = ~n16656 & n16657 ;
  assign n16659 = x53 | n16647 ;
  assign n16660 = n16651 | n16659 ;
  assign n16661 = n16656 | n16660 ;
  assign n16662 = ( ~x53 & n16658 ) | ( ~x53 & n16661 ) | ( n16658 & n16661 ) ;
  assign n16663 = n16645 & n16662 ;
  assign n16664 = ~n16642 & n16661 ;
  assign n16665 = x53 | n16642 ;
  assign n16666 = ( n16658 & n16664 ) | ( n16658 & ~n16665 ) | ( n16664 & ~n16665 ) ;
  assign n16667 = ( n16646 & n16663 ) | ( n16646 & n16666 ) | ( n16663 & n16666 ) ;
  assign n16668 = n16645 | n16662 ;
  assign n16669 = n16642 & ~n16661 ;
  assign n16670 = x53 & n16642 ;
  assign n16671 = ( ~n16658 & n16669 ) | ( ~n16658 & n16670 ) | ( n16669 & n16670 ) ;
  assign n16672 = ( n16646 & n16668 ) | ( n16646 & ~n16671 ) | ( n16668 & ~n16671 ) ;
  assign n16673 = ~n16667 & n16672 ;
  assign n16674 = n16162 | n16165 ;
  assign n16675 = ( n16162 & n16167 ) | ( n16162 & n16674 ) | ( n16167 & n16674 ) ;
  assign n16676 = n16673 & n16675 ;
  assign n16677 = n16673 | n16675 ;
  assign n16678 = ~n16676 & n16677 ;
  assign n16679 = x76 & n11205 ;
  assign n16680 = x75 & n11200 ;
  assign n16681 = x74 & ~n11199 ;
  assign n16682 = n11679 & n16681 ;
  assign n16683 = n16680 | n16682 ;
  assign n16684 = n16679 | n16683 ;
  assign n16685 = n11208 | n16679 ;
  assign n16686 = n16683 | n16685 ;
  assign n16687 = ( n923 & n16684 ) | ( n923 & n16686 ) | ( n16684 & n16686 ) ;
  assign n16688 = x50 & n16686 ;
  assign n16689 = x50 & n16679 ;
  assign n16690 = ( x50 & n16683 ) | ( x50 & n16689 ) | ( n16683 & n16689 ) ;
  assign n16691 = ( n923 & n16688 ) | ( n923 & n16690 ) | ( n16688 & n16690 ) ;
  assign n16692 = x50 & ~n16690 ;
  assign n16693 = x50 & ~n16686 ;
  assign n16694 = ( ~n923 & n16692 ) | ( ~n923 & n16693 ) | ( n16692 & n16693 ) ;
  assign n16695 = ( n16687 & ~n16691 ) | ( n16687 & n16694 ) | ( ~n16691 & n16694 ) ;
  assign n16696 = n16678 | n16695 ;
  assign n16697 = n16678 & n16695 ;
  assign n16698 = n16696 & ~n16697 ;
  assign n16699 = n16189 | n16190 ;
  assign n16700 = ( n16189 & n16191 ) | ( n16189 & n16699 ) | ( n16191 & n16699 ) ;
  assign n16701 = n16698 & n16700 ;
  assign n16702 = n16698 | n16700 ;
  assign n16703 = ~n16701 & n16702 ;
  assign n16704 = x79 & n9933 ;
  assign n16705 = x78 & n9928 ;
  assign n16706 = x77 & ~n9927 ;
  assign n16707 = n10379 & n16706 ;
  assign n16708 = n16705 | n16707 ;
  assign n16709 = n16704 | n16708 ;
  assign n16710 = n9936 | n16704 ;
  assign n16711 = n16708 | n16710 ;
  assign n16712 = ( n1332 & n16709 ) | ( n1332 & n16711 ) | ( n16709 & n16711 ) ;
  assign n16713 = x47 & n16711 ;
  assign n16714 = x47 & n16704 ;
  assign n16715 = ( x47 & n16708 ) | ( x47 & n16714 ) | ( n16708 & n16714 ) ;
  assign n16716 = ( n1332 & n16713 ) | ( n1332 & n16715 ) | ( n16713 & n16715 ) ;
  assign n16717 = x47 & ~n16715 ;
  assign n16718 = x47 & ~n16711 ;
  assign n16719 = ( ~n1332 & n16717 ) | ( ~n1332 & n16718 ) | ( n16717 & n16718 ) ;
  assign n16720 = ( n16712 & ~n16716 ) | ( n16712 & n16719 ) | ( ~n16716 & n16719 ) ;
  assign n16721 = n16703 & n16720 ;
  assign n16722 = n16703 | n16720 ;
  assign n16723 = ~n16721 & n16722 ;
  assign n16724 = n16212 & n16723 ;
  assign n16725 = ( n16216 & n16723 ) | ( n16216 & n16724 ) | ( n16723 & n16724 ) ;
  assign n16726 = n16212 | n16723 ;
  assign n16727 = n16216 | n16726 ;
  assign n16728 = ~n16725 & n16727 ;
  assign n16731 = ( n16602 & n16728 ) | ( n16602 & ~n16730 ) | ( n16728 & ~n16730 ) ;
  assign n16732 = ( ~n16602 & n16730 ) | ( ~n16602 & n16731 ) | ( n16730 & n16731 ) ;
  assign n16733 = x85 & n7566 ;
  assign n16734 = x84 & n7561 ;
  assign n16735 = x83 & ~n7560 ;
  assign n16736 = n7953 & n16735 ;
  assign n16737 = n16734 | n16736 ;
  assign n16738 = n16733 | n16737 ;
  assign n16739 = n7569 | n16733 ;
  assign n16740 = n16737 | n16739 ;
  assign n16741 = ( n2381 & n16738 ) | ( n2381 & n16740 ) | ( n16738 & n16740 ) ;
  assign n16742 = x41 & n16740 ;
  assign n16743 = x41 & n16733 ;
  assign n16744 = ( x41 & n16737 ) | ( x41 & n16743 ) | ( n16737 & n16743 ) ;
  assign n16745 = ( n2381 & n16742 ) | ( n2381 & n16744 ) | ( n16742 & n16744 ) ;
  assign n16746 = x41 & ~n16744 ;
  assign n16747 = x41 & ~n16740 ;
  assign n16748 = ( ~n2381 & n16746 ) | ( ~n2381 & n16747 ) | ( n16746 & n16747 ) ;
  assign n16749 = ( n16741 & ~n16745 ) | ( n16741 & n16748 ) | ( ~n16745 & n16748 ) ;
  assign n16750 = ~n16728 & n16749 ;
  assign n16751 = n16728 & n16749 ;
  assign n16752 = n16602 & n16749 ;
  assign n16753 = ( ~n16730 & n16751 ) | ( ~n16730 & n16752 ) | ( n16751 & n16752 ) ;
  assign n16754 = ( n16732 & n16750 ) | ( n16732 & n16753 ) | ( n16750 & n16753 ) ;
  assign n16755 = n16728 & ~n16749 ;
  assign n16756 = n16728 | n16749 ;
  assign n16757 = n16602 | n16749 ;
  assign n16758 = ( ~n16730 & n16756 ) | ( ~n16730 & n16757 ) | ( n16756 & n16757 ) ;
  assign n16759 = ( n16732 & ~n16755 ) | ( n16732 & n16758 ) | ( ~n16755 & n16758 ) ;
  assign n16760 = ~n16754 & n16759 ;
  assign n16761 = ( n16246 & n16263 ) | ( n16246 & n16273 ) | ( n16263 & n16273 ) ;
  assign n16762 = n16760 | n16761 ;
  assign n16763 = n16760 & n16761 ;
  assign n16764 = n16762 & ~n16763 ;
  assign n16765 = x88 & n6536 ;
  assign n16766 = x87 & n6531 ;
  assign n16767 = x86 & ~n6530 ;
  assign n16768 = n6871 & n16767 ;
  assign n16769 = n16766 | n16768 ;
  assign n16770 = n16765 | n16769 ;
  assign n16771 = n6539 | n16765 ;
  assign n16772 = n16769 | n16771 ;
  assign n16773 = ( ~n3039 & n16770 ) | ( ~n3039 & n16772 ) | ( n16770 & n16772 ) ;
  assign n16774 = n16770 & n16772 ;
  assign n16775 = ( n3023 & n16773 ) | ( n3023 & n16774 ) | ( n16773 & n16774 ) ;
  assign n16776 = x38 & n16772 ;
  assign n16777 = x38 & n16765 ;
  assign n16778 = ( x38 & n16769 ) | ( x38 & n16777 ) | ( n16769 & n16777 ) ;
  assign n16779 = ( ~n3039 & n16776 ) | ( ~n3039 & n16778 ) | ( n16776 & n16778 ) ;
  assign n16780 = n16776 & n16778 ;
  assign n16781 = ( n3023 & n16779 ) | ( n3023 & n16780 ) | ( n16779 & n16780 ) ;
  assign n16782 = x38 & ~n16778 ;
  assign n16783 = x38 & ~n16772 ;
  assign n16784 = ( n3039 & n16782 ) | ( n3039 & n16783 ) | ( n16782 & n16783 ) ;
  assign n16785 = n16782 | n16783 ;
  assign n16786 = ( ~n3023 & n16784 ) | ( ~n3023 & n16785 ) | ( n16784 & n16785 ) ;
  assign n16787 = ( n16775 & ~n16781 ) | ( n16775 & n16786 ) | ( ~n16781 & n16786 ) ;
  assign n16788 = n16764 & n16787 ;
  assign n16789 = n16764 & ~n16788 ;
  assign n16790 = ~n16764 & n16787 ;
  assign n16791 = n16789 | n16790 ;
  assign n16792 = n16294 | n16300 ;
  assign n16793 = n16791 | n16792 ;
  assign n16794 = n16791 & n16792 ;
  assign n16795 = n16793 & ~n16794 ;
  assign n16796 = x91 & n5554 ;
  assign n16797 = x90 & n5549 ;
  assign n16798 = x89 & ~n5548 ;
  assign n16799 = n5893 & n16798 ;
  assign n16800 = n16797 | n16799 ;
  assign n16801 = n16796 | n16800 ;
  assign n16802 = n5557 | n16796 ;
  assign n16803 = n16800 | n16802 ;
  assign n16804 = ( n3768 & n16801 ) | ( n3768 & n16803 ) | ( n16801 & n16803 ) ;
  assign n16805 = x35 & n16803 ;
  assign n16806 = x35 & n16796 ;
  assign n16807 = ( x35 & n16800 ) | ( x35 & n16806 ) | ( n16800 & n16806 ) ;
  assign n16808 = ( n3768 & n16805 ) | ( n3768 & n16807 ) | ( n16805 & n16807 ) ;
  assign n16809 = x35 & ~n16807 ;
  assign n16810 = x35 & ~n16803 ;
  assign n16811 = ( ~n3768 & n16809 ) | ( ~n3768 & n16810 ) | ( n16809 & n16810 ) ;
  assign n16812 = ( n16804 & ~n16808 ) | ( n16804 & n16811 ) | ( ~n16808 & n16811 ) ;
  assign n16813 = n16795 & n16812 ;
  assign n16814 = n16795 & ~n16813 ;
  assign n16815 = ~n16795 & n16812 ;
  assign n16816 = n16814 | n16815 ;
  assign n16817 = n16319 | n16321 ;
  assign n16818 = n16320 | n16817 ;
  assign n16819 = ( n16319 & n16324 ) | ( n16319 & n16818 ) | ( n16324 & n16818 ) ;
  assign n16820 = n16816 | n16819 ;
  assign n16821 = n16816 & n16819 ;
  assign n16822 = n16820 & ~n16821 ;
  assign n16823 = x94 & n4631 ;
  assign n16824 = x93 & n4626 ;
  assign n16825 = x92 & ~n4625 ;
  assign n16826 = n4943 & n16825 ;
  assign n16827 = n16824 | n16826 ;
  assign n16828 = n16823 | n16827 ;
  assign n16829 = n4634 | n16823 ;
  assign n16830 = n16827 | n16829 ;
  assign n16831 = ( n4583 & n16828 ) | ( n4583 & n16830 ) | ( n16828 & n16830 ) ;
  assign n16832 = x32 & n16830 ;
  assign n16833 = x32 & n16823 ;
  assign n16834 = ( x32 & n16827 ) | ( x32 & n16833 ) | ( n16827 & n16833 ) ;
  assign n16835 = ( n4583 & n16832 ) | ( n4583 & n16834 ) | ( n16832 & n16834 ) ;
  assign n16836 = x32 & ~n16834 ;
  assign n16837 = x32 & ~n16830 ;
  assign n16838 = ( ~n4583 & n16836 ) | ( ~n4583 & n16837 ) | ( n16836 & n16837 ) ;
  assign n16839 = ( n16831 & ~n16835 ) | ( n16831 & n16838 ) | ( ~n16835 & n16838 ) ;
  assign n16840 = n16822 | n16839 ;
  assign n16841 = n16822 & n16839 ;
  assign n16842 = n16840 & ~n16841 ;
  assign n16843 = n16345 | n16350 ;
  assign n16844 = ( n16345 & n16347 ) | ( n16345 & n16843 ) | ( n16347 & n16843 ) ;
  assign n16845 = n16842 & n16844 ;
  assign n16846 = n16842 | n16844 ;
  assign n16847 = ~n16845 & n16846 ;
  assign n16848 = x97 & n3816 ;
  assign n16849 = x96 & n3811 ;
  assign n16850 = x95 & ~n3810 ;
  assign n16851 = n4067 & n16850 ;
  assign n16852 = n16849 | n16851 ;
  assign n16853 = n16848 | n16852 ;
  assign n16854 = n3819 | n16848 ;
  assign n16855 = n16852 | n16854 ;
  assign n16856 = ( n5505 & n16853 ) | ( n5505 & n16855 ) | ( n16853 & n16855 ) ;
  assign n16857 = x29 & n16855 ;
  assign n16858 = x29 & n16848 ;
  assign n16859 = ( x29 & n16852 ) | ( x29 & n16858 ) | ( n16852 & n16858 ) ;
  assign n16860 = ( n5505 & n16857 ) | ( n5505 & n16859 ) | ( n16857 & n16859 ) ;
  assign n16861 = x29 & ~n16859 ;
  assign n16862 = x29 & ~n16855 ;
  assign n16863 = ( ~n5505 & n16861 ) | ( ~n5505 & n16862 ) | ( n16861 & n16862 ) ;
  assign n16864 = ( n16856 & ~n16860 ) | ( n16856 & n16863 ) | ( ~n16860 & n16863 ) ;
  assign n16865 = n16847 & n16864 ;
  assign n16866 = n16847 & ~n16865 ;
  assign n16867 = ~n16847 & n16864 ;
  assign n16868 = n16866 | n16867 ;
  assign n16869 = n15815 | n15821 ;
  assign n16870 = n16372 | n16373 ;
  assign n16871 = ( n16372 & n16869 ) | ( n16372 & n16870 ) | ( n16869 & n16870 ) ;
  assign n16872 = ~n16868 & n16871 ;
  assign n16873 = n16868 & ~n16871 ;
  assign n16874 = n16872 | n16873 ;
  assign n16875 = x100 & n3085 ;
  assign n16876 = x99 & n3080 ;
  assign n16877 = x98 & ~n3079 ;
  assign n16878 = n3309 & n16877 ;
  assign n16879 = n16876 | n16878 ;
  assign n16880 = n16875 | n16879 ;
  assign n16881 = n3088 | n16875 ;
  assign n16882 = n16879 | n16881 ;
  assign n16883 = ( n6483 & n16880 ) | ( n6483 & n16882 ) | ( n16880 & n16882 ) ;
  assign n16884 = x26 & n16882 ;
  assign n16885 = x26 & n16875 ;
  assign n16886 = ( x26 & n16879 ) | ( x26 & n16885 ) | ( n16879 & n16885 ) ;
  assign n16887 = ( n6483 & n16884 ) | ( n6483 & n16886 ) | ( n16884 & n16886 ) ;
  assign n16888 = x26 & ~n16886 ;
  assign n16889 = x26 & ~n16882 ;
  assign n16890 = ( ~n6483 & n16888 ) | ( ~n6483 & n16889 ) | ( n16888 & n16889 ) ;
  assign n16891 = ( n16883 & ~n16887 ) | ( n16883 & n16890 ) | ( ~n16887 & n16890 ) ;
  assign n16892 = n16874 & n16891 ;
  assign n16893 = n16874 | n16891 ;
  assign n16894 = ~n16892 & n16893 ;
  assign n16895 = n16396 & n16894 ;
  assign n16896 = ( n16402 & n16894 ) | ( n16402 & n16895 ) | ( n16894 & n16895 ) ;
  assign n16897 = n16396 | n16894 ;
  assign n16898 = n16402 | n16897 ;
  assign n16899 = ~n16896 & n16898 ;
  assign n16900 = x103 & n2429 ;
  assign n16901 = x102 & n2424 ;
  assign n16902 = x101 & ~n2423 ;
  assign n16903 = n2631 & n16902 ;
  assign n16904 = n16901 | n16903 ;
  assign n16905 = n16900 | n16904 ;
  assign n16906 = n2432 | n16900 ;
  assign n16907 = n16904 | n16906 ;
  assign n16908 = ( n7529 & n16905 ) | ( n7529 & n16907 ) | ( n16905 & n16907 ) ;
  assign n16909 = x23 & n16907 ;
  assign n16910 = x23 & n16900 ;
  assign n16911 = ( x23 & n16904 ) | ( x23 & n16910 ) | ( n16904 & n16910 ) ;
  assign n16912 = ( n7529 & n16909 ) | ( n7529 & n16911 ) | ( n16909 & n16911 ) ;
  assign n16913 = x23 & ~n16911 ;
  assign n16914 = x23 & ~n16907 ;
  assign n16915 = ( ~n7529 & n16913 ) | ( ~n7529 & n16914 ) | ( n16913 & n16914 ) ;
  assign n16916 = ( n16908 & ~n16912 ) | ( n16908 & n16915 ) | ( ~n16912 & n16915 ) ;
  assign n16917 = n16899 & n16916 ;
  assign n16918 = n16899 & ~n16917 ;
  assign n16919 = ~n16899 & n16916 ;
  assign n16920 = n16918 | n16919 ;
  assign n16921 = n16421 | n16427 ;
  assign n16922 = n16920 | n16921 ;
  assign n16923 = n16920 & n16921 ;
  assign n16924 = n16922 & ~n16923 ;
  assign n16925 = x106 & n1859 ;
  assign n16926 = x105 & n1854 ;
  assign n16927 = x104 & ~n1853 ;
  assign n16928 = n2037 & n16927 ;
  assign n16929 = n16926 | n16928 ;
  assign n16930 = n16925 | n16929 ;
  assign n16931 = n1862 | n16925 ;
  assign n16932 = n16929 | n16931 ;
  assign n16933 = ( n8656 & n16930 ) | ( n8656 & n16932 ) | ( n16930 & n16932 ) ;
  assign n16934 = x20 & n16932 ;
  assign n16935 = x20 & n16925 ;
  assign n16936 = ( x20 & n16929 ) | ( x20 & n16935 ) | ( n16929 & n16935 ) ;
  assign n16937 = ( n8656 & n16934 ) | ( n8656 & n16936 ) | ( n16934 & n16936 ) ;
  assign n16938 = x20 & ~n16936 ;
  assign n16939 = x20 & ~n16932 ;
  assign n16940 = ( ~n8656 & n16938 ) | ( ~n8656 & n16939 ) | ( n16938 & n16939 ) ;
  assign n16941 = ( n16933 & ~n16937 ) | ( n16933 & n16940 ) | ( ~n16937 & n16940 ) ;
  assign n16942 = n16924 | n16941 ;
  assign n16943 = n16924 & n16941 ;
  assign n16944 = n16942 & ~n16943 ;
  assign n16945 = n16585 & n16944 ;
  assign n16946 = n16585 | n16944 ;
  assign n16947 = ~n16945 & n16946 ;
  assign n16948 = x109 & n1383 ;
  assign n16949 = x108 & n1378 ;
  assign n16950 = x107 & ~n1377 ;
  assign n16951 = n1542 & n16950 ;
  assign n16952 = n16949 | n16951 ;
  assign n16953 = n16948 | n16952 ;
  assign n16954 = n1386 | n16948 ;
  assign n16955 = n16952 | n16954 ;
  assign n16956 = ( n9878 & n16953 ) | ( n9878 & n16955 ) | ( n16953 & n16955 ) ;
  assign n16957 = x17 & n16955 ;
  assign n16958 = x17 & n16948 ;
  assign n16959 = ( x17 & n16952 ) | ( x17 & n16958 ) | ( n16952 & n16958 ) ;
  assign n16960 = ( n9878 & n16957 ) | ( n9878 & n16959 ) | ( n16957 & n16959 ) ;
  assign n16961 = x17 & ~n16959 ;
  assign n16962 = x17 & ~n16955 ;
  assign n16963 = ( ~n9878 & n16961 ) | ( ~n9878 & n16962 ) | ( n16961 & n16962 ) ;
  assign n16964 = ( n16956 & ~n16960 ) | ( n16956 & n16963 ) | ( ~n16960 & n16963 ) ;
  assign n16965 = n16947 & n16964 ;
  assign n16966 = n16947 & ~n16965 ;
  assign n16967 = ( n15922 & n16455 ) | ( n15922 & n16472 ) | ( n16455 & n16472 ) ;
  assign n16968 = n16455 | n16472 ;
  assign n16969 = ( n15927 & n16967 ) | ( n15927 & n16968 ) | ( n16967 & n16968 ) ;
  assign n16970 = ~n16947 & n16964 ;
  assign n16971 = n16969 & n16970 ;
  assign n16972 = ( n16966 & n16969 ) | ( n16966 & n16971 ) | ( n16969 & n16971 ) ;
  assign n16973 = n16969 | n16970 ;
  assign n16974 = n16966 | n16973 ;
  assign n16975 = ~n16972 & n16974 ;
  assign n16976 = x112 & n962 ;
  assign n16977 = x111 & n957 ;
  assign n16978 = x110 & ~n956 ;
  assign n16979 = n1105 & n16978 ;
  assign n16980 = n16977 | n16979 ;
  assign n16981 = n16976 | n16980 ;
  assign n16982 = n965 | n16976 ;
  assign n16983 = n16980 | n16982 ;
  assign n16984 = ( n11172 & n16981 ) | ( n11172 & n16983 ) | ( n16981 & n16983 ) ;
  assign n16985 = x14 & n16983 ;
  assign n16986 = x14 & n16976 ;
  assign n16987 = ( x14 & n16980 ) | ( x14 & n16986 ) | ( n16980 & n16986 ) ;
  assign n16988 = ( n11172 & n16985 ) | ( n11172 & n16987 ) | ( n16985 & n16987 ) ;
  assign n16989 = x14 & ~n16987 ;
  assign n16990 = x14 & ~n16983 ;
  assign n16991 = ( ~n11172 & n16989 ) | ( ~n11172 & n16990 ) | ( n16989 & n16990 ) ;
  assign n16992 = ( n16984 & ~n16988 ) | ( n16984 & n16991 ) | ( ~n16988 & n16991 ) ;
  assign n16993 = n16975 & n16992 ;
  assign n16994 = n16975 & ~n16993 ;
  assign n16995 = ~n16975 & n16992 ;
  assign n16996 = n16994 | n16995 ;
  assign n16997 = n16497 | n16499 ;
  assign n16998 = ( n16497 & n16500 ) | ( n16497 & n16997 ) | ( n16500 & n16997 ) ;
  assign n16999 = n16996 & n16998 ;
  assign n17000 = n16996 | n16998 ;
  assign n17001 = ~n16999 & n17000 ;
  assign n17002 = x115 & n636 ;
  assign n17003 = x114 & n631 ;
  assign n17004 = x113 & ~n630 ;
  assign n17005 = n764 & n17004 ;
  assign n17006 = n17003 | n17005 ;
  assign n17007 = n17002 | n17006 ;
  assign n17008 = n639 | n17002 ;
  assign n17009 = n17006 | n17008 ;
  assign n17010 = ( ~n12550 & n17007 ) | ( ~n12550 & n17009 ) | ( n17007 & n17009 ) ;
  assign n17011 = n17007 & n17009 ;
  assign n17012 = ( n12532 & n17010 ) | ( n12532 & n17011 ) | ( n17010 & n17011 ) ;
  assign n17013 = x11 & n17012 ;
  assign n17014 = x11 & ~n17012 ;
  assign n17015 = ( n17012 & ~n17013 ) | ( n17012 & n17014 ) | ( ~n17013 & n17014 ) ;
  assign n17016 = n17001 & n17015 ;
  assign n17017 = n17001 & ~n17016 ;
  assign n17018 = ~n17001 & n17015 ;
  assign n17019 = n17017 | n17018 ;
  assign n17020 = n16584 & n17019 ;
  assign n17021 = n16584 | n17019 ;
  assign n17022 = ~n17020 & n17021 ;
  assign n17023 = x118 & n389 ;
  assign n17024 = x117 & n384 ;
  assign n17025 = x116 & ~n383 ;
  assign n17026 = n463 & n17025 ;
  assign n17027 = n17024 | n17026 ;
  assign n17028 = n17023 | n17027 ;
  assign n17029 = n392 | n17023 ;
  assign n17030 = n17027 | n17029 ;
  assign n17031 = ( ~n14002 & n17028 ) | ( ~n14002 & n17030 ) | ( n17028 & n17030 ) ;
  assign n17032 = n17028 & n17030 ;
  assign n17033 = ( n13981 & n17031 ) | ( n13981 & n17032 ) | ( n17031 & n17032 ) ;
  assign n17034 = x8 & n17033 ;
  assign n17035 = x8 & ~n17033 ;
  assign n17036 = ( n17033 & ~n17034 ) | ( n17033 & n17035 ) | ( ~n17034 & n17035 ) ;
  assign n17037 = n17022 & n17036 ;
  assign n17038 = n17022 | n17036 ;
  assign n17039 = ~n17037 & n17038 ;
  assign n17040 = n16583 & n17039 ;
  assign n17041 = n16583 | n17039 ;
  assign n17042 = ~n17040 & n17041 ;
  assign n17043 = x121 & n212 ;
  assign n17044 = x120 & n207 ;
  assign n17045 = x119 & ~n206 ;
  assign n17046 = n267 & n17045 ;
  assign n17047 = n17044 | n17046 ;
  assign n17048 = n17043 | n17047 ;
  assign n17049 = n215 | n17043 ;
  assign n17050 = n17047 | n17049 ;
  assign n17051 = ( n15501 & n17048 ) | ( n15501 & n17050 ) | ( n17048 & n17050 ) ;
  assign n17052 = x5 & n17050 ;
  assign n17053 = x5 & n17043 ;
  assign n17054 = ( x5 & n17047 ) | ( x5 & n17053 ) | ( n17047 & n17053 ) ;
  assign n17055 = ( n15501 & n17052 ) | ( n15501 & n17054 ) | ( n17052 & n17054 ) ;
  assign n17056 = x5 & ~n17054 ;
  assign n17057 = x5 & ~n17050 ;
  assign n17058 = ( ~n15501 & n17056 ) | ( ~n15501 & n17057 ) | ( n17056 & n17057 ) ;
  assign n17059 = ( n17051 & ~n17055 ) | ( n17051 & n17058 ) | ( ~n17055 & n17058 ) ;
  assign n17060 = n17042 & n17059 ;
  assign n17061 = n17042 | n17059 ;
  assign n17062 = ~n17060 & n17061 ;
  assign n17063 = x123 | x124 ;
  assign n17064 = x123 & x124 ;
  assign n17065 = n17063 & ~n17064 ;
  assign n17066 = n16026 | n16069 ;
  assign n17067 = ( n16069 & n16070 ) | ( n16069 & n17066 ) | ( n16070 & n17066 ) ;
  assign n17068 = n17065 & n17067 ;
  assign n17069 = n16069 | n16070 ;
  assign n17070 = n17065 & n17069 ;
  assign n17071 = ( n16033 & n17068 ) | ( n16033 & n17070 ) | ( n17068 & n17070 ) ;
  assign n17072 = n16069 & n17065 ;
  assign n17073 = ( n16075 & n17065 ) | ( n16075 & n17072 ) | ( n17065 & n17072 ) ;
  assign n17074 = ( n13965 & n17071 ) | ( n13965 & n17073 ) | ( n17071 & n17073 ) ;
  assign n17075 = n17071 | n17073 ;
  assign n17076 = ( n14002 & n17074 ) | ( n14002 & n17075 ) | ( n17074 & n17075 ) ;
  assign n17077 = n16069 | n16075 ;
  assign n17078 = ( n16033 & n17067 ) | ( n16033 & n17069 ) | ( n17067 & n17069 ) ;
  assign n17079 = n17077 | n17078 ;
  assign n17080 = n17065 | n17079 ;
  assign n17081 = ( n13965 & n17077 ) | ( n13965 & n17078 ) | ( n17077 & n17078 ) ;
  assign n17082 = n17065 | n17081 ;
  assign n17083 = ( n14002 & n17080 ) | ( n14002 & n17082 ) | ( n17080 & n17082 ) ;
  assign n17084 = ~n17076 & n17083 ;
  assign n17085 = x123 & n133 ;
  assign n17086 = x122 & ~n162 ;
  assign n17087 = ( n137 & n17085 ) | ( n137 & n17086 ) | ( n17085 & n17086 ) ;
  assign n17088 = x0 & x124 ;
  assign n17089 = ( ~n137 & n17085 ) | ( ~n137 & n17088 ) | ( n17085 & n17088 ) ;
  assign n17090 = n17087 | n17089 ;
  assign n17091 = n141 | n17090 ;
  assign n17092 = ( n17084 & n17090 ) | ( n17084 & n17091 ) | ( n17090 & n17091 ) ;
  assign n17093 = x2 & n17090 ;
  assign n17094 = ( x2 & n523 ) | ( x2 & n17090 ) | ( n523 & n17090 ) ;
  assign n17095 = ( n17084 & n17093 ) | ( n17084 & n17094 ) | ( n17093 & n17094 ) ;
  assign n17096 = x2 & ~n17094 ;
  assign n17097 = x2 & ~n17090 ;
  assign n17098 = ( ~n17084 & n17096 ) | ( ~n17084 & n17097 ) | ( n17096 & n17097 ) ;
  assign n17099 = ( n17092 & ~n17095 ) | ( n17092 & n17098 ) | ( ~n17095 & n17098 ) ;
  assign n17100 = n17062 & n17099 ;
  assign n17101 = n17062 | n17099 ;
  assign n17102 = ~n17100 & n17101 ;
  assign n17103 = n16547 & n16564 ;
  assign n17104 = n16547 & ~n17103 ;
  assign n17105 = n16101 & ~n16564 ;
  assign n17106 = ( n16101 & n16547 ) | ( n16101 & n17105 ) | ( n16547 & n17105 ) ;
  assign n17107 = ( n16101 & n17103 ) | ( n16101 & ~n17106 ) | ( n17103 & ~n17106 ) ;
  assign n17108 = n16101 | n16564 ;
  assign n17109 = ( n16101 & n16547 ) | ( n16101 & n17108 ) | ( n16547 & n17108 ) ;
  assign n17110 = ( n17104 & n17107 ) | ( n17104 & n17109 ) | ( n17107 & n17109 ) ;
  assign n17111 = n17102 & n17110 ;
  assign n17112 = n17102 | n17110 ;
  assign n17113 = ~n17111 & n17112 ;
  assign n17114 = n16572 | n16580 ;
  assign n17115 = n16572 | n16577 ;
  assign n17116 = ( n16064 & n17114 ) | ( n16064 & n17115 ) | ( n17114 & n17115 ) ;
  assign n17117 = n17113 & n17116 ;
  assign n17118 = n17113 | n17116 ;
  assign n17119 = ~n17117 & n17118 ;
  assign n17120 = n16993 | n16999 ;
  assign n17121 = n16965 | n16972 ;
  assign n17523 = n16943 | n16944 ;
  assign n17524 = ( n16585 & n16943 ) | ( n16585 & n17523 ) | ( n16943 & n17523 ) ;
  assign n17122 = x70 & n14040 ;
  assign n17123 = x69 & ~n14039 ;
  assign n17124 = n14552 & n17123 ;
  assign n17125 = n17122 | n17124 ;
  assign n17126 = x71 & n14045 ;
  assign n17127 = n14048 | n17126 ;
  assign n17128 = n17125 | n17127 ;
  assign n17129 = x56 & ~n17128 ;
  assign n17130 = x56 & ~n17126 ;
  assign n17131 = ~n17125 & n17130 ;
  assign n17132 = ( ~n438 & n17129 ) | ( ~n438 & n17131 ) | ( n17129 & n17131 ) ;
  assign n17133 = ~x56 & n17128 ;
  assign n17134 = ~x56 & n17126 ;
  assign n17135 = ( ~x56 & n17125 ) | ( ~x56 & n17134 ) | ( n17125 & n17134 ) ;
  assign n17136 = ( n438 & n17133 ) | ( n438 & n17135 ) | ( n17133 & n17135 ) ;
  assign n17137 = n17132 | n17136 ;
  assign n17138 = ~x60 & x61 ;
  assign n17139 = x60 & ~x61 ;
  assign n17140 = n17138 | n17139 ;
  assign n17141 = ~n16606 & n17140 ;
  assign n17142 = x64 & n17141 ;
  assign n17143 = ~x61 & x62 ;
  assign n17144 = x61 & ~x62 ;
  assign n17145 = n17143 | n17144 ;
  assign n17146 = n16606 & ~n17145 ;
  assign n17147 = x65 & n17146 ;
  assign n17148 = n17142 | n17147 ;
  assign n17149 = n16606 & n17145 ;
  assign n17150 = x62 | n144 ;
  assign n17151 = ( x62 & n17149 ) | ( x62 & n17150 ) | ( n17149 & n17150 ) ;
  assign n17152 = ~x62 & n17151 ;
  assign n17153 = ( ~x62 & n17148 ) | ( ~x62 & n17152 ) | ( n17148 & n17152 ) ;
  assign n17154 = x62 & ~x64 ;
  assign n17155 = ( x62 & ~n16606 ) | ( x62 & n17154 ) | ( ~n16606 & n17154 ) ;
  assign n17156 = n17151 & n17155 ;
  assign n17157 = ( n17148 & n17155 ) | ( n17148 & n17156 ) | ( n17155 & n17156 ) ;
  assign n17158 = n144 & n17149 ;
  assign n17159 = n17155 & ~n17158 ;
  assign n17160 = ~n17148 & n17159 ;
  assign n17161 = ( n17153 & n17157 ) | ( n17153 & n17160 ) | ( n17157 & n17160 ) ;
  assign n17162 = n17151 | n17155 ;
  assign n17163 = n17148 | n17162 ;
  assign n17164 = ~n17155 & n17158 ;
  assign n17165 = ( n17148 & ~n17155 ) | ( n17148 & n17164 ) | ( ~n17155 & n17164 ) ;
  assign n17166 = ( n17153 & n17163 ) | ( n17153 & ~n17165 ) | ( n17163 & ~n17165 ) ;
  assign n17167 = ~n17161 & n17166 ;
  assign n17168 = n241 & n15555 ;
  assign n17169 = x68 & n15552 ;
  assign n17170 = x67 & n15547 ;
  assign n17171 = x66 & ~n15546 ;
  assign n17172 = n16123 & n17171 ;
  assign n17173 = n17170 | n17172 ;
  assign n17174 = n17169 | n17173 ;
  assign n17175 = n17168 | n17174 ;
  assign n17176 = x59 | n17169 ;
  assign n17177 = n17173 | n17176 ;
  assign n17178 = n17168 | n17177 ;
  assign n17179 = ~x59 & n17177 ;
  assign n17180 = ( ~x59 & n17168 ) | ( ~x59 & n17179 ) | ( n17168 & n17179 ) ;
  assign n17181 = ( ~n17175 & n17178 ) | ( ~n17175 & n17180 ) | ( n17178 & n17180 ) ;
  assign n17182 = n17167 | n17181 ;
  assign n17183 = n17167 & n17181 ;
  assign n17184 = n17182 & ~n17183 ;
  assign n17185 = ( n16137 & n16607 ) | ( n16137 & n16623 ) | ( n16607 & n16623 ) ;
  assign n17186 = n17184 | n17185 ;
  assign n17187 = n17184 & n17185 ;
  assign n17188 = n17186 & ~n17187 ;
  assign n17189 = n17137 | n17188 ;
  assign n17190 = n17137 & n17188 ;
  assign n17191 = n17189 & ~n17190 ;
  assign n17192 = ~n16626 & n16642 ;
  assign n17193 = n16603 & ~n17192 ;
  assign n17194 = n16626 & n16642 ;
  assign n17195 = n16626 & ~n17194 ;
  assign n17196 = ( n16603 & n17194 ) | ( n16603 & n17195 ) | ( n17194 & n17195 ) ;
  assign n17197 = n16603 | n17194 ;
  assign n17198 = ( ~n17193 & n17196 ) | ( ~n17193 & n17197 ) | ( n17196 & n17197 ) ;
  assign n17199 = n17191 & n17198 ;
  assign n17200 = n17191 | n17198 ;
  assign n17201 = ~n17199 & n17200 ;
  assign n17202 = x74 & n12574 ;
  assign n17203 = x73 & n12569 ;
  assign n17204 = x72 & ~n12568 ;
  assign n17205 = n13076 & n17204 ;
  assign n17206 = n17203 | n17205 ;
  assign n17207 = n17202 | n17206 ;
  assign n17208 = n12577 | n17202 ;
  assign n17209 = n17206 | n17208 ;
  assign n17210 = ( n710 & n17207 ) | ( n710 & n17209 ) | ( n17207 & n17209 ) ;
  assign n17211 = x53 & n17209 ;
  assign n17212 = x53 & n17202 ;
  assign n17213 = ( x53 & n17206 ) | ( x53 & n17212 ) | ( n17206 & n17212 ) ;
  assign n17214 = ( n710 & n17211 ) | ( n710 & n17213 ) | ( n17211 & n17213 ) ;
  assign n17215 = x53 & ~n17213 ;
  assign n17216 = x53 & ~n17209 ;
  assign n17217 = ( ~n710 & n17215 ) | ( ~n710 & n17216 ) | ( n17215 & n17216 ) ;
  assign n17218 = ( n17210 & ~n17214 ) | ( n17210 & n17217 ) | ( ~n17214 & n17217 ) ;
  assign n17219 = n17201 & n17218 ;
  assign n17220 = n17201 & ~n17219 ;
  assign n17221 = n16667 | n16673 ;
  assign n17222 = ( n16667 & n16675 ) | ( n16667 & n17221 ) | ( n16675 & n17221 ) ;
  assign n17223 = ~n17201 & n17218 ;
  assign n17224 = n17222 & n17223 ;
  assign n17225 = ( n17220 & n17222 ) | ( n17220 & n17224 ) | ( n17222 & n17224 ) ;
  assign n17226 = n17222 | n17223 ;
  assign n17227 = n17220 | n17226 ;
  assign n17228 = ~n17225 & n17227 ;
  assign n17229 = x77 & n11205 ;
  assign n17230 = x76 & n11200 ;
  assign n17231 = x75 & ~n11199 ;
  assign n17232 = n11679 & n17231 ;
  assign n17233 = n17230 | n17232 ;
  assign n17234 = n17229 | n17233 ;
  assign n17235 = n11208 | n17229 ;
  assign n17236 = n17233 | n17235 ;
  assign n17237 = ( n1059 & n17234 ) | ( n1059 & n17236 ) | ( n17234 & n17236 ) ;
  assign n17238 = x50 & n17236 ;
  assign n17239 = x50 & n17229 ;
  assign n17240 = ( x50 & n17233 ) | ( x50 & n17239 ) | ( n17233 & n17239 ) ;
  assign n17241 = ( n1059 & n17238 ) | ( n1059 & n17240 ) | ( n17238 & n17240 ) ;
  assign n17242 = x50 & ~n17240 ;
  assign n17243 = x50 & ~n17236 ;
  assign n17244 = ( ~n1059 & n17242 ) | ( ~n1059 & n17243 ) | ( n17242 & n17243 ) ;
  assign n17245 = ( n17237 & ~n17241 ) | ( n17237 & n17244 ) | ( ~n17241 & n17244 ) ;
  assign n17246 = n17228 & n17245 ;
  assign n17247 = n17228 | n17245 ;
  assign n17248 = ~n17246 & n17247 ;
  assign n17249 = n16697 | n16698 ;
  assign n17250 = ( n16697 & n16700 ) | ( n16697 & n17249 ) | ( n16700 & n17249 ) ;
  assign n17251 = n17248 & n17250 ;
  assign n17252 = n17250 & ~n17251 ;
  assign n17253 = ( n17248 & ~n17251 ) | ( n17248 & n17252 ) | ( ~n17251 & n17252 ) ;
  assign n17254 = x80 & n9933 ;
  assign n17255 = x79 & n9928 ;
  assign n17256 = x78 & ~n9927 ;
  assign n17257 = n10379 & n17256 ;
  assign n17258 = n17255 | n17257 ;
  assign n17259 = n17254 | n17258 ;
  assign n17260 = n9936 | n17254 ;
  assign n17261 = n17258 | n17260 ;
  assign n17262 = ( n1499 & n17259 ) | ( n1499 & n17261 ) | ( n17259 & n17261 ) ;
  assign n17263 = x47 & n17261 ;
  assign n17264 = x47 & n17254 ;
  assign n17265 = ( x47 & n17258 ) | ( x47 & n17264 ) | ( n17258 & n17264 ) ;
  assign n17266 = ( n1499 & n17263 ) | ( n1499 & n17265 ) | ( n17263 & n17265 ) ;
  assign n17267 = x47 & ~n17265 ;
  assign n17268 = x47 & ~n17261 ;
  assign n17269 = ( ~n1499 & n17267 ) | ( ~n1499 & n17268 ) | ( n17267 & n17268 ) ;
  assign n17270 = ( n17262 & ~n17266 ) | ( n17262 & n17269 ) | ( ~n17266 & n17269 ) ;
  assign n17271 = ~n17251 & n17270 ;
  assign n17272 = n17248 & n17270 ;
  assign n17273 = ( n17252 & n17271 ) | ( n17252 & n17272 ) | ( n17271 & n17272 ) ;
  assign n17274 = n17253 & ~n17273 ;
  assign n17275 = n17251 & n17270 ;
  assign n17276 = ~n17248 & n17270 ;
  assign n17277 = ( ~n17252 & n17275 ) | ( ~n17252 & n17276 ) | ( n17275 & n17276 ) ;
  assign n17278 = n17274 | n17277 ;
  assign n17279 = n16721 | n16725 ;
  assign n17280 = n17278 | n17279 ;
  assign n17281 = n17278 & n17279 ;
  assign n17282 = n17280 & ~n17281 ;
  assign n17283 = x83 & n8724 ;
  assign n17284 = x82 & n8719 ;
  assign n17285 = x81 & ~n8718 ;
  assign n17286 = n9149 & n17285 ;
  assign n17287 = n17284 | n17286 ;
  assign n17288 = n17283 | n17287 ;
  assign n17289 = n8727 | n17283 ;
  assign n17290 = n17287 | n17289 ;
  assign n17291 = ( n2009 & n17288 ) | ( n2009 & n17290 ) | ( n17288 & n17290 ) ;
  assign n17292 = x44 & n17290 ;
  assign n17293 = x44 & n17283 ;
  assign n17294 = ( x44 & n17287 ) | ( x44 & n17293 ) | ( n17287 & n17293 ) ;
  assign n17295 = ( n2009 & n17292 ) | ( n2009 & n17294 ) | ( n17292 & n17294 ) ;
  assign n17296 = x44 & ~n17294 ;
  assign n17297 = x44 & ~n17290 ;
  assign n17298 = ( ~n2009 & n17296 ) | ( ~n2009 & n17297 ) | ( n17296 & n17297 ) ;
  assign n17299 = ( n17291 & ~n17295 ) | ( n17291 & n17298 ) | ( ~n17295 & n17298 ) ;
  assign n17300 = n17282 & n17299 ;
  assign n17301 = n17282 | n17299 ;
  assign n17302 = ~n17300 & n17301 ;
  assign n17303 = n16602 & n16728 ;
  assign n17304 = n16728 & ~n17303 ;
  assign n17305 = n16602 & ~n16728 ;
  assign n17306 = n17304 | n17305 ;
  assign n17307 = n16730 & n17306 ;
  assign n17308 = n17303 | n17307 ;
  assign n17309 = n17302 & n17308 ;
  assign n17310 = n17308 & ~n17309 ;
  assign n17311 = ( n17302 & ~n17309 ) | ( n17302 & n17310 ) | ( ~n17309 & n17310 ) ;
  assign n17312 = x86 & n7566 ;
  assign n17313 = x85 & n7561 ;
  assign n17314 = x84 & ~n7560 ;
  assign n17315 = n7953 & n17314 ;
  assign n17316 = n17313 | n17315 ;
  assign n17317 = n17312 | n17316 ;
  assign n17318 = n7569 | n17312 ;
  assign n17319 = n17316 | n17318 ;
  assign n17320 = ( n2606 & n17317 ) | ( n2606 & n17319 ) | ( n17317 & n17319 ) ;
  assign n17321 = x41 & n17319 ;
  assign n17322 = x41 & n17312 ;
  assign n17323 = ( x41 & n17316 ) | ( x41 & n17322 ) | ( n17316 & n17322 ) ;
  assign n17324 = ( n2606 & n17321 ) | ( n2606 & n17323 ) | ( n17321 & n17323 ) ;
  assign n17325 = x41 & ~n17323 ;
  assign n17326 = x41 & ~n17319 ;
  assign n17327 = ( ~n2606 & n17325 ) | ( ~n2606 & n17326 ) | ( n17325 & n17326 ) ;
  assign n17328 = ( n17320 & ~n17324 ) | ( n17320 & n17327 ) | ( ~n17324 & n17327 ) ;
  assign n17329 = n17302 & n17328 ;
  assign n17330 = ~n17302 & n17328 ;
  assign n17331 = ( ~n17308 & n17328 ) | ( ~n17308 & n17330 ) | ( n17328 & n17330 ) ;
  assign n17332 = ( n17310 & n17329 ) | ( n17310 & n17331 ) | ( n17329 & n17331 ) ;
  assign n17333 = n17311 & ~n17332 ;
  assign n17334 = n17308 & n17329 ;
  assign n17335 = ( ~n17310 & n17330 ) | ( ~n17310 & n17334 ) | ( n17330 & n17334 ) ;
  assign n17336 = n17333 | n17335 ;
  assign n17337 = n16754 | n16763 ;
  assign n17338 = n17336 | n17337 ;
  assign n17339 = n17336 & n17337 ;
  assign n17340 = n17338 & ~n17339 ;
  assign n17341 = x89 & n6536 ;
  assign n17342 = x88 & n6531 ;
  assign n17343 = x87 & ~n6530 ;
  assign n17344 = n6871 & n17343 ;
  assign n17345 = n17342 | n17344 ;
  assign n17346 = n17341 | n17345 ;
  assign n17347 = n6539 | n17341 ;
  assign n17348 = n17345 | n17347 ;
  assign n17349 = ( n3282 & n17346 ) | ( n3282 & n17348 ) | ( n17346 & n17348 ) ;
  assign n17350 = x38 & n17348 ;
  assign n17351 = x38 & n17341 ;
  assign n17352 = ( x38 & n17345 ) | ( x38 & n17351 ) | ( n17345 & n17351 ) ;
  assign n17353 = ( n3282 & n17350 ) | ( n3282 & n17352 ) | ( n17350 & n17352 ) ;
  assign n17354 = x38 & ~n17352 ;
  assign n17355 = x38 & ~n17348 ;
  assign n17356 = ( ~n3282 & n17354 ) | ( ~n3282 & n17355 ) | ( n17354 & n17355 ) ;
  assign n17357 = ( n17349 & ~n17353 ) | ( n17349 & n17356 ) | ( ~n17353 & n17356 ) ;
  assign n17358 = n17340 & n17357 ;
  assign n17359 = n17340 & ~n17358 ;
  assign n17360 = ~n17340 & n17357 ;
  assign n17361 = n17359 | n17360 ;
  assign n17362 = n16788 | n16790 ;
  assign n17363 = n16789 | n17362 ;
  assign n17364 = ( n16788 & n16792 ) | ( n16788 & n17363 ) | ( n16792 & n17363 ) ;
  assign n17365 = n17361 | n17364 ;
  assign n17366 = n17361 & n17364 ;
  assign n17367 = n17365 & ~n17366 ;
  assign n17368 = x92 & n5554 ;
  assign n17369 = x91 & n5549 ;
  assign n17370 = x90 & ~n5548 ;
  assign n17371 = n5893 & n17370 ;
  assign n17372 = n17369 | n17371 ;
  assign n17373 = n17368 | n17372 ;
  assign n17374 = n5557 | n17368 ;
  assign n17375 = n17372 | n17374 ;
  assign n17376 = ( n4040 & n17373 ) | ( n4040 & n17375 ) | ( n17373 & n17375 ) ;
  assign n17377 = x35 & n17375 ;
  assign n17378 = x35 & n17368 ;
  assign n17379 = ( x35 & n17372 ) | ( x35 & n17378 ) | ( n17372 & n17378 ) ;
  assign n17380 = ( n4040 & n17377 ) | ( n4040 & n17379 ) | ( n17377 & n17379 ) ;
  assign n17381 = x35 & ~n17379 ;
  assign n17382 = x35 & ~n17375 ;
  assign n17383 = ( ~n4040 & n17381 ) | ( ~n4040 & n17382 ) | ( n17381 & n17382 ) ;
  assign n17384 = ( n17376 & ~n17380 ) | ( n17376 & n17383 ) | ( ~n17380 & n17383 ) ;
  assign n17385 = n17367 & n17384 ;
  assign n17386 = n17367 & ~n17385 ;
  assign n17387 = ~n17367 & n17384 ;
  assign n17388 = n17386 | n17387 ;
  assign n17389 = n16813 | n16819 ;
  assign n17390 = ( n16813 & n16816 ) | ( n16813 & n17389 ) | ( n16816 & n17389 ) ;
  assign n17391 = n17388 | n17390 ;
  assign n17392 = n17388 & n17390 ;
  assign n17393 = n17391 & ~n17392 ;
  assign n17394 = x95 & n4631 ;
  assign n17395 = x94 & n4626 ;
  assign n17396 = x93 & ~n4625 ;
  assign n17397 = n4943 & n17396 ;
  assign n17398 = n17395 | n17397 ;
  assign n17399 = n17394 | n17398 ;
  assign n17400 = n4634 | n17394 ;
  assign n17401 = n17398 | n17400 ;
  assign n17402 = ( n4897 & n17399 ) | ( n4897 & n17401 ) | ( n17399 & n17401 ) ;
  assign n17403 = x32 & n17401 ;
  assign n17404 = x32 & n17394 ;
  assign n17405 = ( x32 & n17398 ) | ( x32 & n17404 ) | ( n17398 & n17404 ) ;
  assign n17406 = ( n4897 & n17403 ) | ( n4897 & n17405 ) | ( n17403 & n17405 ) ;
  assign n17407 = x32 & ~n17405 ;
  assign n17408 = x32 & ~n17401 ;
  assign n17409 = ( ~n4897 & n17407 ) | ( ~n4897 & n17408 ) | ( n17407 & n17408 ) ;
  assign n17410 = ( n17402 & ~n17406 ) | ( n17402 & n17409 ) | ( ~n17406 & n17409 ) ;
  assign n17411 = n17393 & n17410 ;
  assign n17412 = n17393 & ~n17411 ;
  assign n17413 = ~n17393 & n17410 ;
  assign n17414 = n17412 | n17413 ;
  assign n17415 = n16841 | n16845 ;
  assign n17416 = ~n17414 & n17415 ;
  assign n17417 = n17414 & ~n17415 ;
  assign n17418 = n17416 | n17417 ;
  assign n17419 = x98 & n3816 ;
  assign n17420 = x97 & n3811 ;
  assign n17421 = x96 & ~n3810 ;
  assign n17422 = n4067 & n17421 ;
  assign n17423 = n17420 | n17422 ;
  assign n17424 = n17419 | n17423 ;
  assign n17425 = n3819 | n17419 ;
  assign n17426 = n17423 | n17425 ;
  assign n17427 = ( ~n5850 & n17424 ) | ( ~n5850 & n17426 ) | ( n17424 & n17426 ) ;
  assign n17428 = n17424 & n17426 ;
  assign n17429 = ( n5834 & n17427 ) | ( n5834 & n17428 ) | ( n17427 & n17428 ) ;
  assign n17430 = x29 & n17426 ;
  assign n17431 = x29 & n17419 ;
  assign n17432 = ( x29 & n17423 ) | ( x29 & n17431 ) | ( n17423 & n17431 ) ;
  assign n17433 = ( ~n5850 & n17430 ) | ( ~n5850 & n17432 ) | ( n17430 & n17432 ) ;
  assign n17434 = n17430 & n17432 ;
  assign n17435 = ( n5834 & n17433 ) | ( n5834 & n17434 ) | ( n17433 & n17434 ) ;
  assign n17436 = x29 & ~n17432 ;
  assign n17437 = x29 & ~n17426 ;
  assign n17438 = ( n5850 & n17436 ) | ( n5850 & n17437 ) | ( n17436 & n17437 ) ;
  assign n17439 = n17436 | n17437 ;
  assign n17440 = ( ~n5834 & n17438 ) | ( ~n5834 & n17439 ) | ( n17438 & n17439 ) ;
  assign n17441 = ( n17429 & ~n17435 ) | ( n17429 & n17440 ) | ( ~n17435 & n17440 ) ;
  assign n17442 = n17418 & n17441 ;
  assign n17443 = n17418 | n17441 ;
  assign n17444 = ~n17442 & n17443 ;
  assign n17445 = ( n16847 & n16864 ) | ( n16847 & n16870 ) | ( n16864 & n16870 ) ;
  assign n17446 = ( n16372 & n16847 ) | ( n16372 & n16864 ) | ( n16847 & n16864 ) ;
  assign n17447 = ( n16869 & n17445 ) | ( n16869 & n17446 ) | ( n17445 & n17446 ) ;
  assign n17448 = n17444 | n17447 ;
  assign n17449 = n17444 & n17447 ;
  assign n17450 = n17448 & ~n17449 ;
  assign n17451 = x101 & n3085 ;
  assign n17452 = x100 & n3080 ;
  assign n17453 = x99 & ~n3079 ;
  assign n17454 = n3309 & n17453 ;
  assign n17455 = n17452 | n17454 ;
  assign n17456 = n17451 | n17455 ;
  assign n17457 = n3088 | n17451 ;
  assign n17458 = n17455 | n17457 ;
  assign n17459 = ( n6844 & n17456 ) | ( n6844 & n17458 ) | ( n17456 & n17458 ) ;
  assign n17460 = x26 & n17458 ;
  assign n17461 = x26 & n17451 ;
  assign n17462 = ( x26 & n17455 ) | ( x26 & n17461 ) | ( n17455 & n17461 ) ;
  assign n17463 = ( n6844 & n17460 ) | ( n6844 & n17462 ) | ( n17460 & n17462 ) ;
  assign n17464 = x26 & ~n17462 ;
  assign n17465 = x26 & ~n17458 ;
  assign n17466 = ( ~n6844 & n17464 ) | ( ~n6844 & n17465 ) | ( n17464 & n17465 ) ;
  assign n17467 = ( n17459 & ~n17463 ) | ( n17459 & n17466 ) | ( ~n17463 & n17466 ) ;
  assign n17468 = n17450 & n17467 ;
  assign n17469 = n17450 & ~n17468 ;
  assign n17470 = ~n17450 & n17467 ;
  assign n17471 = n17469 | n17470 ;
  assign n17472 = n16892 | n16896 ;
  assign n17473 = n17471 | n17472 ;
  assign n17474 = n17471 & n17472 ;
  assign n17475 = n17473 & ~n17474 ;
  assign n17476 = x104 & n2429 ;
  assign n17477 = x103 & n2424 ;
  assign n17478 = x102 & ~n2423 ;
  assign n17479 = n2631 & n17478 ;
  assign n17480 = n17477 | n17479 ;
  assign n17481 = n17476 | n17480 ;
  assign n17482 = n2432 | n17476 ;
  assign n17483 = n17480 | n17482 ;
  assign n17484 = ( n7911 & n17481 ) | ( n7911 & n17483 ) | ( n17481 & n17483 ) ;
  assign n17485 = x23 & n17483 ;
  assign n17486 = x23 & n17476 ;
  assign n17487 = ( x23 & n17480 ) | ( x23 & n17486 ) | ( n17480 & n17486 ) ;
  assign n17488 = ( n7911 & n17485 ) | ( n7911 & n17487 ) | ( n17485 & n17487 ) ;
  assign n17489 = x23 & ~n17487 ;
  assign n17490 = x23 & ~n17483 ;
  assign n17491 = ( ~n7911 & n17489 ) | ( ~n7911 & n17490 ) | ( n17489 & n17490 ) ;
  assign n17492 = ( n17484 & ~n17488 ) | ( n17484 & n17491 ) | ( ~n17488 & n17491 ) ;
  assign n17493 = n17475 & n17492 ;
  assign n17494 = n17475 & ~n17493 ;
  assign n17495 = ~n17475 & n17492 ;
  assign n17496 = n17494 | n17495 ;
  assign n17497 = n16917 | n16919 ;
  assign n17498 = n16918 | n17497 ;
  assign n17499 = ( n16917 & n16921 ) | ( n16917 & n17498 ) | ( n16921 & n17498 ) ;
  assign n17500 = n17496 | n17499 ;
  assign n17501 = n17496 & n17499 ;
  assign n17502 = n17500 & ~n17501 ;
  assign n17503 = x107 & n1859 ;
  assign n17504 = x106 & n1854 ;
  assign n17505 = x105 & ~n1853 ;
  assign n17506 = n2037 & n17505 ;
  assign n17507 = n17504 | n17506 ;
  assign n17508 = n17503 | n17507 ;
  assign n17509 = n1862 | n17503 ;
  assign n17510 = n17507 | n17509 ;
  assign n17511 = ( n9084 & n17508 ) | ( n9084 & n17510 ) | ( n17508 & n17510 ) ;
  assign n17512 = x20 & n17510 ;
  assign n17513 = x20 & n17503 ;
  assign n17514 = ( x20 & n17507 ) | ( x20 & n17513 ) | ( n17507 & n17513 ) ;
  assign n17515 = ( n9084 & n17512 ) | ( n9084 & n17514 ) | ( n17512 & n17514 ) ;
  assign n17516 = x20 & ~n17514 ;
  assign n17517 = x20 & ~n17510 ;
  assign n17518 = ( ~n9084 & n17516 ) | ( ~n9084 & n17517 ) | ( n17516 & n17517 ) ;
  assign n17519 = ( n17511 & ~n17515 ) | ( n17511 & n17518 ) | ( ~n17515 & n17518 ) ;
  assign n17520 = n17502 & n17519 ;
  assign n17521 = n17502 | n17519 ;
  assign n17522 = ~n17520 & n17521 ;
  assign n17525 = n17522 & n17524 ;
  assign n17526 = n17524 & ~n17525 ;
  assign n17527 = x110 & n1383 ;
  assign n17528 = x109 & n1378 ;
  assign n17529 = x108 & ~n1377 ;
  assign n17530 = n1542 & n17529 ;
  assign n17531 = n17528 | n17530 ;
  assign n17532 = n17527 | n17531 ;
  assign n17533 = n1386 | n17527 ;
  assign n17534 = n17531 | n17533 ;
  assign n17535 = ( n10330 & n17532 ) | ( n10330 & n17534 ) | ( n17532 & n17534 ) ;
  assign n17536 = x17 & n17534 ;
  assign n17537 = x17 & n17527 ;
  assign n17538 = ( x17 & n17531 ) | ( x17 & n17537 ) | ( n17531 & n17537 ) ;
  assign n17539 = ( n10330 & n17536 ) | ( n10330 & n17538 ) | ( n17536 & n17538 ) ;
  assign n17540 = x17 & ~n17538 ;
  assign n17541 = x17 & ~n17534 ;
  assign n17542 = ( ~n10330 & n17540 ) | ( ~n10330 & n17541 ) | ( n17540 & n17541 ) ;
  assign n17543 = ( n17535 & ~n17539 ) | ( n17535 & n17542 ) | ( ~n17539 & n17542 ) ;
  assign n17544 = n17522 & n17543 ;
  assign n17545 = ~n17522 & n17543 ;
  assign n17546 = ( ~n17524 & n17543 ) | ( ~n17524 & n17545 ) | ( n17543 & n17545 ) ;
  assign n17547 = ( n17526 & n17544 ) | ( n17526 & n17546 ) | ( n17544 & n17546 ) ;
  assign n17548 = n17522 | n17543 ;
  assign n17549 = n17522 & ~n17543 ;
  assign n17550 = n17524 & n17549 ;
  assign n17551 = ( n17526 & n17548 ) | ( n17526 & ~n17550 ) | ( n17548 & ~n17550 ) ;
  assign n17552 = ~n17547 & n17551 ;
  assign n17553 = n17121 & n17552 ;
  assign n17554 = n17121 | n17552 ;
  assign n17555 = ~n17553 & n17554 ;
  assign n17556 = x113 & n962 ;
  assign n17557 = x112 & n957 ;
  assign n17558 = x111 & ~n956 ;
  assign n17559 = n1105 & n17558 ;
  assign n17560 = n17557 | n17559 ;
  assign n17561 = n17556 | n17560 ;
  assign n17562 = n965 | n17556 ;
  assign n17563 = n17560 | n17562 ;
  assign n17564 = ( ~n11642 & n17561 ) | ( ~n11642 & n17563 ) | ( n17561 & n17563 ) ;
  assign n17565 = n17561 & n17563 ;
  assign n17566 = ( n11626 & n17564 ) | ( n11626 & n17565 ) | ( n17564 & n17565 ) ;
  assign n17567 = x14 & n17566 ;
  assign n17568 = x14 & ~n17566 ;
  assign n17569 = ( n17566 & ~n17567 ) | ( n17566 & n17568 ) | ( ~n17567 & n17568 ) ;
  assign n17570 = n17555 | n17569 ;
  assign n17571 = n17555 & n17569 ;
  assign n17572 = n17570 & ~n17571 ;
  assign n17573 = n17120 & n17572 ;
  assign n17574 = n17120 | n17572 ;
  assign n17575 = ~n17573 & n17574 ;
  assign n17576 = x116 & n636 ;
  assign n17577 = x115 & n631 ;
  assign n17578 = x114 & ~n630 ;
  assign n17579 = n764 & n17578 ;
  assign n17580 = n17577 | n17579 ;
  assign n17581 = n17576 | n17580 ;
  assign n17582 = n639 | n17576 ;
  assign n17583 = n17580 | n17582 ;
  assign n17584 = ( ~n13040 & n17581 ) | ( ~n13040 & n17583 ) | ( n17581 & n17583 ) ;
  assign n17585 = n17581 & n17583 ;
  assign n17586 = ( n13022 & n17584 ) | ( n13022 & n17585 ) | ( n17584 & n17585 ) ;
  assign n17587 = x11 & n17586 ;
  assign n17588 = x11 & ~n17586 ;
  assign n17589 = ( n17586 & ~n17587 ) | ( n17586 & n17588 ) | ( ~n17587 & n17588 ) ;
  assign n17590 = n17575 | n17589 ;
  assign n17591 = n17575 & n17589 ;
  assign n17592 = n17590 & ~n17591 ;
  assign n17593 = n17016 | n17018 ;
  assign n17594 = n17017 | n17593 ;
  assign n17595 = ( n16584 & n17016 ) | ( n16584 & n17594 ) | ( n17016 & n17594 ) ;
  assign n17596 = n17592 & n17595 ;
  assign n17597 = n17592 | n17595 ;
  assign n17598 = ~n17596 & n17597 ;
  assign n17599 = x119 & n389 ;
  assign n17600 = x118 & n384 ;
  assign n17601 = x117 & ~n383 ;
  assign n17602 = n463 & n17601 ;
  assign n17603 = n17600 | n17602 ;
  assign n17604 = n17599 | n17603 ;
  assign n17605 = n392 | n17599 ;
  assign n17606 = n17603 | n17605 ;
  assign n17607 = ( n14496 & n17604 ) | ( n14496 & n17606 ) | ( n17604 & n17606 ) ;
  assign n17608 = x8 & n17606 ;
  assign n17609 = x8 & n17599 ;
  assign n17610 = ( x8 & n17603 ) | ( x8 & n17609 ) | ( n17603 & n17609 ) ;
  assign n17611 = ( n14496 & n17608 ) | ( n14496 & n17610 ) | ( n17608 & n17610 ) ;
  assign n17612 = x8 & ~n17610 ;
  assign n17613 = x8 & ~n17606 ;
  assign n17614 = ( ~n14496 & n17612 ) | ( ~n14496 & n17613 ) | ( n17612 & n17613 ) ;
  assign n17615 = ( n17607 & ~n17611 ) | ( n17607 & n17614 ) | ( ~n17611 & n17614 ) ;
  assign n17616 = n17598 & n17615 ;
  assign n17617 = n17598 & ~n17616 ;
  assign n17618 = ~n17598 & n17615 ;
  assign n17619 = n17617 | n17618 ;
  assign n17620 = n17037 | n17039 ;
  assign n17621 = ( n16583 & n17037 ) | ( n16583 & n17620 ) | ( n17037 & n17620 ) ;
  assign n17622 = n17619 | n17621 ;
  assign n17623 = n17619 & n17621 ;
  assign n17624 = n17622 & ~n17623 ;
  assign n17625 = x122 & n212 ;
  assign n17626 = x121 & n207 ;
  assign n17627 = x120 & ~n206 ;
  assign n17628 = n267 & n17627 ;
  assign n17629 = n17626 | n17628 ;
  assign n17630 = n17625 | n17629 ;
  assign n17631 = n215 | n17625 ;
  assign n17632 = n17629 | n17631 ;
  assign n17633 = ( n16043 & n17630 ) | ( n16043 & n17632 ) | ( n17630 & n17632 ) ;
  assign n17634 = x5 & n17632 ;
  assign n17635 = x5 & n17625 ;
  assign n17636 = ( x5 & n17629 ) | ( x5 & n17635 ) | ( n17629 & n17635 ) ;
  assign n17637 = ( n16043 & n17634 ) | ( n16043 & n17636 ) | ( n17634 & n17636 ) ;
  assign n17638 = x5 & ~n17636 ;
  assign n17639 = x5 & ~n17632 ;
  assign n17640 = ( ~n16043 & n17638 ) | ( ~n16043 & n17639 ) | ( n17638 & n17639 ) ;
  assign n17641 = ( n17633 & ~n17637 ) | ( n17633 & n17640 ) | ( ~n17637 & n17640 ) ;
  assign n17642 = n17624 | n17641 ;
  assign n17643 = n17624 & n17641 ;
  assign n17644 = n17642 & ~n17643 ;
  assign n17645 = x124 | x125 ;
  assign n17646 = x124 & x125 ;
  assign n17647 = n17645 & ~n17646 ;
  assign n17648 = n16069 | n17064 ;
  assign n17649 = ( n17064 & n17065 ) | ( n17064 & n17648 ) | ( n17065 & n17648 ) ;
  assign n17650 = n17647 & n17649 ;
  assign n17651 = n17064 | n17065 ;
  assign n17652 = n17647 & n17651 ;
  assign n17653 = ( n16075 & n17650 ) | ( n16075 & n17652 ) | ( n17650 & n17652 ) ;
  assign n17654 = n17064 & n17647 ;
  assign n17655 = ( n17070 & n17647 ) | ( n17070 & n17654 ) | ( n17647 & n17654 ) ;
  assign n17656 = ( n17068 & n17647 ) | ( n17068 & n17654 ) | ( n17647 & n17654 ) ;
  assign n17657 = ( n16033 & n17655 ) | ( n16033 & n17656 ) | ( n17655 & n17656 ) ;
  assign n17658 = ( n13965 & n17653 ) | ( n13965 & n17657 ) | ( n17653 & n17657 ) ;
  assign n17659 = n17653 | n17657 ;
  assign n17660 = ( n14002 & n17658 ) | ( n14002 & n17659 ) | ( n17658 & n17659 ) ;
  assign n17661 = ( n16075 & n17649 ) | ( n16075 & n17651 ) | ( n17649 & n17651 ) ;
  assign n17662 = n17064 | n17070 ;
  assign n17663 = n17064 | n17068 ;
  assign n17664 = ( n16033 & n17662 ) | ( n16033 & n17663 ) | ( n17662 & n17663 ) ;
  assign n17665 = n17661 | n17664 ;
  assign n17666 = n17647 | n17665 ;
  assign n17667 = ( n13965 & n17661 ) | ( n13965 & n17664 ) | ( n17661 & n17664 ) ;
  assign n17668 = n17647 | n17667 ;
  assign n17669 = ( n14002 & n17666 ) | ( n14002 & n17668 ) | ( n17666 & n17668 ) ;
  assign n17670 = ~n17660 & n17669 ;
  assign n17671 = x124 & n133 ;
  assign n17672 = x123 & ~n162 ;
  assign n17673 = ( n137 & n17671 ) | ( n137 & n17672 ) | ( n17671 & n17672 ) ;
  assign n17674 = x0 & x125 ;
  assign n17675 = ( ~n137 & n17671 ) | ( ~n137 & n17674 ) | ( n17671 & n17674 ) ;
  assign n17676 = n17673 | n17675 ;
  assign n17677 = n141 | n17676 ;
  assign n17678 = ( n17670 & n17676 ) | ( n17670 & n17677 ) | ( n17676 & n17677 ) ;
  assign n17679 = x2 & n17676 ;
  assign n17680 = ( x2 & n523 ) | ( x2 & n17676 ) | ( n523 & n17676 ) ;
  assign n17681 = ( n17670 & n17679 ) | ( n17670 & n17680 ) | ( n17679 & n17680 ) ;
  assign n17682 = x2 & ~n17680 ;
  assign n17683 = x2 & ~n17676 ;
  assign n17684 = ( ~n17670 & n17682 ) | ( ~n17670 & n17683 ) | ( n17682 & n17683 ) ;
  assign n17685 = ( n17678 & ~n17681 ) | ( n17678 & n17684 ) | ( ~n17681 & n17684 ) ;
  assign n17686 = ~n17644 & n17685 ;
  assign n17687 = n17059 | n17099 ;
  assign n17688 = ( n17042 & n17099 ) | ( n17042 & n17687 ) | ( n17099 & n17687 ) ;
  assign n17689 = ( n17060 & n17062 ) | ( n17060 & n17688 ) | ( n17062 & n17688 ) ;
  assign n17690 = n17641 | n17685 ;
  assign n17691 = ( n17624 & n17685 ) | ( n17624 & n17690 ) | ( n17685 & n17690 ) ;
  assign n17692 = n17642 & ~n17691 ;
  assign n17693 = n17689 & n17692 ;
  assign n17694 = ( n17686 & n17689 ) | ( n17686 & n17693 ) | ( n17689 & n17693 ) ;
  assign n17695 = n17689 | n17692 ;
  assign n17696 = n17686 | n17695 ;
  assign n17697 = ~n17694 & n17696 ;
  assign n17698 = n17111 | n17113 ;
  assign n17699 = ( n17111 & n17116 ) | ( n17111 & n17698 ) | ( n17116 & n17698 ) ;
  assign n17700 = n17697 & n17699 ;
  assign n17701 = n17697 | n17699 ;
  assign n17702 = ~n17700 & n17701 ;
  assign n17703 = n17616 | n17623 ;
  assign n17704 = n17493 | n17501 ;
  assign n17705 = n17246 | n17251 ;
  assign n17706 = x72 & n14045 ;
  assign n17707 = x71 & n14040 ;
  assign n17708 = x70 & ~n14039 ;
  assign n17709 = n14552 & n17708 ;
  assign n17710 = n17707 | n17709 ;
  assign n17711 = n17706 | n17710 ;
  assign n17712 = ( n513 & n14048 ) | ( n513 & n17711 ) | ( n14048 & n17711 ) ;
  assign n17713 = x56 & n14048 ;
  assign n17714 = ( x56 & n14048 ) | ( x56 & ~n17706 ) | ( n14048 & ~n17706 ) ;
  assign n17715 = ( ~n17710 & n17713 ) | ( ~n17710 & n17714 ) | ( n17713 & n17714 ) ;
  assign n17716 = ( x56 & n513 ) | ( x56 & n17715 ) | ( n513 & n17715 ) ;
  assign n17717 = ~n17712 & n17716 ;
  assign n17718 = n17711 | n17715 ;
  assign n17719 = x56 | n17711 ;
  assign n17720 = ( n513 & n17718 ) | ( n513 & n17719 ) | ( n17718 & n17719 ) ;
  assign n17721 = ( ~x56 & n17717 ) | ( ~x56 & n17720 ) | ( n17717 & n17720 ) ;
  assign n17722 = x66 & n17146 ;
  assign n17723 = x65 & n17141 ;
  assign n17724 = ~n16606 & n17145 ;
  assign n17725 = x64 & ~n17140 ;
  assign n17726 = n17724 & n17725 ;
  assign n17727 = n17723 | n17726 ;
  assign n17728 = n17722 | n17727 ;
  assign n17729 = n159 & n17149 ;
  assign n17730 = n17728 | n17729 ;
  assign n17731 = x62 | n17149 ;
  assign n17732 = ( x62 & n159 ) | ( x62 & n17731 ) | ( n159 & n17731 ) ;
  assign n17733 = n17728 | n17732 ;
  assign n17734 = ~x62 & n17732 ;
  assign n17735 = ( ~x62 & n17728 ) | ( ~x62 & n17734 ) | ( n17728 & n17734 ) ;
  assign n17736 = ( ~n17730 & n17733 ) | ( ~n17730 & n17735 ) | ( n17733 & n17735 ) ;
  assign n17737 = n17161 | n17736 ;
  assign n17738 = n17161 & n17736 ;
  assign n17739 = n17737 & ~n17738 ;
  assign n17740 = n293 & n15555 ;
  assign n17741 = x69 & n15552 ;
  assign n17742 = x68 & n15547 ;
  assign n17743 = x67 & ~n15546 ;
  assign n17744 = n16123 & n17743 ;
  assign n17745 = n17742 | n17744 ;
  assign n17746 = n17741 | n17745 ;
  assign n17747 = n17740 | n17746 ;
  assign n17748 = x59 | n17741 ;
  assign n17749 = n17745 | n17748 ;
  assign n17750 = n17740 | n17749 ;
  assign n17751 = ~x59 & n17749 ;
  assign n17752 = ( ~x59 & n17740 ) | ( ~x59 & n17751 ) | ( n17740 & n17751 ) ;
  assign n17753 = ( ~n17747 & n17750 ) | ( ~n17747 & n17752 ) | ( n17750 & n17752 ) ;
  assign n17754 = n17739 | n17753 ;
  assign n17755 = n17739 & n17753 ;
  assign n17756 = n17754 & ~n17755 ;
  assign n17757 = n17183 | n17185 ;
  assign n17758 = ( n17183 & n17184 ) | ( n17183 & n17757 ) | ( n17184 & n17757 ) ;
  assign n17759 = n17756 & n17758 ;
  assign n17760 = n17756 & ~n17759 ;
  assign n17761 = ~n17756 & n17758 ;
  assign n17762 = n17721 & n17761 ;
  assign n17763 = ( n17721 & n17760 ) | ( n17721 & n17762 ) | ( n17760 & n17762 ) ;
  assign n17764 = n17721 | n17761 ;
  assign n17765 = n17760 | n17764 ;
  assign n17766 = ~n17763 & n17765 ;
  assign n17767 = n17190 | n17191 ;
  assign n17768 = ( n17190 & n17198 ) | ( n17190 & n17767 ) | ( n17198 & n17767 ) ;
  assign n17769 = n17766 & n17768 ;
  assign n17770 = n17766 | n17768 ;
  assign n17771 = ~n17769 & n17770 ;
  assign n17772 = x75 & n12574 ;
  assign n17773 = x74 & n12569 ;
  assign n17774 = x73 & ~n12568 ;
  assign n17775 = n13076 & n17774 ;
  assign n17776 = n17773 | n17775 ;
  assign n17777 = n17772 | n17776 ;
  assign n17778 = n12577 | n17772 ;
  assign n17779 = n17776 | n17778 ;
  assign n17780 = ( n746 & n17777 ) | ( n746 & n17779 ) | ( n17777 & n17779 ) ;
  assign n17781 = x53 & n17779 ;
  assign n17782 = x53 & n17772 ;
  assign n17783 = ( x53 & n17776 ) | ( x53 & n17782 ) | ( n17776 & n17782 ) ;
  assign n17784 = ( n746 & n17781 ) | ( n746 & n17783 ) | ( n17781 & n17783 ) ;
  assign n17785 = x53 & ~n17783 ;
  assign n17786 = x53 & ~n17779 ;
  assign n17787 = ( ~n746 & n17785 ) | ( ~n746 & n17786 ) | ( n17785 & n17786 ) ;
  assign n17788 = ( n17780 & ~n17784 ) | ( n17780 & n17787 ) | ( ~n17784 & n17787 ) ;
  assign n17789 = n17771 | n17788 ;
  assign n17790 = n17771 & n17788 ;
  assign n17791 = n17789 & ~n17790 ;
  assign n17792 = n17219 | n17225 ;
  assign n17793 = n17791 & n17792 ;
  assign n17794 = n17791 | n17792 ;
  assign n17795 = ~n17793 & n17794 ;
  assign n17796 = x78 & n11205 ;
  assign n17797 = x77 & n11200 ;
  assign n17798 = x76 & ~n11199 ;
  assign n17799 = n11679 & n17798 ;
  assign n17800 = n17797 | n17799 ;
  assign n17801 = n17796 | n17800 ;
  assign n17802 = n11208 | n17796 ;
  assign n17803 = n17800 | n17802 ;
  assign n17804 = ( n1192 & n17801 ) | ( n1192 & n17803 ) | ( n17801 & n17803 ) ;
  assign n17805 = x50 & n17803 ;
  assign n17806 = x50 & n17796 ;
  assign n17807 = ( x50 & n17800 ) | ( x50 & n17806 ) | ( n17800 & n17806 ) ;
  assign n17808 = ( n1192 & n17805 ) | ( n1192 & n17807 ) | ( n17805 & n17807 ) ;
  assign n17809 = x50 & ~n17807 ;
  assign n17810 = x50 & ~n17803 ;
  assign n17811 = ( ~n1192 & n17809 ) | ( ~n1192 & n17810 ) | ( n17809 & n17810 ) ;
  assign n17812 = ( n17804 & ~n17808 ) | ( n17804 & n17811 ) | ( ~n17808 & n17811 ) ;
  assign n17813 = n17795 & n17812 ;
  assign n17814 = n17795 & ~n17813 ;
  assign n17815 = ~n17795 & n17812 ;
  assign n17816 = n17814 | n17815 ;
  assign n17817 = n17705 & n17816 ;
  assign n17818 = n17705 | n17816 ;
  assign n17819 = ~n17817 & n17818 ;
  assign n17820 = x81 & n9933 ;
  assign n17821 = x80 & n9928 ;
  assign n17822 = x79 & ~n9927 ;
  assign n17823 = n10379 & n17822 ;
  assign n17824 = n17821 | n17823 ;
  assign n17825 = n17820 | n17824 ;
  assign n17826 = n9936 | n17820 ;
  assign n17827 = n17824 | n17826 ;
  assign n17828 = ( n1651 & n17825 ) | ( n1651 & n17827 ) | ( n17825 & n17827 ) ;
  assign n17829 = x47 & n17827 ;
  assign n17830 = x47 & n17820 ;
  assign n17831 = ( x47 & n17824 ) | ( x47 & n17830 ) | ( n17824 & n17830 ) ;
  assign n17832 = ( n1651 & n17829 ) | ( n1651 & n17831 ) | ( n17829 & n17831 ) ;
  assign n17833 = x47 & ~n17831 ;
  assign n17834 = x47 & ~n17827 ;
  assign n17835 = ( ~n1651 & n17833 ) | ( ~n1651 & n17834 ) | ( n17833 & n17834 ) ;
  assign n17836 = ( n17828 & ~n17832 ) | ( n17828 & n17835 ) | ( ~n17832 & n17835 ) ;
  assign n17837 = n17819 & n17836 ;
  assign n17838 = n17819 & ~n17837 ;
  assign n17839 = ~n17819 & n17836 ;
  assign n17840 = n17838 | n17839 ;
  assign n17841 = n17273 | n17277 ;
  assign n17842 = n17274 | n17841 ;
  assign n17843 = ( n17273 & n17279 ) | ( n17273 & n17842 ) | ( n17279 & n17842 ) ;
  assign n17844 = n17840 & n17843 ;
  assign n17845 = n17840 & ~n17844 ;
  assign n17846 = ~n17840 & n17843 ;
  assign n17847 = n17845 | n17846 ;
  assign n17848 = x84 & n8724 ;
  assign n17849 = x83 & n8719 ;
  assign n17850 = x82 & ~n8718 ;
  assign n17851 = n9149 & n17850 ;
  assign n17852 = n17849 | n17851 ;
  assign n17853 = n17848 | n17852 ;
  assign n17854 = n8727 | n17848 ;
  assign n17855 = n17852 | n17854 ;
  assign n17856 = ( n2194 & n17853 ) | ( n2194 & n17855 ) | ( n17853 & n17855 ) ;
  assign n17857 = x44 & n17855 ;
  assign n17858 = x44 & n17848 ;
  assign n17859 = ( x44 & n17852 ) | ( x44 & n17858 ) | ( n17852 & n17858 ) ;
  assign n17860 = ( n2194 & n17857 ) | ( n2194 & n17859 ) | ( n17857 & n17859 ) ;
  assign n17861 = x44 & ~n17859 ;
  assign n17862 = x44 & ~n17855 ;
  assign n17863 = ( ~n2194 & n17861 ) | ( ~n2194 & n17862 ) | ( n17861 & n17862 ) ;
  assign n17864 = ( n17856 & ~n17860 ) | ( n17856 & n17863 ) | ( ~n17860 & n17863 ) ;
  assign n17865 = n17843 & n17864 ;
  assign n17866 = ~n17840 & n17865 ;
  assign n17867 = ( n17845 & n17864 ) | ( n17845 & n17866 ) | ( n17864 & n17866 ) ;
  assign n17868 = n17847 & ~n17867 ;
  assign n17869 = ~n17843 & n17864 ;
  assign n17870 = ( n17840 & n17864 ) | ( n17840 & n17869 ) | ( n17864 & n17869 ) ;
  assign n17871 = ~n17845 & n17870 ;
  assign n17872 = n17868 | n17871 ;
  assign n17873 = n17300 | n17302 ;
  assign n17874 = ( n17300 & n17308 ) | ( n17300 & n17873 ) | ( n17308 & n17873 ) ;
  assign n17875 = ~n17872 & n17874 ;
  assign n17876 = n17872 & ~n17874 ;
  assign n17877 = n17875 | n17876 ;
  assign n17878 = x87 & n7566 ;
  assign n17879 = x86 & n7561 ;
  assign n17880 = x85 & ~n7560 ;
  assign n17881 = n7953 & n17880 ;
  assign n17882 = n17879 | n17881 ;
  assign n17883 = n17878 | n17882 ;
  assign n17884 = n7569 | n17878 ;
  assign n17885 = n17882 | n17884 ;
  assign n17886 = ( n2816 & n17883 ) | ( n2816 & n17885 ) | ( n17883 & n17885 ) ;
  assign n17887 = x41 & n17885 ;
  assign n17888 = x41 & n17878 ;
  assign n17889 = ( x41 & n17882 ) | ( x41 & n17888 ) | ( n17882 & n17888 ) ;
  assign n17890 = ( n2816 & n17887 ) | ( n2816 & n17889 ) | ( n17887 & n17889 ) ;
  assign n17891 = x41 & ~n17889 ;
  assign n17892 = x41 & ~n17885 ;
  assign n17893 = ( ~n2816 & n17891 ) | ( ~n2816 & n17892 ) | ( n17891 & n17892 ) ;
  assign n17894 = ( n17886 & ~n17890 ) | ( n17886 & n17893 ) | ( ~n17890 & n17893 ) ;
  assign n17895 = n17877 & n17894 ;
  assign n17896 = n17877 | n17894 ;
  assign n17897 = ~n17895 & n17896 ;
  assign n17898 = n17332 | n17337 ;
  assign n17899 = ( n17332 & n17336 ) | ( n17332 & n17898 ) | ( n17336 & n17898 ) ;
  assign n17900 = n17897 | n17899 ;
  assign n17901 = n17897 & n17899 ;
  assign n17902 = n17900 & ~n17901 ;
  assign n17903 = x90 & n6536 ;
  assign n17904 = x89 & n6531 ;
  assign n17905 = x88 & ~n6530 ;
  assign n17906 = n6871 & n17905 ;
  assign n17907 = n17904 | n17906 ;
  assign n17908 = n17903 | n17907 ;
  assign n17909 = n6539 | n17903 ;
  assign n17910 = n17907 | n17909 ;
  assign n17911 = ( n3519 & n17908 ) | ( n3519 & n17910 ) | ( n17908 & n17910 ) ;
  assign n17912 = x38 & n17910 ;
  assign n17913 = x38 & n17903 ;
  assign n17914 = ( x38 & n17907 ) | ( x38 & n17913 ) | ( n17907 & n17913 ) ;
  assign n17915 = ( n3519 & n17912 ) | ( n3519 & n17914 ) | ( n17912 & n17914 ) ;
  assign n17916 = x38 & ~n17914 ;
  assign n17917 = x38 & ~n17910 ;
  assign n17918 = ( ~n3519 & n17916 ) | ( ~n3519 & n17917 ) | ( n17916 & n17917 ) ;
  assign n17919 = ( n17911 & ~n17915 ) | ( n17911 & n17918 ) | ( ~n17915 & n17918 ) ;
  assign n17920 = n17902 & n17919 ;
  assign n17921 = n17902 & ~n17920 ;
  assign n17922 = ~n17902 & n17919 ;
  assign n17923 = n17921 | n17922 ;
  assign n17924 = n17358 | n17364 ;
  assign n17925 = ( n17358 & n17361 ) | ( n17358 & n17924 ) | ( n17361 & n17924 ) ;
  assign n17926 = n17923 | n17925 ;
  assign n17927 = n17923 & n17925 ;
  assign n17928 = n17926 & ~n17927 ;
  assign n17929 = x93 & n5554 ;
  assign n17930 = x92 & n5549 ;
  assign n17931 = x91 & ~n5548 ;
  assign n17932 = n5893 & n17931 ;
  assign n17933 = n17930 | n17932 ;
  assign n17934 = n17929 | n17933 ;
  assign n17935 = n5557 | n17929 ;
  assign n17936 = n17933 | n17935 ;
  assign n17937 = ( n4305 & n17934 ) | ( n4305 & n17936 ) | ( n17934 & n17936 ) ;
  assign n17938 = x35 & n17936 ;
  assign n17939 = x35 & n17929 ;
  assign n17940 = ( x35 & n17933 ) | ( x35 & n17939 ) | ( n17933 & n17939 ) ;
  assign n17941 = ( n4305 & n17938 ) | ( n4305 & n17940 ) | ( n17938 & n17940 ) ;
  assign n17942 = x35 & ~n17940 ;
  assign n17943 = x35 & ~n17936 ;
  assign n17944 = ( ~n4305 & n17942 ) | ( ~n4305 & n17943 ) | ( n17942 & n17943 ) ;
  assign n17945 = ( n17937 & ~n17941 ) | ( n17937 & n17944 ) | ( ~n17941 & n17944 ) ;
  assign n17946 = n17928 & n17945 ;
  assign n17947 = n17928 & ~n17946 ;
  assign n17948 = ~n17928 & n17945 ;
  assign n17949 = n17947 | n17948 ;
  assign n17950 = n17385 | n17390 ;
  assign n17951 = ( n17385 & n17388 ) | ( n17385 & n17950 ) | ( n17388 & n17950 ) ;
  assign n17952 = n17949 | n17951 ;
  assign n17953 = n17949 & n17951 ;
  assign n17954 = n17952 & ~n17953 ;
  assign n17955 = x96 & n4631 ;
  assign n17956 = x95 & n4626 ;
  assign n17957 = x94 & ~n4625 ;
  assign n17958 = n4943 & n17957 ;
  assign n17959 = n17956 | n17958 ;
  assign n17960 = n17955 | n17959 ;
  assign n17961 = n4634 | n17955 ;
  assign n17962 = n17959 | n17961 ;
  assign n17963 = ( n5202 & n17960 ) | ( n5202 & n17962 ) | ( n17960 & n17962 ) ;
  assign n17964 = x32 & n17962 ;
  assign n17965 = x32 & n17955 ;
  assign n17966 = ( x32 & n17959 ) | ( x32 & n17965 ) | ( n17959 & n17965 ) ;
  assign n17967 = ( n5202 & n17964 ) | ( n5202 & n17966 ) | ( n17964 & n17966 ) ;
  assign n17968 = x32 & ~n17966 ;
  assign n17969 = x32 & ~n17962 ;
  assign n17970 = ( ~n5202 & n17968 ) | ( ~n5202 & n17969 ) | ( n17968 & n17969 ) ;
  assign n17971 = ( n17963 & ~n17967 ) | ( n17963 & n17970 ) | ( ~n17967 & n17970 ) ;
  assign n17972 = n17954 & n17971 ;
  assign n17973 = n17954 | n17971 ;
  assign n17974 = ~n17972 & n17973 ;
  assign n17975 = ( n16841 & n17393 ) | ( n16841 & n17410 ) | ( n17393 & n17410 ) ;
  assign n17976 = n17393 | n17410 ;
  assign n17977 = ( n16845 & n17975 ) | ( n16845 & n17976 ) | ( n17975 & n17976 ) ;
  assign n17978 = n17974 & n17977 ;
  assign n17979 = ~n17974 & n17977 ;
  assign n17980 = ( n17974 & ~n17978 ) | ( n17974 & n17979 ) | ( ~n17978 & n17979 ) ;
  assign n17981 = x99 & n3816 ;
  assign n17982 = x98 & n3811 ;
  assign n17983 = x97 & ~n3810 ;
  assign n17984 = n4067 & n17983 ;
  assign n17985 = n17982 | n17984 ;
  assign n17986 = n17981 | n17985 ;
  assign n17987 = n3819 | n17981 ;
  assign n17988 = n17985 | n17987 ;
  assign n17989 = ( n6164 & n17986 ) | ( n6164 & n17988 ) | ( n17986 & n17988 ) ;
  assign n17990 = x29 & n17988 ;
  assign n17991 = x29 & n17981 ;
  assign n17992 = ( x29 & n17985 ) | ( x29 & n17991 ) | ( n17985 & n17991 ) ;
  assign n17993 = ( n6164 & n17990 ) | ( n6164 & n17992 ) | ( n17990 & n17992 ) ;
  assign n17994 = x29 & ~n17992 ;
  assign n17995 = x29 & ~n17988 ;
  assign n17996 = ( ~n6164 & n17994 ) | ( ~n6164 & n17995 ) | ( n17994 & n17995 ) ;
  assign n17997 = ( n17989 & ~n17993 ) | ( n17989 & n17996 ) | ( ~n17993 & n17996 ) ;
  assign n17998 = n17980 & n17997 ;
  assign n17999 = n17980 & ~n17998 ;
  assign n18000 = ~n17980 & n17997 ;
  assign n18001 = n17999 | n18000 ;
  assign n18002 = n17442 | n17447 ;
  assign n18003 = ( n17442 & n17444 ) | ( n17442 & n18002 ) | ( n17444 & n18002 ) ;
  assign n18004 = n18001 | n18003 ;
  assign n18005 = n18001 & n18003 ;
  assign n18006 = n18004 & ~n18005 ;
  assign n18007 = x102 & n3085 ;
  assign n18008 = x101 & n3080 ;
  assign n18009 = x100 & ~n3079 ;
  assign n18010 = n3309 & n18009 ;
  assign n18011 = n18008 | n18010 ;
  assign n18012 = n18007 | n18011 ;
  assign n18013 = n3088 | n18007 ;
  assign n18014 = n18011 | n18013 ;
  assign n18015 = ( n7178 & n18012 ) | ( n7178 & n18014 ) | ( n18012 & n18014 ) ;
  assign n18016 = x26 & n18014 ;
  assign n18017 = x26 & n18007 ;
  assign n18018 = ( x26 & n18011 ) | ( x26 & n18017 ) | ( n18011 & n18017 ) ;
  assign n18019 = ( n7178 & n18016 ) | ( n7178 & n18018 ) | ( n18016 & n18018 ) ;
  assign n18020 = x26 & ~n18018 ;
  assign n18021 = x26 & ~n18014 ;
  assign n18022 = ( ~n7178 & n18020 ) | ( ~n7178 & n18021 ) | ( n18020 & n18021 ) ;
  assign n18023 = ( n18015 & ~n18019 ) | ( n18015 & n18022 ) | ( ~n18019 & n18022 ) ;
  assign n18024 = n18006 & n18023 ;
  assign n18025 = n18006 & ~n18024 ;
  assign n18026 = ~n18006 & n18023 ;
  assign n18027 = n18025 | n18026 ;
  assign n18028 = n17468 | n17474 ;
  assign n18029 = n18027 | n18028 ;
  assign n18030 = n18027 & n18028 ;
  assign n18031 = n18029 & ~n18030 ;
  assign n18032 = x105 & n2429 ;
  assign n18033 = x104 & n2424 ;
  assign n18034 = x103 & ~n2423 ;
  assign n18035 = n2631 & n18034 ;
  assign n18036 = n18033 | n18035 ;
  assign n18037 = n18032 | n18036 ;
  assign n18038 = n2432 | n18032 ;
  assign n18039 = n18036 | n18038 ;
  assign n18040 = ( n8273 & n18037 ) | ( n8273 & n18039 ) | ( n18037 & n18039 ) ;
  assign n18041 = x23 & n18039 ;
  assign n18042 = x23 & n18032 ;
  assign n18043 = ( x23 & n18036 ) | ( x23 & n18042 ) | ( n18036 & n18042 ) ;
  assign n18044 = ( n8273 & n18041 ) | ( n8273 & n18043 ) | ( n18041 & n18043 ) ;
  assign n18045 = x23 & ~n18043 ;
  assign n18046 = x23 & ~n18039 ;
  assign n18047 = ( ~n8273 & n18045 ) | ( ~n8273 & n18046 ) | ( n18045 & n18046 ) ;
  assign n18048 = ( n18040 & ~n18044 ) | ( n18040 & n18047 ) | ( ~n18044 & n18047 ) ;
  assign n18049 = n18031 & n18048 ;
  assign n18050 = n18031 | n18048 ;
  assign n18051 = ~n18049 & n18050 ;
  assign n18052 = n17493 & n18048 ;
  assign n18053 = ( n17493 & n18031 ) | ( n17493 & n18052 ) | ( n18031 & n18052 ) ;
  assign n18054 = ~n18049 & n18053 ;
  assign n18055 = ( n17501 & n18051 ) | ( n17501 & n18054 ) | ( n18051 & n18054 ) ;
  assign n18056 = n17704 & ~n18055 ;
  assign n18057 = x108 & n1859 ;
  assign n18058 = x107 & n1854 ;
  assign n18059 = x106 & ~n1853 ;
  assign n18060 = n2037 & n18059 ;
  assign n18061 = n18058 | n18060 ;
  assign n18062 = n18057 | n18061 ;
  assign n18063 = n1862 | n18057 ;
  assign n18064 = n18061 | n18063 ;
  assign n18065 = ( n9479 & n18062 ) | ( n9479 & n18064 ) | ( n18062 & n18064 ) ;
  assign n18066 = x20 & n18064 ;
  assign n18067 = x20 & n18057 ;
  assign n18068 = ( x20 & n18061 ) | ( x20 & n18067 ) | ( n18061 & n18067 ) ;
  assign n18069 = ( n9479 & n18066 ) | ( n9479 & n18068 ) | ( n18066 & n18068 ) ;
  assign n18070 = x20 & ~n18068 ;
  assign n18071 = x20 & ~n18064 ;
  assign n18072 = ( ~n9479 & n18070 ) | ( ~n9479 & n18071 ) | ( n18070 & n18071 ) ;
  assign n18073 = ( n18065 & ~n18069 ) | ( n18065 & n18072 ) | ( ~n18069 & n18072 ) ;
  assign n18074 = ( n17501 & n18050 ) | ( n17501 & n18053 ) | ( n18050 & n18053 ) ;
  assign n18075 = n18051 & n18073 ;
  assign n18076 = ~n18074 & n18075 ;
  assign n18077 = ( n18056 & n18073 ) | ( n18056 & n18076 ) | ( n18073 & n18076 ) ;
  assign n18078 = n18051 | n18073 ;
  assign n18079 = ( n18073 & ~n18074 ) | ( n18073 & n18078 ) | ( ~n18074 & n18078 ) ;
  assign n18080 = n18056 | n18079 ;
  assign n18081 = ~n18077 & n18080 ;
  assign n18082 = n17520 | n17522 ;
  assign n18083 = ( n17520 & n17524 ) | ( n17520 & n18082 ) | ( n17524 & n18082 ) ;
  assign n18084 = ~n18081 & n18083 ;
  assign n18085 = n18081 & ~n18083 ;
  assign n18086 = n18084 | n18085 ;
  assign n18087 = x111 & n1383 ;
  assign n18088 = x110 & n1378 ;
  assign n18089 = x109 & ~n1377 ;
  assign n18090 = n1542 & n18089 ;
  assign n18091 = n18088 | n18090 ;
  assign n18092 = n18087 | n18091 ;
  assign n18093 = n1386 | n18087 ;
  assign n18094 = n18091 | n18093 ;
  assign n18095 = ( n10749 & n18092 ) | ( n10749 & n18094 ) | ( n18092 & n18094 ) ;
  assign n18096 = x17 & n18094 ;
  assign n18097 = x17 & n18087 ;
  assign n18098 = ( x17 & n18091 ) | ( x17 & n18097 ) | ( n18091 & n18097 ) ;
  assign n18099 = ( n10749 & n18096 ) | ( n10749 & n18098 ) | ( n18096 & n18098 ) ;
  assign n18100 = x17 & ~n18098 ;
  assign n18101 = x17 & ~n18094 ;
  assign n18102 = ( ~n10749 & n18100 ) | ( ~n10749 & n18101 ) | ( n18100 & n18101 ) ;
  assign n18103 = ( n18095 & ~n18099 ) | ( n18095 & n18102 ) | ( ~n18099 & n18102 ) ;
  assign n18104 = n18086 & n18103 ;
  assign n18105 = n18086 | n18103 ;
  assign n18106 = ~n18104 & n18105 ;
  assign n18107 = n17547 | n17552 ;
  assign n18108 = ( n17121 & n17547 ) | ( n17121 & n18107 ) | ( n17547 & n18107 ) ;
  assign n18109 = n18106 & n18108 ;
  assign n18110 = n18106 | n18108 ;
  assign n18111 = ~n18109 & n18110 ;
  assign n18112 = x114 & n962 ;
  assign n18113 = x113 & n957 ;
  assign n18114 = x112 & ~n956 ;
  assign n18115 = n1105 & n18114 ;
  assign n18116 = n18113 | n18115 ;
  assign n18117 = n18112 | n18116 ;
  assign n18118 = n965 | n18112 ;
  assign n18119 = n18116 | n18118 ;
  assign n18120 = ( ~n12095 & n18117 ) | ( ~n12095 & n18119 ) | ( n18117 & n18119 ) ;
  assign n18121 = n18117 & n18119 ;
  assign n18122 = ( n12079 & n18120 ) | ( n12079 & n18121 ) | ( n18120 & n18121 ) ;
  assign n18123 = x14 & n18122 ;
  assign n18124 = x14 & ~n18122 ;
  assign n18125 = ( n18122 & ~n18123 ) | ( n18122 & n18124 ) | ( ~n18123 & n18124 ) ;
  assign n18126 = n18111 & n18125 ;
  assign n18127 = n18111 & ~n18126 ;
  assign n18128 = ~n18111 & n18125 ;
  assign n18129 = n18127 | n18128 ;
  assign n18130 = n17571 | n17572 ;
  assign n18131 = ( n17120 & n17571 ) | ( n17120 & n18130 ) | ( n17571 & n18130 ) ;
  assign n18132 = ~n18129 & n18131 ;
  assign n18133 = n18129 & ~n18131 ;
  assign n18134 = n18132 | n18133 ;
  assign n18135 = x117 & n636 ;
  assign n18136 = x116 & n631 ;
  assign n18137 = x115 & ~n630 ;
  assign n18138 = n764 & n18137 ;
  assign n18139 = n18136 | n18138 ;
  assign n18140 = n18135 | n18139 ;
  assign n18141 = n639 | n18135 ;
  assign n18142 = n18139 | n18141 ;
  assign n18143 = ( ~n13522 & n18140 ) | ( ~n13522 & n18142 ) | ( n18140 & n18142 ) ;
  assign n18144 = n18140 & n18142 ;
  assign n18145 = ( n13503 & n18143 ) | ( n13503 & n18144 ) | ( n18143 & n18144 ) ;
  assign n18146 = x11 & n18145 ;
  assign n18147 = x11 & ~n18145 ;
  assign n18148 = ( n18145 & ~n18146 ) | ( n18145 & n18147 ) | ( ~n18146 & n18147 ) ;
  assign n18149 = n18134 & n18148 ;
  assign n18150 = n18134 | n18148 ;
  assign n18151 = ~n18149 & n18150 ;
  assign n18152 = n17591 | n17592 ;
  assign n18153 = ( n17591 & n17595 ) | ( n17591 & n18152 ) | ( n17595 & n18152 ) ;
  assign n18154 = n18151 & n18153 ;
  assign n18155 = n18151 | n18153 ;
  assign n18156 = ~n18154 & n18155 ;
  assign n18157 = x120 & n389 ;
  assign n18158 = x119 & n384 ;
  assign n18159 = x118 & ~n383 ;
  assign n18160 = n463 & n18159 ;
  assign n18161 = n18158 | n18160 ;
  assign n18162 = n18157 | n18161 ;
  assign n18163 = n392 | n18157 ;
  assign n18164 = n18161 | n18163 ;
  assign n18165 = ( n14991 & n18162 ) | ( n14991 & n18164 ) | ( n18162 & n18164 ) ;
  assign n18166 = x8 & n18164 ;
  assign n18167 = x8 & n18157 ;
  assign n18168 = ( x8 & n18161 ) | ( x8 & n18167 ) | ( n18161 & n18167 ) ;
  assign n18169 = ( n14991 & n18166 ) | ( n14991 & n18168 ) | ( n18166 & n18168 ) ;
  assign n18170 = x8 & ~n18168 ;
  assign n18171 = x8 & ~n18164 ;
  assign n18172 = ( ~n14991 & n18170 ) | ( ~n14991 & n18171 ) | ( n18170 & n18171 ) ;
  assign n18173 = ( n18165 & ~n18169 ) | ( n18165 & n18172 ) | ( ~n18169 & n18172 ) ;
  assign n18174 = n18156 | n18173 ;
  assign n18175 = n18156 & n18173 ;
  assign n18176 = n18174 & ~n18175 ;
  assign n18177 = x123 & n212 ;
  assign n18178 = x122 & n207 ;
  assign n18179 = x121 & ~n206 ;
  assign n18180 = n267 & n18179 ;
  assign n18181 = n18178 | n18180 ;
  assign n18182 = n18177 | n18181 ;
  assign n18183 = n215 | n18177 ;
  assign n18184 = n18181 | n18183 ;
  assign n18185 = ( n16086 & n18182 ) | ( n16086 & n18184 ) | ( n18182 & n18184 ) ;
  assign n18186 = x5 & n18184 ;
  assign n18187 = x5 & n18177 ;
  assign n18188 = ( x5 & n18181 ) | ( x5 & n18187 ) | ( n18181 & n18187 ) ;
  assign n18189 = ( n16086 & n18186 ) | ( n16086 & n18188 ) | ( n18186 & n18188 ) ;
  assign n18190 = x5 & ~n18188 ;
  assign n18191 = x5 & ~n18184 ;
  assign n18192 = ( ~n16086 & n18190 ) | ( ~n16086 & n18191 ) | ( n18190 & n18191 ) ;
  assign n18193 = ( n18185 & ~n18189 ) | ( n18185 & n18192 ) | ( ~n18189 & n18192 ) ;
  assign n18194 = ~n18176 & n18193 ;
  assign n18195 = n17703 & n18194 ;
  assign n18196 = n18173 | n18193 ;
  assign n18197 = ( n18156 & n18193 ) | ( n18156 & n18196 ) | ( n18193 & n18196 ) ;
  assign n18198 = n18174 & ~n18197 ;
  assign n18199 = ( n17703 & n18195 ) | ( n17703 & n18198 ) | ( n18195 & n18198 ) ;
  assign n18200 = x125 | x126 ;
  assign n18201 = x125 & x126 ;
  assign n18202 = n18200 & ~n18201 ;
  assign n18203 = n17646 | n17652 ;
  assign n18204 = n17646 | n17650 ;
  assign n18205 = ( n16075 & n18203 ) | ( n16075 & n18204 ) | ( n18203 & n18204 ) ;
  assign n18206 = n17646 | n17647 ;
  assign n18207 = n17064 | n17646 ;
  assign n18208 = ( n17646 & n17647 ) | ( n17646 & n18207 ) | ( n17647 & n18207 ) ;
  assign n18209 = ( n17070 & n18206 ) | ( n17070 & n18208 ) | ( n18206 & n18208 ) ;
  assign n18210 = ( n17068 & n18206 ) | ( n17068 & n18208 ) | ( n18206 & n18208 ) ;
  assign n18211 = ( n16033 & n18209 ) | ( n16033 & n18210 ) | ( n18209 & n18210 ) ;
  assign n18212 = n18205 | n18211 ;
  assign n18213 = n18202 & n18212 ;
  assign n18214 = ( n13965 & n18205 ) | ( n13965 & n18211 ) | ( n18205 & n18211 ) ;
  assign n18215 = n18202 & n18214 ;
  assign n18216 = ( n14002 & n18213 ) | ( n14002 & n18215 ) | ( n18213 & n18215 ) ;
  assign n18217 = n18202 | n18212 ;
  assign n18218 = n18202 | n18214 ;
  assign n18219 = ( n14002 & n18217 ) | ( n14002 & n18218 ) | ( n18217 & n18218 ) ;
  assign n18220 = ~n18216 & n18219 ;
  assign n18221 = x125 & n133 ;
  assign n18222 = x124 & ~n162 ;
  assign n18223 = ( n137 & n18221 ) | ( n137 & n18222 ) | ( n18221 & n18222 ) ;
  assign n18224 = x0 & x126 ;
  assign n18225 = ( ~n137 & n18221 ) | ( ~n137 & n18224 ) | ( n18221 & n18224 ) ;
  assign n18226 = n18223 | n18225 ;
  assign n18227 = n141 | n18226 ;
  assign n18228 = ( n18220 & n18226 ) | ( n18220 & n18227 ) | ( n18226 & n18227 ) ;
  assign n18229 = x2 & n18226 ;
  assign n18230 = ( x2 & n523 ) | ( x2 & n18226 ) | ( n523 & n18226 ) ;
  assign n18231 = ( n18220 & n18229 ) | ( n18220 & n18230 ) | ( n18229 & n18230 ) ;
  assign n18232 = x2 & ~n18230 ;
  assign n18233 = x2 & ~n18226 ;
  assign n18234 = ( ~n18220 & n18232 ) | ( ~n18220 & n18233 ) | ( n18232 & n18233 ) ;
  assign n18235 = ( n18228 & ~n18231 ) | ( n18228 & n18234 ) | ( ~n18231 & n18234 ) ;
  assign n18236 = n18194 | n18198 ;
  assign n18237 = n17703 | n18236 ;
  assign n18238 = n18235 & n18237 ;
  assign n18239 = ~n18199 & n18238 ;
  assign n18240 = n18235 | n18237 ;
  assign n18241 = ( ~n18199 & n18235 ) | ( ~n18199 & n18240 ) | ( n18235 & n18240 ) ;
  assign n18242 = ~n18239 & n18241 ;
  assign n18243 = ( n17643 & n17644 ) | ( n17643 & n17691 ) | ( n17644 & n17691 ) ;
  assign n18244 = n18242 & n18243 ;
  assign n18245 = n18242 | n18243 ;
  assign n18246 = ~n18244 & n18245 ;
  assign n18247 = n17694 | n17697 ;
  assign n18248 = ( n17694 & n17699 ) | ( n17694 & n18247 ) | ( n17699 & n18247 ) ;
  assign n18249 = n18246 | n18248 ;
  assign n18250 = n18246 & n18247 ;
  assign n18251 = n17694 & n18246 ;
  assign n18252 = ( n17699 & n18250 ) | ( n17699 & n18251 ) | ( n18250 & n18251 ) ;
  assign n18253 = n18249 & ~n18252 ;
  assign n18254 = x124 & n212 ;
  assign n18255 = x123 & n207 ;
  assign n18256 = x122 & ~n206 ;
  assign n18257 = n267 & n18256 ;
  assign n18258 = n18255 | n18257 ;
  assign n18259 = n18254 | n18258 ;
  assign n18260 = n215 | n18254 ;
  assign n18261 = n18258 | n18260 ;
  assign n18262 = ( n17084 & n18259 ) | ( n17084 & n18261 ) | ( n18259 & n18261 ) ;
  assign n18263 = x5 & n18261 ;
  assign n18264 = x5 & n18254 ;
  assign n18265 = ( x5 & n18258 ) | ( x5 & n18264 ) | ( n18258 & n18264 ) ;
  assign n18266 = ( n17084 & n18263 ) | ( n17084 & n18265 ) | ( n18263 & n18265 ) ;
  assign n18267 = x5 & ~n18265 ;
  assign n18268 = x5 & ~n18261 ;
  assign n18269 = ( ~n17084 & n18267 ) | ( ~n17084 & n18268 ) | ( n18267 & n18268 ) ;
  assign n18270 = ( n18262 & ~n18266 ) | ( n18262 & n18269 ) | ( ~n18266 & n18269 ) ;
  assign n18271 = n17755 | n17759 ;
  assign n18272 = x69 & n15547 ;
  assign n18273 = x68 & ~n15546 ;
  assign n18274 = n16123 & n18273 ;
  assign n18275 = n18272 | n18274 ;
  assign n18276 = x70 & n15552 ;
  assign n18277 = n15555 | n18276 ;
  assign n18278 = n18275 | n18277 ;
  assign n18279 = x59 & ~n18278 ;
  assign n18280 = x59 & ~n18276 ;
  assign n18281 = ~n18275 & n18280 ;
  assign n18282 = ( ~n340 & n18279 ) | ( ~n340 & n18281 ) | ( n18279 & n18281 ) ;
  assign n18283 = ~x59 & n18278 ;
  assign n18284 = ~x59 & n18276 ;
  assign n18285 = ( ~x59 & n18275 ) | ( ~x59 & n18284 ) | ( n18275 & n18284 ) ;
  assign n18286 = ( n340 & n18283 ) | ( n340 & n18285 ) | ( n18283 & n18285 ) ;
  assign n18287 = n18282 | n18286 ;
  assign n18288 = x62 & ~x63 ;
  assign n18289 = ~x62 & x63 ;
  assign n18290 = n18288 | n18289 ;
  assign n18291 = x64 & n18290 ;
  assign n18292 = n17161 & n18291 ;
  assign n18293 = n17736 & n18292 ;
  assign n18294 = n17738 & ~n18293 ;
  assign n18295 = x67 & n17146 ;
  assign n18296 = x66 & n17141 ;
  assign n18297 = x65 & ~n17140 ;
  assign n18298 = n17724 & n18297 ;
  assign n18299 = n18296 | n18298 ;
  assign n18300 = n18295 | n18299 ;
  assign n18301 = n186 & n17149 ;
  assign n18302 = n18300 | n18301 ;
  assign n18303 = x62 & ~n18302 ;
  assign n18304 = ~x62 & n18302 ;
  assign n18305 = n18303 | n18304 ;
  assign n18306 = ~n17161 & n18291 ;
  assign n18307 = ( ~n17736 & n18291 ) | ( ~n17736 & n18306 ) | ( n18291 & n18306 ) ;
  assign n18308 = n18305 & n18307 ;
  assign n18309 = ( n18294 & n18305 ) | ( n18294 & n18308 ) | ( n18305 & n18308 ) ;
  assign n18310 = n18305 | n18307 ;
  assign n18311 = n18294 | n18310 ;
  assign n18312 = ~n18309 & n18311 ;
  assign n18313 = n18287 | n18312 ;
  assign n18314 = n18287 & n18312 ;
  assign n18315 = n18313 & ~n18314 ;
  assign n18316 = n18271 & n18315 ;
  assign n18317 = n18271 | n18315 ;
  assign n18318 = ~n18316 & n18317 ;
  assign n18319 = x73 & n14045 ;
  assign n18320 = x72 & n14040 ;
  assign n18321 = x71 & ~n14039 ;
  assign n18322 = n14552 & n18321 ;
  assign n18323 = n18320 | n18322 ;
  assign n18324 = n18319 | n18323 ;
  assign n18325 = ( ~n610 & n14048 ) | ( ~n610 & n18324 ) | ( n14048 & n18324 ) ;
  assign n18326 = n14048 & n18319 ;
  assign n18327 = ( n14048 & n18323 ) | ( n14048 & n18326 ) | ( n18323 & n18326 ) ;
  assign n18328 = ( n598 & n18325 ) | ( n598 & n18327 ) | ( n18325 & n18327 ) ;
  assign n18329 = ( x56 & ~n18324 ) | ( x56 & n18328 ) | ( ~n18324 & n18328 ) ;
  assign n18330 = ~n18328 & n18329 ;
  assign n18331 = x56 | n18319 ;
  assign n18332 = n18323 | n18331 ;
  assign n18333 = n18328 | n18332 ;
  assign n18334 = ( ~x56 & n18330 ) | ( ~x56 & n18333 ) | ( n18330 & n18333 ) ;
  assign n18335 = n18318 & n18334 ;
  assign n18336 = n18318 & ~n18335 ;
  assign n18337 = ~n18318 & n18334 ;
  assign n18338 = n18336 | n18337 ;
  assign n18339 = n17763 | n17766 ;
  assign n18340 = ( n17763 & n17768 ) | ( n17763 & n18339 ) | ( n17768 & n18339 ) ;
  assign n18341 = ~n18338 & n18340 ;
  assign n18342 = n18338 & ~n18340 ;
  assign n18343 = n18341 | n18342 ;
  assign n18344 = x76 & n12574 ;
  assign n18345 = x75 & n12569 ;
  assign n18346 = x74 & ~n12568 ;
  assign n18347 = n13076 & n18346 ;
  assign n18348 = n18345 | n18347 ;
  assign n18349 = n18344 | n18348 ;
  assign n18350 = n12577 | n18344 ;
  assign n18351 = n18348 | n18350 ;
  assign n18352 = ( n923 & n18349 ) | ( n923 & n18351 ) | ( n18349 & n18351 ) ;
  assign n18353 = x53 & n18351 ;
  assign n18354 = x53 & n18344 ;
  assign n18355 = ( x53 & n18348 ) | ( x53 & n18354 ) | ( n18348 & n18354 ) ;
  assign n18356 = ( n923 & n18353 ) | ( n923 & n18355 ) | ( n18353 & n18355 ) ;
  assign n18357 = x53 & ~n18355 ;
  assign n18358 = x53 & ~n18351 ;
  assign n18359 = ( ~n923 & n18357 ) | ( ~n923 & n18358 ) | ( n18357 & n18358 ) ;
  assign n18360 = ( n18352 & ~n18356 ) | ( n18352 & n18359 ) | ( ~n18356 & n18359 ) ;
  assign n18361 = n18343 | n18360 ;
  assign n18362 = n18343 & n18360 ;
  assign n18363 = n18361 & ~n18362 ;
  assign n18364 = n17790 | n17791 ;
  assign n18365 = ( n17790 & n17792 ) | ( n17790 & n18364 ) | ( n17792 & n18364 ) ;
  assign n18366 = n18363 & n18365 ;
  assign n18367 = n18363 | n18365 ;
  assign n18368 = ~n18366 & n18367 ;
  assign n18369 = x79 & n11205 ;
  assign n18370 = x78 & n11200 ;
  assign n18371 = x77 & ~n11199 ;
  assign n18372 = n11679 & n18371 ;
  assign n18373 = n18370 | n18372 ;
  assign n18374 = n18369 | n18373 ;
  assign n18375 = n11208 | n18369 ;
  assign n18376 = n18373 | n18375 ;
  assign n18377 = ( n1332 & n18374 ) | ( n1332 & n18376 ) | ( n18374 & n18376 ) ;
  assign n18378 = x50 & n18376 ;
  assign n18379 = x50 & n18369 ;
  assign n18380 = ( x50 & n18373 ) | ( x50 & n18379 ) | ( n18373 & n18379 ) ;
  assign n18381 = ( n1332 & n18378 ) | ( n1332 & n18380 ) | ( n18378 & n18380 ) ;
  assign n18382 = x50 & ~n18380 ;
  assign n18383 = x50 & ~n18376 ;
  assign n18384 = ( ~n1332 & n18382 ) | ( ~n1332 & n18383 ) | ( n18382 & n18383 ) ;
  assign n18385 = ( n18377 & ~n18381 ) | ( n18377 & n18384 ) | ( ~n18381 & n18384 ) ;
  assign n18386 = n18368 & n18385 ;
  assign n18387 = n18368 & ~n18386 ;
  assign n18388 = ~n18368 & n18385 ;
  assign n18389 = n18387 | n18388 ;
  assign n18390 = n17705 | n17813 ;
  assign n18391 = ( n17813 & n17816 ) | ( n17813 & n18390 ) | ( n17816 & n18390 ) ;
  assign n18392 = n18389 | n18391 ;
  assign n18393 = n18389 & n18391 ;
  assign n18394 = n18392 & ~n18393 ;
  assign n18395 = x82 & n9933 ;
  assign n18396 = x81 & n9928 ;
  assign n18397 = x80 & ~n9927 ;
  assign n18398 = n10379 & n18397 ;
  assign n18399 = n18396 | n18398 ;
  assign n18400 = n18395 | n18399 ;
  assign n18401 = n9936 | n18395 ;
  assign n18402 = n18399 | n18401 ;
  assign n18403 = ( n1811 & n18400 ) | ( n1811 & n18402 ) | ( n18400 & n18402 ) ;
  assign n18404 = x47 & n18402 ;
  assign n18405 = x47 & n18395 ;
  assign n18406 = ( x47 & n18399 ) | ( x47 & n18405 ) | ( n18399 & n18405 ) ;
  assign n18407 = ( n1811 & n18404 ) | ( n1811 & n18406 ) | ( n18404 & n18406 ) ;
  assign n18408 = x47 & ~n18406 ;
  assign n18409 = x47 & ~n18402 ;
  assign n18410 = ( ~n1811 & n18408 ) | ( ~n1811 & n18409 ) | ( n18408 & n18409 ) ;
  assign n18411 = ( n18403 & ~n18407 ) | ( n18403 & n18410 ) | ( ~n18407 & n18410 ) ;
  assign n18412 = n18394 | n18411 ;
  assign n18413 = n18394 & n18411 ;
  assign n18414 = n18412 & ~n18413 ;
  assign n18415 = n17837 | n17843 ;
  assign n18416 = ( n17837 & n17840 ) | ( n17837 & n18415 ) | ( n17840 & n18415 ) ;
  assign n18417 = n18414 & n18416 ;
  assign n18418 = n18414 | n18416 ;
  assign n18419 = ~n18417 & n18418 ;
  assign n18420 = x85 & n8724 ;
  assign n18421 = x84 & n8719 ;
  assign n18422 = x83 & ~n8718 ;
  assign n18423 = n9149 & n18422 ;
  assign n18424 = n18421 | n18423 ;
  assign n18425 = n18420 | n18424 ;
  assign n18426 = n8727 | n18420 ;
  assign n18427 = n18424 | n18426 ;
  assign n18428 = ( n2381 & n18425 ) | ( n2381 & n18427 ) | ( n18425 & n18427 ) ;
  assign n18429 = x44 & n18427 ;
  assign n18430 = x44 & n18420 ;
  assign n18431 = ( x44 & n18424 ) | ( x44 & n18430 ) | ( n18424 & n18430 ) ;
  assign n18432 = ( n2381 & n18429 ) | ( n2381 & n18431 ) | ( n18429 & n18431 ) ;
  assign n18433 = x44 & ~n18431 ;
  assign n18434 = x44 & ~n18427 ;
  assign n18435 = ( ~n2381 & n18433 ) | ( ~n2381 & n18434 ) | ( n18433 & n18434 ) ;
  assign n18436 = ( n18428 & ~n18432 ) | ( n18428 & n18435 ) | ( ~n18432 & n18435 ) ;
  assign n18437 = n18419 & n18436 ;
  assign n18438 = n18419 | n18436 ;
  assign n18439 = ~n18437 & n18438 ;
  assign n18440 = ( n17847 & n17864 ) | ( n17847 & n17874 ) | ( n17864 & n17874 ) ;
  assign n18441 = n18439 | n18440 ;
  assign n18442 = n18439 & n18440 ;
  assign n18443 = n18441 & ~n18442 ;
  assign n18444 = x88 & n7566 ;
  assign n18445 = x87 & n7561 ;
  assign n18446 = x86 & ~n7560 ;
  assign n18447 = n7953 & n18446 ;
  assign n18448 = n18445 | n18447 ;
  assign n18449 = n18444 | n18448 ;
  assign n18450 = n7569 | n18444 ;
  assign n18451 = n18448 | n18450 ;
  assign n18452 = ( ~n3039 & n18449 ) | ( ~n3039 & n18451 ) | ( n18449 & n18451 ) ;
  assign n18453 = n18449 & n18451 ;
  assign n18454 = ( n3023 & n18452 ) | ( n3023 & n18453 ) | ( n18452 & n18453 ) ;
  assign n18455 = x41 & n18451 ;
  assign n18456 = x41 & n18444 ;
  assign n18457 = ( x41 & n18448 ) | ( x41 & n18456 ) | ( n18448 & n18456 ) ;
  assign n18458 = ( ~n3039 & n18455 ) | ( ~n3039 & n18457 ) | ( n18455 & n18457 ) ;
  assign n18459 = n18455 & n18457 ;
  assign n18460 = ( n3023 & n18458 ) | ( n3023 & n18459 ) | ( n18458 & n18459 ) ;
  assign n18461 = x41 & ~n18457 ;
  assign n18462 = x41 & ~n18451 ;
  assign n18463 = ( n3039 & n18461 ) | ( n3039 & n18462 ) | ( n18461 & n18462 ) ;
  assign n18464 = n18461 | n18462 ;
  assign n18465 = ( ~n3023 & n18463 ) | ( ~n3023 & n18464 ) | ( n18463 & n18464 ) ;
  assign n18466 = ( n18454 & ~n18460 ) | ( n18454 & n18465 ) | ( ~n18460 & n18465 ) ;
  assign n18467 = n18443 & n18466 ;
  assign n18468 = n18443 & ~n18467 ;
  assign n18469 = ~n18443 & n18466 ;
  assign n18470 = n18468 | n18469 ;
  assign n18471 = n17895 | n17901 ;
  assign n18472 = n18470 | n18471 ;
  assign n18473 = n18470 & n18471 ;
  assign n18474 = n18472 & ~n18473 ;
  assign n18475 = x91 & n6536 ;
  assign n18476 = x90 & n6531 ;
  assign n18477 = x89 & ~n6530 ;
  assign n18478 = n6871 & n18477 ;
  assign n18479 = n18476 | n18478 ;
  assign n18480 = n18475 | n18479 ;
  assign n18481 = n6539 | n18475 ;
  assign n18482 = n18479 | n18481 ;
  assign n18483 = ( n3768 & n18480 ) | ( n3768 & n18482 ) | ( n18480 & n18482 ) ;
  assign n18484 = x38 & n18482 ;
  assign n18485 = x38 & n18475 ;
  assign n18486 = ( x38 & n18479 ) | ( x38 & n18485 ) | ( n18479 & n18485 ) ;
  assign n18487 = ( n3768 & n18484 ) | ( n3768 & n18486 ) | ( n18484 & n18486 ) ;
  assign n18488 = x38 & ~n18486 ;
  assign n18489 = x38 & ~n18482 ;
  assign n18490 = ( ~n3768 & n18488 ) | ( ~n3768 & n18489 ) | ( n18488 & n18489 ) ;
  assign n18491 = ( n18483 & ~n18487 ) | ( n18483 & n18490 ) | ( ~n18487 & n18490 ) ;
  assign n18492 = n18474 & n18491 ;
  assign n18493 = n18474 & ~n18492 ;
  assign n18494 = ~n18474 & n18491 ;
  assign n18495 = n18493 | n18494 ;
  assign n18496 = n17920 | n17927 ;
  assign n18497 = n18495 | n18496 ;
  assign n18498 = n18495 & n18496 ;
  assign n18499 = n18497 & ~n18498 ;
  assign n18500 = x94 & n5554 ;
  assign n18501 = x93 & n5549 ;
  assign n18502 = x92 & ~n5548 ;
  assign n18503 = n5893 & n18502 ;
  assign n18504 = n18501 | n18503 ;
  assign n18505 = n18500 | n18504 ;
  assign n18506 = n5557 | n18500 ;
  assign n18507 = n18504 | n18506 ;
  assign n18508 = ( n4583 & n18505 ) | ( n4583 & n18507 ) | ( n18505 & n18507 ) ;
  assign n18509 = x35 & n18507 ;
  assign n18510 = x35 & n18500 ;
  assign n18511 = ( x35 & n18504 ) | ( x35 & n18510 ) | ( n18504 & n18510 ) ;
  assign n18512 = ( n4583 & n18509 ) | ( n4583 & n18511 ) | ( n18509 & n18511 ) ;
  assign n18513 = x35 & ~n18511 ;
  assign n18514 = x35 & ~n18507 ;
  assign n18515 = ( ~n4583 & n18513 ) | ( ~n4583 & n18514 ) | ( n18513 & n18514 ) ;
  assign n18516 = ( n18508 & ~n18512 ) | ( n18508 & n18515 ) | ( ~n18512 & n18515 ) ;
  assign n18517 = n18499 | n18516 ;
  assign n18518 = n18499 & n18516 ;
  assign n18519 = n18517 & ~n18518 ;
  assign n18520 = n17946 & n18519 ;
  assign n18521 = ( n17953 & n18519 ) | ( n17953 & n18520 ) | ( n18519 & n18520 ) ;
  assign n18522 = n17946 | n18519 ;
  assign n18523 = n17953 | n18522 ;
  assign n18524 = ~n18521 & n18523 ;
  assign n18525 = x97 & n4631 ;
  assign n18526 = x96 & n4626 ;
  assign n18527 = x95 & ~n4625 ;
  assign n18528 = n4943 & n18527 ;
  assign n18529 = n18526 | n18528 ;
  assign n18530 = n18525 | n18529 ;
  assign n18531 = n4634 | n18525 ;
  assign n18532 = n18529 | n18531 ;
  assign n18533 = ( n5505 & n18530 ) | ( n5505 & n18532 ) | ( n18530 & n18532 ) ;
  assign n18534 = x32 & n18532 ;
  assign n18535 = x32 & n18525 ;
  assign n18536 = ( x32 & n18529 ) | ( x32 & n18535 ) | ( n18529 & n18535 ) ;
  assign n18537 = ( n5505 & n18534 ) | ( n5505 & n18536 ) | ( n18534 & n18536 ) ;
  assign n18538 = x32 & ~n18536 ;
  assign n18539 = x32 & ~n18532 ;
  assign n18540 = ( ~n5505 & n18538 ) | ( ~n5505 & n18539 ) | ( n18538 & n18539 ) ;
  assign n18541 = ( n18533 & ~n18537 ) | ( n18533 & n18540 ) | ( ~n18537 & n18540 ) ;
  assign n18542 = n18524 & n18541 ;
  assign n18543 = n18524 & ~n18542 ;
  assign n18544 = ~n18524 & n18541 ;
  assign n18545 = n17972 | n17977 ;
  assign n18546 = ( n17972 & n17974 ) | ( n17972 & n18545 ) | ( n17974 & n18545 ) ;
  assign n18547 = ~n18544 & n18546 ;
  assign n18548 = ~n18543 & n18547 ;
  assign n18549 = n18544 & ~n18546 ;
  assign n18550 = ( n18543 & ~n18546 ) | ( n18543 & n18549 ) | ( ~n18546 & n18549 ) ;
  assign n18551 = n18548 | n18550 ;
  assign n18552 = x100 & n3816 ;
  assign n18553 = x99 & n3811 ;
  assign n18554 = x98 & ~n3810 ;
  assign n18555 = n4067 & n18554 ;
  assign n18556 = n18553 | n18555 ;
  assign n18557 = n18552 | n18556 ;
  assign n18558 = n3819 | n18552 ;
  assign n18559 = n18556 | n18558 ;
  assign n18560 = ( n6483 & n18557 ) | ( n6483 & n18559 ) | ( n18557 & n18559 ) ;
  assign n18561 = x29 & n18559 ;
  assign n18562 = x29 & n18552 ;
  assign n18563 = ( x29 & n18556 ) | ( x29 & n18562 ) | ( n18556 & n18562 ) ;
  assign n18564 = ( n6483 & n18561 ) | ( n6483 & n18563 ) | ( n18561 & n18563 ) ;
  assign n18565 = x29 & ~n18563 ;
  assign n18566 = x29 & ~n18559 ;
  assign n18567 = ( ~n6483 & n18565 ) | ( ~n6483 & n18566 ) | ( n18565 & n18566 ) ;
  assign n18568 = ( n18560 & ~n18564 ) | ( n18560 & n18567 ) | ( ~n18564 & n18567 ) ;
  assign n18569 = n18551 & n18568 ;
  assign n18570 = n18551 | n18568 ;
  assign n18571 = ~n18569 & n18570 ;
  assign n18572 = n17998 | n18003 ;
  assign n18573 = ( n17998 & n18001 ) | ( n17998 & n18572 ) | ( n18001 & n18572 ) ;
  assign n18574 = n18571 | n18573 ;
  assign n18575 = n18571 & n18573 ;
  assign n18576 = n18574 & ~n18575 ;
  assign n18577 = x103 & n3085 ;
  assign n18578 = x102 & n3080 ;
  assign n18579 = x101 & ~n3079 ;
  assign n18580 = n3309 & n18579 ;
  assign n18581 = n18578 | n18580 ;
  assign n18582 = n18577 | n18581 ;
  assign n18583 = n3088 | n18577 ;
  assign n18584 = n18581 | n18583 ;
  assign n18585 = ( n7529 & n18582 ) | ( n7529 & n18584 ) | ( n18582 & n18584 ) ;
  assign n18586 = x26 & n18584 ;
  assign n18587 = x26 & n18577 ;
  assign n18588 = ( x26 & n18581 ) | ( x26 & n18587 ) | ( n18581 & n18587 ) ;
  assign n18589 = ( n7529 & n18586 ) | ( n7529 & n18588 ) | ( n18586 & n18588 ) ;
  assign n18590 = x26 & ~n18588 ;
  assign n18591 = x26 & ~n18584 ;
  assign n18592 = ( ~n7529 & n18590 ) | ( ~n7529 & n18591 ) | ( n18590 & n18591 ) ;
  assign n18593 = ( n18585 & ~n18589 ) | ( n18585 & n18592 ) | ( ~n18589 & n18592 ) ;
  assign n18594 = n18576 | n18593 ;
  assign n18595 = n18576 & n18593 ;
  assign n18596 = n18594 & ~n18595 ;
  assign n18597 = n18024 & n18596 ;
  assign n18598 = ( n18030 & n18596 ) | ( n18030 & n18597 ) | ( n18596 & n18597 ) ;
  assign n18599 = n18024 | n18596 ;
  assign n18600 = n18030 | n18599 ;
  assign n18601 = ~n18598 & n18600 ;
  assign n18602 = x106 & n2429 ;
  assign n18603 = x105 & n2424 ;
  assign n18604 = x104 & ~n2423 ;
  assign n18605 = n2631 & n18604 ;
  assign n18606 = n18603 | n18605 ;
  assign n18607 = n18602 | n18606 ;
  assign n18608 = n2432 | n18602 ;
  assign n18609 = n18606 | n18608 ;
  assign n18610 = ( n8656 & n18607 ) | ( n8656 & n18609 ) | ( n18607 & n18609 ) ;
  assign n18611 = x23 & n18609 ;
  assign n18612 = x23 & n18602 ;
  assign n18613 = ( x23 & n18606 ) | ( x23 & n18612 ) | ( n18606 & n18612 ) ;
  assign n18614 = ( n8656 & n18611 ) | ( n8656 & n18613 ) | ( n18611 & n18613 ) ;
  assign n18615 = x23 & ~n18613 ;
  assign n18616 = x23 & ~n18609 ;
  assign n18617 = ( ~n8656 & n18615 ) | ( ~n8656 & n18616 ) | ( n18615 & n18616 ) ;
  assign n18618 = ( n18610 & ~n18614 ) | ( n18610 & n18617 ) | ( ~n18614 & n18617 ) ;
  assign n18619 = n18601 & n18618 ;
  assign n18620 = n18601 & ~n18619 ;
  assign n18621 = ~n18601 & n18618 ;
  assign n18622 = n18620 | n18621 ;
  assign n18623 = n18049 | n18053 ;
  assign n18624 = n18049 | n18050 ;
  assign n18625 = ( n17501 & n18623 ) | ( n17501 & n18624 ) | ( n18623 & n18624 ) ;
  assign n18626 = n18622 & n18625 ;
  assign n18627 = n18622 | n18625 ;
  assign n18628 = ~n18626 & n18627 ;
  assign n18629 = x109 & n1859 ;
  assign n18630 = x108 & n1854 ;
  assign n18631 = x107 & ~n1853 ;
  assign n18632 = n2037 & n18631 ;
  assign n18633 = n18630 | n18632 ;
  assign n18634 = n18629 | n18633 ;
  assign n18635 = n1862 | n18629 ;
  assign n18636 = n18633 | n18635 ;
  assign n18637 = ( n9878 & n18634 ) | ( n9878 & n18636 ) | ( n18634 & n18636 ) ;
  assign n18638 = x20 & n18636 ;
  assign n18639 = x20 & n18629 ;
  assign n18640 = ( x20 & n18633 ) | ( x20 & n18639 ) | ( n18633 & n18639 ) ;
  assign n18641 = ( n9878 & n18638 ) | ( n9878 & n18640 ) | ( n18638 & n18640 ) ;
  assign n18642 = x20 & ~n18640 ;
  assign n18643 = x20 & ~n18636 ;
  assign n18644 = ( ~n9878 & n18642 ) | ( ~n9878 & n18643 ) | ( n18642 & n18643 ) ;
  assign n18645 = ( n18637 & ~n18641 ) | ( n18637 & n18644 ) | ( ~n18641 & n18644 ) ;
  assign n18646 = n18628 & n18645 ;
  assign n18647 = n18628 & ~n18646 ;
  assign n18648 = ~n18628 & n18645 ;
  assign n18649 = n18647 | n18648 ;
  assign n18650 = n18077 | n18081 ;
  assign n18651 = ( n18077 & n18083 ) | ( n18077 & n18650 ) | ( n18083 & n18650 ) ;
  assign n18652 = n18649 & n18651 ;
  assign n18653 = n18649 | n18651 ;
  assign n18654 = ~n18652 & n18653 ;
  assign n18655 = x112 & n1383 ;
  assign n18656 = x111 & n1378 ;
  assign n18657 = x110 & ~n1377 ;
  assign n18658 = n1542 & n18657 ;
  assign n18659 = n18656 | n18658 ;
  assign n18660 = n18655 | n18659 ;
  assign n18661 = n1386 | n18655 ;
  assign n18662 = n18659 | n18661 ;
  assign n18663 = ( n11172 & n18660 ) | ( n11172 & n18662 ) | ( n18660 & n18662 ) ;
  assign n18664 = x17 & n18662 ;
  assign n18665 = x17 & n18655 ;
  assign n18666 = ( x17 & n18659 ) | ( x17 & n18665 ) | ( n18659 & n18665 ) ;
  assign n18667 = ( n11172 & n18664 ) | ( n11172 & n18666 ) | ( n18664 & n18666 ) ;
  assign n18668 = x17 & ~n18666 ;
  assign n18669 = x17 & ~n18662 ;
  assign n18670 = ( ~n11172 & n18668 ) | ( ~n11172 & n18669 ) | ( n18668 & n18669 ) ;
  assign n18671 = ( n18663 & ~n18667 ) | ( n18663 & n18670 ) | ( ~n18667 & n18670 ) ;
  assign n18672 = n18654 & n18671 ;
  assign n18673 = n18654 & ~n18672 ;
  assign n18674 = ~n18654 & n18671 ;
  assign n18675 = n18673 | n18674 ;
  assign n18676 = n18104 | n18106 ;
  assign n18677 = ( n18104 & n18108 ) | ( n18104 & n18676 ) | ( n18108 & n18676 ) ;
  assign n18678 = n18675 & n18677 ;
  assign n18679 = n18675 | n18677 ;
  assign n18680 = ~n18678 & n18679 ;
  assign n18681 = x115 & n962 ;
  assign n18682 = x114 & n957 ;
  assign n18683 = x113 & ~n956 ;
  assign n18684 = n1105 & n18683 ;
  assign n18685 = n18682 | n18684 ;
  assign n18686 = n18681 | n18685 ;
  assign n18687 = n965 | n18681 ;
  assign n18688 = n18685 | n18687 ;
  assign n18689 = ( ~n12550 & n18686 ) | ( ~n12550 & n18688 ) | ( n18686 & n18688 ) ;
  assign n18690 = n18686 & n18688 ;
  assign n18691 = ( n12532 & n18689 ) | ( n12532 & n18690 ) | ( n18689 & n18690 ) ;
  assign n18692 = x14 & n18691 ;
  assign n18693 = x14 & ~n18691 ;
  assign n18694 = ( n18691 & ~n18692 ) | ( n18691 & n18693 ) | ( ~n18692 & n18693 ) ;
  assign n18695 = n18680 & n18694 ;
  assign n18696 = n18680 | n18694 ;
  assign n18697 = ~n18695 & n18696 ;
  assign n18698 = ( n18111 & n18125 ) | ( n18111 & n18131 ) | ( n18125 & n18131 ) ;
  assign n18699 = n18697 | n18698 ;
  assign n18700 = n18697 & n18698 ;
  assign n18701 = n18699 & ~n18700 ;
  assign n18702 = x118 & n636 ;
  assign n18703 = x117 & n631 ;
  assign n18704 = x116 & ~n630 ;
  assign n18705 = n764 & n18704 ;
  assign n18706 = n18703 | n18705 ;
  assign n18707 = n18702 | n18706 ;
  assign n18708 = n639 | n18702 ;
  assign n18709 = n18706 | n18708 ;
  assign n18710 = ( ~n14002 & n18707 ) | ( ~n14002 & n18709 ) | ( n18707 & n18709 ) ;
  assign n18711 = n18707 & n18709 ;
  assign n18712 = ( n13981 & n18710 ) | ( n13981 & n18711 ) | ( n18710 & n18711 ) ;
  assign n18713 = x11 & n18712 ;
  assign n18714 = x11 & ~n18712 ;
  assign n18715 = ( n18712 & ~n18713 ) | ( n18712 & n18714 ) | ( ~n18713 & n18714 ) ;
  assign n18716 = n18701 & n18715 ;
  assign n18717 = n18701 & ~n18716 ;
  assign n18718 = ~n18701 & n18715 ;
  assign n18719 = n18717 | n18718 ;
  assign n18720 = n18149 | n18151 ;
  assign n18721 = ( n18149 & n18153 ) | ( n18149 & n18720 ) | ( n18153 & n18720 ) ;
  assign n18722 = n18719 | n18721 ;
  assign n18723 = n18719 & n18721 ;
  assign n18724 = n18722 & ~n18723 ;
  assign n18725 = x121 & n389 ;
  assign n18726 = x120 & n384 ;
  assign n18727 = x119 & ~n383 ;
  assign n18728 = n463 & n18727 ;
  assign n18729 = n18726 | n18728 ;
  assign n18730 = n18725 | n18729 ;
  assign n18731 = n392 | n18725 ;
  assign n18732 = n18729 | n18731 ;
  assign n18733 = ( n15501 & n18730 ) | ( n15501 & n18732 ) | ( n18730 & n18732 ) ;
  assign n18734 = x8 & n18732 ;
  assign n18735 = x8 & n18725 ;
  assign n18736 = ( x8 & n18729 ) | ( x8 & n18735 ) | ( n18729 & n18735 ) ;
  assign n18737 = ( n15501 & n18734 ) | ( n15501 & n18736 ) | ( n18734 & n18736 ) ;
  assign n18738 = x8 & ~n18736 ;
  assign n18739 = x8 & ~n18732 ;
  assign n18740 = ( ~n15501 & n18738 ) | ( ~n15501 & n18739 ) | ( n18738 & n18739 ) ;
  assign n18741 = ( n18733 & ~n18737 ) | ( n18733 & n18740 ) | ( ~n18737 & n18740 ) ;
  assign n18742 = ( n18270 & n18724 ) | ( n18270 & ~n18741 ) | ( n18724 & ~n18741 ) ;
  assign n18743 = ( ~n18724 & n18741 ) | ( ~n18724 & n18742 ) | ( n18741 & n18742 ) ;
  assign n18744 = ( ~n18270 & n18742 ) | ( ~n18270 & n18743 ) | ( n18742 & n18743 ) ;
  assign n18745 = ( n18175 & n18176 ) | ( n18175 & n18197 ) | ( n18176 & n18197 ) ;
  assign n18746 = n18744 | n18745 ;
  assign n18747 = n18744 & n18745 ;
  assign n18748 = n18746 & ~n18747 ;
  assign n18749 = x126 & ~x127 ;
  assign n18750 = ~x126 & x127 ;
  assign n18751 = n18749 | n18750 ;
  assign n18752 = n18201 & n18751 ;
  assign n18753 = ( n18202 & n18751 ) | ( n18202 & n18752 ) | ( n18751 & n18752 ) ;
  assign n18754 = n18751 & n18752 ;
  assign n18755 = ( n18214 & n18753 ) | ( n18214 & n18754 ) | ( n18753 & n18754 ) ;
  assign n18756 = ( n18212 & n18753 ) | ( n18212 & n18754 ) | ( n18753 & n18754 ) ;
  assign n18757 = ( n14002 & n18755 ) | ( n14002 & n18756 ) | ( n18755 & n18756 ) ;
  assign n18758 = n18201 | n18751 ;
  assign n18759 = n18202 | n18758 ;
  assign n18760 = ( n18214 & n18758 ) | ( n18214 & n18759 ) | ( n18758 & n18759 ) ;
  assign n18761 = ( n18212 & n18758 ) | ( n18212 & n18759 ) | ( n18758 & n18759 ) ;
  assign n18762 = ( n14002 & n18760 ) | ( n14002 & n18761 ) | ( n18760 & n18761 ) ;
  assign n18763 = ~n18757 & n18762 ;
  assign n18764 = x126 & n133 ;
  assign n18765 = x125 & ~n162 ;
  assign n18766 = ( n137 & n18764 ) | ( n137 & n18765 ) | ( n18764 & n18765 ) ;
  assign n18767 = x0 & x127 ;
  assign n18768 = ( ~n137 & n18764 ) | ( ~n137 & n18767 ) | ( n18764 & n18767 ) ;
  assign n18769 = n18766 | n18768 ;
  assign n18770 = n141 | n18769 ;
  assign n18771 = ( n18763 & n18769 ) | ( n18763 & n18770 ) | ( n18769 & n18770 ) ;
  assign n18772 = x2 & n18769 ;
  assign n18773 = ( x2 & n523 ) | ( x2 & n18769 ) | ( n523 & n18769 ) ;
  assign n18774 = ( n18763 & n18772 ) | ( n18763 & n18773 ) | ( n18772 & n18773 ) ;
  assign n18775 = x2 & ~n18773 ;
  assign n18776 = x2 & ~n18769 ;
  assign n18777 = ( ~n18763 & n18775 ) | ( ~n18763 & n18776 ) | ( n18775 & n18776 ) ;
  assign n18778 = ( n18771 & ~n18774 ) | ( n18771 & n18777 ) | ( ~n18774 & n18777 ) ;
  assign n18779 = ~n18748 & n18778 ;
  assign n18780 = n18197 | n18778 ;
  assign n18781 = n18175 | n18778 ;
  assign n18782 = ( n18176 & n18780 ) | ( n18176 & n18781 ) | ( n18780 & n18781 ) ;
  assign n18783 = ( n18744 & n18778 ) | ( n18744 & n18782 ) | ( n18778 & n18782 ) ;
  assign n18784 = n18746 & ~n18783 ;
  assign n18785 = n18779 | n18784 ;
  assign n18786 = n18199 | n18239 ;
  assign n18787 = n18785 & n18786 ;
  assign n18788 = n18785 | n18786 ;
  assign n18789 = ~n18787 & n18788 ;
  assign n18790 = n18244 | n18252 ;
  assign n18791 = n18789 | n18790 ;
  assign n18792 = n18244 & n18789 ;
  assign n18793 = ( n18252 & n18789 ) | ( n18252 & n18792 ) | ( n18789 & n18792 ) ;
  assign n18794 = n18791 & ~n18793 ;
  assign n18795 = x107 & n2429 ;
  assign n18796 = x106 & n2424 ;
  assign n18797 = x105 & ~n2423 ;
  assign n18798 = n2631 & n18797 ;
  assign n18799 = n18796 | n18798 ;
  assign n18800 = n18795 | n18799 ;
  assign n18801 = n2432 | n18795 ;
  assign n18802 = n18799 | n18801 ;
  assign n18803 = ( n9084 & n18800 ) | ( n9084 & n18802 ) | ( n18800 & n18802 ) ;
  assign n18804 = x23 & n18802 ;
  assign n18805 = x23 & n18795 ;
  assign n18806 = ( x23 & n18799 ) | ( x23 & n18805 ) | ( n18799 & n18805 ) ;
  assign n18807 = ( n9084 & n18804 ) | ( n9084 & n18806 ) | ( n18804 & n18806 ) ;
  assign n18808 = x23 & ~n18806 ;
  assign n18809 = x23 & ~n18802 ;
  assign n18810 = ( ~n9084 & n18808 ) | ( ~n9084 & n18809 ) | ( n18808 & n18809 ) ;
  assign n18811 = ( n18803 & ~n18807 ) | ( n18803 & n18810 ) | ( ~n18807 & n18810 ) ;
  assign n18812 = n241 & n17149 ;
  assign n18813 = x68 & n17146 ;
  assign n18814 = x67 & n17141 ;
  assign n18815 = x66 & ~n17140 ;
  assign n18816 = n17724 & n18815 ;
  assign n18817 = n18814 | n18816 ;
  assign n18818 = n18813 | n18817 ;
  assign n18819 = n18812 | n18818 ;
  assign n18820 = x62 | n18813 ;
  assign n18821 = n18817 | n18820 ;
  assign n18822 = n18812 | n18821 ;
  assign n18823 = ~x62 & n18821 ;
  assign n18824 = ( ~x62 & n18812 ) | ( ~x62 & n18823 ) | ( n18812 & n18823 ) ;
  assign n18825 = ( ~n18819 & n18822 ) | ( ~n18819 & n18824 ) | ( n18822 & n18824 ) ;
  assign n18826 = x65 & n18290 ;
  assign n18827 = x63 & x64 ;
  assign n18828 = ~n18290 & n18827 ;
  assign n18829 = n18826 | n18828 ;
  assign n18830 = n18821 & n18829 ;
  assign n18831 = ( n18812 & n18829 ) | ( n18812 & n18830 ) | ( n18829 & n18830 ) ;
  assign n18832 = ~n18818 & n18829 ;
  assign n18833 = ~n18812 & n18832 ;
  assign n18834 = ( n18824 & n18831 ) | ( n18824 & n18833 ) | ( n18831 & n18833 ) ;
  assign n18835 = n18825 & ~n18834 ;
  assign n18836 = ~n18821 & n18829 ;
  assign n18837 = ~n18812 & n18836 ;
  assign n18838 = n18818 & n18829 ;
  assign n18839 = ( n18812 & n18829 ) | ( n18812 & n18838 ) | ( n18829 & n18838 ) ;
  assign n18840 = ( ~n18824 & n18837 ) | ( ~n18824 & n18839 ) | ( n18837 & n18839 ) ;
  assign n18841 = n18835 | n18840 ;
  assign n18842 = n18293 | n18309 ;
  assign n18843 = n18841 | n18842 ;
  assign n18844 = n18841 & n18842 ;
  assign n18845 = n18843 & ~n18844 ;
  assign n18846 = x70 & n15547 ;
  assign n18847 = x69 & ~n15546 ;
  assign n18848 = n16123 & n18847 ;
  assign n18849 = n18846 | n18848 ;
  assign n18850 = x71 & n15552 ;
  assign n18851 = n15555 | n18850 ;
  assign n18852 = n18849 | n18851 ;
  assign n18853 = x59 & ~n18852 ;
  assign n18854 = x59 & ~n18850 ;
  assign n18855 = ~n18849 & n18854 ;
  assign n18856 = ( ~n438 & n18853 ) | ( ~n438 & n18855 ) | ( n18853 & n18855 ) ;
  assign n18857 = ~x59 & n18852 ;
  assign n18858 = ~x59 & n18850 ;
  assign n18859 = ( ~x59 & n18849 ) | ( ~x59 & n18858 ) | ( n18849 & n18858 ) ;
  assign n18860 = ( n438 & n18857 ) | ( n438 & n18859 ) | ( n18857 & n18859 ) ;
  assign n18861 = n18856 | n18860 ;
  assign n18862 = n18845 | n18861 ;
  assign n18863 = n18845 & n18861 ;
  assign n18864 = n18862 & ~n18863 ;
  assign n18865 = n18314 | n18316 ;
  assign n18866 = n18864 & n18865 ;
  assign n18867 = n18864 | n18865 ;
  assign n18868 = ~n18866 & n18867 ;
  assign n18869 = x74 & n14045 ;
  assign n18870 = x73 & n14040 ;
  assign n18871 = x72 & ~n14039 ;
  assign n18872 = n14552 & n18871 ;
  assign n18873 = n18870 | n18872 ;
  assign n18874 = n18869 | n18873 ;
  assign n18875 = n14048 | n18869 ;
  assign n18876 = n18873 | n18875 ;
  assign n18877 = ( n710 & n18874 ) | ( n710 & n18876 ) | ( n18874 & n18876 ) ;
  assign n18878 = x56 & n18876 ;
  assign n18879 = x56 & n18869 ;
  assign n18880 = ( x56 & n18873 ) | ( x56 & n18879 ) | ( n18873 & n18879 ) ;
  assign n18881 = ( n710 & n18878 ) | ( n710 & n18880 ) | ( n18878 & n18880 ) ;
  assign n18882 = x56 & ~n18880 ;
  assign n18883 = x56 & ~n18876 ;
  assign n18884 = ( ~n710 & n18882 ) | ( ~n710 & n18883 ) | ( n18882 & n18883 ) ;
  assign n18885 = ( n18877 & ~n18881 ) | ( n18877 & n18884 ) | ( ~n18881 & n18884 ) ;
  assign n18886 = n18868 & n18885 ;
  assign n18887 = n18868 & ~n18886 ;
  assign n18888 = ( n18318 & n18334 ) | ( n18318 & n18340 ) | ( n18334 & n18340 ) ;
  assign n18889 = ~n18868 & n18885 ;
  assign n18890 = n18888 & n18889 ;
  assign n18891 = ( n18887 & n18888 ) | ( n18887 & n18890 ) | ( n18888 & n18890 ) ;
  assign n18892 = n18888 | n18889 ;
  assign n18893 = n18887 | n18892 ;
  assign n18894 = ~n18891 & n18893 ;
  assign n18895 = x77 & n12574 ;
  assign n18896 = x76 & n12569 ;
  assign n18897 = x75 & ~n12568 ;
  assign n18898 = n13076 & n18897 ;
  assign n18899 = n18896 | n18898 ;
  assign n18900 = n18895 | n18899 ;
  assign n18901 = n12577 | n18895 ;
  assign n18902 = n18899 | n18901 ;
  assign n18903 = ( n1059 & n18900 ) | ( n1059 & n18902 ) | ( n18900 & n18902 ) ;
  assign n18904 = x53 & n18902 ;
  assign n18905 = x53 & n18895 ;
  assign n18906 = ( x53 & n18899 ) | ( x53 & n18905 ) | ( n18899 & n18905 ) ;
  assign n18907 = ( n1059 & n18904 ) | ( n1059 & n18906 ) | ( n18904 & n18906 ) ;
  assign n18908 = x53 & ~n18906 ;
  assign n18909 = x53 & ~n18902 ;
  assign n18910 = ( ~n1059 & n18908 ) | ( ~n1059 & n18909 ) | ( n18908 & n18909 ) ;
  assign n18911 = ( n18903 & ~n18907 ) | ( n18903 & n18910 ) | ( ~n18907 & n18910 ) ;
  assign n18912 = n18894 | n18911 ;
  assign n18913 = n18894 & n18911 ;
  assign n18914 = n18912 & ~n18913 ;
  assign n18915 = n18362 | n18366 ;
  assign n18916 = n18914 & n18915 ;
  assign n18917 = n18914 | n18915 ;
  assign n18918 = ~n18916 & n18917 ;
  assign n18919 = x80 & n11205 ;
  assign n18920 = x79 & n11200 ;
  assign n18921 = x78 & ~n11199 ;
  assign n18922 = n11679 & n18921 ;
  assign n18923 = n18920 | n18922 ;
  assign n18924 = n18919 | n18923 ;
  assign n18925 = n11208 | n18919 ;
  assign n18926 = n18923 | n18925 ;
  assign n18927 = ( n1499 & n18924 ) | ( n1499 & n18926 ) | ( n18924 & n18926 ) ;
  assign n18928 = x50 & n18926 ;
  assign n18929 = x50 & n18919 ;
  assign n18930 = ( x50 & n18923 ) | ( x50 & n18929 ) | ( n18923 & n18929 ) ;
  assign n18931 = ( n1499 & n18928 ) | ( n1499 & n18930 ) | ( n18928 & n18930 ) ;
  assign n18932 = x50 & ~n18930 ;
  assign n18933 = x50 & ~n18926 ;
  assign n18934 = ( ~n1499 & n18932 ) | ( ~n1499 & n18933 ) | ( n18932 & n18933 ) ;
  assign n18935 = ( n18927 & ~n18931 ) | ( n18927 & n18934 ) | ( ~n18931 & n18934 ) ;
  assign n18936 = n18918 & n18935 ;
  assign n18937 = n18918 & ~n18936 ;
  assign n18938 = ~n18918 & n18935 ;
  assign n18939 = n18937 | n18938 ;
  assign n18940 = n18386 | n18393 ;
  assign n18941 = n18939 | n18940 ;
  assign n18942 = n18939 & n18940 ;
  assign n18943 = n18941 & ~n18942 ;
  assign n18944 = x83 & n9933 ;
  assign n18945 = x82 & n9928 ;
  assign n18946 = x81 & ~n9927 ;
  assign n18947 = n10379 & n18946 ;
  assign n18948 = n18945 | n18947 ;
  assign n18949 = n18944 | n18948 ;
  assign n18950 = n9936 | n18944 ;
  assign n18951 = n18948 | n18950 ;
  assign n18952 = ( n2009 & n18949 ) | ( n2009 & n18951 ) | ( n18949 & n18951 ) ;
  assign n18953 = x47 & n18951 ;
  assign n18954 = x47 & n18944 ;
  assign n18955 = ( x47 & n18948 ) | ( x47 & n18954 ) | ( n18948 & n18954 ) ;
  assign n18956 = ( n2009 & n18953 ) | ( n2009 & n18955 ) | ( n18953 & n18955 ) ;
  assign n18957 = x47 & ~n18955 ;
  assign n18958 = x47 & ~n18951 ;
  assign n18959 = ( ~n2009 & n18957 ) | ( ~n2009 & n18958 ) | ( n18957 & n18958 ) ;
  assign n18960 = ( n18952 & ~n18956 ) | ( n18952 & n18959 ) | ( ~n18956 & n18959 ) ;
  assign n18961 = n18943 | n18960 ;
  assign n18962 = n18943 & n18960 ;
  assign n18963 = n18961 & ~n18962 ;
  assign n18964 = n18413 | n18414 ;
  assign n18965 = ( n18413 & n18416 ) | ( n18413 & n18964 ) | ( n18416 & n18964 ) ;
  assign n18966 = n18963 & n18965 ;
  assign n18967 = n18963 | n18965 ;
  assign n18968 = ~n18966 & n18967 ;
  assign n18969 = x86 & n8724 ;
  assign n18970 = x85 & n8719 ;
  assign n18971 = x84 & ~n8718 ;
  assign n18972 = n9149 & n18971 ;
  assign n18973 = n18970 | n18972 ;
  assign n18974 = n18969 | n18973 ;
  assign n18975 = n8727 | n18969 ;
  assign n18976 = n18973 | n18975 ;
  assign n18977 = ( n2606 & n18974 ) | ( n2606 & n18976 ) | ( n18974 & n18976 ) ;
  assign n18978 = x44 & n18976 ;
  assign n18979 = x44 & n18969 ;
  assign n18980 = ( x44 & n18973 ) | ( x44 & n18979 ) | ( n18973 & n18979 ) ;
  assign n18981 = ( n2606 & n18978 ) | ( n2606 & n18980 ) | ( n18978 & n18980 ) ;
  assign n18982 = x44 & ~n18980 ;
  assign n18983 = x44 & ~n18976 ;
  assign n18984 = ( ~n2606 & n18982 ) | ( ~n2606 & n18983 ) | ( n18982 & n18983 ) ;
  assign n18985 = ( n18977 & ~n18981 ) | ( n18977 & n18984 ) | ( ~n18981 & n18984 ) ;
  assign n18986 = n18968 & n18985 ;
  assign n18987 = n18968 & ~n18986 ;
  assign n18988 = ~n18968 & n18985 ;
  assign n18989 = n18987 | n18988 ;
  assign n18990 = n18437 | n18442 ;
  assign n18991 = n18989 | n18990 ;
  assign n18992 = n18989 & n18990 ;
  assign n18993 = n18991 & ~n18992 ;
  assign n18994 = x89 & n7566 ;
  assign n18995 = x88 & n7561 ;
  assign n18996 = x87 & ~n7560 ;
  assign n18997 = n7953 & n18996 ;
  assign n18998 = n18995 | n18997 ;
  assign n18999 = n18994 | n18998 ;
  assign n19000 = n7569 | n18994 ;
  assign n19001 = n18998 | n19000 ;
  assign n19002 = ( n3282 & n18999 ) | ( n3282 & n19001 ) | ( n18999 & n19001 ) ;
  assign n19003 = x41 & n19001 ;
  assign n19004 = x41 & n18994 ;
  assign n19005 = ( x41 & n18998 ) | ( x41 & n19004 ) | ( n18998 & n19004 ) ;
  assign n19006 = ( n3282 & n19003 ) | ( n3282 & n19005 ) | ( n19003 & n19005 ) ;
  assign n19007 = x41 & ~n19005 ;
  assign n19008 = x41 & ~n19001 ;
  assign n19009 = ( ~n3282 & n19007 ) | ( ~n3282 & n19008 ) | ( n19007 & n19008 ) ;
  assign n19010 = ( n19002 & ~n19006 ) | ( n19002 & n19009 ) | ( ~n19006 & n19009 ) ;
  assign n19011 = n18993 & n19010 ;
  assign n19012 = n18993 & ~n19011 ;
  assign n19013 = ~n18993 & n19010 ;
  assign n19014 = n19012 | n19013 ;
  assign n19015 = n18467 | n18469 ;
  assign n19016 = n18468 | n19015 ;
  assign n19017 = ( n18467 & n18471 ) | ( n18467 & n19016 ) | ( n18471 & n19016 ) ;
  assign n19018 = n19014 | n19017 ;
  assign n19019 = n19014 & n19017 ;
  assign n19020 = n19018 & ~n19019 ;
  assign n19021 = x92 & n6536 ;
  assign n19022 = x91 & n6531 ;
  assign n19023 = x90 & ~n6530 ;
  assign n19024 = n6871 & n19023 ;
  assign n19025 = n19022 | n19024 ;
  assign n19026 = n19021 | n19025 ;
  assign n19027 = n6539 | n19021 ;
  assign n19028 = n19025 | n19027 ;
  assign n19029 = ( n4040 & n19026 ) | ( n4040 & n19028 ) | ( n19026 & n19028 ) ;
  assign n19030 = x38 & n19028 ;
  assign n19031 = x38 & n19021 ;
  assign n19032 = ( x38 & n19025 ) | ( x38 & n19031 ) | ( n19025 & n19031 ) ;
  assign n19033 = ( n4040 & n19030 ) | ( n4040 & n19032 ) | ( n19030 & n19032 ) ;
  assign n19034 = x38 & ~n19032 ;
  assign n19035 = x38 & ~n19028 ;
  assign n19036 = ( ~n4040 & n19034 ) | ( ~n4040 & n19035 ) | ( n19034 & n19035 ) ;
  assign n19037 = ( n19029 & ~n19033 ) | ( n19029 & n19036 ) | ( ~n19033 & n19036 ) ;
  assign n19038 = n19020 & n19037 ;
  assign n19039 = n19020 & ~n19038 ;
  assign n19040 = ~n19020 & n19037 ;
  assign n19041 = n19039 | n19040 ;
  assign n19042 = n18492 | n18498 ;
  assign n19043 = n19041 | n19042 ;
  assign n19044 = n19041 & n19042 ;
  assign n19045 = n19043 & ~n19044 ;
  assign n19046 = x95 & n5554 ;
  assign n19047 = x94 & n5549 ;
  assign n19048 = x93 & ~n5548 ;
  assign n19049 = n5893 & n19048 ;
  assign n19050 = n19047 | n19049 ;
  assign n19051 = n19046 | n19050 ;
  assign n19052 = n5557 | n19046 ;
  assign n19053 = n19050 | n19052 ;
  assign n19054 = ( n4897 & n19051 ) | ( n4897 & n19053 ) | ( n19051 & n19053 ) ;
  assign n19055 = x35 & n19053 ;
  assign n19056 = x35 & n19046 ;
  assign n19057 = ( x35 & n19050 ) | ( x35 & n19056 ) | ( n19050 & n19056 ) ;
  assign n19058 = ( n4897 & n19055 ) | ( n4897 & n19057 ) | ( n19055 & n19057 ) ;
  assign n19059 = x35 & ~n19057 ;
  assign n19060 = x35 & ~n19053 ;
  assign n19061 = ( ~n4897 & n19059 ) | ( ~n4897 & n19060 ) | ( n19059 & n19060 ) ;
  assign n19062 = ( n19054 & ~n19058 ) | ( n19054 & n19061 ) | ( ~n19058 & n19061 ) ;
  assign n19063 = n19045 | n19062 ;
  assign n19064 = n19045 & n19062 ;
  assign n19065 = n19063 & ~n19064 ;
  assign n19066 = n18518 | n18519 ;
  assign n19067 = n17953 | n18518 ;
  assign n19068 = ( n18520 & n19066 ) | ( n18520 & n19067 ) | ( n19066 & n19067 ) ;
  assign n19069 = n19065 & n19068 ;
  assign n19070 = n19065 | n19068 ;
  assign n19071 = ~n19069 & n19070 ;
  assign n19072 = x98 & n4631 ;
  assign n19073 = x97 & n4626 ;
  assign n19074 = x96 & ~n4625 ;
  assign n19075 = n4943 & n19074 ;
  assign n19076 = n19073 | n19075 ;
  assign n19077 = n19072 | n19076 ;
  assign n19078 = n4634 | n19072 ;
  assign n19079 = n19076 | n19078 ;
  assign n19080 = ( ~n5850 & n19077 ) | ( ~n5850 & n19079 ) | ( n19077 & n19079 ) ;
  assign n19081 = n19077 & n19079 ;
  assign n19082 = ( n5834 & n19080 ) | ( n5834 & n19081 ) | ( n19080 & n19081 ) ;
  assign n19083 = x32 & n19079 ;
  assign n19084 = x32 & n19072 ;
  assign n19085 = ( x32 & n19076 ) | ( x32 & n19084 ) | ( n19076 & n19084 ) ;
  assign n19086 = ( ~n5850 & n19083 ) | ( ~n5850 & n19085 ) | ( n19083 & n19085 ) ;
  assign n19087 = n19083 & n19085 ;
  assign n19088 = ( n5834 & n19086 ) | ( n5834 & n19087 ) | ( n19086 & n19087 ) ;
  assign n19089 = x32 & ~n19085 ;
  assign n19090 = x32 & ~n19079 ;
  assign n19091 = ( n5850 & n19089 ) | ( n5850 & n19090 ) | ( n19089 & n19090 ) ;
  assign n19092 = n19089 | n19090 ;
  assign n19093 = ( ~n5834 & n19091 ) | ( ~n5834 & n19092 ) | ( n19091 & n19092 ) ;
  assign n19094 = ( n19082 & ~n19088 ) | ( n19082 & n19093 ) | ( ~n19088 & n19093 ) ;
  assign n19095 = n19071 & n19094 ;
  assign n19096 = n19071 & ~n19095 ;
  assign n19097 = ( n18524 & n18541 ) | ( n18524 & n18546 ) | ( n18541 & n18546 ) ;
  assign n19098 = ~n19071 & n19094 ;
  assign n19099 = n19097 & n19098 ;
  assign n19100 = ( n19096 & n19097 ) | ( n19096 & n19099 ) | ( n19097 & n19099 ) ;
  assign n19101 = n19097 | n19098 ;
  assign n19102 = n19096 | n19101 ;
  assign n19103 = ~n19100 & n19102 ;
  assign n19104 = x101 & n3816 ;
  assign n19105 = x100 & n3811 ;
  assign n19106 = x99 & ~n3810 ;
  assign n19107 = n4067 & n19106 ;
  assign n19108 = n19105 | n19107 ;
  assign n19109 = n19104 | n19108 ;
  assign n19110 = n3819 | n19104 ;
  assign n19111 = n19108 | n19110 ;
  assign n19112 = ( n6844 & n19109 ) | ( n6844 & n19111 ) | ( n19109 & n19111 ) ;
  assign n19113 = x29 & n19111 ;
  assign n19114 = x29 & n19104 ;
  assign n19115 = ( x29 & n19108 ) | ( x29 & n19114 ) | ( n19108 & n19114 ) ;
  assign n19116 = ( n6844 & n19113 ) | ( n6844 & n19115 ) | ( n19113 & n19115 ) ;
  assign n19117 = x29 & ~n19115 ;
  assign n19118 = x29 & ~n19111 ;
  assign n19119 = ( ~n6844 & n19117 ) | ( ~n6844 & n19118 ) | ( n19117 & n19118 ) ;
  assign n19120 = ( n19112 & ~n19116 ) | ( n19112 & n19119 ) | ( ~n19116 & n19119 ) ;
  assign n19121 = n19103 & n19120 ;
  assign n19122 = n19103 & ~n19121 ;
  assign n19123 = ~n19103 & n19120 ;
  assign n19124 = n19122 | n19123 ;
  assign n19125 = n18569 | n18571 ;
  assign n19126 = ( n18569 & n18573 ) | ( n18569 & n19125 ) | ( n18573 & n19125 ) ;
  assign n19127 = n19124 | n19126 ;
  assign n19128 = n19124 & n19126 ;
  assign n19129 = n19127 & ~n19128 ;
  assign n19130 = x104 & n3085 ;
  assign n19131 = x103 & n3080 ;
  assign n19132 = x102 & ~n3079 ;
  assign n19133 = n3309 & n19132 ;
  assign n19134 = n19131 | n19133 ;
  assign n19135 = n19130 | n19134 ;
  assign n19136 = n3088 | n19130 ;
  assign n19137 = n19134 | n19136 ;
  assign n19138 = ( n7911 & n19135 ) | ( n7911 & n19137 ) | ( n19135 & n19137 ) ;
  assign n19139 = x26 & n19137 ;
  assign n19140 = x26 & n19130 ;
  assign n19141 = ( x26 & n19134 ) | ( x26 & n19140 ) | ( n19134 & n19140 ) ;
  assign n19142 = ( n7911 & n19139 ) | ( n7911 & n19141 ) | ( n19139 & n19141 ) ;
  assign n19143 = x26 & ~n19141 ;
  assign n19144 = x26 & ~n19137 ;
  assign n19145 = ( ~n7911 & n19143 ) | ( ~n7911 & n19144 ) | ( n19143 & n19144 ) ;
  assign n19146 = ( n19138 & ~n19142 ) | ( n19138 & n19145 ) | ( ~n19142 & n19145 ) ;
  assign n19147 = n19129 & n19146 ;
  assign n19148 = n19129 & ~n19147 ;
  assign n19149 = ~n19129 & n19146 ;
  assign n19150 = n19148 | n19149 ;
  assign n19151 = n18595 | n18598 ;
  assign n19152 = n19150 & ~n19151 ;
  assign n19153 = n18811 | n19150 ;
  assign n19154 = n19151 & ~n19153 ;
  assign n19155 = ( ~n18811 & n19152 ) | ( ~n18811 & n19154 ) | ( n19152 & n19154 ) ;
  assign n19156 = n18811 & n19150 ;
  assign n19157 = ( n18811 & ~n19151 ) | ( n18811 & n19156 ) | ( ~n19151 & n19156 ) ;
  assign n19158 = ~n19152 & n19157 ;
  assign n19159 = n19155 | n19158 ;
  assign n19160 = n18619 | n18625 ;
  assign n19161 = ( n18619 & n18622 ) | ( n18619 & n19160 ) | ( n18622 & n19160 ) ;
  assign n19162 = n19159 & n19161 ;
  assign n19163 = n19159 | n19161 ;
  assign n19164 = ~n19162 & n19163 ;
  assign n19165 = x110 & n1859 ;
  assign n19166 = x109 & n1854 ;
  assign n19167 = x108 & ~n1853 ;
  assign n19168 = n2037 & n19167 ;
  assign n19169 = n19166 | n19168 ;
  assign n19170 = n19165 | n19169 ;
  assign n19171 = n1862 | n19165 ;
  assign n19172 = n19169 | n19171 ;
  assign n19173 = ( n10330 & n19170 ) | ( n10330 & n19172 ) | ( n19170 & n19172 ) ;
  assign n19174 = x20 & n19172 ;
  assign n19175 = x20 & n19165 ;
  assign n19176 = ( x20 & n19169 ) | ( x20 & n19175 ) | ( n19169 & n19175 ) ;
  assign n19177 = ( n10330 & n19174 ) | ( n10330 & n19176 ) | ( n19174 & n19176 ) ;
  assign n19178 = x20 & ~n19176 ;
  assign n19179 = x20 & ~n19172 ;
  assign n19180 = ( ~n10330 & n19178 ) | ( ~n10330 & n19179 ) | ( n19178 & n19179 ) ;
  assign n19181 = ( n19173 & ~n19177 ) | ( n19173 & n19180 ) | ( ~n19177 & n19180 ) ;
  assign n19182 = n19164 & n19181 ;
  assign n19183 = n19164 & ~n19182 ;
  assign n19184 = ~n19164 & n19181 ;
  assign n19185 = n19183 | n19184 ;
  assign n19186 = n18646 | n18651 ;
  assign n19187 = ( n18646 & n18649 ) | ( n18646 & n19186 ) | ( n18649 & n19186 ) ;
  assign n19188 = n19185 & n19187 ;
  assign n19189 = n19185 | n19187 ;
  assign n19190 = ~n19188 & n19189 ;
  assign n19191 = x113 & n1383 ;
  assign n19192 = x112 & n1378 ;
  assign n19193 = x111 & ~n1377 ;
  assign n19194 = n1542 & n19193 ;
  assign n19195 = n19192 | n19194 ;
  assign n19196 = n19191 | n19195 ;
  assign n19197 = n1386 | n19191 ;
  assign n19198 = n19195 | n19197 ;
  assign n19199 = ( ~n11642 & n19196 ) | ( ~n11642 & n19198 ) | ( n19196 & n19198 ) ;
  assign n19200 = n19196 & n19198 ;
  assign n19201 = ( n11626 & n19199 ) | ( n11626 & n19200 ) | ( n19199 & n19200 ) ;
  assign n19202 = x17 & n19201 ;
  assign n19203 = x17 & ~n19201 ;
  assign n19204 = ( n19201 & ~n19202 ) | ( n19201 & n19203 ) | ( ~n19202 & n19203 ) ;
  assign n19205 = n19190 & n19204 ;
  assign n19206 = n19190 & ~n19205 ;
  assign n19207 = ~n19190 & n19204 ;
  assign n19208 = n19206 | n19207 ;
  assign n19209 = n18672 | n18677 ;
  assign n19210 = ( n18672 & n18675 ) | ( n18672 & n19209 ) | ( n18675 & n19209 ) ;
  assign n19211 = n19208 & n19210 ;
  assign n19212 = n19208 | n19210 ;
  assign n19213 = ~n19211 & n19212 ;
  assign n19214 = x116 & n962 ;
  assign n19215 = x115 & n957 ;
  assign n19216 = x114 & ~n956 ;
  assign n19217 = n1105 & n19216 ;
  assign n19218 = n19215 | n19217 ;
  assign n19219 = n19214 | n19218 ;
  assign n19220 = n965 | n19214 ;
  assign n19221 = n19218 | n19220 ;
  assign n19222 = ( ~n13040 & n19219 ) | ( ~n13040 & n19221 ) | ( n19219 & n19221 ) ;
  assign n19223 = n19219 & n19221 ;
  assign n19224 = ( n13022 & n19222 ) | ( n13022 & n19223 ) | ( n19222 & n19223 ) ;
  assign n19225 = x14 & n19224 ;
  assign n19226 = x14 & ~n19224 ;
  assign n19227 = ( n19224 & ~n19225 ) | ( n19224 & n19226 ) | ( ~n19225 & n19226 ) ;
  assign n19228 = n19213 & n19227 ;
  assign n19229 = n19213 | n19227 ;
  assign n19230 = ~n19228 & n19229 ;
  assign n19231 = n18695 | n18700 ;
  assign n19232 = n19230 & n19231 ;
  assign n19233 = n19230 | n19231 ;
  assign n19234 = ~n19232 & n19233 ;
  assign n19235 = x119 & n636 ;
  assign n19236 = x118 & n631 ;
  assign n19237 = x117 & ~n630 ;
  assign n19238 = n764 & n19237 ;
  assign n19239 = n19236 | n19238 ;
  assign n19240 = n19235 | n19239 ;
  assign n19241 = n639 | n19235 ;
  assign n19242 = n19239 | n19241 ;
  assign n19243 = ( n14496 & n19240 ) | ( n14496 & n19242 ) | ( n19240 & n19242 ) ;
  assign n19244 = x11 & n19242 ;
  assign n19245 = x11 & n19235 ;
  assign n19246 = ( x11 & n19239 ) | ( x11 & n19245 ) | ( n19239 & n19245 ) ;
  assign n19247 = ( n14496 & n19244 ) | ( n14496 & n19246 ) | ( n19244 & n19246 ) ;
  assign n19248 = x11 & ~n19246 ;
  assign n19249 = x11 & ~n19242 ;
  assign n19250 = ( ~n14496 & n19248 ) | ( ~n14496 & n19249 ) | ( n19248 & n19249 ) ;
  assign n19251 = ( n19243 & ~n19247 ) | ( n19243 & n19250 ) | ( ~n19247 & n19250 ) ;
  assign n19252 = n19234 & n19251 ;
  assign n19253 = n19234 | n19251 ;
  assign n19254 = ~n19252 & n19253 ;
  assign n19255 = n18716 | n18723 ;
  assign n19256 = n19254 & n19255 ;
  assign n19257 = n19254 | n19255 ;
  assign n19258 = ~n19256 & n19257 ;
  assign n19259 = x122 & n389 ;
  assign n19260 = x121 & n384 ;
  assign n19261 = x120 & ~n383 ;
  assign n19262 = n463 & n19261 ;
  assign n19263 = n19260 | n19262 ;
  assign n19264 = n19259 | n19263 ;
  assign n19265 = n392 | n19259 ;
  assign n19266 = n19263 | n19265 ;
  assign n19267 = ( n16043 & n19264 ) | ( n16043 & n19266 ) | ( n19264 & n19266 ) ;
  assign n19268 = x8 & n19266 ;
  assign n19269 = x8 & n19259 ;
  assign n19270 = ( x8 & n19263 ) | ( x8 & n19269 ) | ( n19263 & n19269 ) ;
  assign n19271 = ( n16043 & n19268 ) | ( n16043 & n19270 ) | ( n19268 & n19270 ) ;
  assign n19272 = x8 & ~n19270 ;
  assign n19273 = x8 & ~n19266 ;
  assign n19274 = ( ~n16043 & n19272 ) | ( ~n16043 & n19273 ) | ( n19272 & n19273 ) ;
  assign n19275 = ( n19267 & ~n19271 ) | ( n19267 & n19274 ) | ( ~n19271 & n19274 ) ;
  assign n19276 = x125 & n212 ;
  assign n19277 = x124 & n207 ;
  assign n19278 = x123 & ~n206 ;
  assign n19279 = n267 & n19278 ;
  assign n19280 = n19277 | n19279 ;
  assign n19281 = n19276 | n19280 ;
  assign n19282 = n215 | n19276 ;
  assign n19283 = n19280 | n19282 ;
  assign n19284 = ( n17670 & n19281 ) | ( n17670 & n19283 ) | ( n19281 & n19283 ) ;
  assign n19285 = x5 & n19283 ;
  assign n19286 = x5 & n19276 ;
  assign n19287 = ( x5 & n19280 ) | ( x5 & n19286 ) | ( n19280 & n19286 ) ;
  assign n19288 = ( n17670 & n19285 ) | ( n17670 & n19287 ) | ( n19285 & n19287 ) ;
  assign n19289 = x5 & ~n19287 ;
  assign n19290 = x5 & ~n19283 ;
  assign n19291 = ( ~n17670 & n19289 ) | ( ~n17670 & n19290 ) | ( n19289 & n19290 ) ;
  assign n19292 = ( n19284 & ~n19288 ) | ( n19284 & n19291 ) | ( ~n19288 & n19291 ) ;
  assign n19293 = ( n19258 & ~n19275 ) | ( n19258 & n19292 ) | ( ~n19275 & n19292 ) ;
  assign n19294 = ( ~n19258 & n19275 ) | ( ~n19258 & n19293 ) | ( n19275 & n19293 ) ;
  assign n19295 = n18724 & n18741 ;
  assign n19296 = n18724 & ~n19295 ;
  assign n19297 = n18270 & ~n18741 ;
  assign n19298 = ( n18270 & n18724 ) | ( n18270 & n19297 ) | ( n18724 & n19297 ) ;
  assign n19299 = ( n18270 & n19295 ) | ( n18270 & ~n19298 ) | ( n19295 & ~n19298 ) ;
  assign n19300 = n18270 | n18741 ;
  assign n19301 = ( n18270 & n18724 ) | ( n18270 & n19300 ) | ( n18724 & n19300 ) ;
  assign n19302 = ( n19296 & n19299 ) | ( n19296 & n19301 ) | ( n19299 & n19301 ) ;
  assign n19303 = n19293 & n19302 ;
  assign n19304 = ~n19292 & n19302 ;
  assign n19305 = ( n19294 & n19303 ) | ( n19294 & n19304 ) | ( n19303 & n19304 ) ;
  assign n19306 = n19293 | n19302 ;
  assign n19307 = n19292 & ~n19302 ;
  assign n19308 = ( n19294 & n19306 ) | ( n19294 & ~n19307 ) | ( n19306 & ~n19307 ) ;
  assign n19309 = ~n19305 & n19308 ;
  assign n19310 = x127 & n133 ;
  assign n19311 = x126 & ~n162 ;
  assign n19312 = n137 & n19311 ;
  assign n19313 = n19310 | n19312 ;
  assign n19314 = n18201 & n18749 ;
  assign n19315 = ( n18202 & n18749 ) | ( n18202 & n19314 ) | ( n18749 & n19314 ) ;
  assign n19316 = n18749 & n19314 ;
  assign n19317 = ( n18214 & n19315 ) | ( n18214 & n19316 ) | ( n19315 & n19316 ) ;
  assign n19318 = ( n18212 & n19315 ) | ( n18212 & n19316 ) | ( n19315 & n19316 ) ;
  assign n19319 = ( n14002 & n19317 ) | ( n14002 & n19318 ) | ( n19317 & n19318 ) ;
  assign n19320 = x126 | n18201 ;
  assign n19321 = ( x126 & n18751 ) | ( x126 & n19320 ) | ( n18751 & n19320 ) ;
  assign n19322 = n18202 | n19321 ;
  assign n19323 = x127 & ~n19322 ;
  assign n19324 = x127 & ~n19321 ;
  assign n19325 = ( ~n18212 & n19323 ) | ( ~n18212 & n19324 ) | ( n19323 & n19324 ) ;
  assign n19326 = ( ~n18214 & n19323 ) | ( ~n18214 & n19324 ) | ( n19323 & n19324 ) ;
  assign n19327 = ( ~n14002 & n19325 ) | ( ~n14002 & n19326 ) | ( n19325 & n19326 ) ;
  assign n19328 = n19319 | n19327 ;
  assign n19329 = n141 | n19313 ;
  assign n19330 = ( n19313 & n19328 ) | ( n19313 & n19329 ) | ( n19328 & n19329 ) ;
  assign n19331 = ( x2 & n523 ) | ( x2 & n19313 ) | ( n523 & n19313 ) ;
  assign n19332 = x2 & n19310 ;
  assign n19333 = ( x2 & n19312 ) | ( x2 & n19332 ) | ( n19312 & n19332 ) ;
  assign n19334 = ( n19328 & n19331 ) | ( n19328 & n19333 ) | ( n19331 & n19333 ) ;
  assign n19335 = x2 & ~n19331 ;
  assign n19336 = x2 & ~n19333 ;
  assign n19337 = ( ~n19328 & n19335 ) | ( ~n19328 & n19336 ) | ( n19335 & n19336 ) ;
  assign n19338 = ( n19330 & ~n19334 ) | ( n19330 & n19337 ) | ( ~n19334 & n19337 ) ;
  assign n19339 = n19309 & n19338 ;
  assign n19340 = n19309 | n19338 ;
  assign n19341 = ~n19339 & n19340 ;
  assign n19342 = ( n18747 & n18748 ) | ( n18747 & n18783 ) | ( n18748 & n18783 ) ;
  assign n19343 = n19341 & n19342 ;
  assign n19344 = n19341 | n19342 ;
  assign n19345 = ~n19343 & n19344 ;
  assign n19346 = n18787 | n18789 ;
  assign n19347 = n18244 | n18787 ;
  assign n19348 = ( n18787 & n18789 ) | ( n18787 & n19347 ) | ( n18789 & n19347 ) ;
  assign n19349 = ( n18252 & n19346 ) | ( n18252 & n19348 ) | ( n19346 & n19348 ) ;
  assign n19350 = n19345 | n19349 ;
  assign n19351 = n19345 & n19349 ;
  assign n19352 = n19350 & ~n19351 ;
  assign n19353 = n19182 | n19188 ;
  assign n19354 = n18986 | n18992 ;
  assign n19355 = n18962 | n18966 ;
  assign n19356 = n18886 | n18891 ;
  assign n19357 = n18863 | n18866 ;
  assign n19358 = n293 & n17149 ;
  assign n19359 = x69 & n17146 ;
  assign n19360 = x68 & n17141 ;
  assign n19361 = x67 & ~n17140 ;
  assign n19362 = n17724 & n19361 ;
  assign n19363 = n19360 | n19362 ;
  assign n19364 = n19359 | n19363 ;
  assign n19365 = n19358 | n19364 ;
  assign n19366 = x62 | n19359 ;
  assign n19367 = n19363 | n19366 ;
  assign n19368 = n19358 | n19367 ;
  assign n19369 = ~x62 & n19367 ;
  assign n19370 = ( ~x62 & n19358 ) | ( ~x62 & n19369 ) | ( n19358 & n19369 ) ;
  assign n19371 = ( ~n19365 & n19368 ) | ( ~n19365 & n19370 ) | ( n19368 & n19370 ) ;
  assign n19372 = x66 & n18290 ;
  assign n19373 = x63 & x65 ;
  assign n19374 = ~n18290 & n19373 ;
  assign n19375 = n19372 | n19374 ;
  assign n19376 = n19367 & n19375 ;
  assign n19377 = ( n19358 & n19375 ) | ( n19358 & n19376 ) | ( n19375 & n19376 ) ;
  assign n19378 = ~n19364 & n19375 ;
  assign n19379 = ~n19358 & n19378 ;
  assign n19380 = ( n19370 & n19377 ) | ( n19370 & n19379 ) | ( n19377 & n19379 ) ;
  assign n19381 = n19371 & ~n19380 ;
  assign n19382 = ~n19367 & n19375 ;
  assign n19383 = ~n19358 & n19382 ;
  assign n19384 = n19364 & n19375 ;
  assign n19385 = ( n19358 & n19375 ) | ( n19358 & n19384 ) | ( n19375 & n19384 ) ;
  assign n19386 = ( ~n19370 & n19383 ) | ( ~n19370 & n19385 ) | ( n19383 & n19385 ) ;
  assign n19387 = n19381 | n19386 ;
  assign n19388 = n18834 | n18840 ;
  assign n19389 = n18835 | n19388 ;
  assign n19390 = n19387 | n19389 ;
  assign n19391 = n18834 | n19387 ;
  assign n19392 = ( n18842 & n19390 ) | ( n18842 & n19391 ) | ( n19390 & n19391 ) ;
  assign n19393 = n19387 & n19389 ;
  assign n19394 = n18834 & n19387 ;
  assign n19395 = ( n18842 & n19393 ) | ( n18842 & n19394 ) | ( n19393 & n19394 ) ;
  assign n19396 = n19392 & ~n19395 ;
  assign n19397 = x72 & n15552 ;
  assign n19398 = x71 & n15547 ;
  assign n19399 = x70 & ~n15546 ;
  assign n19400 = n16123 & n19399 ;
  assign n19401 = n19398 | n19400 ;
  assign n19402 = n19397 | n19401 ;
  assign n19403 = ( n513 & n15555 ) | ( n513 & n19402 ) | ( n15555 & n19402 ) ;
  assign n19404 = x59 & n15555 ;
  assign n19405 = ( x59 & n15555 ) | ( x59 & ~n19397 ) | ( n15555 & ~n19397 ) ;
  assign n19406 = ( ~n19401 & n19404 ) | ( ~n19401 & n19405 ) | ( n19404 & n19405 ) ;
  assign n19407 = ( x59 & n513 ) | ( x59 & n19406 ) | ( n513 & n19406 ) ;
  assign n19408 = ~n19403 & n19407 ;
  assign n19409 = n19402 | n19406 ;
  assign n19410 = x59 | n19402 ;
  assign n19411 = ( n513 & n19409 ) | ( n513 & n19410 ) | ( n19409 & n19410 ) ;
  assign n19412 = ( ~x59 & n19408 ) | ( ~x59 & n19411 ) | ( n19408 & n19411 ) ;
  assign n19413 = n19396 & n19412 ;
  assign n19414 = n19396 | n19412 ;
  assign n19415 = ~n19413 & n19414 ;
  assign n19416 = n18863 & n19414 ;
  assign n19417 = ~n19413 & n19416 ;
  assign n19418 = ( n18866 & n19415 ) | ( n18866 & n19417 ) | ( n19415 & n19417 ) ;
  assign n19419 = n19357 & ~n19418 ;
  assign n19420 = x75 & n14045 ;
  assign n19421 = x74 & n14040 ;
  assign n19422 = x73 & ~n14039 ;
  assign n19423 = n14552 & n19422 ;
  assign n19424 = n19421 | n19423 ;
  assign n19425 = n19420 | n19424 ;
  assign n19426 = n14048 | n19420 ;
  assign n19427 = n19424 | n19426 ;
  assign n19428 = ( n746 & n19425 ) | ( n746 & n19427 ) | ( n19425 & n19427 ) ;
  assign n19429 = x56 & n19427 ;
  assign n19430 = x56 & n19420 ;
  assign n19431 = ( x56 & n19424 ) | ( x56 & n19430 ) | ( n19424 & n19430 ) ;
  assign n19432 = ( n746 & n19429 ) | ( n746 & n19431 ) | ( n19429 & n19431 ) ;
  assign n19433 = x56 & ~n19431 ;
  assign n19434 = x56 & ~n19427 ;
  assign n19435 = ( ~n746 & n19433 ) | ( ~n746 & n19434 ) | ( n19433 & n19434 ) ;
  assign n19436 = ( n19428 & ~n19432 ) | ( n19428 & n19435 ) | ( ~n19432 & n19435 ) ;
  assign n19437 = ( n18866 & n19414 ) | ( n18866 & n19416 ) | ( n19414 & n19416 ) ;
  assign n19438 = n19415 & n19436 ;
  assign n19439 = ~n19437 & n19438 ;
  assign n19440 = ( n19419 & n19436 ) | ( n19419 & n19439 ) | ( n19436 & n19439 ) ;
  assign n19441 = n19415 | n19436 ;
  assign n19442 = ( n19436 & ~n19437 ) | ( n19436 & n19441 ) | ( ~n19437 & n19441 ) ;
  assign n19443 = n19419 | n19442 ;
  assign n19444 = ~n19440 & n19443 ;
  assign n19445 = n19356 & n19444 ;
  assign n19446 = n19356 | n19444 ;
  assign n19447 = ~n19445 & n19446 ;
  assign n19448 = x78 & n12574 ;
  assign n19449 = x77 & n12569 ;
  assign n19450 = x76 & ~n12568 ;
  assign n19451 = n13076 & n19450 ;
  assign n19452 = n19449 | n19451 ;
  assign n19453 = n19448 | n19452 ;
  assign n19454 = n12577 | n19448 ;
  assign n19455 = n19452 | n19454 ;
  assign n19456 = ( n1192 & n19453 ) | ( n1192 & n19455 ) | ( n19453 & n19455 ) ;
  assign n19457 = x53 & n19455 ;
  assign n19458 = x53 & n19448 ;
  assign n19459 = ( x53 & n19452 ) | ( x53 & n19458 ) | ( n19452 & n19458 ) ;
  assign n19460 = ( n1192 & n19457 ) | ( n1192 & n19459 ) | ( n19457 & n19459 ) ;
  assign n19461 = x53 & ~n19459 ;
  assign n19462 = x53 & ~n19455 ;
  assign n19463 = ( ~n1192 & n19461 ) | ( ~n1192 & n19462 ) | ( n19461 & n19462 ) ;
  assign n19464 = ( n19456 & ~n19460 ) | ( n19456 & n19463 ) | ( ~n19460 & n19463 ) ;
  assign n19465 = n19447 & n19464 ;
  assign n19466 = n19447 & ~n19465 ;
  assign n19467 = ~n19447 & n19464 ;
  assign n19468 = n19466 | n19467 ;
  assign n19469 = n18913 | n18914 ;
  assign n19470 = ( n18913 & n18915 ) | ( n18913 & n19469 ) | ( n18915 & n19469 ) ;
  assign n19471 = ~n19468 & n19470 ;
  assign n19472 = n19468 & ~n19470 ;
  assign n19473 = n19471 | n19472 ;
  assign n19474 = x81 & n11205 ;
  assign n19475 = x80 & n11200 ;
  assign n19476 = x79 & ~n11199 ;
  assign n19477 = n11679 & n19476 ;
  assign n19478 = n19475 | n19477 ;
  assign n19479 = n19474 | n19478 ;
  assign n19480 = n11208 | n19474 ;
  assign n19481 = n19478 | n19480 ;
  assign n19482 = ( n1651 & n19479 ) | ( n1651 & n19481 ) | ( n19479 & n19481 ) ;
  assign n19483 = x50 & n19481 ;
  assign n19484 = x50 & n19474 ;
  assign n19485 = ( x50 & n19478 ) | ( x50 & n19484 ) | ( n19478 & n19484 ) ;
  assign n19486 = ( n1651 & n19483 ) | ( n1651 & n19485 ) | ( n19483 & n19485 ) ;
  assign n19487 = x50 & ~n19485 ;
  assign n19488 = x50 & ~n19481 ;
  assign n19489 = ( ~n1651 & n19487 ) | ( ~n1651 & n19488 ) | ( n19487 & n19488 ) ;
  assign n19490 = ( n19482 & ~n19486 ) | ( n19482 & n19489 ) | ( ~n19486 & n19489 ) ;
  assign n19491 = n19473 & n19490 ;
  assign n19492 = n19473 | n19490 ;
  assign n19493 = ~n19491 & n19492 ;
  assign n19494 = n18936 | n18942 ;
  assign n19495 = n19493 | n19494 ;
  assign n19496 = n19493 & n19494 ;
  assign n19497 = n19495 & ~n19496 ;
  assign n19498 = x84 & n9933 ;
  assign n19499 = x83 & n9928 ;
  assign n19500 = x82 & ~n9927 ;
  assign n19501 = n10379 & n19500 ;
  assign n19502 = n19499 | n19501 ;
  assign n19503 = n19498 | n19502 ;
  assign n19504 = n9936 | n19498 ;
  assign n19505 = n19502 | n19504 ;
  assign n19506 = ( n2194 & n19503 ) | ( n2194 & n19505 ) | ( n19503 & n19505 ) ;
  assign n19507 = x47 & n19505 ;
  assign n19508 = x47 & n19498 ;
  assign n19509 = ( x47 & n19502 ) | ( x47 & n19508 ) | ( n19502 & n19508 ) ;
  assign n19510 = ( n2194 & n19507 ) | ( n2194 & n19509 ) | ( n19507 & n19509 ) ;
  assign n19511 = x47 & ~n19509 ;
  assign n19512 = x47 & ~n19505 ;
  assign n19513 = ( ~n2194 & n19511 ) | ( ~n2194 & n19512 ) | ( n19511 & n19512 ) ;
  assign n19514 = ( n19506 & ~n19510 ) | ( n19506 & n19513 ) | ( ~n19510 & n19513 ) ;
  assign n19515 = n19497 & n19514 ;
  assign n19516 = n19497 & ~n19515 ;
  assign n19517 = ~n19497 & n19514 ;
  assign n19518 = n19516 | n19517 ;
  assign n19519 = n19355 & ~n19518 ;
  assign n19520 = ~n19355 & n19518 ;
  assign n19521 = n19519 | n19520 ;
  assign n19522 = x87 & n8724 ;
  assign n19523 = x86 & n8719 ;
  assign n19524 = x85 & ~n8718 ;
  assign n19525 = n9149 & n19524 ;
  assign n19526 = n19523 | n19525 ;
  assign n19527 = n19522 | n19526 ;
  assign n19528 = n8727 | n19522 ;
  assign n19529 = n19526 | n19528 ;
  assign n19530 = ( n2816 & n19527 ) | ( n2816 & n19529 ) | ( n19527 & n19529 ) ;
  assign n19531 = x44 & n19529 ;
  assign n19532 = x44 & n19522 ;
  assign n19533 = ( x44 & n19526 ) | ( x44 & n19532 ) | ( n19526 & n19532 ) ;
  assign n19534 = ( n2816 & n19531 ) | ( n2816 & n19533 ) | ( n19531 & n19533 ) ;
  assign n19535 = x44 & ~n19533 ;
  assign n19536 = x44 & ~n19529 ;
  assign n19537 = ( ~n2816 & n19535 ) | ( ~n2816 & n19536 ) | ( n19535 & n19536 ) ;
  assign n19538 = ( n19530 & ~n19534 ) | ( n19530 & n19537 ) | ( ~n19534 & n19537 ) ;
  assign n19539 = n19521 & n19538 ;
  assign n19540 = n19521 | n19538 ;
  assign n19541 = ~n19539 & n19540 ;
  assign n19542 = n19354 | n19541 ;
  assign n19543 = n19354 & n19541 ;
  assign n19544 = n19542 & ~n19543 ;
  assign n19545 = x90 & n7566 ;
  assign n19546 = x89 & n7561 ;
  assign n19547 = x88 & ~n7560 ;
  assign n19548 = n7953 & n19547 ;
  assign n19549 = n19546 | n19548 ;
  assign n19550 = n19545 | n19549 ;
  assign n19551 = n7569 | n19545 ;
  assign n19552 = n19549 | n19551 ;
  assign n19553 = ( n3519 & n19550 ) | ( n3519 & n19552 ) | ( n19550 & n19552 ) ;
  assign n19554 = x41 & n19552 ;
  assign n19555 = x41 & n19545 ;
  assign n19556 = ( x41 & n19549 ) | ( x41 & n19555 ) | ( n19549 & n19555 ) ;
  assign n19557 = ( n3519 & n19554 ) | ( n3519 & n19556 ) | ( n19554 & n19556 ) ;
  assign n19558 = x41 & ~n19556 ;
  assign n19559 = x41 & ~n19552 ;
  assign n19560 = ( ~n3519 & n19558 ) | ( ~n3519 & n19559 ) | ( n19558 & n19559 ) ;
  assign n19561 = ( n19553 & ~n19557 ) | ( n19553 & n19560 ) | ( ~n19557 & n19560 ) ;
  assign n19562 = n19544 & n19561 ;
  assign n19563 = n19544 & ~n19562 ;
  assign n19564 = ~n19544 & n19561 ;
  assign n19565 = n19563 | n19564 ;
  assign n19566 = n19011 | n19019 ;
  assign n19567 = n19565 | n19566 ;
  assign n19568 = n19565 & n19566 ;
  assign n19569 = n19567 & ~n19568 ;
  assign n19570 = x93 & n6536 ;
  assign n19571 = x92 & n6531 ;
  assign n19572 = x91 & ~n6530 ;
  assign n19573 = n6871 & n19572 ;
  assign n19574 = n19571 | n19573 ;
  assign n19575 = n19570 | n19574 ;
  assign n19576 = n6539 | n19570 ;
  assign n19577 = n19574 | n19576 ;
  assign n19578 = ( n4305 & n19575 ) | ( n4305 & n19577 ) | ( n19575 & n19577 ) ;
  assign n19579 = x38 & n19577 ;
  assign n19580 = x38 & n19570 ;
  assign n19581 = ( x38 & n19574 ) | ( x38 & n19580 ) | ( n19574 & n19580 ) ;
  assign n19582 = ( n4305 & n19579 ) | ( n4305 & n19581 ) | ( n19579 & n19581 ) ;
  assign n19583 = x38 & ~n19581 ;
  assign n19584 = x38 & ~n19577 ;
  assign n19585 = ( ~n4305 & n19583 ) | ( ~n4305 & n19584 ) | ( n19583 & n19584 ) ;
  assign n19586 = ( n19578 & ~n19582 ) | ( n19578 & n19585 ) | ( ~n19582 & n19585 ) ;
  assign n19587 = n19569 & n19586 ;
  assign n19588 = n19569 & ~n19587 ;
  assign n19589 = ~n19569 & n19586 ;
  assign n19590 = n19588 | n19589 ;
  assign n19591 = n19038 | n19040 ;
  assign n19592 = n19039 | n19591 ;
  assign n19593 = ( n19038 & n19042 ) | ( n19038 & n19592 ) | ( n19042 & n19592 ) ;
  assign n19594 = n19590 | n19593 ;
  assign n19595 = n19590 & n19593 ;
  assign n19596 = n19594 & ~n19595 ;
  assign n19597 = x96 & n5554 ;
  assign n19598 = x95 & n5549 ;
  assign n19599 = x94 & ~n5548 ;
  assign n19600 = n5893 & n19599 ;
  assign n19601 = n19598 | n19600 ;
  assign n19602 = n19597 | n19601 ;
  assign n19603 = n5557 | n19597 ;
  assign n19604 = n19601 | n19603 ;
  assign n19605 = ( n5202 & n19602 ) | ( n5202 & n19604 ) | ( n19602 & n19604 ) ;
  assign n19606 = x35 & n19604 ;
  assign n19607 = x35 & n19597 ;
  assign n19608 = ( x35 & n19601 ) | ( x35 & n19607 ) | ( n19601 & n19607 ) ;
  assign n19609 = ( n5202 & n19606 ) | ( n5202 & n19608 ) | ( n19606 & n19608 ) ;
  assign n19610 = x35 & ~n19608 ;
  assign n19611 = x35 & ~n19604 ;
  assign n19612 = ( ~n5202 & n19610 ) | ( ~n5202 & n19611 ) | ( n19610 & n19611 ) ;
  assign n19613 = ( n19605 & ~n19609 ) | ( n19605 & n19612 ) | ( ~n19609 & n19612 ) ;
  assign n19614 = n19596 & n19613 ;
  assign n19615 = n19596 | n19613 ;
  assign n19616 = ~n19614 & n19615 ;
  assign n19617 = n19064 | n19065 ;
  assign n19618 = ( n19064 & n19068 ) | ( n19064 & n19617 ) | ( n19068 & n19617 ) ;
  assign n19619 = n19616 & n19618 ;
  assign n19620 = n19618 & ~n19619 ;
  assign n19621 = ( n19616 & ~n19619 ) | ( n19616 & n19620 ) | ( ~n19619 & n19620 ) ;
  assign n19622 = x99 & n4631 ;
  assign n19623 = x98 & n4626 ;
  assign n19624 = x97 & ~n4625 ;
  assign n19625 = n4943 & n19624 ;
  assign n19626 = n19623 | n19625 ;
  assign n19627 = n19622 | n19626 ;
  assign n19628 = n4634 | n19622 ;
  assign n19629 = n19626 | n19628 ;
  assign n19630 = ( n6164 & n19627 ) | ( n6164 & n19629 ) | ( n19627 & n19629 ) ;
  assign n19631 = x32 & n19629 ;
  assign n19632 = x32 & n19622 ;
  assign n19633 = ( x32 & n19626 ) | ( x32 & n19632 ) | ( n19626 & n19632 ) ;
  assign n19634 = ( n6164 & n19631 ) | ( n6164 & n19633 ) | ( n19631 & n19633 ) ;
  assign n19635 = x32 & ~n19633 ;
  assign n19636 = x32 & ~n19629 ;
  assign n19637 = ( ~n6164 & n19635 ) | ( ~n6164 & n19636 ) | ( n19635 & n19636 ) ;
  assign n19638 = ( n19630 & ~n19634 ) | ( n19630 & n19637 ) | ( ~n19634 & n19637 ) ;
  assign n19639 = n19616 & n19638 ;
  assign n19640 = ~n19616 & n19638 ;
  assign n19641 = ( ~n19618 & n19638 ) | ( ~n19618 & n19640 ) | ( n19638 & n19640 ) ;
  assign n19642 = ( n19620 & n19639 ) | ( n19620 & n19641 ) | ( n19639 & n19641 ) ;
  assign n19643 = n19621 & ~n19642 ;
  assign n19644 = n19618 & n19639 ;
  assign n19645 = ( ~n19620 & n19640 ) | ( ~n19620 & n19644 ) | ( n19640 & n19644 ) ;
  assign n19646 = n19643 | n19645 ;
  assign n19647 = n19095 | n19100 ;
  assign n19648 = n19646 | n19647 ;
  assign n19649 = n19646 & n19647 ;
  assign n19650 = n19648 & ~n19649 ;
  assign n19651 = x102 & n3816 ;
  assign n19652 = x101 & n3811 ;
  assign n19653 = x100 & ~n3810 ;
  assign n19654 = n4067 & n19653 ;
  assign n19655 = n19652 | n19654 ;
  assign n19656 = n19651 | n19655 ;
  assign n19657 = n3819 | n19651 ;
  assign n19658 = n19655 | n19657 ;
  assign n19659 = ( n7178 & n19656 ) | ( n7178 & n19658 ) | ( n19656 & n19658 ) ;
  assign n19660 = x29 & n19658 ;
  assign n19661 = x29 & n19651 ;
  assign n19662 = ( x29 & n19655 ) | ( x29 & n19661 ) | ( n19655 & n19661 ) ;
  assign n19663 = ( n7178 & n19660 ) | ( n7178 & n19662 ) | ( n19660 & n19662 ) ;
  assign n19664 = x29 & ~n19662 ;
  assign n19665 = x29 & ~n19658 ;
  assign n19666 = ( ~n7178 & n19664 ) | ( ~n7178 & n19665 ) | ( n19664 & n19665 ) ;
  assign n19667 = ( n19659 & ~n19663 ) | ( n19659 & n19666 ) | ( ~n19663 & n19666 ) ;
  assign n19668 = n19650 & n19667 ;
  assign n19669 = n19650 & ~n19668 ;
  assign n19670 = ~n19650 & n19667 ;
  assign n19671 = n19669 | n19670 ;
  assign n19672 = n19121 | n19128 ;
  assign n19673 = n19671 | n19672 ;
  assign n19674 = n19671 & n19672 ;
  assign n19675 = n19673 & ~n19674 ;
  assign n19676 = x105 & n3085 ;
  assign n19677 = x104 & n3080 ;
  assign n19678 = x103 & ~n3079 ;
  assign n19679 = n3309 & n19678 ;
  assign n19680 = n19677 | n19679 ;
  assign n19681 = n19676 | n19680 ;
  assign n19682 = n3088 | n19676 ;
  assign n19683 = n19680 | n19682 ;
  assign n19684 = ( n8273 & n19681 ) | ( n8273 & n19683 ) | ( n19681 & n19683 ) ;
  assign n19685 = x26 & n19683 ;
  assign n19686 = x26 & n19676 ;
  assign n19687 = ( x26 & n19680 ) | ( x26 & n19686 ) | ( n19680 & n19686 ) ;
  assign n19688 = ( n8273 & n19685 ) | ( n8273 & n19687 ) | ( n19685 & n19687 ) ;
  assign n19689 = x26 & ~n19687 ;
  assign n19690 = x26 & ~n19683 ;
  assign n19691 = ( ~n8273 & n19689 ) | ( ~n8273 & n19690 ) | ( n19689 & n19690 ) ;
  assign n19692 = ( n19684 & ~n19688 ) | ( n19684 & n19691 ) | ( ~n19688 & n19691 ) ;
  assign n19693 = n19675 & n19692 ;
  assign n19694 = n19675 | n19692 ;
  assign n19695 = ~n19693 & n19694 ;
  assign n19696 = n19147 | n19150 ;
  assign n19697 = ( n19147 & n19151 ) | ( n19147 & n19696 ) | ( n19151 & n19696 ) ;
  assign n19698 = n19695 & n19697 ;
  assign n19699 = n19697 & ~n19698 ;
  assign n19700 = ( n19695 & ~n19698 ) | ( n19695 & n19699 ) | ( ~n19698 & n19699 ) ;
  assign n19701 = x108 & n2429 ;
  assign n19702 = x107 & n2424 ;
  assign n19703 = x106 & ~n2423 ;
  assign n19704 = n2631 & n19703 ;
  assign n19705 = n19702 | n19704 ;
  assign n19706 = n19701 | n19705 ;
  assign n19707 = n2432 | n19701 ;
  assign n19708 = n19705 | n19707 ;
  assign n19709 = ( n9479 & n19706 ) | ( n9479 & n19708 ) | ( n19706 & n19708 ) ;
  assign n19710 = x23 & n19708 ;
  assign n19711 = x23 & n19701 ;
  assign n19712 = ( x23 & n19705 ) | ( x23 & n19711 ) | ( n19705 & n19711 ) ;
  assign n19713 = ( n9479 & n19710 ) | ( n9479 & n19712 ) | ( n19710 & n19712 ) ;
  assign n19714 = x23 & ~n19712 ;
  assign n19715 = x23 & ~n19708 ;
  assign n19716 = ( ~n9479 & n19714 ) | ( ~n9479 & n19715 ) | ( n19714 & n19715 ) ;
  assign n19717 = ( n19709 & ~n19713 ) | ( n19709 & n19716 ) | ( ~n19713 & n19716 ) ;
  assign n19718 = ~n19698 & n19717 ;
  assign n19719 = n19695 & n19717 ;
  assign n19720 = ( n19699 & n19718 ) | ( n19699 & n19719 ) | ( n19718 & n19719 ) ;
  assign n19721 = n19700 & ~n19720 ;
  assign n19722 = ~n19150 & n19151 ;
  assign n19723 = n19152 | n19722 ;
  assign n19724 = ( n18619 & n18811 ) | ( n18619 & n19723 ) | ( n18811 & n19723 ) ;
  assign n19725 = n18811 | n19723 ;
  assign n19726 = ( n18626 & n19724 ) | ( n18626 & n19725 ) | ( n19724 & n19725 ) ;
  assign n19727 = n19698 & n19717 ;
  assign n19728 = ~n19695 & n19717 ;
  assign n19729 = ( ~n19699 & n19727 ) | ( ~n19699 & n19728 ) | ( n19727 & n19728 ) ;
  assign n19730 = n19726 & n19729 ;
  assign n19731 = ( n19721 & n19726 ) | ( n19721 & n19730 ) | ( n19726 & n19730 ) ;
  assign n19732 = n19726 | n19729 ;
  assign n19733 = n19721 | n19732 ;
  assign n19734 = ~n19731 & n19733 ;
  assign n19735 = x111 & n1859 ;
  assign n19736 = x110 & n1854 ;
  assign n19737 = x109 & ~n1853 ;
  assign n19738 = n2037 & n19737 ;
  assign n19739 = n19736 | n19738 ;
  assign n19740 = n19735 | n19739 ;
  assign n19741 = n1862 | n19735 ;
  assign n19742 = n19739 | n19741 ;
  assign n19743 = ( n10749 & n19740 ) | ( n10749 & n19742 ) | ( n19740 & n19742 ) ;
  assign n19744 = x20 & n19742 ;
  assign n19745 = x20 & n19735 ;
  assign n19746 = ( x20 & n19739 ) | ( x20 & n19745 ) | ( n19739 & n19745 ) ;
  assign n19747 = ( n10749 & n19744 ) | ( n10749 & n19746 ) | ( n19744 & n19746 ) ;
  assign n19748 = x20 & ~n19746 ;
  assign n19749 = x20 & ~n19742 ;
  assign n19750 = ( ~n10749 & n19748 ) | ( ~n10749 & n19749 ) | ( n19748 & n19749 ) ;
  assign n19751 = ( n19743 & ~n19747 ) | ( n19743 & n19750 ) | ( ~n19747 & n19750 ) ;
  assign n19752 = n19734 & n19751 ;
  assign n19753 = n19734 & ~n19752 ;
  assign n19754 = ~n19734 & n19751 ;
  assign n19755 = n19753 | n19754 ;
  assign n19756 = n19353 & n19755 ;
  assign n19757 = n19353 & ~n19756 ;
  assign n19758 = x114 & n1383 ;
  assign n19759 = x113 & n1378 ;
  assign n19760 = x112 & ~n1377 ;
  assign n19761 = n1542 & n19760 ;
  assign n19762 = n19759 | n19761 ;
  assign n19763 = n19758 | n19762 ;
  assign n19764 = n1386 | n19758 ;
  assign n19765 = n19762 | n19764 ;
  assign n19766 = ( ~n12095 & n19763 ) | ( ~n12095 & n19765 ) | ( n19763 & n19765 ) ;
  assign n19767 = n19763 & n19765 ;
  assign n19768 = ( n12079 & n19766 ) | ( n12079 & n19767 ) | ( n19766 & n19767 ) ;
  assign n19769 = x17 & n19768 ;
  assign n19770 = x17 & ~n19768 ;
  assign n19771 = ( n19768 & ~n19769 ) | ( n19768 & n19770 ) | ( ~n19769 & n19770 ) ;
  assign n19772 = ~n19353 & n19755 ;
  assign n19773 = n19771 | n19772 ;
  assign n19774 = n19757 | n19773 ;
  assign n19775 = n19771 & n19772 ;
  assign n19776 = ( n19757 & n19771 ) | ( n19757 & n19775 ) | ( n19771 & n19775 ) ;
  assign n19777 = n19774 & ~n19776 ;
  assign n19778 = n19205 | n19210 ;
  assign n19779 = ( n19205 & n19208 ) | ( n19205 & n19778 ) | ( n19208 & n19778 ) ;
  assign n19780 = n19777 & n19779 ;
  assign n19781 = n19777 | n19779 ;
  assign n19782 = ~n19780 & n19781 ;
  assign n19783 = x117 & n962 ;
  assign n19784 = x116 & n957 ;
  assign n19785 = x115 & ~n956 ;
  assign n19786 = n1105 & n19785 ;
  assign n19787 = n19784 | n19786 ;
  assign n19788 = n19783 | n19787 ;
  assign n19789 = n965 | n19783 ;
  assign n19790 = n19787 | n19789 ;
  assign n19791 = ( ~n13522 & n19788 ) | ( ~n13522 & n19790 ) | ( n19788 & n19790 ) ;
  assign n19792 = n19788 & n19790 ;
  assign n19793 = ( n13503 & n19791 ) | ( n13503 & n19792 ) | ( n19791 & n19792 ) ;
  assign n19794 = x14 & n19793 ;
  assign n19795 = x14 & ~n19793 ;
  assign n19796 = ( n19793 & ~n19794 ) | ( n19793 & n19795 ) | ( ~n19794 & n19795 ) ;
  assign n19797 = n19782 & n19796 ;
  assign n19798 = n19782 & ~n19797 ;
  assign n19799 = ~n19782 & n19796 ;
  assign n19800 = n19798 | n19799 ;
  assign n19801 = n19228 | n19230 ;
  assign n19802 = ( n19228 & n19231 ) | ( n19228 & n19801 ) | ( n19231 & n19801 ) ;
  assign n19803 = n19800 | n19802 ;
  assign n19804 = n19800 & n19802 ;
  assign n19805 = n19803 & ~n19804 ;
  assign n19806 = x120 & n636 ;
  assign n19807 = x119 & n631 ;
  assign n19808 = x118 & ~n630 ;
  assign n19809 = n764 & n19808 ;
  assign n19810 = n19807 | n19809 ;
  assign n19811 = n19806 | n19810 ;
  assign n19812 = n639 | n19806 ;
  assign n19813 = n19810 | n19812 ;
  assign n19814 = ( n14991 & n19811 ) | ( n14991 & n19813 ) | ( n19811 & n19813 ) ;
  assign n19815 = x11 & n19813 ;
  assign n19816 = x11 & n19806 ;
  assign n19817 = ( x11 & n19810 ) | ( x11 & n19816 ) | ( n19810 & n19816 ) ;
  assign n19818 = ( n14991 & n19815 ) | ( n14991 & n19817 ) | ( n19815 & n19817 ) ;
  assign n19819 = x11 & ~n19817 ;
  assign n19820 = x11 & ~n19813 ;
  assign n19821 = ( ~n14991 & n19819 ) | ( ~n14991 & n19820 ) | ( n19819 & n19820 ) ;
  assign n19822 = ( n19814 & ~n19818 ) | ( n19814 & n19821 ) | ( ~n19818 & n19821 ) ;
  assign n19823 = n19805 | n19822 ;
  assign n19824 = n19805 & n19822 ;
  assign n19825 = n19823 & ~n19824 ;
  assign n19826 = x123 & n389 ;
  assign n19827 = x122 & n384 ;
  assign n19828 = x121 & ~n383 ;
  assign n19829 = n463 & n19828 ;
  assign n19830 = n19827 | n19829 ;
  assign n19831 = n19826 | n19830 ;
  assign n19832 = n392 | n19826 ;
  assign n19833 = n19830 | n19832 ;
  assign n19834 = ( n16086 & n19831 ) | ( n16086 & n19833 ) | ( n19831 & n19833 ) ;
  assign n19835 = x8 & n19833 ;
  assign n19836 = x8 & n19826 ;
  assign n19837 = ( x8 & n19830 ) | ( x8 & n19836 ) | ( n19830 & n19836 ) ;
  assign n19838 = ( n16086 & n19835 ) | ( n16086 & n19837 ) | ( n19835 & n19837 ) ;
  assign n19839 = x8 & ~n19837 ;
  assign n19840 = x8 & ~n19833 ;
  assign n19841 = ( ~n16086 & n19839 ) | ( ~n16086 & n19840 ) | ( n19839 & n19840 ) ;
  assign n19842 = ( n19834 & ~n19838 ) | ( n19834 & n19841 ) | ( ~n19838 & n19841 ) ;
  assign n19843 = ~n19825 & n19842 ;
  assign n19844 = n19252 | n19254 ;
  assign n19845 = ( n19252 & n19255 ) | ( n19252 & n19844 ) | ( n19255 & n19844 ) ;
  assign n19846 = n19822 | n19842 ;
  assign n19847 = ( n19805 & n19842 ) | ( n19805 & n19846 ) | ( n19842 & n19846 ) ;
  assign n19848 = n19823 & ~n19847 ;
  assign n19849 = n19845 & n19848 ;
  assign n19850 = ( n19843 & n19845 ) | ( n19843 & n19849 ) | ( n19845 & n19849 ) ;
  assign n19851 = n19845 | n19848 ;
  assign n19852 = n19843 | n19851 ;
  assign n19853 = ~n19850 & n19852 ;
  assign n19854 = x126 & n212 ;
  assign n19855 = x125 & n207 ;
  assign n19856 = x124 & ~n206 ;
  assign n19857 = n267 & n19856 ;
  assign n19858 = n19855 | n19857 ;
  assign n19859 = n19854 | n19858 ;
  assign n19860 = n215 | n19854 ;
  assign n19861 = n19858 | n19860 ;
  assign n19862 = ( n18220 & n19859 ) | ( n18220 & n19861 ) | ( n19859 & n19861 ) ;
  assign n19863 = x5 & n19861 ;
  assign n19864 = x5 & n19854 ;
  assign n19865 = ( x5 & n19858 ) | ( x5 & n19864 ) | ( n19858 & n19864 ) ;
  assign n19866 = ( n18220 & n19863 ) | ( n18220 & n19865 ) | ( n19863 & n19865 ) ;
  assign n19867 = x5 & ~n19865 ;
  assign n19868 = x5 & ~n19861 ;
  assign n19869 = ( ~n18220 & n19867 ) | ( ~n18220 & n19868 ) | ( n19867 & n19868 ) ;
  assign n19870 = ( n19862 & ~n19866 ) | ( n19862 & n19869 ) | ( ~n19866 & n19869 ) ;
  assign n19871 = n19853 & n19870 ;
  assign n19872 = n19853 & ~n19871 ;
  assign n19873 = ~n19853 & n19870 ;
  assign n19874 = n19872 | n19873 ;
  assign n19875 = n19258 & n19275 ;
  assign n19876 = n19258 & ~n19875 ;
  assign n19877 = x127 & n19321 ;
  assign n19878 = n141 & n19877 ;
  assign n19879 = x126 & x127 ;
  assign n19880 = ( x127 & n18751 ) | ( x127 & n19879 ) | ( n18751 & n19879 ) ;
  assign n19881 = n141 & n19880 ;
  assign n19882 = n19878 & n19881 ;
  assign n19883 = x2 | n19882 ;
  assign n19884 = ( n18202 & n19878 ) | ( n18202 & n19881 ) | ( n19878 & n19881 ) ;
  assign n19885 = x2 | n19884 ;
  assign n19886 = ( n18212 & n19883 ) | ( n18212 & n19885 ) | ( n19883 & n19885 ) ;
  assign n19887 = ( n18214 & n19883 ) | ( n18214 & n19885 ) | ( n19883 & n19885 ) ;
  assign n19888 = ( n14002 & n19886 ) | ( n14002 & n19887 ) | ( n19886 & n19887 ) ;
  assign n19889 = x127 & ~n162 ;
  assign n19890 = n137 & n19889 ;
  assign n19891 = n19881 | n19890 ;
  assign n19892 = n141 | n19890 ;
  assign n19893 = ( n19877 & n19890 ) | ( n19877 & n19892 ) | ( n19890 & n19892 ) ;
  assign n19894 = n19891 & n19893 ;
  assign n19895 = x2 & n19894 ;
  assign n19896 = ( n18202 & n19891 ) | ( n18202 & n19893 ) | ( n19891 & n19893 ) ;
  assign n19897 = x2 & n19896 ;
  assign n19898 = ( n18212 & n19895 ) | ( n18212 & n19897 ) | ( n19895 & n19897 ) ;
  assign n19899 = ( n18214 & n19895 ) | ( n18214 & n19897 ) | ( n19895 & n19897 ) ;
  assign n19900 = ( n14002 & n19898 ) | ( n14002 & n19899 ) | ( n19898 & n19899 ) ;
  assign n19901 = n19888 & ~n19900 ;
  assign n19902 = n19275 & n19292 ;
  assign n19903 = ~n19258 & n19902 ;
  assign n19904 = n19275 & n19901 ;
  assign n19905 = n19258 & n19904 ;
  assign n19906 = ( n19901 & n19903 ) | ( n19901 & n19905 ) | ( n19903 & n19905 ) ;
  assign n19907 = ( n19292 & n19901 ) | ( n19292 & n19904 ) | ( n19901 & n19904 ) ;
  assign n19908 = n19292 & n19901 ;
  assign n19909 = ( n19258 & n19907 ) | ( n19258 & n19908 ) | ( n19907 & n19908 ) ;
  assign n19910 = ( n19876 & n19906 ) | ( n19876 & n19909 ) | ( n19906 & n19909 ) ;
  assign n19911 = n19275 | n19901 ;
  assign n19912 = ( n19258 & n19901 ) | ( n19258 & n19911 ) | ( n19901 & n19911 ) ;
  assign n19913 = n19903 | n19912 ;
  assign n19914 = n19292 | n19911 ;
  assign n19915 = n19292 | n19901 ;
  assign n19916 = ( n19258 & n19914 ) | ( n19258 & n19915 ) | ( n19914 & n19915 ) ;
  assign n19917 = ( n19876 & n19913 ) | ( n19876 & n19916 ) | ( n19913 & n19916 ) ;
  assign n19918 = ~n19910 & n19917 ;
  assign n19919 = n19874 & n19918 ;
  assign n19920 = n19874 | n19918 ;
  assign n19921 = ~n19919 & n19920 ;
  assign n19922 = n19305 | n19338 ;
  assign n19923 = ( n19305 & n19309 ) | ( n19305 & n19922 ) | ( n19309 & n19922 ) ;
  assign n19924 = n19921 | n19923 ;
  assign n19925 = n19921 & n19923 ;
  assign n19926 = n19924 & ~n19925 ;
  assign n19927 = n19343 | n19345 ;
  assign n19928 = ( n19343 & n19349 ) | ( n19343 & n19927 ) | ( n19349 & n19927 ) ;
  assign n19929 = n19926 | n19928 ;
  assign n19930 = n19926 & n19927 ;
  assign n19931 = n19343 & n19926 ;
  assign n19932 = ( n19349 & n19930 ) | ( n19349 & n19931 ) | ( n19930 & n19931 ) ;
  assign n19933 = n19929 & ~n19932 ;
  assign n19951 = n19850 | n19870 ;
  assign n19952 = ( n19850 & n19853 ) | ( n19850 & n19951 ) | ( n19853 & n19951 ) ;
  assign n19934 = x127 & n212 ;
  assign n19935 = x126 & n207 ;
  assign n19936 = x125 & ~n206 ;
  assign n19937 = n267 & n19936 ;
  assign n19938 = n19935 | n19937 ;
  assign n19939 = n19934 | n19938 ;
  assign n19940 = n215 | n19934 ;
  assign n19941 = n19938 | n19940 ;
  assign n19942 = ( n18763 & n19939 ) | ( n18763 & n19941 ) | ( n19939 & n19941 ) ;
  assign n19943 = x5 & n19941 ;
  assign n19944 = x5 & n19934 ;
  assign n19945 = ( x5 & n19938 ) | ( x5 & n19944 ) | ( n19938 & n19944 ) ;
  assign n19946 = ( n18763 & n19943 ) | ( n18763 & n19945 ) | ( n19943 & n19945 ) ;
  assign n19947 = x5 & ~n19945 ;
  assign n19948 = x5 & ~n19941 ;
  assign n19949 = ( ~n18763 & n19947 ) | ( ~n18763 & n19948 ) | ( n19947 & n19948 ) ;
  assign n19950 = ( n19942 & ~n19946 ) | ( n19942 & n19949 ) | ( ~n19946 & n19949 ) ;
  assign n19953 = n19950 & n19952 ;
  assign n19954 = n19952 & ~n19953 ;
  assign n19955 = x121 & n636 ;
  assign n19956 = x120 & n631 ;
  assign n19957 = x119 & ~n630 ;
  assign n19958 = n764 & n19957 ;
  assign n19959 = n19956 | n19958 ;
  assign n19960 = n19955 | n19959 ;
  assign n19961 = n639 | n19955 ;
  assign n19962 = n19959 | n19961 ;
  assign n19963 = ( n15501 & n19960 ) | ( n15501 & n19962 ) | ( n19960 & n19962 ) ;
  assign n19964 = x11 & n19962 ;
  assign n19965 = x11 & n19955 ;
  assign n19966 = ( x11 & n19959 ) | ( x11 & n19965 ) | ( n19959 & n19965 ) ;
  assign n19967 = ( n15501 & n19964 ) | ( n15501 & n19966 ) | ( n19964 & n19966 ) ;
  assign n19968 = x11 & ~n19966 ;
  assign n19969 = x11 & ~n19962 ;
  assign n19970 = ( ~n15501 & n19968 ) | ( ~n15501 & n19969 ) | ( n19968 & n19969 ) ;
  assign n19971 = ( n19963 & ~n19967 ) | ( n19963 & n19970 ) | ( ~n19967 & n19970 ) ;
  assign n19972 = n19796 | n19971 ;
  assign n19973 = ( n19782 & n19971 ) | ( n19782 & n19972 ) | ( n19971 & n19972 ) ;
  assign n19974 = n19802 | n19973 ;
  assign n19975 = ( n19800 & n19973 ) | ( n19800 & n19974 ) | ( n19973 & n19974 ) ;
  assign n19976 = n19796 & n19971 ;
  assign n19977 = n19782 & n19976 ;
  assign n19978 = ( n19802 & n19971 ) | ( n19802 & n19977 ) | ( n19971 & n19977 ) ;
  assign n19979 = n19971 & n19977 ;
  assign n19980 = ( n19800 & n19978 ) | ( n19800 & n19979 ) | ( n19978 & n19979 ) ;
  assign n19981 = n19975 & ~n19980 ;
  assign n19983 = x117 & n957 ;
  assign n19984 = x116 & ~n956 ;
  assign n19985 = n1105 & n19984 ;
  assign n19986 = n19983 | n19985 ;
  assign n19982 = x118 & n962 ;
  assign n19988 = n965 | n19982 ;
  assign n19989 = n19986 | n19988 ;
  assign n19987 = n19982 | n19986 ;
  assign n19990 = n19987 & n19989 ;
  assign n19991 = ( ~n14002 & n19989 ) | ( ~n14002 & n19990 ) | ( n19989 & n19990 ) ;
  assign n19992 = n19989 & n19990 ;
  assign n19993 = ( n13981 & n19991 ) | ( n13981 & n19992 ) | ( n19991 & n19992 ) ;
  assign n19994 = x14 & n19993 ;
  assign n19995 = x14 & ~n19993 ;
  assign n19996 = ( n19993 & ~n19994 ) | ( n19993 & n19995 ) | ( ~n19994 & n19995 ) ;
  assign n19997 = n19776 & n19996 ;
  assign n19998 = ( n19777 & n19996 ) | ( n19777 & n19997 ) | ( n19996 & n19997 ) ;
  assign n19999 = n19996 & n19997 ;
  assign n20000 = ( n19779 & n19998 ) | ( n19779 & n19999 ) | ( n19998 & n19999 ) ;
  assign n20001 = ( n19776 & n19780 ) | ( n19776 & ~n20000 ) | ( n19780 & ~n20000 ) ;
  assign n20003 = x102 & n3811 ;
  assign n20004 = x101 & ~n3810 ;
  assign n20005 = n4067 & n20004 ;
  assign n20006 = n20003 | n20005 ;
  assign n20002 = x103 & n3816 ;
  assign n20008 = n3819 | n20002 ;
  assign n20009 = n20006 | n20008 ;
  assign n20007 = n20002 | n20006 ;
  assign n20010 = n20007 & n20009 ;
  assign n20011 = ( n7529 & n20009 ) | ( n7529 & n20010 ) | ( n20009 & n20010 ) ;
  assign n20012 = x29 & n20010 ;
  assign n20013 = x29 & n20009 ;
  assign n20014 = ( n7529 & n20012 ) | ( n7529 & n20013 ) | ( n20012 & n20013 ) ;
  assign n20015 = x29 & ~n20010 ;
  assign n20016 = x29 & ~n20009 ;
  assign n20017 = ( ~n7529 & n20015 ) | ( ~n7529 & n20016 ) | ( n20015 & n20016 ) ;
  assign n20018 = ( n20011 & ~n20014 ) | ( n20011 & n20017 ) | ( ~n20014 & n20017 ) ;
  assign n20019 = n19641 & n20018 ;
  assign n20020 = n19639 & n20018 ;
  assign n20021 = ( n19620 & n20019 ) | ( n19620 & n20020 ) | ( n20019 & n20020 ) ;
  assign n20022 = ( n19647 & n20018 ) | ( n19647 & n20021 ) | ( n20018 & n20021 ) ;
  assign n20023 = n20018 & n20021 ;
  assign n20024 = ( n19646 & n20022 ) | ( n19646 & n20023 ) | ( n20022 & n20023 ) ;
  assign n20025 = n19641 | n20018 ;
  assign n20026 = n19639 | n20018 ;
  assign n20027 = ( n19620 & n20025 ) | ( n19620 & n20026 ) | ( n20025 & n20026 ) ;
  assign n20028 = n19647 | n20027 ;
  assign n20029 = ( n19646 & n20027 ) | ( n19646 & n20028 ) | ( n20027 & n20028 ) ;
  assign n20030 = ~n20024 & n20029 ;
  assign n20032 = x99 & n4626 ;
  assign n20033 = x98 & ~n4625 ;
  assign n20034 = n4943 & n20033 ;
  assign n20035 = n20032 | n20034 ;
  assign n20031 = x100 & n4631 ;
  assign n20037 = n4634 | n20031 ;
  assign n20038 = n20035 | n20037 ;
  assign n20036 = n20031 | n20035 ;
  assign n20039 = n20036 & n20038 ;
  assign n20040 = ( n6483 & n20038 ) | ( n6483 & n20039 ) | ( n20038 & n20039 ) ;
  assign n20041 = x32 & n20039 ;
  assign n20042 = x32 & n20038 ;
  assign n20043 = ( n6483 & n20041 ) | ( n6483 & n20042 ) | ( n20041 & n20042 ) ;
  assign n20044 = x32 & ~n20039 ;
  assign n20045 = x32 & ~n20038 ;
  assign n20046 = ( ~n6483 & n20044 ) | ( ~n6483 & n20045 ) | ( n20044 & n20045 ) ;
  assign n20047 = ( n20040 & ~n20043 ) | ( n20040 & n20046 ) | ( ~n20043 & n20046 ) ;
  assign n20048 = n19613 & n20047 ;
  assign n20049 = n19596 & n20048 ;
  assign n20050 = ( n19616 & n20047 ) | ( n19616 & n20049 ) | ( n20047 & n20049 ) ;
  assign n20051 = n20047 & n20048 ;
  assign n20052 = n19596 & n20051 ;
  assign n20053 = ( n19618 & n20050 ) | ( n19618 & n20052 ) | ( n20050 & n20052 ) ;
  assign n20054 = n19614 | n19616 ;
  assign n20055 = ( n19614 & n19618 ) | ( n19614 & n20054 ) | ( n19618 & n20054 ) ;
  assign n20056 = ~n20053 & n20055 ;
  assign n20057 = ( n18834 & n18842 ) | ( n18834 & n19389 ) | ( n18842 & n19389 ) ;
  assign n20058 = x67 & n18290 ;
  assign n20059 = x63 & x66 ;
  assign n20060 = ~n18290 & n20059 ;
  assign n20061 = n20058 | n20060 ;
  assign n20062 = x2 & n20061 ;
  assign n20063 = x2 | n20061 ;
  assign n20064 = ~n20062 & n20063 ;
  assign n20065 = x69 & n17141 ;
  assign n20066 = x68 & ~n17140 ;
  assign n20067 = n17724 & n20066 ;
  assign n20068 = n20065 | n20067 ;
  assign n20069 = x70 & n17146 ;
  assign n20070 = n17149 | n20069 ;
  assign n20071 = n20068 | n20070 ;
  assign n20072 = x62 & ~n20071 ;
  assign n20073 = n20068 | n20069 ;
  assign n20074 = x62 & ~n20073 ;
  assign n20075 = ( ~n340 & n20072 ) | ( ~n340 & n20074 ) | ( n20072 & n20074 ) ;
  assign n20076 = ~x62 & n20071 ;
  assign n20077 = ~x62 & n20073 ;
  assign n20078 = ( n340 & n20076 ) | ( n340 & n20077 ) | ( n20076 & n20077 ) ;
  assign n20079 = n20075 | n20078 ;
  assign n20080 = n20064 & n20079 ;
  assign n20081 = n20064 | n20079 ;
  assign n20082 = ~n20080 & n20081 ;
  assign n20083 = n19380 | n19386 ;
  assign n20084 = n19381 | n20083 ;
  assign n20085 = n20082 & n20084 ;
  assign n20086 = n19380 & n20082 ;
  assign n20087 = ( n20057 & n20085 ) | ( n20057 & n20086 ) | ( n20085 & n20086 ) ;
  assign n20088 = n20082 | n20084 ;
  assign n20089 = n19380 | n20082 ;
  assign n20090 = ( n20057 & n20088 ) | ( n20057 & n20089 ) | ( n20088 & n20089 ) ;
  assign n20091 = ~n20087 & n20090 ;
  assign n20092 = x73 & n15552 ;
  assign n20093 = x72 & n15547 ;
  assign n20094 = x71 & ~n15546 ;
  assign n20095 = n16123 & n20094 ;
  assign n20096 = n20093 | n20095 ;
  assign n20097 = n20092 | n20096 ;
  assign n20098 = ( ~n610 & n15555 ) | ( ~n610 & n20097 ) | ( n15555 & n20097 ) ;
  assign n20099 = n15555 & n20092 ;
  assign n20100 = ( n15555 & n20096 ) | ( n15555 & n20099 ) | ( n20096 & n20099 ) ;
  assign n20101 = ( n598 & n20098 ) | ( n598 & n20100 ) | ( n20098 & n20100 ) ;
  assign n20102 = ( x59 & ~n20097 ) | ( x59 & n20101 ) | ( ~n20097 & n20101 ) ;
  assign n20103 = ~n20101 & n20102 ;
  assign n20104 = x59 | n20092 ;
  assign n20105 = n20096 | n20104 ;
  assign n20106 = n20101 | n20105 ;
  assign n20107 = ( ~x59 & n20103 ) | ( ~x59 & n20106 ) | ( n20103 & n20106 ) ;
  assign n20108 = n20091 & ~n20107 ;
  assign n20109 = n20091 | n20107 ;
  assign n20110 = ( ~n20091 & n20108 ) | ( ~n20091 & n20109 ) | ( n20108 & n20109 ) ;
  assign n20111 = n19413 & ~n20110 ;
  assign n20112 = ( n19437 & ~n20110 ) | ( n19437 & n20111 ) | ( ~n20110 & n20111 ) ;
  assign n20113 = ~n19413 & n20110 ;
  assign n20114 = ~n19437 & n20113 ;
  assign n20115 = n20112 | n20114 ;
  assign n20116 = x76 & n14045 ;
  assign n20117 = x75 & n14040 ;
  assign n20118 = x74 & ~n14039 ;
  assign n20119 = n14552 & n20118 ;
  assign n20120 = n20117 | n20119 ;
  assign n20121 = n20116 | n20120 ;
  assign n20122 = n14048 | n20116 ;
  assign n20123 = n20120 | n20122 ;
  assign n20124 = ( n923 & n20121 ) | ( n923 & n20123 ) | ( n20121 & n20123 ) ;
  assign n20125 = x56 & n20123 ;
  assign n20126 = x56 & n20116 ;
  assign n20127 = ( x56 & n20120 ) | ( x56 & n20126 ) | ( n20120 & n20126 ) ;
  assign n20128 = ( n923 & n20125 ) | ( n923 & n20127 ) | ( n20125 & n20127 ) ;
  assign n20129 = x56 & ~n20127 ;
  assign n20130 = x56 & ~n20123 ;
  assign n20131 = ( ~n923 & n20129 ) | ( ~n923 & n20130 ) | ( n20129 & n20130 ) ;
  assign n20132 = ( n20124 & ~n20128 ) | ( n20124 & n20131 ) | ( ~n20128 & n20131 ) ;
  assign n20133 = n20115 | n20132 ;
  assign n20134 = n20115 & n20132 ;
  assign n20135 = n20133 & ~n20134 ;
  assign n20136 = n19440 & n20135 ;
  assign n20137 = ( n19445 & n20135 ) | ( n19445 & n20136 ) | ( n20135 & n20136 ) ;
  assign n20138 = n19440 | n20135 ;
  assign n20139 = n19445 | n20138 ;
  assign n20140 = ~n20137 & n20139 ;
  assign n20141 = x79 & n12574 ;
  assign n20142 = x78 & n12569 ;
  assign n20143 = x77 & ~n12568 ;
  assign n20144 = n13076 & n20143 ;
  assign n20145 = n20142 | n20144 ;
  assign n20146 = n20141 | n20145 ;
  assign n20147 = n12577 | n20141 ;
  assign n20148 = n20145 | n20147 ;
  assign n20149 = ( n1332 & n20146 ) | ( n1332 & n20148 ) | ( n20146 & n20148 ) ;
  assign n20150 = x53 & n20148 ;
  assign n20151 = x53 & n20141 ;
  assign n20152 = ( x53 & n20145 ) | ( x53 & n20151 ) | ( n20145 & n20151 ) ;
  assign n20153 = ( n1332 & n20150 ) | ( n1332 & n20152 ) | ( n20150 & n20152 ) ;
  assign n20154 = x53 & ~n20152 ;
  assign n20155 = x53 & ~n20148 ;
  assign n20156 = ( ~n1332 & n20154 ) | ( ~n1332 & n20155 ) | ( n20154 & n20155 ) ;
  assign n20157 = ( n20149 & ~n20153 ) | ( n20149 & n20156 ) | ( ~n20153 & n20156 ) ;
  assign n20158 = n20140 & ~n20157 ;
  assign n20159 = n20140 | n20157 ;
  assign n20160 = ( ~n20140 & n20158 ) | ( ~n20140 & n20159 ) | ( n20158 & n20159 ) ;
  assign n20161 = ( n19447 & n19464 ) | ( n19447 & n19470 ) | ( n19464 & n19470 ) ;
  assign n20162 = n20160 | n20161 ;
  assign n20163 = n20160 & n20161 ;
  assign n20164 = n20162 & ~n20163 ;
  assign n20165 = x82 & n11205 ;
  assign n20166 = x81 & n11200 ;
  assign n20167 = x80 & ~n11199 ;
  assign n20168 = n11679 & n20167 ;
  assign n20169 = n20166 | n20168 ;
  assign n20170 = n20165 | n20169 ;
  assign n20171 = n11208 | n20165 ;
  assign n20172 = n20169 | n20171 ;
  assign n20173 = ( n1811 & n20170 ) | ( n1811 & n20172 ) | ( n20170 & n20172 ) ;
  assign n20174 = x50 & n20172 ;
  assign n20175 = x50 & n20165 ;
  assign n20176 = ( x50 & n20169 ) | ( x50 & n20175 ) | ( n20169 & n20175 ) ;
  assign n20177 = ( n1811 & n20174 ) | ( n1811 & n20176 ) | ( n20174 & n20176 ) ;
  assign n20178 = x50 & ~n20176 ;
  assign n20179 = x50 & ~n20172 ;
  assign n20180 = ( ~n1811 & n20178 ) | ( ~n1811 & n20179 ) | ( n20178 & n20179 ) ;
  assign n20181 = ( n20173 & ~n20177 ) | ( n20173 & n20180 ) | ( ~n20177 & n20180 ) ;
  assign n20182 = ~n20164 & n20181 ;
  assign n20183 = n20163 | n20181 ;
  assign n20184 = n20162 & ~n20183 ;
  assign n20185 = n20182 | n20184 ;
  assign n20186 = n19491 | n19493 ;
  assign n20187 = ( n19491 & n19494 ) | ( n19491 & n20186 ) | ( n19494 & n20186 ) ;
  assign n20188 = n20185 | n20187 ;
  assign n20189 = n20185 & n20187 ;
  assign n20190 = n20188 & ~n20189 ;
  assign n20191 = x85 & n9933 ;
  assign n20192 = x84 & n9928 ;
  assign n20193 = x83 & ~n9927 ;
  assign n20194 = n10379 & n20193 ;
  assign n20195 = n20192 | n20194 ;
  assign n20196 = n20191 | n20195 ;
  assign n20197 = n9936 | n20191 ;
  assign n20198 = n20195 | n20197 ;
  assign n20199 = ( n2381 & n20196 ) | ( n2381 & n20198 ) | ( n20196 & n20198 ) ;
  assign n20200 = x47 & n20198 ;
  assign n20201 = x47 & n20191 ;
  assign n20202 = ( x47 & n20195 ) | ( x47 & n20201 ) | ( n20195 & n20201 ) ;
  assign n20203 = ( n2381 & n20200 ) | ( n2381 & n20202 ) | ( n20200 & n20202 ) ;
  assign n20204 = x47 & ~n20202 ;
  assign n20205 = x47 & ~n20198 ;
  assign n20206 = ( ~n2381 & n20204 ) | ( ~n2381 & n20205 ) | ( n20204 & n20205 ) ;
  assign n20207 = ( n20199 & ~n20203 ) | ( n20199 & n20206 ) | ( ~n20203 & n20206 ) ;
  assign n20208 = n20190 | n20207 ;
  assign n20209 = n20190 & n20207 ;
  assign n20210 = n20208 & ~n20209 ;
  assign n20211 = ( n18962 & n19497 ) | ( n18962 & n19514 ) | ( n19497 & n19514 ) ;
  assign n20212 = n19497 | n19514 ;
  assign n20213 = ( n18966 & n20211 ) | ( n18966 & n20212 ) | ( n20211 & n20212 ) ;
  assign n20214 = n20210 & n20213 ;
  assign n20215 = n20210 | n20213 ;
  assign n20216 = ~n20214 & n20215 ;
  assign n20217 = x88 & n8724 ;
  assign n20218 = x87 & n8719 ;
  assign n20219 = x86 & ~n8718 ;
  assign n20220 = n9149 & n20219 ;
  assign n20221 = n20218 | n20220 ;
  assign n20222 = n20217 | n20221 ;
  assign n20223 = n8727 | n20217 ;
  assign n20224 = n20221 | n20223 ;
  assign n20225 = ( ~n3039 & n20222 ) | ( ~n3039 & n20224 ) | ( n20222 & n20224 ) ;
  assign n20226 = n20222 & n20224 ;
  assign n20227 = ( n3023 & n20225 ) | ( n3023 & n20226 ) | ( n20225 & n20226 ) ;
  assign n20228 = x44 & n20224 ;
  assign n20229 = x44 & n20217 ;
  assign n20230 = ( x44 & n20221 ) | ( x44 & n20229 ) | ( n20221 & n20229 ) ;
  assign n20231 = ( ~n3039 & n20228 ) | ( ~n3039 & n20230 ) | ( n20228 & n20230 ) ;
  assign n20232 = n20228 & n20230 ;
  assign n20233 = ( n3023 & n20231 ) | ( n3023 & n20232 ) | ( n20231 & n20232 ) ;
  assign n20234 = x44 & ~n20230 ;
  assign n20235 = x44 & ~n20224 ;
  assign n20236 = ( n3039 & n20234 ) | ( n3039 & n20235 ) | ( n20234 & n20235 ) ;
  assign n20237 = n20234 | n20235 ;
  assign n20238 = ( ~n3023 & n20236 ) | ( ~n3023 & n20237 ) | ( n20236 & n20237 ) ;
  assign n20239 = ( n20227 & ~n20233 ) | ( n20227 & n20238 ) | ( ~n20233 & n20238 ) ;
  assign n20240 = n20216 & ~n20239 ;
  assign n20241 = n20216 | n20239 ;
  assign n20242 = ( ~n20216 & n20240 ) | ( ~n20216 & n20241 ) | ( n20240 & n20241 ) ;
  assign n20243 = n19539 & n20242 ;
  assign n20244 = ( n19543 & n20242 ) | ( n19543 & n20243 ) | ( n20242 & n20243 ) ;
  assign n20245 = n19539 | n20242 ;
  assign n20246 = n19543 | n20245 ;
  assign n20247 = ~n20244 & n20246 ;
  assign n20248 = x91 & n7566 ;
  assign n20249 = x90 & n7561 ;
  assign n20250 = x89 & ~n7560 ;
  assign n20251 = n7953 & n20250 ;
  assign n20252 = n20249 | n20251 ;
  assign n20253 = n20248 | n20252 ;
  assign n20254 = n7569 | n20248 ;
  assign n20255 = n20252 | n20254 ;
  assign n20256 = ( n3768 & n20253 ) | ( n3768 & n20255 ) | ( n20253 & n20255 ) ;
  assign n20257 = x41 & n20255 ;
  assign n20258 = x41 & n20248 ;
  assign n20259 = ( x41 & n20252 ) | ( x41 & n20258 ) | ( n20252 & n20258 ) ;
  assign n20260 = ( n3768 & n20257 ) | ( n3768 & n20259 ) | ( n20257 & n20259 ) ;
  assign n20261 = x41 & ~n20259 ;
  assign n20262 = x41 & ~n20255 ;
  assign n20263 = ( ~n3768 & n20261 ) | ( ~n3768 & n20262 ) | ( n20261 & n20262 ) ;
  assign n20264 = ( n20256 & ~n20260 ) | ( n20256 & n20263 ) | ( ~n20260 & n20263 ) ;
  assign n20265 = ~n20247 & n20264 ;
  assign n20266 = n20244 | n20264 ;
  assign n20267 = n20246 & ~n20266 ;
  assign n20268 = n20265 | n20267 ;
  assign n20269 = n19562 & n20268 ;
  assign n20270 = ( n19568 & n20268 ) | ( n19568 & n20269 ) | ( n20268 & n20269 ) ;
  assign n20271 = n19562 | n20268 ;
  assign n20272 = n19568 | n20271 ;
  assign n20273 = ~n20270 & n20272 ;
  assign n20274 = x94 & n6536 ;
  assign n20275 = x93 & n6531 ;
  assign n20276 = x92 & ~n6530 ;
  assign n20277 = n6871 & n20276 ;
  assign n20278 = n20275 | n20277 ;
  assign n20279 = n20274 | n20278 ;
  assign n20280 = n6539 | n20274 ;
  assign n20281 = n20278 | n20280 ;
  assign n20282 = ( n4583 & n20279 ) | ( n4583 & n20281 ) | ( n20279 & n20281 ) ;
  assign n20283 = x38 & n20281 ;
  assign n20284 = x38 & n20274 ;
  assign n20285 = ( x38 & n20278 ) | ( x38 & n20284 ) | ( n20278 & n20284 ) ;
  assign n20286 = ( n4583 & n20283 ) | ( n4583 & n20285 ) | ( n20283 & n20285 ) ;
  assign n20287 = x38 & ~n20285 ;
  assign n20288 = x38 & ~n20281 ;
  assign n20289 = ( ~n4583 & n20287 ) | ( ~n4583 & n20288 ) | ( n20287 & n20288 ) ;
  assign n20290 = ( n20282 & ~n20286 ) | ( n20282 & n20289 ) | ( ~n20286 & n20289 ) ;
  assign n20291 = n20273 | n20290 ;
  assign n20292 = n20273 & n20290 ;
  assign n20293 = n20291 & ~n20292 ;
  assign n20294 = n19587 & n20293 ;
  assign n20295 = ( n19595 & n20293 ) | ( n19595 & n20294 ) | ( n20293 & n20294 ) ;
  assign n20296 = n19587 | n20293 ;
  assign n20297 = n19595 | n20296 ;
  assign n20298 = ~n20295 & n20297 ;
  assign n20299 = x97 & n5554 ;
  assign n20300 = x96 & n5549 ;
  assign n20301 = x95 & ~n5548 ;
  assign n20302 = n5893 & n20301 ;
  assign n20303 = n20300 | n20302 ;
  assign n20304 = n20299 | n20303 ;
  assign n20305 = n5557 | n20299 ;
  assign n20306 = n20303 | n20305 ;
  assign n20307 = ( n5505 & n20304 ) | ( n5505 & n20306 ) | ( n20304 & n20306 ) ;
  assign n20308 = x35 & n20306 ;
  assign n20309 = x35 & n20299 ;
  assign n20310 = ( x35 & n20303 ) | ( x35 & n20309 ) | ( n20303 & n20309 ) ;
  assign n20311 = ( n5505 & n20308 ) | ( n5505 & n20310 ) | ( n20308 & n20310 ) ;
  assign n20312 = x35 & ~n20310 ;
  assign n20313 = x35 & ~n20306 ;
  assign n20314 = ( ~n5505 & n20312 ) | ( ~n5505 & n20313 ) | ( n20312 & n20313 ) ;
  assign n20315 = ( n20307 & ~n20311 ) | ( n20307 & n20314 ) | ( ~n20311 & n20314 ) ;
  assign n20316 = n20298 & ~n20315 ;
  assign n20317 = n20298 | n20315 ;
  assign n20318 = ( ~n20298 & n20316 ) | ( ~n20298 & n20317 ) | ( n20316 & n20317 ) ;
  assign n20319 = n20047 & ~n20048 ;
  assign n20320 = ( ~n19596 & n20047 ) | ( ~n19596 & n20319 ) | ( n20047 & n20319 ) ;
  assign n20321 = ~n19616 & n20320 ;
  assign n20322 = ( ~n19618 & n20320 ) | ( ~n19618 & n20321 ) | ( n20320 & n20321 ) ;
  assign n20323 = n20318 & n20322 ;
  assign n20324 = ( n20056 & n20318 ) | ( n20056 & n20323 ) | ( n20318 & n20323 ) ;
  assign n20325 = n20318 | n20322 ;
  assign n20326 = n20056 | n20325 ;
  assign n20327 = ~n20324 & n20326 ;
  assign n20328 = n20030 & ~n20327 ;
  assign n20329 = n20030 | n20327 ;
  assign n20330 = ( ~n20030 & n20328 ) | ( ~n20030 & n20329 ) | ( n20328 & n20329 ) ;
  assign n20331 = x106 & n3085 ;
  assign n20332 = x105 & n3080 ;
  assign n20333 = x104 & ~n3079 ;
  assign n20334 = n3309 & n20333 ;
  assign n20335 = n20332 | n20334 ;
  assign n20336 = n20331 | n20335 ;
  assign n20337 = n3088 | n20331 ;
  assign n20338 = n20335 | n20337 ;
  assign n20339 = ( n8656 & n20336 ) | ( n8656 & n20338 ) | ( n20336 & n20338 ) ;
  assign n20340 = x26 & n20338 ;
  assign n20341 = x26 & n20331 ;
  assign n20342 = ( x26 & n20335 ) | ( x26 & n20341 ) | ( n20335 & n20341 ) ;
  assign n20343 = ( n8656 & n20340 ) | ( n8656 & n20342 ) | ( n20340 & n20342 ) ;
  assign n20344 = x26 & ~n20342 ;
  assign n20345 = x26 & ~n20338 ;
  assign n20346 = ( ~n8656 & n20344 ) | ( ~n8656 & n20345 ) | ( n20344 & n20345 ) ;
  assign n20347 = ( n20339 & ~n20343 ) | ( n20339 & n20346 ) | ( ~n20343 & n20346 ) ;
  assign n20348 = n19667 | n20347 ;
  assign n20349 = ( n19650 & n20347 ) | ( n19650 & n20348 ) | ( n20347 & n20348 ) ;
  assign n20350 = n19672 | n20349 ;
  assign n20351 = ( n19671 & n20349 ) | ( n19671 & n20350 ) | ( n20349 & n20350 ) ;
  assign n20352 = n19667 & n20347 ;
  assign n20353 = n19650 & n20352 ;
  assign n20354 = ( n19672 & n20347 ) | ( n19672 & n20353 ) | ( n20347 & n20353 ) ;
  assign n20355 = n20347 & n20353 ;
  assign n20356 = ( n19671 & n20354 ) | ( n19671 & n20355 ) | ( n20354 & n20355 ) ;
  assign n20357 = n20351 & ~n20356 ;
  assign n20358 = n19693 | n19695 ;
  assign n20359 = ( n19693 & n19697 ) | ( n19693 & n20358 ) | ( n19697 & n20358 ) ;
  assign n20360 = x109 & n2429 ;
  assign n20361 = x108 & n2424 ;
  assign n20362 = x107 & ~n2423 ;
  assign n20363 = n2631 & n20362 ;
  assign n20364 = n20361 | n20363 ;
  assign n20365 = n20360 | n20364 ;
  assign n20366 = n2432 | n20360 ;
  assign n20367 = n20364 | n20366 ;
  assign n20368 = ( n9878 & n20365 ) | ( n9878 & n20367 ) | ( n20365 & n20367 ) ;
  assign n20369 = x23 & n20367 ;
  assign n20370 = x23 & n20360 ;
  assign n20371 = ( x23 & n20364 ) | ( x23 & n20370 ) | ( n20364 & n20370 ) ;
  assign n20372 = ( n9878 & n20369 ) | ( n9878 & n20371 ) | ( n20369 & n20371 ) ;
  assign n20373 = x23 & ~n20371 ;
  assign n20374 = x23 & ~n20367 ;
  assign n20375 = ( ~n9878 & n20373 ) | ( ~n9878 & n20374 ) | ( n20373 & n20374 ) ;
  assign n20376 = ( n20368 & ~n20372 ) | ( n20368 & n20375 ) | ( ~n20372 & n20375 ) ;
  assign n20377 = n19697 | n20376 ;
  assign n20378 = n19693 | n20376 ;
  assign n20379 = ( n20358 & n20377 ) | ( n20358 & n20378 ) | ( n20377 & n20378 ) ;
  assign n20380 = n19697 & ~n20376 ;
  assign n20381 = n19693 & ~n20376 ;
  assign n20382 = ( n20358 & n20380 ) | ( n20358 & n20381 ) | ( n20380 & n20381 ) ;
  assign n20383 = ( ~n20359 & n20379 ) | ( ~n20359 & n20382 ) | ( n20379 & n20382 ) ;
  assign n20384 = ( n20330 & ~n20357 ) | ( n20330 & n20383 ) | ( ~n20357 & n20383 ) ;
  assign n20385 = ( n20357 & ~n20383 ) | ( n20357 & n20384 ) | ( ~n20383 & n20384 ) ;
  assign n20386 = ( ~n20330 & n20384 ) | ( ~n20330 & n20385 ) | ( n20384 & n20385 ) ;
  assign n20387 = x115 & n1383 ;
  assign n20388 = x114 & n1378 ;
  assign n20389 = x113 & ~n1377 ;
  assign n20390 = n1542 & n20389 ;
  assign n20391 = n20388 | n20390 ;
  assign n20392 = n20387 | n20391 ;
  assign n20393 = n1386 | n20387 ;
  assign n20394 = n20391 | n20393 ;
  assign n20395 = ( ~n12550 & n20392 ) | ( ~n12550 & n20394 ) | ( n20392 & n20394 ) ;
  assign n20396 = n20392 & n20394 ;
  assign n20397 = ( n12532 & n20395 ) | ( n12532 & n20396 ) | ( n20395 & n20396 ) ;
  assign n20398 = x17 & n20397 ;
  assign n20399 = x17 & ~n20397 ;
  assign n20400 = ( n20397 & ~n20398 ) | ( n20397 & n20399 ) | ( ~n20398 & n20399 ) ;
  assign n20401 = n19751 & n20400 ;
  assign n20402 = n19734 & n20401 ;
  assign n20403 = ( n19754 & n20400 ) | ( n19754 & n20402 ) | ( n20400 & n20402 ) ;
  assign n20404 = n20400 | n20402 ;
  assign n20405 = ( n19753 & n20403 ) | ( n19753 & n20404 ) | ( n20403 & n20404 ) ;
  assign n20406 = n20400 & n20401 ;
  assign n20407 = n19734 & n20406 ;
  assign n20408 = ( n19353 & n20405 ) | ( n19353 & n20407 ) | ( n20405 & n20407 ) ;
  assign n20409 = n19751 | n20400 ;
  assign n20410 = ( n19734 & n20400 ) | ( n19734 & n20409 ) | ( n20400 & n20409 ) ;
  assign n20411 = n19754 | n20410 ;
  assign n20412 = n19753 | n20411 ;
  assign n20413 = ( n19353 & n20410 ) | ( n19353 & n20412 ) | ( n20410 & n20412 ) ;
  assign n20414 = ~n20408 & n20413 ;
  assign n20415 = x112 & n1859 ;
  assign n20416 = x111 & n1854 ;
  assign n20417 = x110 & ~n1853 ;
  assign n20418 = n2037 & n20417 ;
  assign n20419 = n20416 | n20418 ;
  assign n20420 = n20415 | n20419 ;
  assign n20421 = n1862 | n20415 ;
  assign n20422 = n20419 | n20421 ;
  assign n20423 = ( n11172 & n20420 ) | ( n11172 & n20422 ) | ( n20420 & n20422 ) ;
  assign n20424 = x20 & n20422 ;
  assign n20425 = x20 & n20415 ;
  assign n20426 = ( x20 & n20419 ) | ( x20 & n20425 ) | ( n20419 & n20425 ) ;
  assign n20427 = ( n11172 & n20424 ) | ( n11172 & n20426 ) | ( n20424 & n20426 ) ;
  assign n20428 = x20 & ~n20426 ;
  assign n20429 = x20 & ~n20422 ;
  assign n20430 = ( ~n11172 & n20428 ) | ( ~n11172 & n20429 ) | ( n20428 & n20429 ) ;
  assign n20431 = ( n20423 & ~n20427 ) | ( n20423 & n20430 ) | ( ~n20427 & n20430 ) ;
  assign n20432 = n19720 | n20431 ;
  assign n20433 = n19726 | n20432 ;
  assign n20434 = n19721 | n20432 ;
  assign n20435 = ( n19730 & n20433 ) | ( n19730 & n20434 ) | ( n20433 & n20434 ) ;
  assign n20436 = n19720 & n20431 ;
  assign n20437 = ( n19726 & n20431 ) | ( n19726 & n20436 ) | ( n20431 & n20436 ) ;
  assign n20438 = ( n19721 & n20431 ) | ( n19721 & n20436 ) | ( n20431 & n20436 ) ;
  assign n20439 = ( n19730 & n20437 ) | ( n19730 & n20438 ) | ( n20437 & n20438 ) ;
  assign n20440 = n20435 & ~n20439 ;
  assign n20441 = ( n20386 & n20414 ) | ( n20386 & ~n20440 ) | ( n20414 & ~n20440 ) ;
  assign n20442 = ( ~n20414 & n20440 ) | ( ~n20414 & n20441 ) | ( n20440 & n20441 ) ;
  assign n20443 = ( ~n20386 & n20441 ) | ( ~n20386 & n20442 ) | ( n20441 & n20442 ) ;
  assign n20444 = ~n19776 & n19996 ;
  assign n20445 = ~n19777 & n20444 ;
  assign n20446 = ( ~n19779 & n20444 ) | ( ~n19779 & n20445 ) | ( n20444 & n20445 ) ;
  assign n20447 = n20443 & n20446 ;
  assign n20448 = ( n20001 & n20443 ) | ( n20001 & n20447 ) | ( n20443 & n20447 ) ;
  assign n20449 = n20443 | n20446 ;
  assign n20450 = n20001 | n20449 ;
  assign n20451 = ~n20448 & n20450 ;
  assign n20452 = ~n19981 & n20451 ;
  assign n20453 = n19977 | n20451 ;
  assign n20454 = n19971 | n20451 ;
  assign n20455 = ( n19804 & n20453 ) | ( n19804 & n20454 ) | ( n20453 & n20454 ) ;
  assign n20456 = n19975 & ~n20455 ;
  assign n20457 = n20452 | n20456 ;
  assign n20458 = ( n19824 & n19825 ) | ( n19824 & n19847 ) | ( n19825 & n19847 ) ;
  assign n20459 = x124 & n389 ;
  assign n20460 = x123 & n384 ;
  assign n20461 = x122 & ~n383 ;
  assign n20462 = n463 & n20461 ;
  assign n20463 = n20460 | n20462 ;
  assign n20464 = n20459 | n20463 ;
  assign n20465 = n392 | n20459 ;
  assign n20466 = n20463 | n20465 ;
  assign n20467 = ( n17084 & n20464 ) | ( n17084 & n20466 ) | ( n20464 & n20466 ) ;
  assign n20468 = x8 & n20466 ;
  assign n20469 = x8 & n20459 ;
  assign n20470 = ( x8 & n20463 ) | ( x8 & n20469 ) | ( n20463 & n20469 ) ;
  assign n20471 = ( n17084 & n20468 ) | ( n17084 & n20470 ) | ( n20468 & n20470 ) ;
  assign n20472 = x8 & ~n20470 ;
  assign n20473 = x8 & ~n20466 ;
  assign n20474 = ( ~n17084 & n20472 ) | ( ~n17084 & n20473 ) | ( n20472 & n20473 ) ;
  assign n20475 = ( n20467 & ~n20471 ) | ( n20467 & n20474 ) | ( ~n20471 & n20474 ) ;
  assign n20476 = n19847 & n20475 ;
  assign n20477 = n19824 & n20475 ;
  assign n20478 = ( n19825 & n20476 ) | ( n19825 & n20477 ) | ( n20476 & n20477 ) ;
  assign n20479 = n20458 & ~n20478 ;
  assign n20480 = ~n19847 & n20475 ;
  assign n20481 = ~n19824 & n20475 ;
  assign n20482 = ( ~n19825 & n20480 ) | ( ~n19825 & n20481 ) | ( n20480 & n20481 ) ;
  assign n20483 = n20457 & n20482 ;
  assign n20484 = ( n20457 & n20479 ) | ( n20457 & n20483 ) | ( n20479 & n20483 ) ;
  assign n20485 = n20457 | n20482 ;
  assign n20486 = n20479 | n20485 ;
  assign n20487 = ~n20484 & n20486 ;
  assign n20488 = n19950 & ~n19952 ;
  assign n20489 = n20487 & n20488 ;
  assign n20490 = ( n19954 & n20487 ) | ( n19954 & n20489 ) | ( n20487 & n20489 ) ;
  assign n20491 = n20487 | n20488 ;
  assign n20492 = n19954 | n20491 ;
  assign n20493 = ~n20490 & n20492 ;
  assign n20494 = n19910 | n19918 ;
  assign n20495 = ( n19874 & n19910 ) | ( n19874 & n20494 ) | ( n19910 & n20494 ) ;
  assign n20496 = n20493 | n20495 ;
  assign n20497 = n20493 & n20495 ;
  assign n20498 = n20496 & ~n20497 ;
  assign n20499 = n19925 | n19932 ;
  assign n20500 = n20498 | n20499 ;
  assign n20501 = n19925 & n20498 ;
  assign n20502 = ( n19932 & n20498 ) | ( n19932 & n20501 ) | ( n20498 & n20501 ) ;
  assign n20503 = n20500 & ~n20502 ;
  assign n20504 = n19953 | n20490 ;
  assign n20505 = n20478 | n20484 ;
  assign n20506 = x127 & n207 ;
  assign n20507 = x126 & ~n206 ;
  assign n20508 = n267 & n20507 ;
  assign n20509 = n20506 | n20508 ;
  assign n20510 = n215 | n20509 ;
  assign n20511 = ( n19328 & n20509 ) | ( n19328 & n20510 ) | ( n20509 & n20510 ) ;
  assign n20512 = x5 & n20509 ;
  assign n20513 = x5 & n215 ;
  assign n20514 = ( x5 & n20509 ) | ( x5 & n20513 ) | ( n20509 & n20513 ) ;
  assign n20515 = ( n19328 & n20512 ) | ( n19328 & n20514 ) | ( n20512 & n20514 ) ;
  assign n20516 = x5 & ~n20513 ;
  assign n20517 = ~n20509 & n20516 ;
  assign n20518 = x5 & ~n20509 ;
  assign n20519 = ( ~n19328 & n20517 ) | ( ~n19328 & n20518 ) | ( n20517 & n20518 ) ;
  assign n20520 = ( n20511 & ~n20515 ) | ( n20511 & n20519 ) | ( ~n20515 & n20519 ) ;
  assign n20521 = n20475 & n20520 ;
  assign n20522 = n19847 & n20521 ;
  assign n20523 = n19824 & n20521 ;
  assign n20524 = ( n19825 & n20522 ) | ( n19825 & n20523 ) | ( n20522 & n20523 ) ;
  assign n20525 = ( n20484 & n20520 ) | ( n20484 & n20524 ) | ( n20520 & n20524 ) ;
  assign n20526 = n20505 & ~n20525 ;
  assign n20527 = n20520 & ~n20521 ;
  assign n20528 = ( ~n19847 & n20520 ) | ( ~n19847 & n20527 ) | ( n20520 & n20527 ) ;
  assign n20529 = ( ~n19824 & n20520 ) | ( ~n19824 & n20527 ) | ( n20520 & n20527 ) ;
  assign n20530 = ( ~n19825 & n20528 ) | ( ~n19825 & n20529 ) | ( n20528 & n20529 ) ;
  assign n20531 = ~n20484 & n20530 ;
  assign n20549 = n19980 | n20451 ;
  assign n20550 = ( n19980 & n19981 ) | ( n19980 & n20549 ) | ( n19981 & n20549 ) ;
  assign n20533 = x124 & n384 ;
  assign n20534 = x123 & ~n383 ;
  assign n20535 = n463 & n20534 ;
  assign n20536 = n20533 | n20535 ;
  assign n20532 = x125 & n389 ;
  assign n20538 = n392 | n20532 ;
  assign n20539 = n20536 | n20538 ;
  assign n20537 = n20532 | n20536 ;
  assign n20540 = n20537 & n20539 ;
  assign n20541 = ( n17670 & n20539 ) | ( n17670 & n20540 ) | ( n20539 & n20540 ) ;
  assign n20542 = x8 & n20540 ;
  assign n20543 = x8 & n20539 ;
  assign n20544 = ( n17670 & n20542 ) | ( n17670 & n20543 ) | ( n20542 & n20543 ) ;
  assign n20545 = x8 & ~n20540 ;
  assign n20546 = x8 & ~n20539 ;
  assign n20547 = ( ~n17670 & n20545 ) | ( ~n17670 & n20546 ) | ( n20545 & n20546 ) ;
  assign n20548 = ( n20541 & ~n20544 ) | ( n20541 & n20547 ) | ( ~n20544 & n20547 ) ;
  assign n20551 = n20548 & n20550 ;
  assign n20552 = n20550 & ~n20551 ;
  assign n20553 = x119 & n962 ;
  assign n20554 = x118 & n957 ;
  assign n20555 = x117 & ~n956 ;
  assign n20556 = n1105 & n20555 ;
  assign n20557 = n20554 | n20556 ;
  assign n20558 = n20553 | n20557 ;
  assign n20559 = n965 | n20553 ;
  assign n20560 = n20557 | n20559 ;
  assign n20561 = ( n14496 & n20558 ) | ( n14496 & n20560 ) | ( n20558 & n20560 ) ;
  assign n20562 = x14 & n20560 ;
  assign n20563 = x14 & n20553 ;
  assign n20564 = ( x14 & n20557 ) | ( x14 & n20563 ) | ( n20557 & n20563 ) ;
  assign n20565 = ( n14496 & n20562 ) | ( n14496 & n20564 ) | ( n20562 & n20564 ) ;
  assign n20566 = x14 & ~n20564 ;
  assign n20567 = x14 & ~n20560 ;
  assign n20568 = ( ~n14496 & n20566 ) | ( ~n14496 & n20567 ) | ( n20566 & n20567 ) ;
  assign n20569 = ( n20561 & ~n20565 ) | ( n20561 & n20568 ) | ( ~n20565 & n20568 ) ;
  assign n20570 = n20386 & n20440 ;
  assign n20571 = n20386 | n20440 ;
  assign n20572 = ~n20570 & n20571 ;
  assign n20573 = n20408 | n20572 ;
  assign n20574 = ( n20408 & n20414 ) | ( n20408 & n20573 ) | ( n20414 & n20573 ) ;
  assign n20575 = n20569 | n20574 ;
  assign n20576 = n20569 & n20574 ;
  assign n20577 = n20575 & ~n20576 ;
  assign n20578 = x113 & n1859 ;
  assign n20579 = x112 & n1854 ;
  assign n20580 = x111 & ~n1853 ;
  assign n20581 = n2037 & n20580 ;
  assign n20582 = n20579 | n20581 ;
  assign n20583 = n20578 | n20582 ;
  assign n20584 = n1862 | n20578 ;
  assign n20585 = n20582 | n20584 ;
  assign n20586 = ( ~n11642 & n20583 ) | ( ~n11642 & n20585 ) | ( n20583 & n20585 ) ;
  assign n20587 = n20583 & n20585 ;
  assign n20588 = ( n11626 & n20586 ) | ( n11626 & n20587 ) | ( n20586 & n20587 ) ;
  assign n20589 = x20 & n20588 ;
  assign n20590 = x20 & ~n20588 ;
  assign n20591 = ( n20588 & ~n20589 ) | ( n20588 & n20590 ) | ( ~n20589 & n20590 ) ;
  assign n20592 = n19692 & n20376 ;
  assign n20593 = n19675 & n20592 ;
  assign n20594 = ( n19695 & n20376 ) | ( n19695 & n20593 ) | ( n20376 & n20593 ) ;
  assign n20595 = n20330 & n20357 ;
  assign n20596 = n20330 | n20357 ;
  assign n20597 = ~n20595 & n20596 ;
  assign n20598 = n19697 | n20597 ;
  assign n20599 = n20376 & n20592 ;
  assign n20600 = n19675 & n20599 ;
  assign n20601 = n20597 | n20600 ;
  assign n20602 = ( n20594 & n20598 ) | ( n20594 & n20601 ) | ( n20598 & n20601 ) ;
  assign n20603 = n20591 | n20602 ;
  assign n20604 = n19697 | n20591 ;
  assign n20605 = n20591 | n20600 ;
  assign n20606 = ( n20594 & n20604 ) | ( n20594 & n20605 ) | ( n20604 & n20605 ) ;
  assign n20607 = ( n20383 & n20603 ) | ( n20383 & n20606 ) | ( n20603 & n20606 ) ;
  assign n20608 = n20591 & n20602 ;
  assign n20609 = n19697 & n20591 ;
  assign n20610 = n20591 & n20600 ;
  assign n20611 = ( n20594 & n20609 ) | ( n20594 & n20610 ) | ( n20609 & n20610 ) ;
  assign n20612 = ( n20383 & n20608 ) | ( n20383 & n20611 ) | ( n20608 & n20611 ) ;
  assign n20613 = n20607 & ~n20612 ;
  assign n20614 = x107 & n3085 ;
  assign n20615 = x106 & n3080 ;
  assign n20616 = x105 & ~n3079 ;
  assign n20617 = n3309 & n20616 ;
  assign n20618 = n20615 | n20617 ;
  assign n20619 = n20614 | n20618 ;
  assign n20620 = n3088 | n20614 ;
  assign n20621 = n20618 | n20620 ;
  assign n20622 = ( n9084 & n20619 ) | ( n9084 & n20621 ) | ( n20619 & n20621 ) ;
  assign n20623 = x26 & n20621 ;
  assign n20624 = x26 & n20614 ;
  assign n20625 = ( x26 & n20618 ) | ( x26 & n20624 ) | ( n20618 & n20624 ) ;
  assign n20626 = ( n9084 & n20623 ) | ( n9084 & n20625 ) | ( n20623 & n20625 ) ;
  assign n20627 = x26 & ~n20625 ;
  assign n20628 = x26 & ~n20621 ;
  assign n20629 = ( ~n9084 & n20627 ) | ( ~n9084 & n20628 ) | ( n20627 & n20628 ) ;
  assign n20630 = ( n20622 & ~n20626 ) | ( n20622 & n20629 ) | ( ~n20626 & n20629 ) ;
  assign n20631 = n20024 | n20327 ;
  assign n20632 = ( n20024 & n20030 ) | ( n20024 & n20631 ) | ( n20030 & n20631 ) ;
  assign n20633 = n20630 | n20632 ;
  assign n20634 = n20630 & n20632 ;
  assign n20635 = n20633 & ~n20634 ;
  assign n20637 = x100 & n4626 ;
  assign n20638 = x99 & ~n4625 ;
  assign n20639 = n4943 & n20638 ;
  assign n20640 = n20637 | n20639 ;
  assign n20636 = x101 & n4631 ;
  assign n20642 = n4634 | n20636 ;
  assign n20643 = n20640 | n20642 ;
  assign n20641 = n20636 | n20640 ;
  assign n20644 = n20641 & n20643 ;
  assign n20645 = ( n6844 & n20643 ) | ( n6844 & n20644 ) | ( n20643 & n20644 ) ;
  assign n20646 = x32 & n20644 ;
  assign n20647 = x32 & n20643 ;
  assign n20648 = ( n6844 & n20646 ) | ( n6844 & n20647 ) | ( n20646 & n20647 ) ;
  assign n20649 = x32 & ~n20644 ;
  assign n20650 = x32 & ~n20643 ;
  assign n20651 = ( ~n6844 & n20649 ) | ( ~n6844 & n20650 ) | ( n20649 & n20650 ) ;
  assign n20652 = ( n20645 & ~n20648 ) | ( n20645 & n20651 ) | ( ~n20648 & n20651 ) ;
  assign n20653 = n20295 | n20315 ;
  assign n20654 = ( n20295 & n20298 ) | ( n20295 & n20653 ) | ( n20298 & n20653 ) ;
  assign n20655 = n20652 & n20654 ;
  assign n20656 = n20652 | n20654 ;
  assign n20657 = ~n20655 & n20656 ;
  assign n20901 = n20270 | n20290 ;
  assign n20902 = ( n20270 & n20273 ) | ( n20270 & n20901 ) | ( n20273 & n20901 ) ;
  assign n20658 = n20185 | n20207 ;
  assign n20659 = ( n20187 & n20207 ) | ( n20187 & n20658 ) | ( n20207 & n20658 ) ;
  assign n20660 = ( n20189 & n20190 ) | ( n20189 & n20659 ) | ( n20190 & n20659 ) ;
  assign n20661 = x70 & n17141 ;
  assign n20662 = x69 & ~n17140 ;
  assign n20663 = n17724 & n20662 ;
  assign n20664 = n20661 | n20663 ;
  assign n20665 = x71 & n17146 ;
  assign n20666 = n17149 | n20665 ;
  assign n20667 = n20664 | n20666 ;
  assign n20668 = x62 & ~n20667 ;
  assign n20669 = x62 & ~n20665 ;
  assign n20670 = ~n20664 & n20669 ;
  assign n20671 = ( ~n438 & n20668 ) | ( ~n438 & n20670 ) | ( n20668 & n20670 ) ;
  assign n20672 = ~x62 & n20667 ;
  assign n20673 = ~x62 & n20665 ;
  assign n20674 = ( ~x62 & n20664 ) | ( ~x62 & n20673 ) | ( n20664 & n20673 ) ;
  assign n20675 = ( n438 & n20672 ) | ( n438 & n20674 ) | ( n20672 & n20674 ) ;
  assign n20676 = n20671 | n20675 ;
  assign n20677 = x68 & n18290 ;
  assign n20678 = x63 & x67 ;
  assign n20679 = ~n18290 & n20678 ;
  assign n20680 = n20677 | n20679 ;
  assign n20681 = x2 & n20680 ;
  assign n20682 = n20680 & ~n20681 ;
  assign n20683 = x2 & ~n20680 ;
  assign n20684 = n20682 | n20683 ;
  assign n20685 = n20676 & n20684 ;
  assign n20686 = n20676 | n20684 ;
  assign n20687 = ~n20685 & n20686 ;
  assign n20688 = n20062 | n20064 ;
  assign n20689 = ( n20062 & n20079 ) | ( n20062 & n20688 ) | ( n20079 & n20688 ) ;
  assign n20690 = n20687 | n20689 ;
  assign n20691 = n20687 & n20689 ;
  assign n20692 = n20690 & ~n20691 ;
  assign n20693 = x74 & n15552 ;
  assign n20694 = x73 & n15547 ;
  assign n20695 = x72 & ~n15546 ;
  assign n20696 = n16123 & n20695 ;
  assign n20697 = n20694 | n20696 ;
  assign n20698 = n20693 | n20697 ;
  assign n20699 = n15555 | n20693 ;
  assign n20700 = n20697 | n20699 ;
  assign n20701 = ( n710 & n20698 ) | ( n710 & n20700 ) | ( n20698 & n20700 ) ;
  assign n20702 = x59 & n20700 ;
  assign n20703 = x59 & n20693 ;
  assign n20704 = ( x59 & n20697 ) | ( x59 & n20703 ) | ( n20697 & n20703 ) ;
  assign n20705 = ( n710 & n20702 ) | ( n710 & n20704 ) | ( n20702 & n20704 ) ;
  assign n20706 = x59 & ~n20704 ;
  assign n20707 = x59 & ~n20700 ;
  assign n20708 = ( ~n710 & n20706 ) | ( ~n710 & n20707 ) | ( n20706 & n20707 ) ;
  assign n20709 = ( n20701 & ~n20705 ) | ( n20701 & n20708 ) | ( ~n20705 & n20708 ) ;
  assign n20710 = ~n20692 & n20709 ;
  assign n20711 = n20689 | n20709 ;
  assign n20712 = ( n20687 & n20709 ) | ( n20687 & n20711 ) | ( n20709 & n20711 ) ;
  assign n20713 = n20690 & ~n20712 ;
  assign n20714 = n20710 | n20713 ;
  assign n20715 = n20086 | n20107 ;
  assign n20716 = n20085 | n20107 ;
  assign n20717 = ( n20057 & n20715 ) | ( n20057 & n20716 ) | ( n20715 & n20716 ) ;
  assign n20718 = ( n20087 & n20091 ) | ( n20087 & n20717 ) | ( n20091 & n20717 ) ;
  assign n20719 = n20714 | n20718 ;
  assign n20720 = n20714 & n20718 ;
  assign n20721 = n20719 & ~n20720 ;
  assign n20722 = x77 & n14045 ;
  assign n20723 = x76 & n14040 ;
  assign n20724 = x75 & ~n14039 ;
  assign n20725 = n14552 & n20724 ;
  assign n20726 = n20723 | n20725 ;
  assign n20727 = n20722 | n20726 ;
  assign n20728 = n14048 | n20722 ;
  assign n20729 = n20726 | n20728 ;
  assign n20730 = ( n1059 & n20727 ) | ( n1059 & n20729 ) | ( n20727 & n20729 ) ;
  assign n20731 = x56 & n20729 ;
  assign n20732 = x56 & n20722 ;
  assign n20733 = ( x56 & n20726 ) | ( x56 & n20732 ) | ( n20726 & n20732 ) ;
  assign n20734 = ( n1059 & n20731 ) | ( n1059 & n20733 ) | ( n20731 & n20733 ) ;
  assign n20735 = x56 & ~n20733 ;
  assign n20736 = x56 & ~n20729 ;
  assign n20737 = ( ~n1059 & n20735 ) | ( ~n1059 & n20736 ) | ( n20735 & n20736 ) ;
  assign n20738 = ( n20730 & ~n20734 ) | ( n20730 & n20737 ) | ( ~n20734 & n20737 ) ;
  assign n20739 = n20721 | n20738 ;
  assign n20740 = n20721 & n20738 ;
  assign n20741 = n20739 & ~n20740 ;
  assign n20742 = ( n19413 & n20110 ) | ( n19413 & n20132 ) | ( n20110 & n20132 ) ;
  assign n20743 = n20110 | n20132 ;
  assign n20744 = ( n19437 & n20742 ) | ( n19437 & n20743 ) | ( n20742 & n20743 ) ;
  assign n20745 = n20741 | n20744 ;
  assign n20746 = n20741 & n20744 ;
  assign n20747 = n20745 & ~n20746 ;
  assign n20748 = x80 & n12574 ;
  assign n20749 = x79 & n12569 ;
  assign n20750 = x78 & ~n12568 ;
  assign n20751 = n13076 & n20750 ;
  assign n20752 = n20749 | n20751 ;
  assign n20753 = n20748 | n20752 ;
  assign n20754 = n12577 | n20748 ;
  assign n20755 = n20752 | n20754 ;
  assign n20756 = ( n1499 & n20753 ) | ( n1499 & n20755 ) | ( n20753 & n20755 ) ;
  assign n20757 = x53 & n20755 ;
  assign n20758 = x53 & n20748 ;
  assign n20759 = ( x53 & n20752 ) | ( x53 & n20758 ) | ( n20752 & n20758 ) ;
  assign n20760 = ( n1499 & n20757 ) | ( n1499 & n20759 ) | ( n20757 & n20759 ) ;
  assign n20761 = x53 & ~n20759 ;
  assign n20762 = x53 & ~n20755 ;
  assign n20763 = ( ~n1499 & n20761 ) | ( ~n1499 & n20762 ) | ( n20761 & n20762 ) ;
  assign n20764 = ( n20756 & ~n20760 ) | ( n20756 & n20763 ) | ( ~n20760 & n20763 ) ;
  assign n20765 = n20747 & ~n20764 ;
  assign n20766 = n20747 | n20764 ;
  assign n20767 = ( ~n20747 & n20765 ) | ( ~n20747 & n20766 ) | ( n20765 & n20766 ) ;
  assign n20768 = n20137 | n20157 ;
  assign n20769 = ( n20137 & n20140 ) | ( n20137 & n20768 ) | ( n20140 & n20768 ) ;
  assign n20770 = n20767 | n20769 ;
  assign n20771 = n20767 & n20769 ;
  assign n20772 = n20770 & ~n20771 ;
  assign n20773 = x83 & n11205 ;
  assign n20774 = x82 & n11200 ;
  assign n20775 = x81 & ~n11199 ;
  assign n20776 = n11679 & n20775 ;
  assign n20777 = n20774 | n20776 ;
  assign n20778 = n20773 | n20777 ;
  assign n20779 = n11208 | n20773 ;
  assign n20780 = n20777 | n20779 ;
  assign n20781 = ( n2009 & n20778 ) | ( n2009 & n20780 ) | ( n20778 & n20780 ) ;
  assign n20782 = x50 & n20780 ;
  assign n20783 = x50 & n20773 ;
  assign n20784 = ( x50 & n20777 ) | ( x50 & n20783 ) | ( n20777 & n20783 ) ;
  assign n20785 = ( n2009 & n20782 ) | ( n2009 & n20784 ) | ( n20782 & n20784 ) ;
  assign n20786 = x50 & ~n20784 ;
  assign n20787 = x50 & ~n20780 ;
  assign n20788 = ( ~n2009 & n20786 ) | ( ~n2009 & n20787 ) | ( n20786 & n20787 ) ;
  assign n20789 = ( n20781 & ~n20785 ) | ( n20781 & n20788 ) | ( ~n20785 & n20788 ) ;
  assign n20790 = ~n20772 & n20789 ;
  assign n20791 = n20767 | n20789 ;
  assign n20792 = ( n20769 & n20789 ) | ( n20769 & n20791 ) | ( n20789 & n20791 ) ;
  assign n20793 = n20770 & ~n20792 ;
  assign n20794 = n20790 | n20793 ;
  assign n20795 = ( n20163 & n20164 ) | ( n20163 & n20183 ) | ( n20164 & n20183 ) ;
  assign n20796 = n20794 | n20795 ;
  assign n20797 = n20794 & n20795 ;
  assign n20798 = n20796 & ~n20797 ;
  assign n20799 = x86 & n9933 ;
  assign n20800 = x85 & n9928 ;
  assign n20801 = x84 & ~n9927 ;
  assign n20802 = n10379 & n20801 ;
  assign n20803 = n20800 | n20802 ;
  assign n20804 = n20799 | n20803 ;
  assign n20805 = n9936 | n20799 ;
  assign n20806 = n20803 | n20805 ;
  assign n20807 = ( n2606 & n20804 ) | ( n2606 & n20806 ) | ( n20804 & n20806 ) ;
  assign n20808 = x47 & n20806 ;
  assign n20809 = x47 & n20799 ;
  assign n20810 = ( x47 & n20803 ) | ( x47 & n20809 ) | ( n20803 & n20809 ) ;
  assign n20811 = ( n2606 & n20808 ) | ( n2606 & n20810 ) | ( n20808 & n20810 ) ;
  assign n20812 = x47 & ~n20810 ;
  assign n20813 = x47 & ~n20806 ;
  assign n20814 = ( ~n2606 & n20812 ) | ( ~n2606 & n20813 ) | ( n20812 & n20813 ) ;
  assign n20815 = ( n20807 & ~n20811 ) | ( n20807 & n20814 ) | ( ~n20811 & n20814 ) ;
  assign n20816 = ~n20798 & n20815 ;
  assign n20817 = n20797 | n20815 ;
  assign n20818 = n20796 & ~n20817 ;
  assign n20819 = n20816 | n20818 ;
  assign n20820 = n20659 & n20819 ;
  assign n20821 = n20189 & n20819 ;
  assign n20822 = ( n20190 & n20820 ) | ( n20190 & n20821 ) | ( n20820 & n20821 ) ;
  assign n20823 = n20660 & ~n20822 ;
  assign n20824 = x89 & n8724 ;
  assign n20825 = x88 & n8719 ;
  assign n20826 = x87 & ~n8718 ;
  assign n20827 = n9149 & n20826 ;
  assign n20828 = n20825 | n20827 ;
  assign n20829 = n20824 | n20828 ;
  assign n20830 = n8727 | n20824 ;
  assign n20831 = n20828 | n20830 ;
  assign n20832 = ( n3282 & n20829 ) | ( n3282 & n20831 ) | ( n20829 & n20831 ) ;
  assign n20833 = x44 & n20831 ;
  assign n20834 = x44 & n20824 ;
  assign n20835 = ( x44 & n20828 ) | ( x44 & n20834 ) | ( n20828 & n20834 ) ;
  assign n20836 = ( n3282 & n20833 ) | ( n3282 & n20835 ) | ( n20833 & n20835 ) ;
  assign n20837 = x44 & ~n20835 ;
  assign n20838 = x44 & ~n20831 ;
  assign n20839 = ( ~n3282 & n20837 ) | ( ~n3282 & n20838 ) | ( n20837 & n20838 ) ;
  assign n20840 = ( n20832 & ~n20836 ) | ( n20832 & n20839 ) | ( ~n20836 & n20839 ) ;
  assign n20841 = ~n20659 & n20819 ;
  assign n20842 = ~n20189 & n20819 ;
  assign n20843 = ( ~n20190 & n20841 ) | ( ~n20190 & n20842 ) | ( n20841 & n20842 ) ;
  assign n20844 = n20840 & ~n20843 ;
  assign n20845 = ~n20823 & n20844 ;
  assign n20846 = ~n20840 & n20843 ;
  assign n20847 = ( n20823 & ~n20840 ) | ( n20823 & n20846 ) | ( ~n20840 & n20846 ) ;
  assign n20848 = n20845 | n20847 ;
  assign n20849 = n20213 | n20239 ;
  assign n20850 = ( n20210 & n20239 ) | ( n20210 & n20849 ) | ( n20239 & n20849 ) ;
  assign n20851 = ( n20214 & n20216 ) | ( n20214 & n20850 ) | ( n20216 & n20850 ) ;
  assign n20852 = n20848 | n20851 ;
  assign n20853 = n20848 & n20851 ;
  assign n20854 = n20852 & ~n20853 ;
  assign n20855 = x92 & n7566 ;
  assign n20856 = x91 & n7561 ;
  assign n20857 = x90 & ~n7560 ;
  assign n20858 = n7953 & n20857 ;
  assign n20859 = n20856 | n20858 ;
  assign n20860 = n20855 | n20859 ;
  assign n20861 = n7569 | n20855 ;
  assign n20862 = n20859 | n20861 ;
  assign n20863 = ( n4040 & n20860 ) | ( n4040 & n20862 ) | ( n20860 & n20862 ) ;
  assign n20864 = x41 & n20862 ;
  assign n20865 = x41 & n20855 ;
  assign n20866 = ( x41 & n20859 ) | ( x41 & n20865 ) | ( n20859 & n20865 ) ;
  assign n20867 = ( n4040 & n20864 ) | ( n4040 & n20866 ) | ( n20864 & n20866 ) ;
  assign n20868 = x41 & ~n20866 ;
  assign n20869 = x41 & ~n20862 ;
  assign n20870 = ( ~n4040 & n20868 ) | ( ~n4040 & n20869 ) | ( n20868 & n20869 ) ;
  assign n20871 = ( n20863 & ~n20867 ) | ( n20863 & n20870 ) | ( ~n20867 & n20870 ) ;
  assign n20872 = ~n20854 & n20871 ;
  assign n20873 = n20848 | n20871 ;
  assign n20874 = ( n20851 & n20871 ) | ( n20851 & n20873 ) | ( n20871 & n20873 ) ;
  assign n20875 = n20852 & ~n20874 ;
  assign n20876 = n20872 | n20875 ;
  assign n20877 = ( n20244 & n20247 ) | ( n20244 & n20266 ) | ( n20247 & n20266 ) ;
  assign n20878 = n20876 | n20877 ;
  assign n20879 = n20876 & n20877 ;
  assign n20880 = n20878 & ~n20879 ;
  assign n20881 = x95 & n6536 ;
  assign n20882 = x94 & n6531 ;
  assign n20883 = x93 & ~n6530 ;
  assign n20884 = n6871 & n20883 ;
  assign n20885 = n20882 | n20884 ;
  assign n20886 = n20881 | n20885 ;
  assign n20887 = n6539 | n20881 ;
  assign n20888 = n20885 | n20887 ;
  assign n20889 = ( n4897 & n20886 ) | ( n4897 & n20888 ) | ( n20886 & n20888 ) ;
  assign n20890 = x38 & n20888 ;
  assign n20891 = x38 & n20881 ;
  assign n20892 = ( x38 & n20885 ) | ( x38 & n20891 ) | ( n20885 & n20891 ) ;
  assign n20893 = ( n4897 & n20890 ) | ( n4897 & n20892 ) | ( n20890 & n20892 ) ;
  assign n20894 = x38 & ~n20892 ;
  assign n20895 = x38 & ~n20888 ;
  assign n20896 = ( ~n4897 & n20894 ) | ( ~n4897 & n20895 ) | ( n20894 & n20895 ) ;
  assign n20897 = ( n20889 & ~n20893 ) | ( n20889 & n20896 ) | ( ~n20893 & n20896 ) ;
  assign n20898 = n20880 | n20897 ;
  assign n20899 = n20880 & n20897 ;
  assign n20900 = n20898 & ~n20899 ;
  assign n20903 = n20900 & n20902 ;
  assign n20904 = n20902 & ~n20903 ;
  assign n20905 = x98 & n5554 ;
  assign n20906 = x97 & n5549 ;
  assign n20907 = x96 & ~n5548 ;
  assign n20908 = n5893 & n20907 ;
  assign n20909 = n20906 | n20908 ;
  assign n20910 = n20905 | n20909 ;
  assign n20911 = n5557 | n20905 ;
  assign n20912 = n20909 | n20911 ;
  assign n20913 = ( ~n5850 & n20910 ) | ( ~n5850 & n20912 ) | ( n20910 & n20912 ) ;
  assign n20914 = n20910 & n20912 ;
  assign n20915 = ( n5834 & n20913 ) | ( n5834 & n20914 ) | ( n20913 & n20914 ) ;
  assign n20916 = x35 & n20912 ;
  assign n20917 = x35 & n20905 ;
  assign n20918 = ( x35 & n20909 ) | ( x35 & n20917 ) | ( n20909 & n20917 ) ;
  assign n20919 = ( ~n5850 & n20916 ) | ( ~n5850 & n20918 ) | ( n20916 & n20918 ) ;
  assign n20920 = n20916 & n20918 ;
  assign n20921 = ( n5834 & n20919 ) | ( n5834 & n20920 ) | ( n20919 & n20920 ) ;
  assign n20922 = x35 & ~n20918 ;
  assign n20923 = x35 & ~n20912 ;
  assign n20924 = ( n5850 & n20922 ) | ( n5850 & n20923 ) | ( n20922 & n20923 ) ;
  assign n20925 = n20922 | n20923 ;
  assign n20926 = ( ~n5834 & n20924 ) | ( ~n5834 & n20925 ) | ( n20924 & n20925 ) ;
  assign n20927 = ( n20915 & ~n20921 ) | ( n20915 & n20926 ) | ( ~n20921 & n20926 ) ;
  assign n20928 = ~n20900 & n20927 ;
  assign n20929 = ( n20902 & n20927 ) | ( n20902 & n20928 ) | ( n20927 & n20928 ) ;
  assign n20930 = ~n20904 & n20929 ;
  assign n20931 = n20900 & ~n20927 ;
  assign n20932 = ~n20902 & n20931 ;
  assign n20933 = ( n20904 & ~n20927 ) | ( n20904 & n20932 ) | ( ~n20927 & n20932 ) ;
  assign n20934 = n20930 | n20933 ;
  assign n20935 = n20657 | n20934 ;
  assign n20936 = n20657 & n20934 ;
  assign n20937 = n20935 & ~n20936 ;
  assign n20938 = n20053 | n20324 ;
  assign n20940 = x103 & n3811 ;
  assign n20941 = x102 & ~n3810 ;
  assign n20942 = n4067 & n20941 ;
  assign n20943 = n20940 | n20942 ;
  assign n20939 = x104 & n3816 ;
  assign n20945 = n3819 | n20939 ;
  assign n20946 = n20943 | n20945 ;
  assign n20944 = n20939 | n20943 ;
  assign n20947 = n20944 & n20946 ;
  assign n20948 = ( n7911 & n20946 ) | ( n7911 & n20947 ) | ( n20946 & n20947 ) ;
  assign n20949 = x29 & n20947 ;
  assign n20950 = x29 & n20946 ;
  assign n20951 = ( n7911 & n20949 ) | ( n7911 & n20950 ) | ( n20949 & n20950 ) ;
  assign n20952 = x29 & ~n20947 ;
  assign n20953 = x29 & ~n20946 ;
  assign n20954 = ( ~n7911 & n20952 ) | ( ~n7911 & n20953 ) | ( n20952 & n20953 ) ;
  assign n20955 = ( n20948 & ~n20951 ) | ( n20948 & n20954 ) | ( ~n20951 & n20954 ) ;
  assign n20956 = n20053 & n20955 ;
  assign n20957 = ( n20324 & n20955 ) | ( n20324 & n20956 ) | ( n20955 & n20956 ) ;
  assign n20958 = n20938 & ~n20957 ;
  assign n20959 = ~n20053 & n20955 ;
  assign n20960 = ~n20324 & n20959 ;
  assign n20961 = n20937 & n20960 ;
  assign n20962 = ( n20937 & n20958 ) | ( n20937 & n20961 ) | ( n20958 & n20961 ) ;
  assign n20963 = n20937 | n20960 ;
  assign n20964 = n20958 | n20963 ;
  assign n20965 = ~n20962 & n20964 ;
  assign n20966 = ~n20635 & n20965 ;
  assign n20967 = n20630 | n20965 ;
  assign n20968 = ( n20632 & n20965 ) | ( n20632 & n20967 ) | ( n20965 & n20967 ) ;
  assign n20969 = n20633 & ~n20968 ;
  assign n20970 = n20966 | n20969 ;
  assign n20971 = x110 & n2429 ;
  assign n20972 = x109 & n2424 ;
  assign n20973 = x108 & ~n2423 ;
  assign n20974 = n2631 & n20973 ;
  assign n20975 = n20972 | n20974 ;
  assign n20976 = n20971 | n20975 ;
  assign n20977 = n2432 | n20971 ;
  assign n20978 = n20975 | n20977 ;
  assign n20979 = ( n10330 & n20976 ) | ( n10330 & n20978 ) | ( n20976 & n20978 ) ;
  assign n20980 = x23 & n20978 ;
  assign n20981 = x23 & n20971 ;
  assign n20982 = ( x23 & n20975 ) | ( x23 & n20981 ) | ( n20975 & n20981 ) ;
  assign n20983 = ( n10330 & n20980 ) | ( n10330 & n20982 ) | ( n20980 & n20982 ) ;
  assign n20984 = x23 & ~n20982 ;
  assign n20985 = x23 & ~n20978 ;
  assign n20986 = ( ~n10330 & n20984 ) | ( ~n10330 & n20985 ) | ( n20984 & n20985 ) ;
  assign n20987 = ( n20979 & ~n20983 ) | ( n20979 & n20986 ) | ( ~n20983 & n20986 ) ;
  assign n20988 = n20330 | n20356 ;
  assign n20989 = ( n20356 & n20357 ) | ( n20356 & n20988 ) | ( n20357 & n20988 ) ;
  assign n20990 = ( n20970 & n20987 ) | ( n20970 & ~n20989 ) | ( n20987 & ~n20989 ) ;
  assign n20991 = ( ~n20987 & n20989 ) | ( ~n20987 & n20990 ) | ( n20989 & n20990 ) ;
  assign n20992 = ( ~n20970 & n20990 ) | ( ~n20970 & n20991 ) | ( n20990 & n20991 ) ;
  assign n20993 = ~n20613 & n20992 ;
  assign n20994 = n20612 | n20992 ;
  assign n20995 = n20607 & ~n20994 ;
  assign n20996 = n20993 | n20995 ;
  assign n20997 = x116 & n1383 ;
  assign n20998 = x115 & n1378 ;
  assign n20999 = x114 & ~n1377 ;
  assign n21000 = n1542 & n20999 ;
  assign n21001 = n20998 | n21000 ;
  assign n21002 = n20997 | n21001 ;
  assign n21003 = n1386 | n20997 ;
  assign n21004 = n21001 | n21003 ;
  assign n21005 = ( ~n13040 & n21002 ) | ( ~n13040 & n21004 ) | ( n21002 & n21004 ) ;
  assign n21006 = n21002 & n21004 ;
  assign n21007 = ( n13022 & n21005 ) | ( n13022 & n21006 ) | ( n21005 & n21006 ) ;
  assign n21008 = x17 & n21007 ;
  assign n21009 = x17 & ~n21007 ;
  assign n21010 = ( n21007 & ~n21008 ) | ( n21007 & n21009 ) | ( ~n21008 & n21009 ) ;
  assign n21011 = n20386 | n20439 ;
  assign n21012 = ( n20439 & n20440 ) | ( n20439 & n21011 ) | ( n20440 & n21011 ) ;
  assign n21013 = ( n20996 & n21010 ) | ( n20996 & ~n21012 ) | ( n21010 & ~n21012 ) ;
  assign n21014 = ( ~n21010 & n21012 ) | ( ~n21010 & n21013 ) | ( n21012 & n21013 ) ;
  assign n21015 = ( ~n20996 & n21013 ) | ( ~n20996 & n21014 ) | ( n21013 & n21014 ) ;
  assign n21016 = ~n20577 & n21015 ;
  assign n21017 = n20569 | n21013 ;
  assign n21018 = ~n20569 & n20996 ;
  assign n21019 = ( n21014 & n21017 ) | ( n21014 & ~n21018 ) | ( n21017 & ~n21018 ) ;
  assign n21020 = ( n20574 & n21015 ) | ( n20574 & n21019 ) | ( n21015 & n21019 ) ;
  assign n21021 = n20575 & ~n21020 ;
  assign n21022 = n21016 | n21021 ;
  assign n21023 = n20000 | n20448 ;
  assign n21025 = x121 & n631 ;
  assign n21026 = x120 & ~n630 ;
  assign n21027 = n764 & n21026 ;
  assign n21028 = n21025 | n21027 ;
  assign n21024 = x122 & n636 ;
  assign n21030 = n639 | n21024 ;
  assign n21031 = n21028 | n21030 ;
  assign n21029 = n21024 | n21028 ;
  assign n21032 = n21029 & n21031 ;
  assign n21033 = ( n16043 & n21031 ) | ( n16043 & n21032 ) | ( n21031 & n21032 ) ;
  assign n21034 = x11 & n21032 ;
  assign n21035 = x11 & n21031 ;
  assign n21036 = ( n16043 & n21034 ) | ( n16043 & n21035 ) | ( n21034 & n21035 ) ;
  assign n21037 = x11 & ~n21032 ;
  assign n21038 = x11 & ~n21031 ;
  assign n21039 = ( ~n16043 & n21037 ) | ( ~n16043 & n21038 ) | ( n21037 & n21038 ) ;
  assign n21040 = ( n21033 & ~n21036 ) | ( n21033 & n21039 ) | ( ~n21036 & n21039 ) ;
  assign n21041 = n19996 & n21040 ;
  assign n21042 = n19776 & n21041 ;
  assign n21043 = ( n19777 & n21041 ) | ( n19777 & n21042 ) | ( n21041 & n21042 ) ;
  assign n21044 = n21041 & n21042 ;
  assign n21045 = ( n19779 & n21043 ) | ( n19779 & n21044 ) | ( n21043 & n21044 ) ;
  assign n21046 = ( n20448 & n21040 ) | ( n20448 & n21045 ) | ( n21040 & n21045 ) ;
  assign n21047 = n21023 & ~n21046 ;
  assign n21048 = n21040 & ~n21045 ;
  assign n21049 = n21022 & n21048 ;
  assign n21050 = ~n20448 & n21049 ;
  assign n21051 = ( n21022 & n21047 ) | ( n21022 & n21050 ) | ( n21047 & n21050 ) ;
  assign n21052 = n21022 | n21048 ;
  assign n21053 = ( ~n20448 & n21022 ) | ( ~n20448 & n21052 ) | ( n21022 & n21052 ) ;
  assign n21054 = n21047 | n21053 ;
  assign n21055 = ~n21051 & n21054 ;
  assign n21056 = n20548 & n21055 ;
  assign n21057 = ~n20550 & n21056 ;
  assign n21058 = ( n20552 & n21055 ) | ( n20552 & n21057 ) | ( n21055 & n21057 ) ;
  assign n21059 = n20548 | n21055 ;
  assign n21060 = ( ~n20550 & n21055 ) | ( ~n20550 & n21059 ) | ( n21055 & n21059 ) ;
  assign n21061 = n20552 | n21060 ;
  assign n21062 = ~n21058 & n21061 ;
  assign n21063 = n20531 | n21062 ;
  assign n21064 = n20526 | n21063 ;
  assign n21065 = n20531 & n21062 ;
  assign n21066 = ( n20526 & n21062 ) | ( n20526 & n21065 ) | ( n21062 & n21065 ) ;
  assign n21067 = n21064 & ~n21066 ;
  assign n21068 = ~n20504 & n21067 ;
  assign n21069 = n20497 | n20502 ;
  assign n21070 = ( n20504 & ~n21067 ) | ( n20504 & n21069 ) | ( ~n21067 & n21069 ) ;
  assign n21071 = n20504 & n21067 ;
  assign n21072 = n20504 & ~n21071 ;
  assign n21073 = n21068 | n21072 ;
  assign n21074 = n20497 & n21068 ;
  assign n21075 = ( n20497 & n21072 ) | ( n20497 & n21074 ) | ( n21072 & n21074 ) ;
  assign n21076 = ( n20501 & n21073 ) | ( n20501 & n21075 ) | ( n21073 & n21075 ) ;
  assign n21077 = ( n20498 & n21073 ) | ( n20498 & n21075 ) | ( n21073 & n21075 ) ;
  assign n21078 = ( n19932 & n21076 ) | ( n19932 & n21077 ) | ( n21076 & n21077 ) ;
  assign n21079 = ( n21068 & n21070 ) | ( n21068 & ~n21078 ) | ( n21070 & ~n21078 ) ;
  assign n21080 = n20525 | n21066 ;
  assign n21081 = n20551 | n21057 ;
  assign n21082 = n20551 | n21055 ;
  assign n21083 = ( n20552 & n21081 ) | ( n20552 & n21082 ) | ( n21081 & n21082 ) ;
  assign n21084 = x127 & ~n206 ;
  assign n21085 = n267 & n21084 ;
  assign n21086 = n215 & n19877 ;
  assign n21087 = n21085 | n21086 ;
  assign n21088 = n215 & n19880 ;
  assign n21089 = n21085 | n21088 ;
  assign n21090 = ( n18202 & n21087 ) | ( n18202 & n21089 ) | ( n21087 & n21089 ) ;
  assign n21091 = n21087 & n21089 ;
  assign n21092 = ( n18212 & n21090 ) | ( n18212 & n21091 ) | ( n21090 & n21091 ) ;
  assign n21093 = ( n18214 & n21090 ) | ( n18214 & n21091 ) | ( n21090 & n21091 ) ;
  assign n21094 = ( n14002 & n21092 ) | ( n14002 & n21093 ) | ( n21092 & n21093 ) ;
  assign n21095 = x5 & n21092 ;
  assign n21096 = x5 & n21093 ;
  assign n21097 = ( n14002 & n21095 ) | ( n14002 & n21096 ) | ( n21095 & n21096 ) ;
  assign n21098 = x5 & ~n21096 ;
  assign n21099 = x5 & ~n21095 ;
  assign n21100 = ( ~n14002 & n21098 ) | ( ~n14002 & n21099 ) | ( n21098 & n21099 ) ;
  assign n21101 = ( n21094 & ~n21097 ) | ( n21094 & n21100 ) | ( ~n21097 & n21100 ) ;
  assign n21102 = n20548 & n21101 ;
  assign n21103 = n20550 & n21102 ;
  assign n21104 = ( n21057 & n21101 ) | ( n21057 & n21103 ) | ( n21101 & n21103 ) ;
  assign n21105 = ( n21055 & n21101 ) | ( n21055 & n21103 ) | ( n21101 & n21103 ) ;
  assign n21106 = ( n20552 & n21104 ) | ( n20552 & n21105 ) | ( n21104 & n21105 ) ;
  assign n21107 = n21083 & ~n21106 ;
  assign n21108 = n21046 | n21050 ;
  assign n21109 = n21022 | n21046 ;
  assign n21110 = ( n21047 & n21108 ) | ( n21047 & n21109 ) | ( n21108 & n21109 ) ;
  assign n21112 = x125 & n384 ;
  assign n21113 = x124 & ~n383 ;
  assign n21114 = n463 & n21113 ;
  assign n21115 = n21112 | n21114 ;
  assign n21111 = x126 & n389 ;
  assign n21117 = n392 | n21111 ;
  assign n21118 = n21115 | n21117 ;
  assign n21116 = n21111 | n21115 ;
  assign n21119 = n21116 & n21118 ;
  assign n21120 = ( n18220 & n21118 ) | ( n18220 & n21119 ) | ( n21118 & n21119 ) ;
  assign n21121 = x8 & n21119 ;
  assign n21122 = x8 & n21118 ;
  assign n21123 = ( n18220 & n21121 ) | ( n18220 & n21122 ) | ( n21121 & n21122 ) ;
  assign n21124 = x8 & ~n21119 ;
  assign n21125 = x8 & ~n21118 ;
  assign n21126 = ( ~n18220 & n21124 ) | ( ~n18220 & n21125 ) | ( n21124 & n21125 ) ;
  assign n21127 = ( n21120 & ~n21123 ) | ( n21120 & n21126 ) | ( ~n21123 & n21126 ) ;
  assign n21128 = n21045 & n21127 ;
  assign n21129 = n21040 & n21127 ;
  assign n21130 = ( n20448 & n21128 ) | ( n20448 & n21129 ) | ( n21128 & n21129 ) ;
  assign n21131 = ( n21050 & n21127 ) | ( n21050 & n21130 ) | ( n21127 & n21130 ) ;
  assign n21132 = ( n21022 & n21127 ) | ( n21022 & n21130 ) | ( n21127 & n21130 ) ;
  assign n21133 = ( n21047 & n21131 ) | ( n21047 & n21132 ) | ( n21131 & n21132 ) ;
  assign n21134 = n21110 & ~n21133 ;
  assign n21135 = x123 & n636 ;
  assign n21136 = x122 & n631 ;
  assign n21137 = x121 & ~n630 ;
  assign n21138 = n764 & n21137 ;
  assign n21139 = n21136 | n21138 ;
  assign n21140 = n21135 | n21139 ;
  assign n21141 = n639 | n21135 ;
  assign n21142 = n21139 | n21141 ;
  assign n21143 = ( n16086 & n21140 ) | ( n16086 & n21142 ) | ( n21140 & n21142 ) ;
  assign n21144 = x11 & n21142 ;
  assign n21145 = x11 & n21135 ;
  assign n21146 = ( x11 & n21139 ) | ( x11 & n21145 ) | ( n21139 & n21145 ) ;
  assign n21147 = ( n16086 & n21144 ) | ( n16086 & n21146 ) | ( n21144 & n21146 ) ;
  assign n21148 = x11 & ~n21146 ;
  assign n21149 = x11 & ~n21142 ;
  assign n21150 = ( ~n16086 & n21148 ) | ( ~n16086 & n21149 ) | ( n21148 & n21149 ) ;
  assign n21151 = ( n21143 & ~n21147 ) | ( n21143 & n21150 ) | ( ~n21147 & n21150 ) ;
  assign n21152 = n21020 | n21151 ;
  assign n21153 = n20576 | n21151 ;
  assign n21154 = ( n20577 & n21152 ) | ( n20577 & n21153 ) | ( n21152 & n21153 ) ;
  assign n21155 = n21020 & n21151 ;
  assign n21156 = n20576 & n21151 ;
  assign n21157 = ( n20577 & n21155 ) | ( n20577 & n21156 ) | ( n21155 & n21156 ) ;
  assign n21158 = n21154 & ~n21157 ;
  assign n21159 = x120 & n962 ;
  assign n21160 = x119 & n957 ;
  assign n21161 = x118 & ~n956 ;
  assign n21162 = n1105 & n21161 ;
  assign n21163 = n21160 | n21162 ;
  assign n21164 = n21159 | n21163 ;
  assign n21165 = n965 | n21159 ;
  assign n21166 = n21163 | n21165 ;
  assign n21167 = ( n14991 & n21164 ) | ( n14991 & n21166 ) | ( n21164 & n21166 ) ;
  assign n21168 = x14 & n21166 ;
  assign n21169 = x14 & n21159 ;
  assign n21170 = ( x14 & n21163 ) | ( x14 & n21169 ) | ( n21163 & n21169 ) ;
  assign n21171 = ( n14991 & n21168 ) | ( n14991 & n21170 ) | ( n21168 & n21170 ) ;
  assign n21172 = x14 & ~n21170 ;
  assign n21173 = x14 & ~n21166 ;
  assign n21174 = ( ~n14991 & n21172 ) | ( ~n14991 & n21173 ) | ( n21172 & n21173 ) ;
  assign n21175 = ( n21167 & ~n21171 ) | ( n21167 & n21174 ) | ( ~n21171 & n21174 ) ;
  assign n21177 = x116 & n1378 ;
  assign n21178 = x115 & ~n1377 ;
  assign n21179 = n1542 & n21178 ;
  assign n21180 = n21177 | n21179 ;
  assign n21176 = x117 & n1383 ;
  assign n21182 = n1386 | n21176 ;
  assign n21183 = n21180 | n21182 ;
  assign n21181 = n21176 | n21180 ;
  assign n21184 = n21181 & n21183 ;
  assign n21185 = ( ~n13522 & n21183 ) | ( ~n13522 & n21184 ) | ( n21183 & n21184 ) ;
  assign n21186 = n21183 & n21184 ;
  assign n21187 = ( n13503 & n21185 ) | ( n13503 & n21186 ) | ( n21185 & n21186 ) ;
  assign n21188 = x17 & n21187 ;
  assign n21189 = x17 & ~n21187 ;
  assign n21190 = ( n21187 & ~n21188 ) | ( n21187 & n21189 ) | ( ~n21188 & n21189 ) ;
  assign n21191 = ( n20612 & n20613 ) | ( n20612 & n20994 ) | ( n20613 & n20994 ) ;
  assign n21192 = n21190 & n21191 ;
  assign n21193 = n21190 | n21191 ;
  assign n21194 = ~n21192 & n21193 ;
  assign n21195 = x114 & n1859 ;
  assign n21196 = x113 & n1854 ;
  assign n21197 = x112 & ~n1853 ;
  assign n21198 = n2037 & n21197 ;
  assign n21199 = n21196 | n21198 ;
  assign n21200 = n21195 | n21199 ;
  assign n21201 = n1862 | n21195 ;
  assign n21202 = n21199 | n21201 ;
  assign n21203 = ( ~n12095 & n21200 ) | ( ~n12095 & n21202 ) | ( n21200 & n21202 ) ;
  assign n21204 = n21200 & n21202 ;
  assign n21205 = ( n12079 & n21203 ) | ( n12079 & n21204 ) | ( n21203 & n21204 ) ;
  assign n21206 = x20 & n21205 ;
  assign n21207 = x20 & ~n21205 ;
  assign n21208 = ( n21205 & ~n21206 ) | ( n21205 & n21207 ) | ( ~n21206 & n21207 ) ;
  assign n21209 = x111 & n2429 ;
  assign n21210 = x110 & n2424 ;
  assign n21211 = x109 & ~n2423 ;
  assign n21212 = n2631 & n21211 ;
  assign n21213 = n21210 | n21212 ;
  assign n21214 = n21209 | n21213 ;
  assign n21215 = n2432 | n21209 ;
  assign n21216 = n21213 | n21215 ;
  assign n21217 = ( n10749 & n21214 ) | ( n10749 & n21216 ) | ( n21214 & n21216 ) ;
  assign n21218 = x23 & n21216 ;
  assign n21219 = x23 & n21209 ;
  assign n21220 = ( x23 & n21213 ) | ( x23 & n21219 ) | ( n21213 & n21219 ) ;
  assign n21221 = ( n10749 & n21218 ) | ( n10749 & n21220 ) | ( n21218 & n21220 ) ;
  assign n21222 = x23 & ~n21220 ;
  assign n21223 = x23 & ~n21216 ;
  assign n21224 = ( ~n10749 & n21222 ) | ( ~n10749 & n21223 ) | ( n21222 & n21223 ) ;
  assign n21225 = ( n21217 & ~n21221 ) | ( n21217 & n21224 ) | ( ~n21221 & n21224 ) ;
  assign n21226 = n20968 | n21225 ;
  assign n21227 = n20634 | n21225 ;
  assign n21228 = ( n20635 & n21226 ) | ( n20635 & n21227 ) | ( n21226 & n21227 ) ;
  assign n21229 = n20968 & n21225 ;
  assign n21230 = n20634 & n21225 ;
  assign n21231 = ( n20635 & n21229 ) | ( n20635 & n21230 ) | ( n21229 & n21230 ) ;
  assign n21232 = n21228 & ~n21231 ;
  assign n21233 = x105 & n3816 ;
  assign n21234 = x104 & n3811 ;
  assign n21235 = x103 & ~n3810 ;
  assign n21236 = n4067 & n21235 ;
  assign n21237 = n21234 | n21236 ;
  assign n21238 = n21233 | n21237 ;
  assign n21239 = n3819 | n21233 ;
  assign n21240 = n21237 | n21239 ;
  assign n21241 = ( n8273 & n21238 ) | ( n8273 & n21240 ) | ( n21238 & n21240 ) ;
  assign n21242 = x29 & n21240 ;
  assign n21243 = x29 & n21233 ;
  assign n21244 = ( x29 & n21237 ) | ( x29 & n21243 ) | ( n21237 & n21243 ) ;
  assign n21245 = ( n8273 & n21242 ) | ( n8273 & n21244 ) | ( n21242 & n21244 ) ;
  assign n21246 = x29 & ~n21244 ;
  assign n21247 = x29 & ~n21240 ;
  assign n21248 = ( ~n8273 & n21246 ) | ( ~n8273 & n21247 ) | ( n21246 & n21247 ) ;
  assign n21249 = ( n21241 & ~n21245 ) | ( n21241 & n21248 ) | ( ~n21245 & n21248 ) ;
  assign n21250 = n20652 | n20934 ;
  assign n21251 = ( n20654 & n20934 ) | ( n20654 & n21250 ) | ( n20934 & n21250 ) ;
  assign n21252 = n21249 | n21251 ;
  assign n21253 = n20655 | n21249 ;
  assign n21254 = ( n20657 & n21252 ) | ( n20657 & n21253 ) | ( n21252 & n21253 ) ;
  assign n21255 = n21249 & n21251 ;
  assign n21256 = n20655 & n21249 ;
  assign n21257 = ( n20657 & n21255 ) | ( n20657 & n21256 ) | ( n21255 & n21256 ) ;
  assign n21258 = n21254 & ~n21257 ;
  assign n21260 = x101 & n4626 ;
  assign n21261 = x100 & ~n4625 ;
  assign n21262 = n4943 & n21261 ;
  assign n21263 = n21260 | n21262 ;
  assign n21259 = x102 & n4631 ;
  assign n21265 = n4634 | n21259 ;
  assign n21266 = n21263 | n21265 ;
  assign n21264 = n21259 | n21263 ;
  assign n21267 = n21264 & n21266 ;
  assign n21268 = ( n7178 & n21266 ) | ( n7178 & n21267 ) | ( n21266 & n21267 ) ;
  assign n21269 = x32 & n21267 ;
  assign n21270 = x32 & n21266 ;
  assign n21271 = ( n7178 & n21269 ) | ( n7178 & n21270 ) | ( n21269 & n21270 ) ;
  assign n21272 = x32 & ~n21267 ;
  assign n21273 = x32 & ~n21266 ;
  assign n21274 = ( ~n7178 & n21272 ) | ( ~n7178 & n21273 ) | ( n21272 & n21273 ) ;
  assign n21275 = ( n21268 & ~n21271 ) | ( n21268 & n21274 ) | ( ~n21271 & n21274 ) ;
  assign n21276 = n20900 & ~n20902 ;
  assign n21277 = n20900 | n20927 ;
  assign n21278 = ( n20902 & n20927 ) | ( n20902 & n21277 ) | ( n20927 & n21277 ) ;
  assign n21279 = ( n20903 & n21276 ) | ( n20903 & n21278 ) | ( n21276 & n21278 ) ;
  assign n21280 = n20903 | n21278 ;
  assign n21281 = ( n20904 & n21279 ) | ( n20904 & n21280 ) | ( n21279 & n21280 ) ;
  assign n21282 = n21275 & n21281 ;
  assign n21283 = n21275 | n21281 ;
  assign n21284 = ~n21282 & n21283 ;
  assign n21285 = n20840 & n20843 ;
  assign n21286 = ( n20823 & n20840 ) | ( n20823 & n21285 ) | ( n20840 & n21285 ) ;
  assign n21287 = n20681 | n20683 ;
  assign n21288 = n20682 | n21287 ;
  assign n21289 = ( n20676 & n20681 ) | ( n20676 & n21288 ) | ( n20681 & n21288 ) ;
  assign n21290 = x72 & n17146 ;
  assign n21291 = x71 & n17141 ;
  assign n21292 = x70 & ~n17140 ;
  assign n21293 = n17724 & n21292 ;
  assign n21294 = n21291 | n21293 ;
  assign n21295 = n21290 | n21294 ;
  assign n21296 = ( n513 & n17149 ) | ( n513 & n21295 ) | ( n17149 & n21295 ) ;
  assign n21297 = ( x62 & n17149 ) | ( x62 & ~n21290 ) | ( n17149 & ~n21290 ) ;
  assign n21298 = x62 & n17149 ;
  assign n21299 = ( ~n21294 & n21297 ) | ( ~n21294 & n21298 ) | ( n21297 & n21298 ) ;
  assign n21300 = ( x62 & n513 ) | ( x62 & n21299 ) | ( n513 & n21299 ) ;
  assign n21301 = ~n21296 & n21300 ;
  assign n21302 = x69 & n18290 ;
  assign n21303 = x63 & x68 ;
  assign n21304 = ~n18290 & n21303 ;
  assign n21305 = n21302 | n21304 ;
  assign n21306 = x2 & n21305 ;
  assign n21307 = n21305 & ~n21306 ;
  assign n21308 = x2 & ~n21305 ;
  assign n21309 = n21307 | n21308 ;
  assign n21310 = n21295 | n21299 ;
  assign n21311 = x62 | n21295 ;
  assign n21312 = ( n513 & n21310 ) | ( n513 & n21311 ) | ( n21310 & n21311 ) ;
  assign n21313 = n21309 & ~n21312 ;
  assign n21314 = x62 & n21309 ;
  assign n21315 = ( ~n21301 & n21313 ) | ( ~n21301 & n21314 ) | ( n21313 & n21314 ) ;
  assign n21316 = n21289 & n21315 ;
  assign n21317 = ~n21309 & n21312 ;
  assign n21318 = x62 | n21309 ;
  assign n21319 = ( n21301 & n21317 ) | ( n21301 & ~n21318 ) | ( n21317 & ~n21318 ) ;
  assign n21320 = ( n21289 & n21316 ) | ( n21289 & n21319 ) | ( n21316 & n21319 ) ;
  assign n21321 = n21289 | n21315 ;
  assign n21322 = n21319 | n21321 ;
  assign n21323 = ~n21320 & n21322 ;
  assign n21324 = x75 & n15552 ;
  assign n21325 = x74 & n15547 ;
  assign n21326 = x73 & ~n15546 ;
  assign n21327 = n16123 & n21326 ;
  assign n21328 = n21325 | n21327 ;
  assign n21329 = n21324 | n21328 ;
  assign n21330 = n15555 | n21324 ;
  assign n21331 = n21328 | n21330 ;
  assign n21332 = ( n746 & n21329 ) | ( n746 & n21331 ) | ( n21329 & n21331 ) ;
  assign n21333 = x59 & n21331 ;
  assign n21334 = x59 & n21324 ;
  assign n21335 = ( x59 & n21328 ) | ( x59 & n21334 ) | ( n21328 & n21334 ) ;
  assign n21336 = ( n746 & n21333 ) | ( n746 & n21335 ) | ( n21333 & n21335 ) ;
  assign n21337 = x59 & ~n21335 ;
  assign n21338 = x59 & ~n21331 ;
  assign n21339 = ( ~n746 & n21337 ) | ( ~n746 & n21338 ) | ( n21337 & n21338 ) ;
  assign n21340 = ( n21332 & ~n21336 ) | ( n21332 & n21339 ) | ( ~n21336 & n21339 ) ;
  assign n21341 = n21323 | n21340 ;
  assign n21342 = n21323 & n21340 ;
  assign n21343 = n21341 & ~n21342 ;
  assign n21344 = ( n20691 & n20692 ) | ( n20691 & n20712 ) | ( n20692 & n20712 ) ;
  assign n21345 = n21343 & n21344 ;
  assign n21346 = n21343 | n21344 ;
  assign n21347 = ~n21345 & n21346 ;
  assign n21348 = x78 & n14045 ;
  assign n21349 = x77 & n14040 ;
  assign n21350 = x76 & ~n14039 ;
  assign n21351 = n14552 & n21350 ;
  assign n21352 = n21349 | n21351 ;
  assign n21353 = n21348 | n21352 ;
  assign n21354 = n14048 | n21348 ;
  assign n21355 = n21352 | n21354 ;
  assign n21356 = ( n1192 & n21353 ) | ( n1192 & n21355 ) | ( n21353 & n21355 ) ;
  assign n21357 = x56 & n21355 ;
  assign n21358 = x56 & n21348 ;
  assign n21359 = ( x56 & n21352 ) | ( x56 & n21358 ) | ( n21352 & n21358 ) ;
  assign n21360 = ( n1192 & n21357 ) | ( n1192 & n21359 ) | ( n21357 & n21359 ) ;
  assign n21361 = x56 & ~n21359 ;
  assign n21362 = x56 & ~n21355 ;
  assign n21363 = ( ~n1192 & n21361 ) | ( ~n1192 & n21362 ) | ( n21361 & n21362 ) ;
  assign n21364 = ( n21356 & ~n21360 ) | ( n21356 & n21363 ) | ( ~n21360 & n21363 ) ;
  assign n21365 = n21347 & ~n21364 ;
  assign n21366 = n21347 | n21364 ;
  assign n21367 = ( ~n21347 & n21365 ) | ( ~n21347 & n21366 ) | ( n21365 & n21366 ) ;
  assign n21368 = n20714 | n20738 ;
  assign n21369 = ( n20718 & n20738 ) | ( n20718 & n21368 ) | ( n20738 & n21368 ) ;
  assign n21370 = ( n20720 & n20721 ) | ( n20720 & n21369 ) | ( n20721 & n21369 ) ;
  assign n21371 = n21367 & n21370 ;
  assign n21372 = n21367 & ~n21371 ;
  assign n21373 = x81 & n12574 ;
  assign n21374 = x80 & n12569 ;
  assign n21375 = x79 & ~n12568 ;
  assign n21376 = n13076 & n21375 ;
  assign n21377 = n21374 | n21376 ;
  assign n21378 = n21373 | n21377 ;
  assign n21379 = n12577 | n21373 ;
  assign n21380 = n21377 | n21379 ;
  assign n21381 = ( n1651 & n21378 ) | ( n1651 & n21380 ) | ( n21378 & n21380 ) ;
  assign n21382 = x53 & n21380 ;
  assign n21383 = x53 & n21373 ;
  assign n21384 = ( x53 & n21377 ) | ( x53 & n21383 ) | ( n21377 & n21383 ) ;
  assign n21385 = ( n1651 & n21382 ) | ( n1651 & n21384 ) | ( n21382 & n21384 ) ;
  assign n21386 = x53 & ~n21384 ;
  assign n21387 = x53 & ~n21380 ;
  assign n21388 = ( ~n1651 & n21386 ) | ( ~n1651 & n21387 ) | ( n21386 & n21387 ) ;
  assign n21389 = ( n21381 & ~n21385 ) | ( n21381 & n21388 ) | ( ~n21385 & n21388 ) ;
  assign n21390 = ~n21367 & n21370 ;
  assign n21391 = n21389 & n21390 ;
  assign n21392 = ( n21372 & n21389 ) | ( n21372 & n21391 ) | ( n21389 & n21391 ) ;
  assign n21393 = n21389 | n21390 ;
  assign n21394 = n21372 | n21393 ;
  assign n21395 = ~n21392 & n21394 ;
  assign n21396 = n20744 | n20764 ;
  assign n21397 = ( n20741 & n20764 ) | ( n20741 & n21396 ) | ( n20764 & n21396 ) ;
  assign n21398 = ( n20746 & n20747 ) | ( n20746 & n21397 ) | ( n20747 & n21397 ) ;
  assign n21399 = n21395 | n21398 ;
  assign n21400 = n21395 & n21398 ;
  assign n21401 = n21399 & ~n21400 ;
  assign n21402 = x84 & n11205 ;
  assign n21403 = x83 & n11200 ;
  assign n21404 = x82 & ~n11199 ;
  assign n21405 = n11679 & n21404 ;
  assign n21406 = n21403 | n21405 ;
  assign n21407 = n21402 | n21406 ;
  assign n21408 = n11208 | n21402 ;
  assign n21409 = n21406 | n21408 ;
  assign n21410 = ( n2194 & n21407 ) | ( n2194 & n21409 ) | ( n21407 & n21409 ) ;
  assign n21411 = x50 & n21409 ;
  assign n21412 = x50 & n21402 ;
  assign n21413 = ( x50 & n21406 ) | ( x50 & n21412 ) | ( n21406 & n21412 ) ;
  assign n21414 = ( n2194 & n21411 ) | ( n2194 & n21413 ) | ( n21411 & n21413 ) ;
  assign n21415 = x50 & ~n21413 ;
  assign n21416 = x50 & ~n21409 ;
  assign n21417 = ( ~n2194 & n21415 ) | ( ~n2194 & n21416 ) | ( n21415 & n21416 ) ;
  assign n21418 = ( n21410 & ~n21414 ) | ( n21410 & n21417 ) | ( ~n21414 & n21417 ) ;
  assign n21419 = n21401 | n21418 ;
  assign n21420 = n21401 & n21418 ;
  assign n21421 = n21419 & ~n21420 ;
  assign n21422 = n20792 & n21421 ;
  assign n21423 = n20771 & n21421 ;
  assign n21424 = ( n20772 & n21422 ) | ( n20772 & n21423 ) | ( n21422 & n21423 ) ;
  assign n21425 = n20792 | n21421 ;
  assign n21426 = n20771 | n21421 ;
  assign n21427 = ( n20772 & n21425 ) | ( n20772 & n21426 ) | ( n21425 & n21426 ) ;
  assign n21428 = ~n21424 & n21427 ;
  assign n21429 = x87 & n9933 ;
  assign n21430 = x86 & n9928 ;
  assign n21431 = x85 & ~n9927 ;
  assign n21432 = n10379 & n21431 ;
  assign n21433 = n21430 | n21432 ;
  assign n21434 = n21429 | n21433 ;
  assign n21435 = n9936 | n21429 ;
  assign n21436 = n21433 | n21435 ;
  assign n21437 = ( n2816 & n21434 ) | ( n2816 & n21436 ) | ( n21434 & n21436 ) ;
  assign n21438 = x47 & n21436 ;
  assign n21439 = x47 & n21429 ;
  assign n21440 = ( x47 & n21433 ) | ( x47 & n21439 ) | ( n21433 & n21439 ) ;
  assign n21441 = ( n2816 & n21438 ) | ( n2816 & n21440 ) | ( n21438 & n21440 ) ;
  assign n21442 = x47 & ~n21440 ;
  assign n21443 = x47 & ~n21436 ;
  assign n21444 = ( ~n2816 & n21442 ) | ( ~n2816 & n21443 ) | ( n21442 & n21443 ) ;
  assign n21445 = ( n21437 & ~n21441 ) | ( n21437 & n21444 ) | ( ~n21441 & n21444 ) ;
  assign n21446 = n21428 & ~n21445 ;
  assign n21447 = n21428 | n21445 ;
  assign n21448 = ( ~n21428 & n21446 ) | ( ~n21428 & n21447 ) | ( n21446 & n21447 ) ;
  assign n21449 = ( n20797 & n20798 ) | ( n20797 & n20817 ) | ( n20798 & n20817 ) ;
  assign n21450 = n21448 | n21449 ;
  assign n21451 = n21448 & n21449 ;
  assign n21452 = n21450 & ~n21451 ;
  assign n21453 = x90 & n8724 ;
  assign n21454 = x89 & n8719 ;
  assign n21455 = x88 & ~n8718 ;
  assign n21456 = n9149 & n21455 ;
  assign n21457 = n21454 | n21456 ;
  assign n21458 = n21453 | n21457 ;
  assign n21459 = n8727 | n21453 ;
  assign n21460 = n21457 | n21459 ;
  assign n21461 = ( n3519 & n21458 ) | ( n3519 & n21460 ) | ( n21458 & n21460 ) ;
  assign n21462 = x44 & n21460 ;
  assign n21463 = x44 & n21453 ;
  assign n21464 = ( x44 & n21457 ) | ( x44 & n21463 ) | ( n21457 & n21463 ) ;
  assign n21465 = ( n3519 & n21462 ) | ( n3519 & n21464 ) | ( n21462 & n21464 ) ;
  assign n21466 = x44 & ~n21464 ;
  assign n21467 = x44 & ~n21460 ;
  assign n21468 = ( ~n3519 & n21466 ) | ( ~n3519 & n21467 ) | ( n21466 & n21467 ) ;
  assign n21469 = ( n21461 & ~n21465 ) | ( n21461 & n21468 ) | ( ~n21465 & n21468 ) ;
  assign n21470 = ~n21452 & n21469 ;
  assign n21471 = n21448 | n21469 ;
  assign n21472 = ( n21449 & n21469 ) | ( n21449 & n21471 ) | ( n21469 & n21471 ) ;
  assign n21473 = n21450 & ~n21472 ;
  assign n21474 = n21470 | n21473 ;
  assign n21475 = n20822 | n21474 ;
  assign n21476 = n21286 | n21475 ;
  assign n21477 = n20822 & n21474 ;
  assign n21478 = ( n21286 & n21474 ) | ( n21286 & n21477 ) | ( n21474 & n21477 ) ;
  assign n21479 = n21476 & ~n21478 ;
  assign n21480 = x93 & n7566 ;
  assign n21481 = x92 & n7561 ;
  assign n21482 = x91 & ~n7560 ;
  assign n21483 = n7953 & n21482 ;
  assign n21484 = n21481 | n21483 ;
  assign n21485 = n21480 | n21484 ;
  assign n21486 = n7569 | n21480 ;
  assign n21487 = n21484 | n21486 ;
  assign n21488 = ( n4305 & n21485 ) | ( n4305 & n21487 ) | ( n21485 & n21487 ) ;
  assign n21489 = x41 & n21487 ;
  assign n21490 = x41 & n21480 ;
  assign n21491 = ( x41 & n21484 ) | ( x41 & n21490 ) | ( n21484 & n21490 ) ;
  assign n21492 = ( n4305 & n21489 ) | ( n4305 & n21491 ) | ( n21489 & n21491 ) ;
  assign n21493 = x41 & ~n21491 ;
  assign n21494 = x41 & ~n21487 ;
  assign n21495 = ( ~n4305 & n21493 ) | ( ~n4305 & n21494 ) | ( n21493 & n21494 ) ;
  assign n21496 = ( n21488 & ~n21492 ) | ( n21488 & n21495 ) | ( ~n21492 & n21495 ) ;
  assign n21497 = ~n21479 & n21496 ;
  assign n21498 = n20822 | n21496 ;
  assign n21499 = ( n21474 & n21496 ) | ( n21474 & n21498 ) | ( n21496 & n21498 ) ;
  assign n21500 = n21473 | n21496 ;
  assign n21501 = n21470 | n21500 ;
  assign n21502 = ( n21286 & n21499 ) | ( n21286 & n21501 ) | ( n21499 & n21501 ) ;
  assign n21503 = n21476 & ~n21502 ;
  assign n21504 = n21497 | n21503 ;
  assign n21505 = ( n20853 & n20854 ) | ( n20853 & n20874 ) | ( n20854 & n20874 ) ;
  assign n21506 = n21504 | n21505 ;
  assign n21507 = n21504 & n21505 ;
  assign n21508 = n21506 & ~n21507 ;
  assign n21509 = x96 & n6536 ;
  assign n21510 = x95 & n6531 ;
  assign n21511 = x94 & ~n6530 ;
  assign n21512 = n6871 & n21511 ;
  assign n21513 = n21510 | n21512 ;
  assign n21514 = n21509 | n21513 ;
  assign n21515 = n6539 | n21509 ;
  assign n21516 = n21513 | n21515 ;
  assign n21517 = ( n5202 & n21514 ) | ( n5202 & n21516 ) | ( n21514 & n21516 ) ;
  assign n21518 = x38 & n21516 ;
  assign n21519 = x38 & n21509 ;
  assign n21520 = ( x38 & n21513 ) | ( x38 & n21519 ) | ( n21513 & n21519 ) ;
  assign n21521 = ( n5202 & n21518 ) | ( n5202 & n21520 ) | ( n21518 & n21520 ) ;
  assign n21522 = x38 & ~n21520 ;
  assign n21523 = x38 & ~n21516 ;
  assign n21524 = ( ~n5202 & n21522 ) | ( ~n5202 & n21523 ) | ( n21522 & n21523 ) ;
  assign n21525 = ( n21517 & ~n21521 ) | ( n21517 & n21524 ) | ( ~n21521 & n21524 ) ;
  assign n21526 = n21508 | n21525 ;
  assign n21527 = n21508 & n21525 ;
  assign n21528 = n21526 & ~n21527 ;
  assign n21529 = n20876 | n20897 ;
  assign n21530 = ( n20877 & n20897 ) | ( n20877 & n21529 ) | ( n20897 & n21529 ) ;
  assign n21531 = ( n20879 & n20880 ) | ( n20879 & n21530 ) | ( n20880 & n21530 ) ;
  assign n21532 = n21528 & n21531 ;
  assign n21533 = n21528 | n21531 ;
  assign n21534 = ~n21532 & n21533 ;
  assign n21535 = x99 & n5554 ;
  assign n21536 = x98 & n5549 ;
  assign n21537 = x97 & ~n5548 ;
  assign n21538 = n5893 & n21537 ;
  assign n21539 = n21536 | n21538 ;
  assign n21540 = n21535 | n21539 ;
  assign n21541 = n5557 | n21535 ;
  assign n21542 = n21539 | n21541 ;
  assign n21543 = ( n6164 & n21540 ) | ( n6164 & n21542 ) | ( n21540 & n21542 ) ;
  assign n21544 = x35 & n21542 ;
  assign n21545 = x35 & n21535 ;
  assign n21546 = ( x35 & n21539 ) | ( x35 & n21545 ) | ( n21539 & n21545 ) ;
  assign n21547 = ( n6164 & n21544 ) | ( n6164 & n21546 ) | ( n21544 & n21546 ) ;
  assign n21548 = x35 & ~n21546 ;
  assign n21549 = x35 & ~n21542 ;
  assign n21550 = ( ~n6164 & n21548 ) | ( ~n6164 & n21549 ) | ( n21548 & n21549 ) ;
  assign n21551 = ( n21543 & ~n21547 ) | ( n21543 & n21550 ) | ( ~n21547 & n21550 ) ;
  assign n21552 = n21534 & ~n21551 ;
  assign n21553 = n21534 | n21551 ;
  assign n21554 = ( ~n21534 & n21552 ) | ( ~n21534 & n21553 ) | ( n21552 & n21553 ) ;
  assign n21555 = n21284 & ~n21554 ;
  assign n21556 = n21284 | n21554 ;
  assign n21557 = ( ~n21284 & n21555 ) | ( ~n21284 & n21556 ) | ( n21555 & n21556 ) ;
  assign n21558 = ~n21258 & n21557 ;
  assign n21559 = ( n20655 & n20657 ) | ( n20655 & n21251 ) | ( n20657 & n21251 ) ;
  assign n21560 = n21249 | n21557 ;
  assign n21561 = ( n21557 & n21559 ) | ( n21557 & n21560 ) | ( n21559 & n21560 ) ;
  assign n21562 = n21254 & ~n21561 ;
  assign n21563 = n21558 | n21562 ;
  assign n21564 = n20957 | n20962 ;
  assign n21566 = x107 & n3080 ;
  assign n21567 = x106 & ~n3079 ;
  assign n21568 = n3309 & n21567 ;
  assign n21569 = n21566 | n21568 ;
  assign n21565 = x108 & n3085 ;
  assign n21571 = n3088 | n21565 ;
  assign n21572 = n21569 | n21571 ;
  assign n21570 = n21565 | n21569 ;
  assign n21573 = n21570 & n21572 ;
  assign n21574 = ( n9479 & n21572 ) | ( n9479 & n21573 ) | ( n21572 & n21573 ) ;
  assign n21575 = x26 & n21573 ;
  assign n21576 = x26 & n21572 ;
  assign n21577 = ( n9479 & n21575 ) | ( n9479 & n21576 ) | ( n21575 & n21576 ) ;
  assign n21578 = x26 & ~n21573 ;
  assign n21579 = x26 & ~n21572 ;
  assign n21580 = ( ~n9479 & n21578 ) | ( ~n9479 & n21579 ) | ( n21578 & n21579 ) ;
  assign n21581 = ( n21574 & ~n21577 ) | ( n21574 & n21580 ) | ( ~n21577 & n21580 ) ;
  assign n21582 = n20955 & n21581 ;
  assign n21583 = n20053 & n21582 ;
  assign n21584 = ( n20324 & n21582 ) | ( n20324 & n21583 ) | ( n21582 & n21583 ) ;
  assign n21585 = ( n20962 & n21581 ) | ( n20962 & n21584 ) | ( n21581 & n21584 ) ;
  assign n21586 = n21564 & ~n21585 ;
  assign n21587 = n21581 & ~n21583 ;
  assign n21588 = n21581 & ~n21582 ;
  assign n21589 = ( ~n20324 & n21587 ) | ( ~n20324 & n21588 ) | ( n21587 & n21588 ) ;
  assign n21590 = n21563 & n21589 ;
  assign n21591 = ~n20962 & n21590 ;
  assign n21592 = ( n21563 & n21586 ) | ( n21563 & n21591 ) | ( n21586 & n21591 ) ;
  assign n21593 = n21563 | n21589 ;
  assign n21594 = ( ~n20962 & n21563 ) | ( ~n20962 & n21593 ) | ( n21563 & n21593 ) ;
  assign n21595 = n21586 | n21594 ;
  assign n21596 = ~n21592 & n21595 ;
  assign n21597 = ~n21232 & n21596 ;
  assign n21598 = ( n20634 & n20635 ) | ( n20634 & n20968 ) | ( n20635 & n20968 ) ;
  assign n21599 = n21225 | n21596 ;
  assign n21600 = ( n21596 & n21598 ) | ( n21596 & n21599 ) | ( n21598 & n21599 ) ;
  assign n21601 = n21228 & ~n21600 ;
  assign n21602 = n21597 | n21601 ;
  assign n21603 = n20987 & n20989 ;
  assign n21604 = n20989 & ~n21603 ;
  assign n21605 = n20969 & n20987 ;
  assign n21606 = ( n20966 & n20987 ) | ( n20966 & n21605 ) | ( n20987 & n21605 ) ;
  assign n21607 = ~n20989 & n21606 ;
  assign n21608 = n21603 | n21607 ;
  assign n21609 = n20970 | n20987 ;
  assign n21610 = ( n20970 & n20989 ) | ( n20970 & n21609 ) | ( n20989 & n21609 ) ;
  assign n21611 = ( n21604 & n21608 ) | ( n21604 & n21610 ) | ( n21608 & n21610 ) ;
  assign n21612 = ( n21208 & n21602 ) | ( n21208 & ~n21611 ) | ( n21602 & ~n21611 ) ;
  assign n21613 = ( ~n21602 & n21611 ) | ( ~n21602 & n21612 ) | ( n21611 & n21612 ) ;
  assign n21614 = ( ~n21208 & n21612 ) | ( ~n21208 & n21613 ) | ( n21612 & n21613 ) ;
  assign n21615 = n21194 & ~n21614 ;
  assign n21616 = n21194 | n21614 ;
  assign n21617 = ( ~n21194 & n21615 ) | ( ~n21194 & n21616 ) | ( n21615 & n21616 ) ;
  assign n21618 = n21010 & n21012 ;
  assign n21619 = n21012 & ~n21618 ;
  assign n21620 = n20996 & n21010 ;
  assign n21621 = ~n21012 & n21620 ;
  assign n21622 = n21618 | n21621 ;
  assign n21623 = n20996 | n21010 ;
  assign n21624 = ( n20996 & n21012 ) | ( n20996 & n21623 ) | ( n21012 & n21623 ) ;
  assign n21625 = ( n21619 & n21622 ) | ( n21619 & n21624 ) | ( n21622 & n21624 ) ;
  assign n21626 = ( n21175 & n21617 ) | ( n21175 & ~n21625 ) | ( n21617 & ~n21625 ) ;
  assign n21627 = ( ~n21617 & n21625 ) | ( ~n21617 & n21626 ) | ( n21625 & n21626 ) ;
  assign n21628 = ( ~n21175 & n21626 ) | ( ~n21175 & n21627 ) | ( n21626 & n21627 ) ;
  assign n21629 = ~n21158 & n21628 ;
  assign n21630 = n21151 | n21626 ;
  assign n21631 = ~n21151 & n21175 ;
  assign n21632 = ( n21627 & n21630 ) | ( n21627 & ~n21631 ) | ( n21630 & ~n21631 ) ;
  assign n21633 = ( n21020 & n21628 ) | ( n21020 & n21632 ) | ( n21628 & n21632 ) ;
  assign n21634 = ( n20576 & n21628 ) | ( n20576 & n21632 ) | ( n21628 & n21632 ) ;
  assign n21635 = ( n20577 & n21633 ) | ( n20577 & n21634 ) | ( n21633 & n21634 ) ;
  assign n21636 = n21154 & ~n21635 ;
  assign n21637 = n21629 | n21636 ;
  assign n21638 = n21127 & ~n21129 ;
  assign n21639 = ~n21045 & n21127 ;
  assign n21640 = ( ~n20448 & n21638 ) | ( ~n20448 & n21639 ) | ( n21638 & n21639 ) ;
  assign n21641 = n21637 | n21640 ;
  assign n21642 = ( ~n21051 & n21637 ) | ( ~n21051 & n21641 ) | ( n21637 & n21641 ) ;
  assign n21643 = n21134 | n21642 ;
  assign n21644 = n21637 & n21640 ;
  assign n21645 = ~n21051 & n21644 ;
  assign n21646 = ( n21134 & n21637 ) | ( n21134 & n21645 ) | ( n21637 & n21645 ) ;
  assign n21647 = n21643 & ~n21646 ;
  assign n21648 = ~n20548 & n21101 ;
  assign n21649 = ( ~n20550 & n21101 ) | ( ~n20550 & n21648 ) | ( n21101 & n21648 ) ;
  assign n21650 = n21647 & n21649 ;
  assign n21651 = ~n21058 & n21650 ;
  assign n21652 = ( n21107 & n21647 ) | ( n21107 & n21651 ) | ( n21647 & n21651 ) ;
  assign n21653 = n21647 | n21649 ;
  assign n21654 = ( ~n21058 & n21647 ) | ( ~n21058 & n21653 ) | ( n21647 & n21653 ) ;
  assign n21655 = n21107 | n21654 ;
  assign n21656 = ~n21652 & n21655 ;
  assign n21657 = n20525 & n21656 ;
  assign n21658 = ( n21066 & n21656 ) | ( n21066 & n21657 ) | ( n21656 & n21657 ) ;
  assign n21659 = n21080 & ~n21658 ;
  assign n21660 = ~n20525 & n21656 ;
  assign n21661 = ~n21066 & n21660 ;
  assign n21662 = n21659 | n21661 ;
  assign n21663 = n21071 | n21078 ;
  assign n21664 = n21662 | n21663 ;
  assign n21665 = ~n21663 & n21664 ;
  assign n21666 = ( ~n21662 & n21664 ) | ( ~n21662 & n21665 ) | ( n21664 & n21665 ) ;
  assign n21667 = x127 & n389 ;
  assign n21668 = x126 & n384 ;
  assign n21669 = x125 & ~n383 ;
  assign n21670 = n463 & n21669 ;
  assign n21671 = n21668 | n21670 ;
  assign n21672 = n21667 | n21671 ;
  assign n21673 = n392 | n21667 ;
  assign n21674 = n21671 | n21673 ;
  assign n21675 = ( n18763 & n21672 ) | ( n18763 & n21674 ) | ( n21672 & n21674 ) ;
  assign n21676 = x8 & n21674 ;
  assign n21677 = x8 & n21667 ;
  assign n21678 = ( x8 & n21671 ) | ( x8 & n21677 ) | ( n21671 & n21677 ) ;
  assign n21679 = ( n18763 & n21676 ) | ( n18763 & n21678 ) | ( n21676 & n21678 ) ;
  assign n21680 = x8 & ~n21678 ;
  assign n21681 = x8 & ~n21674 ;
  assign n21682 = ( ~n18763 & n21680 ) | ( ~n18763 & n21681 ) | ( n21680 & n21681 ) ;
  assign n21683 = ( n21675 & ~n21679 ) | ( n21675 & n21682 ) | ( ~n21679 & n21682 ) ;
  assign n22210 = n21133 | n21645 ;
  assign n21684 = x124 & n636 ;
  assign n21685 = x123 & n631 ;
  assign n21686 = x122 & ~n630 ;
  assign n21687 = n764 & n21686 ;
  assign n21688 = n21685 | n21687 ;
  assign n21689 = n21684 | n21688 ;
  assign n21690 = n639 | n21684 ;
  assign n21691 = n21688 | n21690 ;
  assign n21692 = ( n17084 & n21689 ) | ( n17084 & n21691 ) | ( n21689 & n21691 ) ;
  assign n21693 = x11 & n21691 ;
  assign n21694 = x11 & n21684 ;
  assign n21695 = ( x11 & n21688 ) | ( x11 & n21694 ) | ( n21688 & n21694 ) ;
  assign n21696 = ( n17084 & n21693 ) | ( n17084 & n21695 ) | ( n21693 & n21695 ) ;
  assign n21697 = x11 & ~n21695 ;
  assign n21698 = x11 & ~n21691 ;
  assign n21699 = ( ~n17084 & n21697 ) | ( ~n17084 & n21698 ) | ( n21697 & n21698 ) ;
  assign n21700 = ( n21692 & ~n21696 ) | ( n21692 & n21699 ) | ( ~n21696 & n21699 ) ;
  assign n21701 = n21635 | n21700 ;
  assign n21702 = n21157 | n21700 ;
  assign n21703 = ( n21158 & n21701 ) | ( n21158 & n21702 ) | ( n21701 & n21702 ) ;
  assign n21704 = n21635 & n21700 ;
  assign n21705 = n21157 & n21700 ;
  assign n21706 = ( n21158 & n21704 ) | ( n21158 & n21705 ) | ( n21704 & n21705 ) ;
  assign n21707 = n21703 & ~n21706 ;
  assign n21708 = n21010 & n21175 ;
  assign n21709 = n21012 & n21708 ;
  assign n21710 = ( n21175 & n21621 ) | ( n21175 & n21709 ) | ( n21621 & n21709 ) ;
  assign n21711 = ( n20996 & n21175 ) | ( n20996 & n21708 ) | ( n21175 & n21708 ) ;
  assign n21712 = n20996 & n21175 ;
  assign n21713 = ( n21012 & n21711 ) | ( n21012 & n21712 ) | ( n21711 & n21712 ) ;
  assign n21714 = ( n21619 & n21710 ) | ( n21619 & n21713 ) | ( n21710 & n21713 ) ;
  assign n21715 = n21625 & ~n21714 ;
  assign n21716 = n21175 & ~n21708 ;
  assign n21717 = ( ~n21012 & n21175 ) | ( ~n21012 & n21716 ) | ( n21175 & n21716 ) ;
  assign n21718 = ~n21621 & n21717 ;
  assign n21719 = ~n20996 & n21716 ;
  assign n21720 = ~n20996 & n21175 ;
  assign n21721 = ( ~n21012 & n21719 ) | ( ~n21012 & n21720 ) | ( n21719 & n21720 ) ;
  assign n21722 = ( ~n21619 & n21718 ) | ( ~n21619 & n21721 ) | ( n21718 & n21721 ) ;
  assign n21723 = n21617 & n21722 ;
  assign n21724 = ( n21617 & n21715 ) | ( n21617 & n21723 ) | ( n21715 & n21723 ) ;
  assign n21725 = x121 & n962 ;
  assign n21726 = x120 & n957 ;
  assign n21727 = x119 & ~n956 ;
  assign n21728 = n1105 & n21727 ;
  assign n21729 = n21726 | n21728 ;
  assign n21730 = n21725 | n21729 ;
  assign n21731 = n965 | n21725 ;
  assign n21732 = n21729 | n21731 ;
  assign n21733 = ( n15501 & n21730 ) | ( n15501 & n21732 ) | ( n21730 & n21732 ) ;
  assign n21734 = x14 & n21732 ;
  assign n21735 = x14 & n21725 ;
  assign n21736 = ( x14 & n21729 ) | ( x14 & n21735 ) | ( n21729 & n21735 ) ;
  assign n21737 = ( n15501 & n21734 ) | ( n15501 & n21736 ) | ( n21734 & n21736 ) ;
  assign n21738 = x14 & ~n21736 ;
  assign n21739 = x14 & ~n21732 ;
  assign n21740 = ( ~n15501 & n21738 ) | ( ~n15501 & n21739 ) | ( n21738 & n21739 ) ;
  assign n21741 = ( n21733 & ~n21737 ) | ( n21733 & n21740 ) | ( ~n21737 & n21740 ) ;
  assign n21742 = n21714 & n21741 ;
  assign n21743 = ( n21724 & n21741 ) | ( n21724 & n21742 ) | ( n21741 & n21742 ) ;
  assign n21744 = n21714 | n21741 ;
  assign n21745 = n21724 | n21744 ;
  assign n21746 = ~n21743 & n21745 ;
  assign n21747 = n21190 | n21614 ;
  assign n21748 = ( n21191 & n21614 ) | ( n21191 & n21747 ) | ( n21614 & n21747 ) ;
  assign n21749 = ( n21192 & n21194 ) | ( n21192 & n21748 ) | ( n21194 & n21748 ) ;
  assign n21750 = x118 & n1383 ;
  assign n21751 = x117 & n1378 ;
  assign n21752 = x116 & ~n1377 ;
  assign n21753 = n1542 & n21752 ;
  assign n21754 = n21751 | n21753 ;
  assign n21755 = n21750 | n21754 ;
  assign n21756 = n1386 | n21750 ;
  assign n21757 = n21754 | n21756 ;
  assign n21758 = ( ~n14002 & n21755 ) | ( ~n14002 & n21757 ) | ( n21755 & n21757 ) ;
  assign n21759 = n21755 & n21757 ;
  assign n21760 = ( n13981 & n21758 ) | ( n13981 & n21759 ) | ( n21758 & n21759 ) ;
  assign n21761 = x17 & n21760 ;
  assign n21762 = x17 & ~n21760 ;
  assign n21763 = ( n21760 & ~n21761 ) | ( n21760 & n21762 ) | ( ~n21761 & n21762 ) ;
  assign n21764 = n21748 & n21763 ;
  assign n21765 = n21192 & n21763 ;
  assign n21766 = ( n21194 & n21764 ) | ( n21194 & n21765 ) | ( n21764 & n21765 ) ;
  assign n21767 = n21749 & ~n21766 ;
  assign n21768 = n20987 & n21208 ;
  assign n21769 = n20989 & n21768 ;
  assign n21770 = ( n21208 & n21607 ) | ( n21208 & n21769 ) | ( n21607 & n21769 ) ;
  assign n21771 = ( n20970 & n21208 ) | ( n20970 & n21768 ) | ( n21208 & n21768 ) ;
  assign n21772 = n20970 & n21208 ;
  assign n21773 = ( n20989 & n21771 ) | ( n20989 & n21772 ) | ( n21771 & n21772 ) ;
  assign n21774 = ( n21604 & n21770 ) | ( n21604 & n21773 ) | ( n21770 & n21773 ) ;
  assign n21775 = n21611 & ~n21774 ;
  assign n21776 = n21208 & ~n21768 ;
  assign n21777 = ( ~n20989 & n21208 ) | ( ~n20989 & n21776 ) | ( n21208 & n21776 ) ;
  assign n21778 = ~n21607 & n21777 ;
  assign n21779 = ~n20970 & n21776 ;
  assign n21780 = ~n20970 & n21208 ;
  assign n21781 = ( ~n20989 & n21779 ) | ( ~n20989 & n21780 ) | ( n21779 & n21780 ) ;
  assign n21782 = ( ~n21604 & n21778 ) | ( ~n21604 & n21781 ) | ( n21778 & n21781 ) ;
  assign n21783 = n21602 & n21782 ;
  assign n21784 = ( n21602 & n21775 ) | ( n21602 & n21783 ) | ( n21775 & n21783 ) ;
  assign n21785 = x115 & n1859 ;
  assign n21786 = x114 & n1854 ;
  assign n21787 = x113 & ~n1853 ;
  assign n21788 = n2037 & n21787 ;
  assign n21789 = n21786 | n21788 ;
  assign n21790 = n21785 | n21789 ;
  assign n21791 = n1862 | n21785 ;
  assign n21792 = n21789 | n21791 ;
  assign n21793 = ( ~n12550 & n21790 ) | ( ~n12550 & n21792 ) | ( n21790 & n21792 ) ;
  assign n21794 = n21790 & n21792 ;
  assign n21795 = ( n12532 & n21793 ) | ( n12532 & n21794 ) | ( n21793 & n21794 ) ;
  assign n21796 = x20 & n21795 ;
  assign n21797 = x20 & ~n21795 ;
  assign n21798 = ( n21795 & ~n21796 ) | ( n21795 & n21797 ) | ( ~n21796 & n21797 ) ;
  assign n21799 = n21774 & n21798 ;
  assign n21800 = ( n21784 & n21798 ) | ( n21784 & n21799 ) | ( n21798 & n21799 ) ;
  assign n21801 = n21774 | n21798 ;
  assign n21802 = n21784 | n21801 ;
  assign n21803 = ~n21800 & n21802 ;
  assign n21804 = x112 & n2429 ;
  assign n21805 = x111 & n2424 ;
  assign n21806 = x110 & ~n2423 ;
  assign n21807 = n2631 & n21806 ;
  assign n21808 = n21805 | n21807 ;
  assign n21809 = n21804 | n21808 ;
  assign n21810 = n2432 | n21804 ;
  assign n21811 = n21808 | n21810 ;
  assign n21812 = ( n11172 & n21809 ) | ( n11172 & n21811 ) | ( n21809 & n21811 ) ;
  assign n21813 = x23 & n21811 ;
  assign n21814 = x23 & n21804 ;
  assign n21815 = ( x23 & n21808 ) | ( x23 & n21814 ) | ( n21808 & n21814 ) ;
  assign n21816 = ( n11172 & n21813 ) | ( n11172 & n21815 ) | ( n21813 & n21815 ) ;
  assign n21817 = x23 & ~n21815 ;
  assign n21818 = x23 & ~n21811 ;
  assign n21819 = ( ~n11172 & n21817 ) | ( ~n11172 & n21818 ) | ( n21817 & n21818 ) ;
  assign n21820 = ( n21812 & ~n21816 ) | ( n21812 & n21819 ) | ( ~n21816 & n21819 ) ;
  assign n21821 = ( n21231 & n21232 ) | ( n21231 & n21600 ) | ( n21232 & n21600 ) ;
  assign n21822 = n21820 | n21821 ;
  assign n21823 = n21820 & n21821 ;
  assign n21824 = n21822 & ~n21823 ;
  assign n21825 = x109 & n3085 ;
  assign n21826 = x108 & n3080 ;
  assign n21827 = x107 & ~n3079 ;
  assign n21828 = n3309 & n21827 ;
  assign n21829 = n21826 | n21828 ;
  assign n21830 = n21825 | n21829 ;
  assign n21831 = n3088 | n21825 ;
  assign n21832 = n21829 | n21831 ;
  assign n21833 = ( n9878 & n21830 ) | ( n9878 & n21832 ) | ( n21830 & n21832 ) ;
  assign n21834 = x26 & n21832 ;
  assign n21835 = x26 & n21825 ;
  assign n21836 = ( x26 & n21829 ) | ( x26 & n21835 ) | ( n21829 & n21835 ) ;
  assign n21837 = ( n9878 & n21834 ) | ( n9878 & n21836 ) | ( n21834 & n21836 ) ;
  assign n21838 = x26 & ~n21836 ;
  assign n21839 = x26 & ~n21832 ;
  assign n21840 = ( ~n9878 & n21838 ) | ( ~n9878 & n21839 ) | ( n21838 & n21839 ) ;
  assign n21841 = ( n21833 & ~n21837 ) | ( n21833 & n21840 ) | ( ~n21837 & n21840 ) ;
  assign n21842 = x106 & n3816 ;
  assign n21843 = x105 & n3811 ;
  assign n21844 = x104 & ~n3810 ;
  assign n21845 = n4067 & n21844 ;
  assign n21846 = n21843 | n21845 ;
  assign n21847 = n21842 | n21846 ;
  assign n21848 = n3819 | n21842 ;
  assign n21849 = n21846 | n21848 ;
  assign n21850 = ( n8656 & n21847 ) | ( n8656 & n21849 ) | ( n21847 & n21849 ) ;
  assign n21851 = x29 & n21849 ;
  assign n21852 = x29 & n21842 ;
  assign n21853 = ( x29 & n21846 ) | ( x29 & n21852 ) | ( n21846 & n21852 ) ;
  assign n21854 = ( n8656 & n21851 ) | ( n8656 & n21853 ) | ( n21851 & n21853 ) ;
  assign n21855 = x29 & ~n21853 ;
  assign n21856 = x29 & ~n21849 ;
  assign n21857 = ( ~n8656 & n21855 ) | ( ~n8656 & n21856 ) | ( n21855 & n21856 ) ;
  assign n21858 = ( n21850 & ~n21854 ) | ( n21850 & n21857 ) | ( ~n21854 & n21857 ) ;
  assign n21859 = ( n21257 & n21258 ) | ( n21257 & n21561 ) | ( n21258 & n21561 ) ;
  assign n21860 = n21858 | n21859 ;
  assign n21861 = n21858 & n21859 ;
  assign n21862 = n21860 & ~n21861 ;
  assign n21863 = x70 & n18290 ;
  assign n21864 = x63 & x69 ;
  assign n21865 = ~n18290 & n21864 ;
  assign n21866 = n21863 | n21865 ;
  assign n21867 = x2 & ~x5 ;
  assign n21868 = ~x2 & x5 ;
  assign n21869 = n21867 | n21868 ;
  assign n21870 = n21866 & n21869 ;
  assign n21871 = n21866 | n21869 ;
  assign n21872 = ~n21870 & n21871 ;
  assign n21873 = n21306 | n21308 ;
  assign n21874 = n21307 | n21873 ;
  assign n21875 = n21872 & n21874 ;
  assign n21876 = n21306 & n21872 ;
  assign n21877 = ( n21312 & n21875 ) | ( n21312 & n21876 ) | ( n21875 & n21876 ) ;
  assign n21878 = ( ~x62 & n21875 ) | ( ~x62 & n21876 ) | ( n21875 & n21876 ) ;
  assign n21879 = ( n21301 & n21877 ) | ( n21301 & n21878 ) | ( n21877 & n21878 ) ;
  assign n21880 = n21872 | n21874 ;
  assign n21881 = n21306 | n21872 ;
  assign n21882 = ( n21312 & n21880 ) | ( n21312 & n21881 ) | ( n21880 & n21881 ) ;
  assign n21883 = ( ~x62 & n21880 ) | ( ~x62 & n21881 ) | ( n21880 & n21881 ) ;
  assign n21884 = ( n21301 & n21882 ) | ( n21301 & n21883 ) | ( n21882 & n21883 ) ;
  assign n21885 = ~n21879 & n21884 ;
  assign n21886 = x73 & n17146 ;
  assign n21887 = x72 & n17141 ;
  assign n21888 = x71 & ~n17140 ;
  assign n21889 = n17724 & n21888 ;
  assign n21890 = n21887 | n21889 ;
  assign n21891 = n21886 | n21890 ;
  assign n21892 = ( ~n610 & n17149 ) | ( ~n610 & n21891 ) | ( n17149 & n21891 ) ;
  assign n21893 = n17149 & n21886 ;
  assign n21894 = ( n17149 & n21890 ) | ( n17149 & n21893 ) | ( n21890 & n21893 ) ;
  assign n21895 = ( n598 & n21892 ) | ( n598 & n21894 ) | ( n21892 & n21894 ) ;
  assign n21896 = ( x62 & ~n21891 ) | ( x62 & n21895 ) | ( ~n21891 & n21895 ) ;
  assign n21897 = ~n21895 & n21896 ;
  assign n21898 = x62 | n21886 ;
  assign n21899 = n21890 | n21898 ;
  assign n21900 = n21895 | n21899 ;
  assign n21901 = ( ~x62 & n21897 ) | ( ~x62 & n21900 ) | ( n21897 & n21900 ) ;
  assign n21902 = n21885 | n21901 ;
  assign n21903 = n21885 & n21901 ;
  assign n21904 = n21902 & ~n21903 ;
  assign n21905 = x76 & n15552 ;
  assign n21906 = x75 & n15547 ;
  assign n21907 = x74 & ~n15546 ;
  assign n21908 = n16123 & n21907 ;
  assign n21909 = n21906 | n21908 ;
  assign n21910 = n21905 | n21909 ;
  assign n21911 = n15555 | n21905 ;
  assign n21912 = n21909 | n21911 ;
  assign n21913 = ( n923 & n21910 ) | ( n923 & n21912 ) | ( n21910 & n21912 ) ;
  assign n21914 = x59 & n21912 ;
  assign n21915 = x59 & n21905 ;
  assign n21916 = ( x59 & n21909 ) | ( x59 & n21915 ) | ( n21909 & n21915 ) ;
  assign n21917 = ( n923 & n21914 ) | ( n923 & n21916 ) | ( n21914 & n21916 ) ;
  assign n21918 = x59 & ~n21916 ;
  assign n21919 = x59 & ~n21912 ;
  assign n21920 = ( ~n923 & n21918 ) | ( ~n923 & n21919 ) | ( n21918 & n21919 ) ;
  assign n21921 = ( n21913 & ~n21917 ) | ( n21913 & n21920 ) | ( ~n21917 & n21920 ) ;
  assign n21922 = n21904 & n21921 ;
  assign n21923 = n21904 & ~n21922 ;
  assign n21924 = n21319 | n21340 ;
  assign n21925 = n21289 | n21340 ;
  assign n21926 = ( n21316 & n21924 ) | ( n21316 & n21925 ) | ( n21924 & n21925 ) ;
  assign n21927 = ( n21320 & n21323 ) | ( n21320 & n21926 ) | ( n21323 & n21926 ) ;
  assign n21928 = ~n21904 & n21921 ;
  assign n21929 = n21927 & n21928 ;
  assign n21930 = ( n21923 & n21927 ) | ( n21923 & n21929 ) | ( n21927 & n21929 ) ;
  assign n21931 = n21927 | n21928 ;
  assign n21932 = n21923 | n21931 ;
  assign n21933 = ~n21930 & n21932 ;
  assign n21934 = x79 & n14045 ;
  assign n21935 = x78 & n14040 ;
  assign n21936 = x77 & ~n14039 ;
  assign n21937 = n14552 & n21936 ;
  assign n21938 = n21935 | n21937 ;
  assign n21939 = n21934 | n21938 ;
  assign n21940 = n14048 | n21934 ;
  assign n21941 = n21938 | n21940 ;
  assign n21942 = ( n1332 & n21939 ) | ( n1332 & n21941 ) | ( n21939 & n21941 ) ;
  assign n21943 = x56 & n21941 ;
  assign n21944 = x56 & n21934 ;
  assign n21945 = ( x56 & n21938 ) | ( x56 & n21944 ) | ( n21938 & n21944 ) ;
  assign n21946 = ( n1332 & n21943 ) | ( n1332 & n21945 ) | ( n21943 & n21945 ) ;
  assign n21947 = x56 & ~n21945 ;
  assign n21948 = x56 & ~n21941 ;
  assign n21949 = ( ~n1332 & n21947 ) | ( ~n1332 & n21948 ) | ( n21947 & n21948 ) ;
  assign n21950 = ( n21942 & ~n21946 ) | ( n21942 & n21949 ) | ( ~n21946 & n21949 ) ;
  assign n21951 = n21933 & n21950 ;
  assign n21952 = n21933 & ~n21951 ;
  assign n21954 = n21344 | n21364 ;
  assign n21955 = ( n21343 & n21364 ) | ( n21343 & n21954 ) | ( n21364 & n21954 ) ;
  assign n21956 = ( n21345 & n21347 ) | ( n21345 & n21955 ) | ( n21347 & n21955 ) ;
  assign n21953 = ~n21933 & n21950 ;
  assign n21957 = n21953 & n21956 ;
  assign n21958 = ( n21952 & n21956 ) | ( n21952 & n21957 ) | ( n21956 & n21957 ) ;
  assign n21959 = n21953 | n21956 ;
  assign n21960 = n21952 | n21959 ;
  assign n21961 = ~n21958 & n21960 ;
  assign n21962 = x82 & n12574 ;
  assign n21963 = x81 & n12569 ;
  assign n21964 = x80 & ~n12568 ;
  assign n21965 = n13076 & n21964 ;
  assign n21966 = n21963 | n21965 ;
  assign n21967 = n21962 | n21966 ;
  assign n21968 = n12577 | n21962 ;
  assign n21969 = n21966 | n21968 ;
  assign n21970 = ( n1811 & n21967 ) | ( n1811 & n21969 ) | ( n21967 & n21969 ) ;
  assign n21971 = x53 & n21969 ;
  assign n21972 = x53 & n21962 ;
  assign n21973 = ( x53 & n21966 ) | ( x53 & n21972 ) | ( n21966 & n21972 ) ;
  assign n21974 = ( n1811 & n21971 ) | ( n1811 & n21973 ) | ( n21971 & n21973 ) ;
  assign n21975 = x53 & ~n21973 ;
  assign n21976 = x53 & ~n21969 ;
  assign n21977 = ( ~n1811 & n21975 ) | ( ~n1811 & n21976 ) | ( n21975 & n21976 ) ;
  assign n21978 = ( n21970 & ~n21974 ) | ( n21970 & n21977 ) | ( ~n21974 & n21977 ) ;
  assign n21979 = n21961 & n21978 ;
  assign n21980 = n21961 & ~n21979 ;
  assign n21981 = ~n21961 & n21978 ;
  assign n21982 = n21980 | n21981 ;
  assign n21983 = n21371 | n21392 ;
  assign n21984 = n21982 | n21983 ;
  assign n21985 = n21982 & n21983 ;
  assign n21986 = n21984 & ~n21985 ;
  assign n21987 = x85 & n11205 ;
  assign n21988 = x84 & n11200 ;
  assign n21989 = x83 & ~n11199 ;
  assign n21990 = n11679 & n21989 ;
  assign n21991 = n21988 | n21990 ;
  assign n21992 = n21987 | n21991 ;
  assign n21993 = n11208 | n21987 ;
  assign n21994 = n21991 | n21993 ;
  assign n21995 = ( n2381 & n21992 ) | ( n2381 & n21994 ) | ( n21992 & n21994 ) ;
  assign n21996 = x50 & n21994 ;
  assign n21997 = x50 & n21987 ;
  assign n21998 = ( x50 & n21991 ) | ( x50 & n21997 ) | ( n21991 & n21997 ) ;
  assign n21999 = ( n2381 & n21996 ) | ( n2381 & n21998 ) | ( n21996 & n21998 ) ;
  assign n22000 = x50 & ~n21998 ;
  assign n22001 = x50 & ~n21994 ;
  assign n22002 = ( ~n2381 & n22000 ) | ( ~n2381 & n22001 ) | ( n22000 & n22001 ) ;
  assign n22003 = ( n21995 & ~n21999 ) | ( n21995 & n22002 ) | ( ~n21999 & n22002 ) ;
  assign n22004 = n21400 | n21418 ;
  assign n22005 = ( n21400 & n21401 ) | ( n21400 & n22004 ) | ( n21401 & n22004 ) ;
  assign n22006 = ( n21986 & ~n22003 ) | ( n21986 & n22005 ) | ( ~n22003 & n22005 ) ;
  assign n22007 = ( ~n21986 & n22003 ) | ( ~n21986 & n22006 ) | ( n22003 & n22006 ) ;
  assign n22008 = x88 & n9933 ;
  assign n22009 = x87 & n9928 ;
  assign n22010 = x86 & ~n9927 ;
  assign n22011 = n10379 & n22010 ;
  assign n22012 = n22009 | n22011 ;
  assign n22013 = n22008 | n22012 ;
  assign n22014 = n9936 | n22008 ;
  assign n22015 = n22012 | n22014 ;
  assign n22016 = ( ~n3039 & n22013 ) | ( ~n3039 & n22015 ) | ( n22013 & n22015 ) ;
  assign n22017 = n22013 & n22015 ;
  assign n22018 = ( n3023 & n22016 ) | ( n3023 & n22017 ) | ( n22016 & n22017 ) ;
  assign n22019 = x47 & n22015 ;
  assign n22020 = x47 & n22008 ;
  assign n22021 = ( x47 & n22012 ) | ( x47 & n22020 ) | ( n22012 & n22020 ) ;
  assign n22022 = ( ~n3039 & n22019 ) | ( ~n3039 & n22021 ) | ( n22019 & n22021 ) ;
  assign n22023 = n22019 & n22021 ;
  assign n22024 = ( n3023 & n22022 ) | ( n3023 & n22023 ) | ( n22022 & n22023 ) ;
  assign n22025 = x47 & ~n22021 ;
  assign n22026 = x47 & ~n22015 ;
  assign n22027 = ( n3039 & n22025 ) | ( n3039 & n22026 ) | ( n22025 & n22026 ) ;
  assign n22028 = n22025 | n22026 ;
  assign n22029 = ( ~n3023 & n22027 ) | ( ~n3023 & n22028 ) | ( n22027 & n22028 ) ;
  assign n22030 = ( n22018 & ~n22024 ) | ( n22018 & n22029 ) | ( ~n22024 & n22029 ) ;
  assign n22031 = n22006 & n22030 ;
  assign n22032 = ~n22005 & n22030 ;
  assign n22033 = ( n22007 & n22031 ) | ( n22007 & n22032 ) | ( n22031 & n22032 ) ;
  assign n22034 = n22006 | n22030 ;
  assign n22035 = n22005 & ~n22030 ;
  assign n22036 = ( n22007 & n22034 ) | ( n22007 & ~n22035 ) | ( n22034 & ~n22035 ) ;
  assign n22037 = ~n22033 & n22036 ;
  assign n22038 = n21424 | n21445 ;
  assign n22039 = ( n21424 & n21428 ) | ( n21424 & n22038 ) | ( n21428 & n22038 ) ;
  assign n22040 = n22037 | n22039 ;
  assign n22041 = n22037 & n22039 ;
  assign n22042 = n22040 & ~n22041 ;
  assign n22043 = x91 & n8724 ;
  assign n22044 = x90 & n8719 ;
  assign n22045 = x89 & ~n8718 ;
  assign n22046 = n9149 & n22045 ;
  assign n22047 = n22044 | n22046 ;
  assign n22048 = n22043 | n22047 ;
  assign n22049 = n8727 | n22043 ;
  assign n22050 = n22047 | n22049 ;
  assign n22051 = ( n3768 & n22048 ) | ( n3768 & n22050 ) | ( n22048 & n22050 ) ;
  assign n22052 = x44 & n22050 ;
  assign n22053 = x44 & n22043 ;
  assign n22054 = ( x44 & n22047 ) | ( x44 & n22053 ) | ( n22047 & n22053 ) ;
  assign n22055 = ( n3768 & n22052 ) | ( n3768 & n22054 ) | ( n22052 & n22054 ) ;
  assign n22056 = x44 & ~n22054 ;
  assign n22057 = x44 & ~n22050 ;
  assign n22058 = ( ~n3768 & n22056 ) | ( ~n3768 & n22057 ) | ( n22056 & n22057 ) ;
  assign n22059 = ( n22051 & ~n22055 ) | ( n22051 & n22058 ) | ( ~n22055 & n22058 ) ;
  assign n22060 = n22042 & n22059 ;
  assign n22061 = n22042 & ~n22060 ;
  assign n22062 = ~n22042 & n22059 ;
  assign n22063 = n22061 | n22062 ;
  assign n22064 = ( n21451 & n21452 ) | ( n21451 & n21472 ) | ( n21452 & n21472 ) ;
  assign n22065 = n22063 | n22064 ;
  assign n22066 = n22063 & n22064 ;
  assign n22067 = n22065 & ~n22066 ;
  assign n22068 = x94 & n7566 ;
  assign n22069 = x93 & n7561 ;
  assign n22070 = x92 & ~n7560 ;
  assign n22071 = n7953 & n22070 ;
  assign n22072 = n22069 | n22071 ;
  assign n22073 = n22068 | n22072 ;
  assign n22074 = n7569 | n22068 ;
  assign n22075 = n22072 | n22074 ;
  assign n22076 = ( n4583 & n22073 ) | ( n4583 & n22075 ) | ( n22073 & n22075 ) ;
  assign n22077 = x41 & n22075 ;
  assign n22078 = x41 & n22068 ;
  assign n22079 = ( x41 & n22072 ) | ( x41 & n22078 ) | ( n22072 & n22078 ) ;
  assign n22080 = ( n4583 & n22077 ) | ( n4583 & n22079 ) | ( n22077 & n22079 ) ;
  assign n22081 = x41 & ~n22079 ;
  assign n22082 = x41 & ~n22075 ;
  assign n22083 = ( ~n4583 & n22081 ) | ( ~n4583 & n22082 ) | ( n22081 & n22082 ) ;
  assign n22084 = ( n22076 & ~n22080 ) | ( n22076 & n22083 ) | ( ~n22080 & n22083 ) ;
  assign n22085 = n22067 & n22084 ;
  assign n22086 = n22067 | n22084 ;
  assign n22087 = ~n22085 & n22086 ;
  assign n22088 = n21478 | n21496 ;
  assign n22089 = ( n21478 & n21479 ) | ( n21478 & n22088 ) | ( n21479 & n22088 ) ;
  assign n22090 = n22087 & ~n22089 ;
  assign n22091 = ~n22087 & n22089 ;
  assign n22092 = n22090 | n22091 ;
  assign n22093 = x97 & n6536 ;
  assign n22094 = x96 & n6531 ;
  assign n22095 = x95 & ~n6530 ;
  assign n22096 = n6871 & n22095 ;
  assign n22097 = n22094 | n22096 ;
  assign n22098 = n22093 | n22097 ;
  assign n22099 = n6539 | n22093 ;
  assign n22100 = n22097 | n22099 ;
  assign n22101 = ( n5505 & n22098 ) | ( n5505 & n22100 ) | ( n22098 & n22100 ) ;
  assign n22102 = x38 & n22100 ;
  assign n22103 = x38 & n22093 ;
  assign n22104 = ( x38 & n22097 ) | ( x38 & n22103 ) | ( n22097 & n22103 ) ;
  assign n22105 = ( n5505 & n22102 ) | ( n5505 & n22104 ) | ( n22102 & n22104 ) ;
  assign n22106 = x38 & ~n22104 ;
  assign n22107 = x38 & ~n22100 ;
  assign n22108 = ( ~n5505 & n22106 ) | ( ~n5505 & n22107 ) | ( n22106 & n22107 ) ;
  assign n22109 = ( n22101 & ~n22105 ) | ( n22101 & n22108 ) | ( ~n22105 & n22108 ) ;
  assign n22110 = n22092 & n22109 ;
  assign n22111 = n22092 | n22109 ;
  assign n22112 = ~n22110 & n22111 ;
  assign n22113 = n21504 | n21525 ;
  assign n22114 = ( n21505 & n21525 ) | ( n21505 & n22113 ) | ( n21525 & n22113 ) ;
  assign n22115 = ( n21507 & n21508 ) | ( n21507 & n22114 ) | ( n21508 & n22114 ) ;
  assign n22116 = ~n22112 & n22115 ;
  assign n22117 = n22112 & ~n22115 ;
  assign n22118 = n22116 | n22117 ;
  assign n22119 = x100 & n5554 ;
  assign n22120 = x99 & n5549 ;
  assign n22121 = x98 & ~n5548 ;
  assign n22122 = n5893 & n22121 ;
  assign n22123 = n22120 | n22122 ;
  assign n22124 = n22119 | n22123 ;
  assign n22125 = n5557 | n22119 ;
  assign n22126 = n22123 | n22125 ;
  assign n22127 = ( n6483 & n22124 ) | ( n6483 & n22126 ) | ( n22124 & n22126 ) ;
  assign n22128 = x35 & n22126 ;
  assign n22129 = x35 & n22119 ;
  assign n22130 = ( x35 & n22123 ) | ( x35 & n22129 ) | ( n22123 & n22129 ) ;
  assign n22131 = ( n6483 & n22128 ) | ( n6483 & n22130 ) | ( n22128 & n22130 ) ;
  assign n22132 = x35 & ~n22130 ;
  assign n22133 = x35 & ~n22126 ;
  assign n22134 = ( ~n6483 & n22132 ) | ( ~n6483 & n22133 ) | ( n22132 & n22133 ) ;
  assign n22135 = ( n22127 & ~n22131 ) | ( n22127 & n22134 ) | ( ~n22131 & n22134 ) ;
  assign n22136 = n22118 & n22135 ;
  assign n22137 = n22118 | n22135 ;
  assign n22138 = ~n22136 & n22137 ;
  assign n22139 = n21528 | n21551 ;
  assign n22140 = ( n21531 & n21551 ) | ( n21531 & n22139 ) | ( n21551 & n22139 ) ;
  assign n22141 = ( n21532 & n21534 ) | ( n21532 & n22140 ) | ( n21534 & n22140 ) ;
  assign n22142 = n22138 | n22141 ;
  assign n22143 = n22138 & n22141 ;
  assign n22144 = n22142 & ~n22143 ;
  assign n22145 = x103 & n4631 ;
  assign n22146 = x102 & n4626 ;
  assign n22147 = x101 & ~n4625 ;
  assign n22148 = n4943 & n22147 ;
  assign n22149 = n22146 | n22148 ;
  assign n22150 = n22145 | n22149 ;
  assign n22151 = n4634 | n22145 ;
  assign n22152 = n22149 | n22151 ;
  assign n22153 = ( n7529 & n22150 ) | ( n7529 & n22152 ) | ( n22150 & n22152 ) ;
  assign n22154 = x32 & n22152 ;
  assign n22155 = x32 & n22145 ;
  assign n22156 = ( x32 & n22149 ) | ( x32 & n22155 ) | ( n22149 & n22155 ) ;
  assign n22157 = ( n7529 & n22154 ) | ( n7529 & n22156 ) | ( n22154 & n22156 ) ;
  assign n22158 = x32 & ~n22156 ;
  assign n22159 = x32 & ~n22152 ;
  assign n22160 = ( ~n7529 & n22158 ) | ( ~n7529 & n22159 ) | ( n22158 & n22159 ) ;
  assign n22161 = ( n22153 & ~n22157 ) | ( n22153 & n22160 ) | ( ~n22157 & n22160 ) ;
  assign n22162 = n21275 | n21554 ;
  assign n22163 = ( n21281 & n21554 ) | ( n21281 & n22162 ) | ( n21554 & n22162 ) ;
  assign n22164 = n22161 | n22163 ;
  assign n22165 = n21282 | n22161 ;
  assign n22166 = ( n21284 & n22164 ) | ( n21284 & n22165 ) | ( n22164 & n22165 ) ;
  assign n22167 = n22161 & n22163 ;
  assign n22168 = n21282 & n22161 ;
  assign n22169 = ( n21284 & n22167 ) | ( n21284 & n22168 ) | ( n22167 & n22168 ) ;
  assign n22170 = n22166 & ~n22169 ;
  assign n22171 = n22144 & n22170 ;
  assign n22172 = n22144 | n22170 ;
  assign n22173 = ~n22171 & n22172 ;
  assign n22174 = n21862 & n22173 ;
  assign n22175 = n21862 | n22173 ;
  assign n22176 = ~n22174 & n22175 ;
  assign n22177 = n21585 | n21591 ;
  assign n22178 = n21563 | n21585 ;
  assign n22179 = ( n21586 & n22177 ) | ( n21586 & n22178 ) | ( n22177 & n22178 ) ;
  assign n22180 = ( n21841 & n22176 ) | ( n21841 & ~n22179 ) | ( n22176 & ~n22179 ) ;
  assign n22181 = ( ~n22176 & n22179 ) | ( ~n22176 & n22180 ) | ( n22179 & n22180 ) ;
  assign n22182 = ( ~n21841 & n22180 ) | ( ~n21841 & n22181 ) | ( n22180 & n22181 ) ;
  assign n22183 = ~n21824 & n22182 ;
  assign n22184 = n21820 | n22180 ;
  assign n22185 = ~n21820 & n21841 ;
  assign n22186 = ( n22181 & n22184 ) | ( n22181 & ~n22185 ) | ( n22184 & ~n22185 ) ;
  assign n22187 = ( n21821 & n22182 ) | ( n21821 & n22186 ) | ( n22182 & n22186 ) ;
  assign n22188 = n21822 & ~n22187 ;
  assign n22189 = n22183 | n22188 ;
  assign n22190 = n21803 & ~n22189 ;
  assign n22191 = n21803 | n22189 ;
  assign n22192 = ( ~n21803 & n22190 ) | ( ~n21803 & n22191 ) | ( n22190 & n22191 ) ;
  assign n22193 = ~n21748 & n21763 ;
  assign n22194 = ~n21192 & n21763 ;
  assign n22195 = ( ~n21194 & n22193 ) | ( ~n21194 & n22194 ) | ( n22193 & n22194 ) ;
  assign n22196 = n22192 & n22195 ;
  assign n22197 = ( n21767 & n22192 ) | ( n21767 & n22196 ) | ( n22192 & n22196 ) ;
  assign n22198 = n22192 | n22195 ;
  assign n22199 = n21767 | n22198 ;
  assign n22200 = ~n22197 & n22199 ;
  assign n22201 = n21746 & ~n22200 ;
  assign n22202 = n21746 | n22200 ;
  assign n22203 = ( ~n21746 & n22201 ) | ( ~n21746 & n22202 ) | ( n22201 & n22202 ) ;
  assign n22204 = ~n21707 & n22203 ;
  assign n22205 = ( n21157 & n21158 ) | ( n21157 & n21635 ) | ( n21158 & n21635 ) ;
  assign n22206 = n21700 | n22203 ;
  assign n22207 = ( n22203 & n22205 ) | ( n22203 & n22206 ) | ( n22205 & n22206 ) ;
  assign n22208 = n21703 & ~n22207 ;
  assign n22209 = n22204 | n22208 ;
  assign n22211 = n21133 | n21637 ;
  assign n22213 = ( n21683 & n22209 ) | ( n21683 & ~n22211 ) | ( n22209 & ~n22211 ) ;
  assign n22214 = ( ~n21134 & n21683 ) | ( ~n21134 & n22209 ) | ( n21683 & n22209 ) ;
  assign n22215 = ( ~n22210 & n22213 ) | ( ~n22210 & n22214 ) | ( n22213 & n22214 ) ;
  assign n22212 = ( n21134 & n22210 ) | ( n21134 & n22211 ) | ( n22210 & n22211 ) ;
  assign n22216 = ( ~n22209 & n22212 ) | ( ~n22209 & n22215 ) | ( n22212 & n22215 ) ;
  assign n22217 = ( ~n21683 & n22215 ) | ( ~n21683 & n22216 ) | ( n22215 & n22216 ) ;
  assign n22218 = n21106 & n22217 ;
  assign n22219 = ( n21652 & n22217 ) | ( n21652 & n22218 ) | ( n22217 & n22218 ) ;
  assign n22220 = n21106 | n22217 ;
  assign n22221 = n21652 | n22220 ;
  assign n22222 = ~n22219 & n22221 ;
  assign n22223 = n21658 | n21661 ;
  assign n22224 = n21659 | n22223 ;
  assign n22225 = ( n21658 & n21663 ) | ( n21658 & n22224 ) | ( n21663 & n22224 ) ;
  assign n22226 = n22222 | n22225 ;
  assign n22227 = n22222 & n22224 ;
  assign n22228 = n21658 & n22222 ;
  assign n22229 = ( n21663 & n22227 ) | ( n21663 & n22228 ) | ( n22227 & n22228 ) ;
  assign n22230 = n22226 & ~n22229 ;
  assign n22759 = n21127 & n21683 ;
  assign n22760 = n21128 & n21683 ;
  assign n22761 = n21129 & n21683 ;
  assign n22762 = ( n20448 & n22760 ) | ( n20448 & n22761 ) | ( n22760 & n22761 ) ;
  assign n22763 = ( n21050 & n22759 ) | ( n21050 & n22762 ) | ( n22759 & n22762 ) ;
  assign n22764 = ( n21022 & n22759 ) | ( n21022 & n22762 ) | ( n22759 & n22762 ) ;
  assign n22765 = ( n21047 & n22763 ) | ( n21047 & n22764 ) | ( n22763 & n22764 ) ;
  assign n22766 = ( n21645 & n21683 ) | ( n21645 & n22765 ) | ( n21683 & n22765 ) ;
  assign n22767 = ( n21637 & n21683 ) | ( n21637 & n22765 ) | ( n21683 & n22765 ) ;
  assign n22768 = ( n21134 & n22766 ) | ( n21134 & n22767 ) | ( n22766 & n22767 ) ;
  assign n22769 = n22212 & ~n22768 ;
  assign n22770 = n21683 & ~n22762 ;
  assign n22771 = n21683 & ~n22759 ;
  assign n22772 = ( ~n21051 & n22770 ) | ( ~n21051 & n22771 ) | ( n22770 & n22771 ) ;
  assign n22773 = ~n21645 & n22772 ;
  assign n22774 = ~n21637 & n22770 ;
  assign n22775 = ~n21637 & n22771 ;
  assign n22776 = ( ~n21051 & n22774 ) | ( ~n21051 & n22775 ) | ( n22774 & n22775 ) ;
  assign n22777 = n22209 & ~n22776 ;
  assign n22778 = n21134 & n22209 ;
  assign n22779 = ( ~n22773 & n22777 ) | ( ~n22773 & n22778 ) | ( n22777 & n22778 ) ;
  assign n22780 = ( n22209 & n22768 ) | ( n22209 & ~n22779 ) | ( n22768 & ~n22779 ) ;
  assign n22781 = n22209 | n22768 ;
  assign n22782 = ( n22769 & n22780 ) | ( n22769 & n22781 ) | ( n22780 & n22781 ) ;
  assign n22231 = x116 & n1859 ;
  assign n22232 = x115 & n1854 ;
  assign n22233 = x114 & ~n1853 ;
  assign n22234 = n2037 & n22233 ;
  assign n22235 = n22232 | n22234 ;
  assign n22236 = n22231 | n22235 ;
  assign n22237 = n1862 | n22231 ;
  assign n22238 = n22235 | n22237 ;
  assign n22239 = ( ~n13040 & n22236 ) | ( ~n13040 & n22238 ) | ( n22236 & n22238 ) ;
  assign n22240 = n22236 & n22238 ;
  assign n22241 = ( n13022 & n22239 ) | ( n13022 & n22240 ) | ( n22239 & n22240 ) ;
  assign n22242 = x20 & n22241 ;
  assign n22243 = x20 & ~n22241 ;
  assign n22244 = ( n22241 & ~n22242 ) | ( n22241 & n22243 ) | ( ~n22242 & n22243 ) ;
  assign n22245 = n22187 & n22244 ;
  assign n22246 = n21823 & n22244 ;
  assign n22247 = ( n21824 & n22245 ) | ( n21824 & n22246 ) | ( n22245 & n22246 ) ;
  assign n22248 = n22187 | n22244 ;
  assign n22249 = n21823 | n22244 ;
  assign n22250 = ( n21824 & n22248 ) | ( n21824 & n22249 ) | ( n22248 & n22249 ) ;
  assign n22251 = ~n22247 & n22250 ;
  assign n22252 = x113 & n2429 ;
  assign n22253 = x112 & n2424 ;
  assign n22254 = x111 & ~n2423 ;
  assign n22255 = n2631 & n22254 ;
  assign n22256 = n22253 | n22255 ;
  assign n22257 = n22252 | n22256 ;
  assign n22258 = n2432 | n22252 ;
  assign n22259 = n22256 | n22258 ;
  assign n22260 = ( ~n11642 & n22257 ) | ( ~n11642 & n22259 ) | ( n22257 & n22259 ) ;
  assign n22261 = n22257 & n22259 ;
  assign n22262 = ( n11626 & n22260 ) | ( n11626 & n22261 ) | ( n22260 & n22261 ) ;
  assign n22263 = x23 & n22262 ;
  assign n22264 = x23 & ~n22262 ;
  assign n22265 = ( n22262 & ~n22263 ) | ( n22262 & n22264 ) | ( ~n22263 & n22264 ) ;
  assign n22266 = n21581 & n21841 ;
  assign n22267 = n21583 & n21841 ;
  assign n22268 = n21582 & n21841 ;
  assign n22269 = ( n20324 & n22267 ) | ( n20324 & n22268 ) | ( n22267 & n22268 ) ;
  assign n22270 = ( n20962 & n22266 ) | ( n20962 & n22269 ) | ( n22266 & n22269 ) ;
  assign n22271 = ( n21591 & n21841 ) | ( n21591 & n22270 ) | ( n21841 & n22270 ) ;
  assign n22272 = ( n21563 & n21841 ) | ( n21563 & n22270 ) | ( n21841 & n22270 ) ;
  assign n22273 = ( n21586 & n22271 ) | ( n21586 & n22272 ) | ( n22271 & n22272 ) ;
  assign n22274 = n22179 & ~n22273 ;
  assign n22275 = n21841 & ~n22269 ;
  assign n22276 = n21841 & ~n22266 ;
  assign n22277 = ( ~n20962 & n22275 ) | ( ~n20962 & n22276 ) | ( n22275 & n22276 ) ;
  assign n22278 = ~n21591 & n22277 ;
  assign n22279 = ~n21563 & n22277 ;
  assign n22280 = ( ~n21586 & n22278 ) | ( ~n21586 & n22279 ) | ( n22278 & n22279 ) ;
  assign n22281 = n22176 & n22280 ;
  assign n22282 = ( n22176 & n22274 ) | ( n22176 & n22281 ) | ( n22274 & n22281 ) ;
  assign n22285 = x109 & n3080 ;
  assign n22286 = x108 & ~n3079 ;
  assign n22287 = n3309 & n22286 ;
  assign n22288 = n22285 | n22287 ;
  assign n22284 = x110 & n3085 ;
  assign n22290 = n3088 | n22284 ;
  assign n22291 = n22288 | n22290 ;
  assign n22289 = n22284 | n22288 ;
  assign n22292 = n22289 & n22291 ;
  assign n22293 = ( n10330 & n22291 ) | ( n10330 & n22292 ) | ( n22291 & n22292 ) ;
  assign n22294 = x26 & n22292 ;
  assign n22295 = x26 & n22291 ;
  assign n22296 = ( n10330 & n22294 ) | ( n10330 & n22295 ) | ( n22294 & n22295 ) ;
  assign n22297 = x26 & ~n22292 ;
  assign n22298 = x26 & ~n22291 ;
  assign n22299 = ( ~n10330 & n22297 ) | ( ~n10330 & n22298 ) | ( n22297 & n22298 ) ;
  assign n22300 = ( n22293 & ~n22296 ) | ( n22293 & n22299 ) | ( ~n22296 & n22299 ) ;
  assign n22301 = n21858 | n22173 ;
  assign n22302 = ( n21859 & n22173 ) | ( n21859 & n22301 ) | ( n22173 & n22301 ) ;
  assign n22303 = n22300 & n22302 ;
  assign n22304 = n21861 & n22300 ;
  assign n22305 = ( n21862 & n22303 ) | ( n21862 & n22304 ) | ( n22303 & n22304 ) ;
  assign n22306 = n22300 | n22302 ;
  assign n22307 = n21861 | n22300 ;
  assign n22308 = ( n21862 & n22306 ) | ( n21862 & n22307 ) | ( n22306 & n22307 ) ;
  assign n22309 = ~n22305 & n22308 ;
  assign n22310 = x104 & n4631 ;
  assign n22311 = x103 & n4626 ;
  assign n22312 = x102 & ~n4625 ;
  assign n22313 = n4943 & n22312 ;
  assign n22314 = n22311 | n22313 ;
  assign n22315 = n22310 | n22314 ;
  assign n22316 = n4634 | n22310 ;
  assign n22317 = n22314 | n22316 ;
  assign n22318 = ( n7911 & n22315 ) | ( n7911 & n22317 ) | ( n22315 & n22317 ) ;
  assign n22319 = x32 & n22317 ;
  assign n22320 = x32 & n22310 ;
  assign n22321 = ( x32 & n22314 ) | ( x32 & n22320 ) | ( n22314 & n22320 ) ;
  assign n22322 = ( n7911 & n22319 ) | ( n7911 & n22321 ) | ( n22319 & n22321 ) ;
  assign n22323 = x32 & ~n22321 ;
  assign n22324 = x32 & ~n22317 ;
  assign n22325 = ( ~n7911 & n22323 ) | ( ~n7911 & n22324 ) | ( n22323 & n22324 ) ;
  assign n22326 = ( n22318 & ~n22322 ) | ( n22318 & n22325 ) | ( ~n22322 & n22325 ) ;
  assign n22327 = n22136 | n22138 ;
  assign n22328 = ( n22136 & n22141 ) | ( n22136 & n22327 ) | ( n22141 & n22327 ) ;
  assign n22329 = n22326 | n22328 ;
  assign n22330 = n22326 & n22328 ;
  assign n22331 = n22329 & ~n22330 ;
  assign n22332 = n22112 & n22115 ;
  assign n22333 = n21922 | n21930 ;
  assign n22334 = x74 & n17146 ;
  assign n22335 = x73 & n17141 ;
  assign n22336 = x72 & ~n17140 ;
  assign n22337 = n17724 & n22336 ;
  assign n22338 = n22335 | n22337 ;
  assign n22339 = n22334 | n22338 ;
  assign n22340 = n17149 | n22334 ;
  assign n22341 = n22338 | n22340 ;
  assign n22342 = n22339 & n22341 ;
  assign n22343 = x62 & n22342 ;
  assign n22344 = x62 & n22341 ;
  assign n22345 = ( n710 & n22343 ) | ( n710 & n22344 ) | ( n22343 & n22344 ) ;
  assign n22346 = x62 & ~n22345 ;
  assign n22347 = x71 & n18290 ;
  assign n22348 = x63 & x70 ;
  assign n22349 = ~n18290 & n22348 ;
  assign n22350 = n22347 | n22349 ;
  assign n22351 = ( x2 & x5 ) | ( x2 & ~n21866 ) | ( x5 & ~n21866 ) ;
  assign n22352 = n22350 | n22351 ;
  assign n22353 = n22350 & n22351 ;
  assign n22354 = n22352 & ~n22353 ;
  assign n22355 = ~n22345 & n22354 ;
  assign n22356 = n22342 & n22354 ;
  assign n22357 = n22341 & n22354 ;
  assign n22358 = ( n710 & n22356 ) | ( n710 & n22357 ) | ( n22356 & n22357 ) ;
  assign n22359 = ( n22346 & n22355 ) | ( n22346 & n22358 ) | ( n22355 & n22358 ) ;
  assign n22360 = n22345 & ~n22354 ;
  assign n22361 = n22342 | n22354 ;
  assign n22362 = n22341 | n22354 ;
  assign n22363 = ( n710 & n22361 ) | ( n710 & n22362 ) | ( n22361 & n22362 ) ;
  assign n22364 = ( n22346 & ~n22360 ) | ( n22346 & n22363 ) | ( ~n22360 & n22363 ) ;
  assign n22365 = ~n22359 & n22364 ;
  assign n22366 = n21879 | n21901 ;
  assign n22367 = ( n21879 & n21885 ) | ( n21879 & n22366 ) | ( n21885 & n22366 ) ;
  assign n22368 = n22365 & n22367 ;
  assign n22369 = n22365 | n22367 ;
  assign n22370 = ~n22368 & n22369 ;
  assign n22371 = x77 & n15552 ;
  assign n22372 = x76 & n15547 ;
  assign n22373 = x75 & ~n15546 ;
  assign n22374 = n16123 & n22373 ;
  assign n22375 = n22372 | n22374 ;
  assign n22376 = n22371 | n22375 ;
  assign n22377 = n15555 | n22371 ;
  assign n22378 = n22375 | n22377 ;
  assign n22379 = ( n1059 & n22376 ) | ( n1059 & n22378 ) | ( n22376 & n22378 ) ;
  assign n22380 = x59 & n22378 ;
  assign n22381 = x59 & n22371 ;
  assign n22382 = ( x59 & n22375 ) | ( x59 & n22381 ) | ( n22375 & n22381 ) ;
  assign n22383 = ( n1059 & n22380 ) | ( n1059 & n22382 ) | ( n22380 & n22382 ) ;
  assign n22384 = x59 & ~n22382 ;
  assign n22385 = x59 & ~n22378 ;
  assign n22386 = ( ~n1059 & n22384 ) | ( ~n1059 & n22385 ) | ( n22384 & n22385 ) ;
  assign n22387 = ( n22379 & ~n22383 ) | ( n22379 & n22386 ) | ( ~n22383 & n22386 ) ;
  assign n22388 = n22370 & ~n22387 ;
  assign n22389 = n22370 | n22387 ;
  assign n22390 = ( ~n22370 & n22388 ) | ( ~n22370 & n22389 ) | ( n22388 & n22389 ) ;
  assign n22391 = n22333 | n22390 ;
  assign n22392 = n22333 & n22390 ;
  assign n22393 = n22391 & ~n22392 ;
  assign n22394 = x80 & n14045 ;
  assign n22395 = x79 & n14040 ;
  assign n22396 = x78 & ~n14039 ;
  assign n22397 = n14552 & n22396 ;
  assign n22398 = n22395 | n22397 ;
  assign n22399 = n22394 | n22398 ;
  assign n22400 = n14048 | n22394 ;
  assign n22401 = n22398 | n22400 ;
  assign n22402 = ( n1499 & n22399 ) | ( n1499 & n22401 ) | ( n22399 & n22401 ) ;
  assign n22403 = x56 & n22401 ;
  assign n22404 = x56 & n22394 ;
  assign n22405 = ( x56 & n22398 ) | ( x56 & n22404 ) | ( n22398 & n22404 ) ;
  assign n22406 = ( n1499 & n22403 ) | ( n1499 & n22405 ) | ( n22403 & n22405 ) ;
  assign n22407 = x56 & ~n22405 ;
  assign n22408 = x56 & ~n22401 ;
  assign n22409 = ( ~n1499 & n22407 ) | ( ~n1499 & n22408 ) | ( n22407 & n22408 ) ;
  assign n22410 = ( n22402 & ~n22406 ) | ( n22402 & n22409 ) | ( ~n22406 & n22409 ) ;
  assign n22411 = ~n22393 & n22410 ;
  assign n22412 = n22390 | n22410 ;
  assign n22413 = ( n22333 & n22410 ) | ( n22333 & n22412 ) | ( n22410 & n22412 ) ;
  assign n22414 = n22391 & ~n22413 ;
  assign n22415 = n22411 | n22414 ;
  assign n22416 = n21951 | n21958 ;
  assign n22417 = n22415 | n22416 ;
  assign n22418 = n22415 & n22416 ;
  assign n22419 = n22417 & ~n22418 ;
  assign n22420 = x83 & n12574 ;
  assign n22421 = x82 & n12569 ;
  assign n22422 = x81 & ~n12568 ;
  assign n22423 = n13076 & n22422 ;
  assign n22424 = n22421 | n22423 ;
  assign n22425 = n22420 | n22424 ;
  assign n22426 = n12577 | n22420 ;
  assign n22427 = n22424 | n22426 ;
  assign n22428 = ( n2009 & n22425 ) | ( n2009 & n22427 ) | ( n22425 & n22427 ) ;
  assign n22429 = x53 & n22427 ;
  assign n22430 = x53 & n22420 ;
  assign n22431 = ( x53 & n22424 ) | ( x53 & n22430 ) | ( n22424 & n22430 ) ;
  assign n22432 = ( n2009 & n22429 ) | ( n2009 & n22431 ) | ( n22429 & n22431 ) ;
  assign n22433 = x53 & ~n22431 ;
  assign n22434 = x53 & ~n22427 ;
  assign n22435 = ( ~n2009 & n22433 ) | ( ~n2009 & n22434 ) | ( n22433 & n22434 ) ;
  assign n22436 = ( n22428 & ~n22432 ) | ( n22428 & n22435 ) | ( ~n22432 & n22435 ) ;
  assign n22437 = ~n22419 & n22436 ;
  assign n22438 = n22418 | n22436 ;
  assign n22439 = n22417 & ~n22438 ;
  assign n22440 = n22437 | n22439 ;
  assign n22441 = n21979 | n21983 ;
  assign n22442 = ( n21979 & n21982 ) | ( n21979 & n22441 ) | ( n21982 & n22441 ) ;
  assign n22443 = n22440 | n22442 ;
  assign n22444 = n22440 & n22442 ;
  assign n22445 = n22443 & ~n22444 ;
  assign n22446 = x86 & n11205 ;
  assign n22447 = x85 & n11200 ;
  assign n22448 = x84 & ~n11199 ;
  assign n22449 = n11679 & n22448 ;
  assign n22450 = n22447 | n22449 ;
  assign n22451 = n22446 | n22450 ;
  assign n22452 = n11208 | n22446 ;
  assign n22453 = n22450 | n22452 ;
  assign n22454 = ( n2606 & n22451 ) | ( n2606 & n22453 ) | ( n22451 & n22453 ) ;
  assign n22455 = x50 & n22453 ;
  assign n22456 = x50 & n22446 ;
  assign n22457 = ( x50 & n22450 ) | ( x50 & n22456 ) | ( n22450 & n22456 ) ;
  assign n22458 = ( n2606 & n22455 ) | ( n2606 & n22457 ) | ( n22455 & n22457 ) ;
  assign n22459 = x50 & ~n22457 ;
  assign n22460 = x50 & ~n22453 ;
  assign n22461 = ( ~n2606 & n22459 ) | ( ~n2606 & n22460 ) | ( n22459 & n22460 ) ;
  assign n22462 = ( n22454 & ~n22458 ) | ( n22454 & n22461 ) | ( ~n22458 & n22461 ) ;
  assign n22463 = ~n22445 & n22462 ;
  assign n22464 = n22444 | n22462 ;
  assign n22465 = n22443 & ~n22464 ;
  assign n22466 = n22463 | n22465 ;
  assign n22467 = n21986 & n22003 ;
  assign n22468 = n21986 & ~n22467 ;
  assign n22469 = ~n21986 & n22003 ;
  assign n22470 = n22005 & ~n22469 ;
  assign n22471 = ~n22468 & n22470 ;
  assign n22472 = ( n22005 & n22467 ) | ( n22005 & ~n22471 ) | ( n22467 & ~n22471 ) ;
  assign n22473 = n22466 | n22472 ;
  assign n22474 = n22466 & n22472 ;
  assign n22475 = n22473 & ~n22474 ;
  assign n22476 = x89 & n9933 ;
  assign n22477 = x88 & n9928 ;
  assign n22478 = x87 & ~n9927 ;
  assign n22479 = n10379 & n22478 ;
  assign n22480 = n22477 | n22479 ;
  assign n22481 = n22476 | n22480 ;
  assign n22482 = n9936 | n22476 ;
  assign n22483 = n22480 | n22482 ;
  assign n22484 = ( n3282 & n22481 ) | ( n3282 & n22483 ) | ( n22481 & n22483 ) ;
  assign n22485 = x47 & n22483 ;
  assign n22486 = x47 & n22476 ;
  assign n22487 = ( x47 & n22480 ) | ( x47 & n22486 ) | ( n22480 & n22486 ) ;
  assign n22488 = ( n3282 & n22485 ) | ( n3282 & n22487 ) | ( n22485 & n22487 ) ;
  assign n22489 = x47 & ~n22487 ;
  assign n22490 = x47 & ~n22483 ;
  assign n22491 = ( ~n3282 & n22489 ) | ( ~n3282 & n22490 ) | ( n22489 & n22490 ) ;
  assign n22492 = ( n22484 & ~n22488 ) | ( n22484 & n22491 ) | ( ~n22488 & n22491 ) ;
  assign n22493 = ~n22475 & n22492 ;
  assign n22494 = n22033 | n22037 ;
  assign n22495 = ( n22033 & n22039 ) | ( n22033 & n22494 ) | ( n22039 & n22494 ) ;
  assign n22496 = n22466 | n22492 ;
  assign n22497 = ( n22472 & n22492 ) | ( n22472 & n22496 ) | ( n22492 & n22496 ) ;
  assign n22498 = n22473 & ~n22497 ;
  assign n22499 = n22495 & n22498 ;
  assign n22500 = ( n22493 & n22495 ) | ( n22493 & n22499 ) | ( n22495 & n22499 ) ;
  assign n22501 = n22495 | n22498 ;
  assign n22502 = n22493 | n22501 ;
  assign n22503 = ~n22500 & n22502 ;
  assign n22504 = x92 & n8724 ;
  assign n22505 = x91 & n8719 ;
  assign n22506 = x90 & ~n8718 ;
  assign n22507 = n9149 & n22506 ;
  assign n22508 = n22505 | n22507 ;
  assign n22509 = n22504 | n22508 ;
  assign n22510 = n8727 | n22504 ;
  assign n22511 = n22508 | n22510 ;
  assign n22512 = ( n4040 & n22509 ) | ( n4040 & n22511 ) | ( n22509 & n22511 ) ;
  assign n22513 = x44 & n22511 ;
  assign n22514 = x44 & n22504 ;
  assign n22515 = ( x44 & n22508 ) | ( x44 & n22514 ) | ( n22508 & n22514 ) ;
  assign n22516 = ( n4040 & n22513 ) | ( n4040 & n22515 ) | ( n22513 & n22515 ) ;
  assign n22517 = x44 & ~n22515 ;
  assign n22518 = x44 & ~n22511 ;
  assign n22519 = ( ~n4040 & n22517 ) | ( ~n4040 & n22518 ) | ( n22517 & n22518 ) ;
  assign n22520 = ( n22512 & ~n22516 ) | ( n22512 & n22519 ) | ( ~n22516 & n22519 ) ;
  assign n22521 = n22503 & ~n22520 ;
  assign n22522 = n22503 | n22520 ;
  assign n22523 = ( ~n22503 & n22521 ) | ( ~n22503 & n22522 ) | ( n22521 & n22522 ) ;
  assign n22524 = n21472 | n22060 ;
  assign n22525 = n21451 | n22060 ;
  assign n22526 = ( n21452 & n22524 ) | ( n21452 & n22525 ) | ( n22524 & n22525 ) ;
  assign n22527 = ( n22060 & n22063 ) | ( n22060 & n22526 ) | ( n22063 & n22526 ) ;
  assign n22528 = n22523 | n22527 ;
  assign n22529 = n22523 & n22527 ;
  assign n22530 = n22528 & ~n22529 ;
  assign n22531 = x95 & n7566 ;
  assign n22532 = x94 & n7561 ;
  assign n22533 = x93 & ~n7560 ;
  assign n22534 = n7953 & n22533 ;
  assign n22535 = n22532 | n22534 ;
  assign n22536 = n22531 | n22535 ;
  assign n22537 = n7569 | n22531 ;
  assign n22538 = n22535 | n22537 ;
  assign n22539 = ( n4897 & n22536 ) | ( n4897 & n22538 ) | ( n22536 & n22538 ) ;
  assign n22540 = x41 & n22538 ;
  assign n22541 = x41 & n22531 ;
  assign n22542 = ( x41 & n22535 ) | ( x41 & n22541 ) | ( n22535 & n22541 ) ;
  assign n22543 = ( n4897 & n22540 ) | ( n4897 & n22542 ) | ( n22540 & n22542 ) ;
  assign n22544 = x41 & ~n22542 ;
  assign n22545 = x41 & ~n22538 ;
  assign n22546 = ( ~n4897 & n22544 ) | ( ~n4897 & n22545 ) | ( n22544 & n22545 ) ;
  assign n22547 = ( n22539 & ~n22543 ) | ( n22539 & n22546 ) | ( ~n22543 & n22546 ) ;
  assign n22548 = n22530 | n22547 ;
  assign n22549 = n22530 & n22547 ;
  assign n22550 = n22548 & ~n22549 ;
  assign n22551 = n22085 | n22087 ;
  assign n22552 = ( n22085 & n22089 ) | ( n22085 & n22551 ) | ( n22089 & n22551 ) ;
  assign n22553 = n22550 & n22552 ;
  assign n22554 = n22550 | n22552 ;
  assign n22555 = ~n22553 & n22554 ;
  assign n22556 = x98 & n6536 ;
  assign n22557 = x97 & n6531 ;
  assign n22558 = x96 & ~n6530 ;
  assign n22559 = n6871 & n22558 ;
  assign n22560 = n22557 | n22559 ;
  assign n22561 = n22556 | n22560 ;
  assign n22562 = n6539 | n22556 ;
  assign n22563 = n22560 | n22562 ;
  assign n22564 = ( ~n5850 & n22561 ) | ( ~n5850 & n22563 ) | ( n22561 & n22563 ) ;
  assign n22565 = n22561 & n22563 ;
  assign n22566 = ( n5834 & n22564 ) | ( n5834 & n22565 ) | ( n22564 & n22565 ) ;
  assign n22567 = x38 & n22563 ;
  assign n22568 = x38 & n22556 ;
  assign n22569 = ( x38 & n22560 ) | ( x38 & n22568 ) | ( n22560 & n22568 ) ;
  assign n22570 = ( ~n5850 & n22567 ) | ( ~n5850 & n22569 ) | ( n22567 & n22569 ) ;
  assign n22571 = n22567 & n22569 ;
  assign n22572 = ( n5834 & n22570 ) | ( n5834 & n22571 ) | ( n22570 & n22571 ) ;
  assign n22573 = x38 & ~n22569 ;
  assign n22574 = x38 & ~n22563 ;
  assign n22575 = ( n5850 & n22573 ) | ( n5850 & n22574 ) | ( n22573 & n22574 ) ;
  assign n22576 = n22573 | n22574 ;
  assign n22577 = ( ~n5834 & n22575 ) | ( ~n5834 & n22576 ) | ( n22575 & n22576 ) ;
  assign n22578 = ( n22566 & ~n22572 ) | ( n22566 & n22577 ) | ( ~n22572 & n22577 ) ;
  assign n22579 = n22555 & n22578 ;
  assign n22580 = n22555 | n22578 ;
  assign n22581 = ~n22579 & n22580 ;
  assign n22582 = n22110 & n22581 ;
  assign n22583 = ( n22332 & n22581 ) | ( n22332 & n22582 ) | ( n22581 & n22582 ) ;
  assign n22584 = n22110 | n22581 ;
  assign n22585 = n22332 | n22584 ;
  assign n22586 = ~n22583 & n22585 ;
  assign n22587 = x101 & n5554 ;
  assign n22588 = x100 & n5549 ;
  assign n22589 = x99 & ~n5548 ;
  assign n22590 = n5893 & n22589 ;
  assign n22591 = n22588 | n22590 ;
  assign n22592 = n22587 | n22591 ;
  assign n22593 = n5557 | n22587 ;
  assign n22594 = n22591 | n22593 ;
  assign n22595 = ( n6844 & n22592 ) | ( n6844 & n22594 ) | ( n22592 & n22594 ) ;
  assign n22596 = x35 & n22594 ;
  assign n22597 = x35 & n22587 ;
  assign n22598 = ( x35 & n22591 ) | ( x35 & n22597 ) | ( n22591 & n22597 ) ;
  assign n22599 = ( n6844 & n22596 ) | ( n6844 & n22598 ) | ( n22596 & n22598 ) ;
  assign n22600 = x35 & ~n22598 ;
  assign n22601 = x35 & ~n22594 ;
  assign n22602 = ( ~n6844 & n22600 ) | ( ~n6844 & n22601 ) | ( n22600 & n22601 ) ;
  assign n22603 = ( n22595 & ~n22599 ) | ( n22595 & n22602 ) | ( ~n22599 & n22602 ) ;
  assign n22604 = n22586 & ~n22603 ;
  assign n22605 = n22586 | n22603 ;
  assign n22606 = ( ~n22586 & n22604 ) | ( ~n22586 & n22605 ) | ( n22604 & n22605 ) ;
  assign n22607 = ~n22331 & n22606 ;
  assign n22608 = n22326 | n22606 ;
  assign n22609 = ( n22328 & n22606 ) | ( n22328 & n22608 ) | ( n22606 & n22608 ) ;
  assign n22610 = n22329 & ~n22609 ;
  assign n22611 = n22607 | n22610 ;
  assign n22612 = x107 & n3816 ;
  assign n22613 = x106 & n3811 ;
  assign n22614 = x105 & ~n3810 ;
  assign n22615 = n4067 & n22614 ;
  assign n22616 = n22613 | n22615 ;
  assign n22617 = n22612 | n22616 ;
  assign n22618 = n3819 | n22612 ;
  assign n22619 = n22616 | n22618 ;
  assign n22620 = ( n9084 & n22617 ) | ( n9084 & n22619 ) | ( n22617 & n22619 ) ;
  assign n22621 = x29 & n22619 ;
  assign n22622 = x29 & n22612 ;
  assign n22623 = ( x29 & n22616 ) | ( x29 & n22622 ) | ( n22616 & n22622 ) ;
  assign n22624 = ( n9084 & n22621 ) | ( n9084 & n22623 ) | ( n22621 & n22623 ) ;
  assign n22625 = x29 & ~n22623 ;
  assign n22626 = x29 & ~n22619 ;
  assign n22627 = ( ~n9084 & n22625 ) | ( ~n9084 & n22626 ) | ( n22625 & n22626 ) ;
  assign n22628 = ( n22620 & ~n22624 ) | ( n22620 & n22627 ) | ( ~n22624 & n22627 ) ;
  assign n22629 = n22144 | n22169 ;
  assign n22630 = ( n22169 & n22170 ) | ( n22169 & n22629 ) | ( n22170 & n22629 ) ;
  assign n22631 = ( n22611 & n22628 ) | ( n22611 & ~n22630 ) | ( n22628 & ~n22630 ) ;
  assign n22632 = ( ~n22628 & n22630 ) | ( ~n22628 & n22631 ) | ( n22630 & n22631 ) ;
  assign n22633 = ( ~n22611 & n22631 ) | ( ~n22611 & n22632 ) | ( n22631 & n22632 ) ;
  assign n22634 = n22309 & ~n22633 ;
  assign n22635 = n22309 | n22633 ;
  assign n22636 = ( ~n22309 & n22634 ) | ( ~n22309 & n22635 ) | ( n22634 & n22635 ) ;
  assign n22637 = ( n22265 & ~n22273 ) | ( n22265 & n22636 ) | ( ~n22273 & n22636 ) ;
  assign n22638 = n22265 & n22636 ;
  assign n22639 = ( ~n22282 & n22637 ) | ( ~n22282 & n22638 ) | ( n22637 & n22638 ) ;
  assign n22283 = n22273 | n22282 ;
  assign n22640 = ( n22283 & ~n22636 ) | ( n22283 & n22639 ) | ( ~n22636 & n22639 ) ;
  assign n22641 = ( ~n22265 & n22639 ) | ( ~n22265 & n22640 ) | ( n22639 & n22640 ) ;
  assign n22642 = ~n22251 & n22641 ;
  assign n22643 = n22244 | n22639 ;
  assign n22644 = ~n22244 & n22265 ;
  assign n22645 = ( n22640 & n22643 ) | ( n22640 & ~n22644 ) | ( n22643 & ~n22644 ) ;
  assign n22646 = ( n22187 & n22641 ) | ( n22187 & n22645 ) | ( n22641 & n22645 ) ;
  assign n22647 = ( n21823 & n22641 ) | ( n21823 & n22645 ) | ( n22641 & n22645 ) ;
  assign n22648 = ( n21824 & n22646 ) | ( n21824 & n22647 ) | ( n22646 & n22647 ) ;
  assign n22649 = n22250 & ~n22648 ;
  assign n22650 = n22642 | n22649 ;
  assign n22652 = x121 & n957 ;
  assign n22653 = x120 & ~n956 ;
  assign n22654 = n1105 & n22653 ;
  assign n22655 = n22652 | n22654 ;
  assign n22651 = x122 & n962 ;
  assign n22657 = n965 | n22651 ;
  assign n22658 = n22655 | n22657 ;
  assign n22656 = n22651 | n22655 ;
  assign n22659 = n22656 & n22658 ;
  assign n22660 = ( n16043 & n22658 ) | ( n16043 & n22659 ) | ( n22658 & n22659 ) ;
  assign n22661 = x14 & n22659 ;
  assign n22662 = x14 & n22658 ;
  assign n22663 = ( n16043 & n22661 ) | ( n16043 & n22662 ) | ( n22661 & n22662 ) ;
  assign n22664 = x14 & ~n22659 ;
  assign n22665 = x14 & ~n22658 ;
  assign n22666 = ( ~n16043 & n22664 ) | ( ~n16043 & n22665 ) | ( n22664 & n22665 ) ;
  assign n22667 = ( n22660 & ~n22663 ) | ( n22660 & n22666 ) | ( ~n22663 & n22666 ) ;
  assign n22668 = n21763 & n22667 ;
  assign n22669 = n21748 & n22668 ;
  assign n22670 = n21192 & n22668 ;
  assign n22671 = ( n21194 & n22669 ) | ( n21194 & n22670 ) | ( n22669 & n22670 ) ;
  assign n22672 = ( n22197 & n22667 ) | ( n22197 & n22671 ) | ( n22667 & n22671 ) ;
  assign n22673 = n21763 | n22667 ;
  assign n22674 = ( n21748 & n22667 ) | ( n21748 & n22673 ) | ( n22667 & n22673 ) ;
  assign n22675 = ( n21192 & n22667 ) | ( n21192 & n22673 ) | ( n22667 & n22673 ) ;
  assign n22676 = ( n21194 & n22674 ) | ( n21194 & n22675 ) | ( n22674 & n22675 ) ;
  assign n22677 = n22197 | n22676 ;
  assign n22678 = ~n22672 & n22677 ;
  assign n22679 = x119 & n1383 ;
  assign n22680 = x118 & n1378 ;
  assign n22681 = x117 & ~n1377 ;
  assign n22682 = n1542 & n22681 ;
  assign n22683 = n22680 | n22682 ;
  assign n22684 = n22679 | n22683 ;
  assign n22685 = n1386 | n22679 ;
  assign n22686 = n22683 | n22685 ;
  assign n22687 = ( n14496 & n22684 ) | ( n14496 & n22686 ) | ( n22684 & n22686 ) ;
  assign n22688 = x17 & n22686 ;
  assign n22689 = x17 & n22679 ;
  assign n22690 = ( x17 & n22683 ) | ( x17 & n22689 ) | ( n22683 & n22689 ) ;
  assign n22691 = ( n14496 & n22688 ) | ( n14496 & n22690 ) | ( n22688 & n22690 ) ;
  assign n22692 = x17 & ~n22690 ;
  assign n22693 = x17 & ~n22686 ;
  assign n22694 = ( ~n14496 & n22692 ) | ( ~n14496 & n22693 ) | ( n22692 & n22693 ) ;
  assign n22695 = ( n22687 & ~n22691 ) | ( n22687 & n22694 ) | ( ~n22691 & n22694 ) ;
  assign n22696 = n21799 | n22189 ;
  assign n22697 = n21798 | n22189 ;
  assign n22698 = ( n21784 & n22696 ) | ( n21784 & n22697 ) | ( n22696 & n22697 ) ;
  assign n22699 = n22695 | n22698 ;
  assign n22700 = n21800 | n22695 ;
  assign n22701 = ( n21803 & n22699 ) | ( n21803 & n22700 ) | ( n22699 & n22700 ) ;
  assign n22702 = n22695 & n22698 ;
  assign n22703 = n21800 & n22695 ;
  assign n22704 = ( n21803 & n22702 ) | ( n21803 & n22703 ) | ( n22702 & n22703 ) ;
  assign n22705 = n22701 & ~n22704 ;
  assign n22706 = ( n22650 & n22678 ) | ( n22650 & ~n22705 ) | ( n22678 & ~n22705 ) ;
  assign n22707 = ( ~n22678 & n22705 ) | ( ~n22678 & n22706 ) | ( n22705 & n22706 ) ;
  assign n22708 = ( ~n22650 & n22706 ) | ( ~n22650 & n22707 ) | ( n22706 & n22707 ) ;
  assign n22709 = x127 & n384 ;
  assign n22710 = x126 & ~n383 ;
  assign n22711 = n463 & n22710 ;
  assign n22712 = n22709 | n22711 ;
  assign n22713 = n392 | n22712 ;
  assign n22714 = ( n19328 & n22712 ) | ( n19328 & n22713 ) | ( n22712 & n22713 ) ;
  assign n22715 = x8 & n22712 ;
  assign n22716 = x8 & n392 ;
  assign n22717 = ( x8 & n22712 ) | ( x8 & n22716 ) | ( n22712 & n22716 ) ;
  assign n22718 = ( n19328 & n22715 ) | ( n19328 & n22717 ) | ( n22715 & n22717 ) ;
  assign n22719 = x8 & ~n22716 ;
  assign n22720 = ~n22712 & n22719 ;
  assign n22721 = x8 & ~n22712 ;
  assign n22722 = ( ~n19328 & n22720 ) | ( ~n19328 & n22721 ) | ( n22720 & n22721 ) ;
  assign n22723 = ( n22714 & ~n22718 ) | ( n22714 & n22722 ) | ( ~n22718 & n22722 ) ;
  assign n22724 = n21706 | n22203 ;
  assign n22725 = ( n21706 & n21707 ) | ( n21706 & n22724 ) | ( n21707 & n22724 ) ;
  assign n22726 = n22723 & n22725 ;
  assign n22727 = n22723 | n22725 ;
  assign n22728 = ~n22726 & n22727 ;
  assign n22729 = x125 & n636 ;
  assign n22730 = x124 & n631 ;
  assign n22731 = x123 & ~n630 ;
  assign n22732 = n764 & n22731 ;
  assign n22733 = n22730 | n22732 ;
  assign n22734 = n22729 | n22733 ;
  assign n22735 = n639 | n22729 ;
  assign n22736 = n22733 | n22735 ;
  assign n22737 = ( n17670 & n22734 ) | ( n17670 & n22736 ) | ( n22734 & n22736 ) ;
  assign n22738 = x11 & n22736 ;
  assign n22739 = x11 & n22729 ;
  assign n22740 = ( x11 & n22733 ) | ( x11 & n22739 ) | ( n22733 & n22739 ) ;
  assign n22741 = ( n17670 & n22738 ) | ( n17670 & n22740 ) | ( n22738 & n22740 ) ;
  assign n22742 = x11 & ~n22740 ;
  assign n22743 = x11 & ~n22736 ;
  assign n22744 = ( ~n17670 & n22742 ) | ( ~n17670 & n22743 ) | ( n22742 & n22743 ) ;
  assign n22745 = ( n22737 & ~n22741 ) | ( n22737 & n22744 ) | ( ~n22741 & n22744 ) ;
  assign n22746 = n21742 | n22200 ;
  assign n22747 = n21741 | n22200 ;
  assign n22748 = ( n21724 & n22746 ) | ( n21724 & n22747 ) | ( n22746 & n22747 ) ;
  assign n22749 = n22745 | n22748 ;
  assign n22750 = n21743 | n22745 ;
  assign n22751 = ( n21746 & n22749 ) | ( n21746 & n22750 ) | ( n22749 & n22750 ) ;
  assign n22752 = n22745 & n22748 ;
  assign n22753 = n21743 & n22745 ;
  assign n22754 = ( n21746 & n22752 ) | ( n21746 & n22753 ) | ( n22752 & n22753 ) ;
  assign n22755 = n22751 & ~n22754 ;
  assign n22756 = ( n22708 & n22728 ) | ( n22708 & ~n22755 ) | ( n22728 & ~n22755 ) ;
  assign n22757 = ( ~n22728 & n22755 ) | ( ~n22728 & n22756 ) | ( n22755 & n22756 ) ;
  assign n22758 = ( ~n22708 & n22756 ) | ( ~n22708 & n22757 ) | ( n22756 & n22757 ) ;
  assign n22783 = n22758 & n22782 ;
  assign n22784 = n22782 & ~n22783 ;
  assign n22785 = n22758 & ~n22782 ;
  assign n22786 = n22784 | n22785 ;
  assign n22787 = n22219 | n22222 ;
  assign n22788 = ( n22219 & n22224 ) | ( n22219 & n22787 ) | ( n22224 & n22787 ) ;
  assign n22789 = ( n21658 & n22219 ) | ( n21658 & n22787 ) | ( n22219 & n22787 ) ;
  assign n22790 = ( n21071 & n22788 ) | ( n21071 & n22789 ) | ( n22788 & n22789 ) ;
  assign n22791 = n22787 | n22789 ;
  assign n22792 = n22219 | n22789 ;
  assign n22793 = ( n22224 & n22791 ) | ( n22224 & n22792 ) | ( n22791 & n22792 ) ;
  assign n22794 = ( n21078 & n22790 ) | ( n21078 & n22793 ) | ( n22790 & n22793 ) ;
  assign n22795 = n22786 | n22794 ;
  assign n22796 = n22786 & n22794 ;
  assign n22797 = n22795 & ~n22796 ;
  assign n22816 = n22708 | n22754 ;
  assign n22817 = ( n22754 & n22755 ) | ( n22754 & n22816 ) | ( n22755 & n22816 ) ;
  assign n22798 = x127 & ~n383 ;
  assign n22799 = n463 & n22798 ;
  assign n22800 = n392 & n19877 ;
  assign n22801 = n22799 | n22800 ;
  assign n22802 = n392 & n19880 ;
  assign n22803 = n22799 | n22802 ;
  assign n22804 = ( n18202 & n22801 ) | ( n18202 & n22803 ) | ( n22801 & n22803 ) ;
  assign n22805 = n22801 & n22803 ;
  assign n22806 = ( n18212 & n22804 ) | ( n18212 & n22805 ) | ( n22804 & n22805 ) ;
  assign n22807 = ( n18214 & n22804 ) | ( n18214 & n22805 ) | ( n22804 & n22805 ) ;
  assign n22808 = ( n14002 & n22806 ) | ( n14002 & n22807 ) | ( n22806 & n22807 ) ;
  assign n22809 = x8 & n22806 ;
  assign n22810 = x8 & n22807 ;
  assign n22811 = ( n14002 & n22809 ) | ( n14002 & n22810 ) | ( n22809 & n22810 ) ;
  assign n22812 = x8 & ~n22810 ;
  assign n22813 = x8 & ~n22809 ;
  assign n22814 = ( ~n14002 & n22812 ) | ( ~n14002 & n22813 ) | ( n22812 & n22813 ) ;
  assign n22815 = ( n22808 & ~n22811 ) | ( n22808 & n22814 ) | ( ~n22811 & n22814 ) ;
  assign n22818 = n22815 & n22817 ;
  assign n22819 = n22817 & ~n22818 ;
  assign n22820 = n22650 & n22705 ;
  assign n22821 = n22650 | n22705 ;
  assign n22822 = ~n22820 & n22821 ;
  assign n22823 = n22671 | n22822 ;
  assign n22824 = n22667 | n22822 ;
  assign n22825 = ( n22197 & n22823 ) | ( n22197 & n22824 ) | ( n22823 & n22824 ) ;
  assign n22826 = ( n22672 & n22678 ) | ( n22672 & n22825 ) | ( n22678 & n22825 ) ;
  assign n22828 = x125 & n631 ;
  assign n22829 = x124 & ~n630 ;
  assign n22830 = n764 & n22829 ;
  assign n22831 = n22828 | n22830 ;
  assign n22827 = x126 & n636 ;
  assign n22833 = n639 | n22827 ;
  assign n22834 = n22831 | n22833 ;
  assign n22832 = n22827 | n22831 ;
  assign n22835 = n22832 & n22834 ;
  assign n22836 = ( n18220 & n22834 ) | ( n18220 & n22835 ) | ( n22834 & n22835 ) ;
  assign n22837 = x11 & n22835 ;
  assign n22838 = x11 & n22834 ;
  assign n22839 = ( n18220 & n22837 ) | ( n18220 & n22838 ) | ( n22837 & n22838 ) ;
  assign n22840 = x11 & ~n22835 ;
  assign n22841 = x11 & ~n22834 ;
  assign n22842 = ( ~n18220 & n22840 ) | ( ~n18220 & n22841 ) | ( n22840 & n22841 ) ;
  assign n22843 = ( n22836 & ~n22839 ) | ( n22836 & n22842 ) | ( ~n22839 & n22842 ) ;
  assign n22844 = n22825 & n22843 ;
  assign n22845 = n22672 & n22843 ;
  assign n22846 = ( n22678 & n22844 ) | ( n22678 & n22845 ) | ( n22844 & n22845 ) ;
  assign n22847 = n22826 & ~n22846 ;
  assign n22848 = x120 & n1383 ;
  assign n22849 = x119 & n1378 ;
  assign n22850 = x118 & ~n1377 ;
  assign n22851 = n1542 & n22850 ;
  assign n22852 = n22849 | n22851 ;
  assign n22853 = n22848 | n22852 ;
  assign n22854 = n1386 | n22848 ;
  assign n22855 = n22852 | n22854 ;
  assign n22856 = ( n14991 & n22853 ) | ( n14991 & n22855 ) | ( n22853 & n22855 ) ;
  assign n22857 = x17 & n22855 ;
  assign n22858 = x17 & n22848 ;
  assign n22859 = ( x17 & n22852 ) | ( x17 & n22858 ) | ( n22852 & n22858 ) ;
  assign n22860 = ( n14991 & n22857 ) | ( n14991 & n22859 ) | ( n22857 & n22859 ) ;
  assign n22861 = x17 & ~n22859 ;
  assign n22862 = x17 & ~n22855 ;
  assign n22863 = ( ~n14991 & n22861 ) | ( ~n14991 & n22862 ) | ( n22861 & n22862 ) ;
  assign n22864 = ( n22856 & ~n22860 ) | ( n22856 & n22863 ) | ( ~n22860 & n22863 ) ;
  assign n22865 = n22648 & n22864 ;
  assign n22866 = n22247 & n22864 ;
  assign n22867 = ( n22251 & n22865 ) | ( n22251 & n22866 ) | ( n22865 & n22866 ) ;
  assign n22868 = n22648 | n22864 ;
  assign n22869 = n22247 | n22864 ;
  assign n22870 = ( n22251 & n22868 ) | ( n22251 & n22869 ) | ( n22868 & n22869 ) ;
  assign n22871 = ~n22867 & n22870 ;
  assign n22872 = x114 & n2429 ;
  assign n22873 = x113 & n2424 ;
  assign n22874 = x112 & ~n2423 ;
  assign n22875 = n2631 & n22874 ;
  assign n22876 = n22873 | n22875 ;
  assign n22877 = n22872 | n22876 ;
  assign n22878 = n2432 | n22872 ;
  assign n22879 = n22876 | n22878 ;
  assign n22880 = ( ~n12095 & n22877 ) | ( ~n12095 & n22879 ) | ( n22877 & n22879 ) ;
  assign n22881 = n22877 & n22879 ;
  assign n22882 = ( n12079 & n22880 ) | ( n12079 & n22881 ) | ( n22880 & n22881 ) ;
  assign n22883 = x23 & n22882 ;
  assign n22884 = x23 & ~n22882 ;
  assign n22885 = ( n22882 & ~n22883 ) | ( n22882 & n22884 ) | ( ~n22883 & n22884 ) ;
  assign n22886 = n22305 | n22633 ;
  assign n22887 = ( n22305 & n22309 ) | ( n22305 & n22886 ) | ( n22309 & n22886 ) ;
  assign n22888 = n22885 | n22887 ;
  assign n22889 = n22885 & n22887 ;
  assign n22890 = n22888 & ~n22889 ;
  assign n22891 = n22628 & n22630 ;
  assign n22892 = n22630 & ~n22891 ;
  assign n22893 = n22610 & n22628 ;
  assign n22894 = ( n22607 & n22628 ) | ( n22607 & n22893 ) | ( n22628 & n22893 ) ;
  assign n22895 = ~n22630 & n22894 ;
  assign n22896 = n22891 | n22895 ;
  assign n22897 = n22611 | n22628 ;
  assign n22898 = ( n22611 & n22630 ) | ( n22611 & n22897 ) | ( n22630 & n22897 ) ;
  assign n22899 = ( n22892 & n22896 ) | ( n22892 & n22898 ) | ( n22896 & n22898 ) ;
  assign n22900 = x111 & n3085 ;
  assign n22901 = x110 & n3080 ;
  assign n22902 = x109 & ~n3079 ;
  assign n22903 = n3309 & n22902 ;
  assign n22904 = n22901 | n22903 ;
  assign n22905 = n22900 | n22904 ;
  assign n22906 = n3088 | n22900 ;
  assign n22907 = n22904 | n22906 ;
  assign n22908 = ( n10749 & n22905 ) | ( n10749 & n22907 ) | ( n22905 & n22907 ) ;
  assign n22909 = x26 & n22907 ;
  assign n22910 = x26 & n22900 ;
  assign n22911 = ( x26 & n22904 ) | ( x26 & n22910 ) | ( n22904 & n22910 ) ;
  assign n22912 = ( n10749 & n22909 ) | ( n10749 & n22911 ) | ( n22909 & n22911 ) ;
  assign n22913 = x26 & ~n22911 ;
  assign n22914 = x26 & ~n22907 ;
  assign n22915 = ( ~n10749 & n22913 ) | ( ~n10749 & n22914 ) | ( n22913 & n22914 ) ;
  assign n22916 = ( n22908 & ~n22912 ) | ( n22908 & n22915 ) | ( ~n22912 & n22915 ) ;
  assign n22917 = n22628 & n22916 ;
  assign n22918 = n22630 & n22917 ;
  assign n22919 = ( n22895 & n22916 ) | ( n22895 & n22918 ) | ( n22916 & n22918 ) ;
  assign n22920 = ( n22611 & n22916 ) | ( n22611 & n22917 ) | ( n22916 & n22917 ) ;
  assign n22921 = n22611 & n22916 ;
  assign n22922 = ( n22630 & n22920 ) | ( n22630 & n22921 ) | ( n22920 & n22921 ) ;
  assign n22923 = ( n22892 & n22919 ) | ( n22892 & n22922 ) | ( n22919 & n22922 ) ;
  assign n22924 = n22899 & ~n22923 ;
  assign n22925 = ( n22330 & n22331 ) | ( n22330 & n22609 ) | ( n22331 & n22609 ) ;
  assign n22927 = x107 & n3811 ;
  assign n22928 = x106 & ~n3810 ;
  assign n22929 = n4067 & n22928 ;
  assign n22930 = n22927 | n22929 ;
  assign n22926 = x108 & n3816 ;
  assign n22932 = n3819 | n22926 ;
  assign n22933 = n22930 | n22932 ;
  assign n22931 = n22926 | n22930 ;
  assign n22934 = n22931 & n22933 ;
  assign n22935 = ( n9479 & n22933 ) | ( n9479 & n22934 ) | ( n22933 & n22934 ) ;
  assign n22936 = x29 & n22934 ;
  assign n22937 = x29 & n22933 ;
  assign n22938 = ( n9479 & n22936 ) | ( n9479 & n22937 ) | ( n22936 & n22937 ) ;
  assign n22939 = x29 & ~n22934 ;
  assign n22940 = x29 & ~n22933 ;
  assign n22941 = ( ~n9479 & n22939 ) | ( ~n9479 & n22940 ) | ( n22939 & n22940 ) ;
  assign n22942 = ( n22935 & ~n22938 ) | ( n22935 & n22941 ) | ( ~n22938 & n22941 ) ;
  assign n22943 = n22609 & n22942 ;
  assign n22944 = n22330 & n22942 ;
  assign n22945 = ( n22331 & n22943 ) | ( n22331 & n22944 ) | ( n22943 & n22944 ) ;
  assign n22946 = n22925 & ~n22945 ;
  assign n22947 = x102 & n5554 ;
  assign n22948 = x101 & n5549 ;
  assign n22949 = x100 & ~n5548 ;
  assign n22950 = n5893 & n22949 ;
  assign n22951 = n22948 | n22950 ;
  assign n22952 = n22947 | n22951 ;
  assign n22953 = n5557 | n22947 ;
  assign n22954 = n22951 | n22953 ;
  assign n22955 = ( n7178 & n22952 ) | ( n7178 & n22954 ) | ( n22952 & n22954 ) ;
  assign n22956 = x35 & n22954 ;
  assign n22957 = x35 & n22947 ;
  assign n22958 = ( x35 & n22951 ) | ( x35 & n22957 ) | ( n22951 & n22957 ) ;
  assign n22959 = ( n7178 & n22956 ) | ( n7178 & n22958 ) | ( n22956 & n22958 ) ;
  assign n22960 = x35 & ~n22958 ;
  assign n22961 = x35 & ~n22954 ;
  assign n22962 = ( ~n7178 & n22960 ) | ( ~n7178 & n22961 ) | ( n22960 & n22961 ) ;
  assign n22963 = ( n22955 & ~n22959 ) | ( n22955 & n22962 ) | ( ~n22959 & n22962 ) ;
  assign n22964 = x105 & n4631 ;
  assign n22965 = x104 & n4626 ;
  assign n22966 = x103 & ~n4625 ;
  assign n22967 = n4943 & n22966 ;
  assign n22968 = n22965 | n22967 ;
  assign n22969 = n22964 | n22968 ;
  assign n22970 = n4634 | n22964 ;
  assign n22971 = n22968 | n22970 ;
  assign n22972 = ( n8273 & n22969 ) | ( n8273 & n22971 ) | ( n22969 & n22971 ) ;
  assign n22973 = x32 & n22971 ;
  assign n22974 = x32 & n22964 ;
  assign n22975 = ( x32 & n22968 ) | ( x32 & n22974 ) | ( n22968 & n22974 ) ;
  assign n22976 = ( n8273 & n22973 ) | ( n8273 & n22975 ) | ( n22973 & n22975 ) ;
  assign n22977 = x32 & ~n22975 ;
  assign n22978 = x32 & ~n22971 ;
  assign n22979 = ( ~n8273 & n22977 ) | ( ~n8273 & n22978 ) | ( n22977 & n22978 ) ;
  assign n22980 = ( n22972 & ~n22976 ) | ( n22972 & n22979 ) | ( ~n22976 & n22979 ) ;
  assign n22981 = n22583 | n22603 ;
  assign n22982 = ( n22583 & n22586 ) | ( n22583 & n22981 ) | ( n22586 & n22981 ) ;
  assign n22983 = n22980 | n22982 ;
  assign n22984 = n22980 & n22982 ;
  assign n22985 = n22983 & ~n22984 ;
  assign n23116 = ( n22418 & n22419 ) | ( n22418 & n22438 ) | ( n22419 & n22438 ) ;
  assign n22986 = x72 & n18290 ;
  assign n22987 = x63 & x71 ;
  assign n22988 = ~n18290 & n22987 ;
  assign n22989 = n22986 | n22988 ;
  assign n22990 = ~n22350 & n22989 ;
  assign n22991 = n22350 & ~n22989 ;
  assign n22992 = n22352 | n22991 ;
  assign n22993 = ( ~n22354 & n22991 ) | ( ~n22354 & n22992 ) | ( n22991 & n22992 ) ;
  assign n22994 = n22990 | n22993 ;
  assign n22995 = n22990 | n22991 ;
  assign n22996 = n22352 | n22995 ;
  assign n22997 = ( n22345 & n22994 ) | ( n22345 & n22996 ) | ( n22994 & n22996 ) ;
  assign n22998 = ( n710 & n22341 ) | ( n710 & n22342 ) | ( n22341 & n22342 ) ;
  assign n22999 = ( n22994 & n22996 ) | ( n22994 & ~n22998 ) | ( n22996 & ~n22998 ) ;
  assign n23000 = ( ~n22346 & n22997 ) | ( ~n22346 & n22999 ) | ( n22997 & n22999 ) ;
  assign n23001 = ( ~n22352 & n22359 ) | ( ~n22352 & n23000 ) | ( n22359 & n23000 ) ;
  assign n23002 = ~n22995 & n23000 ;
  assign n23003 = n23001 | n23002 ;
  assign n23004 = x75 & n17146 ;
  assign n23005 = x74 & n17141 ;
  assign n23006 = x73 & ~n17140 ;
  assign n23007 = n17724 & n23006 ;
  assign n23008 = n23005 | n23007 ;
  assign n23009 = n23004 | n23008 ;
  assign n23010 = n17149 | n23004 ;
  assign n23011 = n23008 | n23010 ;
  assign n23012 = ( n746 & n23009 ) | ( n746 & n23011 ) | ( n23009 & n23011 ) ;
  assign n23013 = x62 & n23011 ;
  assign n23014 = x62 & n23004 ;
  assign n23015 = ( x62 & n23008 ) | ( x62 & n23014 ) | ( n23008 & n23014 ) ;
  assign n23016 = ( n746 & n23013 ) | ( n746 & n23015 ) | ( n23013 & n23015 ) ;
  assign n23017 = x62 & ~n23015 ;
  assign n23018 = x62 & ~n23011 ;
  assign n23019 = ( ~n746 & n23017 ) | ( ~n746 & n23018 ) | ( n23017 & n23018 ) ;
  assign n23020 = ( n23012 & ~n23016 ) | ( n23012 & n23019 ) | ( ~n23016 & n23019 ) ;
  assign n23021 = n23003 & ~n23020 ;
  assign n23022 = ~n23003 & n23020 ;
  assign n23023 = n23021 | n23022 ;
  assign n23024 = x78 & n15552 ;
  assign n23025 = x77 & n15547 ;
  assign n23026 = x76 & ~n15546 ;
  assign n23027 = n16123 & n23026 ;
  assign n23028 = n23025 | n23027 ;
  assign n23029 = n23024 | n23028 ;
  assign n23030 = n15555 | n23024 ;
  assign n23031 = n23028 | n23030 ;
  assign n23032 = ( n1192 & n23029 ) | ( n1192 & n23031 ) | ( n23029 & n23031 ) ;
  assign n23033 = x59 & n23031 ;
  assign n23034 = x59 & n23024 ;
  assign n23035 = ( x59 & n23028 ) | ( x59 & n23034 ) | ( n23028 & n23034 ) ;
  assign n23036 = ( n1192 & n23033 ) | ( n1192 & n23035 ) | ( n23033 & n23035 ) ;
  assign n23037 = x59 & ~n23035 ;
  assign n23038 = x59 & ~n23031 ;
  assign n23039 = ( ~n1192 & n23037 ) | ( ~n1192 & n23038 ) | ( n23037 & n23038 ) ;
  assign n23040 = ( n23032 & ~n23036 ) | ( n23032 & n23039 ) | ( ~n23036 & n23039 ) ;
  assign n23041 = n23023 & n23040 ;
  assign n23042 = n23023 | n23040 ;
  assign n23043 = ~n23041 & n23042 ;
  assign n23044 = n22365 | n22387 ;
  assign n23045 = ( n22367 & n22387 ) | ( n22367 & n23044 ) | ( n22387 & n23044 ) ;
  assign n23046 = ( n22368 & n22370 ) | ( n22368 & n23045 ) | ( n22370 & n23045 ) ;
  assign n23047 = n23043 | n23046 ;
  assign n23048 = n23043 & n23046 ;
  assign n23049 = n23047 & ~n23048 ;
  assign n23050 = x81 & n14045 ;
  assign n23051 = x80 & n14040 ;
  assign n23052 = x79 & ~n14039 ;
  assign n23053 = n14552 & n23052 ;
  assign n23054 = n23051 | n23053 ;
  assign n23055 = n23050 | n23054 ;
  assign n23056 = n14048 | n23050 ;
  assign n23057 = n23054 | n23056 ;
  assign n23058 = ( n1651 & n23055 ) | ( n1651 & n23057 ) | ( n23055 & n23057 ) ;
  assign n23059 = x56 & n23057 ;
  assign n23060 = x56 & n23050 ;
  assign n23061 = ( x56 & n23054 ) | ( x56 & n23060 ) | ( n23054 & n23060 ) ;
  assign n23062 = ( n1651 & n23059 ) | ( n1651 & n23061 ) | ( n23059 & n23061 ) ;
  assign n23063 = x56 & ~n23061 ;
  assign n23064 = x56 & ~n23057 ;
  assign n23065 = ( ~n1651 & n23063 ) | ( ~n1651 & n23064 ) | ( n23063 & n23064 ) ;
  assign n23066 = ( n23058 & ~n23062 ) | ( n23058 & n23065 ) | ( ~n23062 & n23065 ) ;
  assign n23067 = ~n23049 & n23066 ;
  assign n23068 = n23045 | n23066 ;
  assign n23069 = n22368 | n23066 ;
  assign n23070 = ( n22370 & n23068 ) | ( n22370 & n23069 ) | ( n23068 & n23069 ) ;
  assign n23071 = ( n23043 & n23066 ) | ( n23043 & n23070 ) | ( n23066 & n23070 ) ;
  assign n23072 = n23047 & ~n23071 ;
  assign n23073 = n23067 | n23072 ;
  assign n23074 = n22392 | n22410 ;
  assign n23075 = ( n22392 & n22393 ) | ( n22392 & n23074 ) | ( n22393 & n23074 ) ;
  assign n23076 = n23073 | n23075 ;
  assign n23077 = n23073 & n23075 ;
  assign n23078 = n23076 & ~n23077 ;
  assign n23079 = x84 & n12574 ;
  assign n23080 = x83 & n12569 ;
  assign n23081 = x82 & ~n12568 ;
  assign n23082 = n13076 & n23081 ;
  assign n23083 = n23080 | n23082 ;
  assign n23084 = n23079 | n23083 ;
  assign n23085 = n12577 | n23079 ;
  assign n23086 = n23083 | n23085 ;
  assign n23087 = ( n2194 & n23084 ) | ( n2194 & n23086 ) | ( n23084 & n23086 ) ;
  assign n23088 = x53 & n23086 ;
  assign n23089 = x53 & n23079 ;
  assign n23090 = ( x53 & n23083 ) | ( x53 & n23089 ) | ( n23083 & n23089 ) ;
  assign n23091 = ( n2194 & n23088 ) | ( n2194 & n23090 ) | ( n23088 & n23090 ) ;
  assign n23092 = x53 & ~n23090 ;
  assign n23093 = x53 & ~n23086 ;
  assign n23094 = ( ~n2194 & n23092 ) | ( ~n2194 & n23093 ) | ( n23092 & n23093 ) ;
  assign n23095 = ( n23087 & ~n23091 ) | ( n23087 & n23094 ) | ( ~n23091 & n23094 ) ;
  assign n23096 = n23078 | n23095 ;
  assign n23097 = n23078 & n23095 ;
  assign n23098 = n23096 & ~n23097 ;
  assign n23099 = x87 & n11205 ;
  assign n23100 = x86 & n11200 ;
  assign n23101 = x85 & ~n11199 ;
  assign n23102 = n11679 & n23101 ;
  assign n23103 = n23100 | n23102 ;
  assign n23104 = n23099 | n23103 ;
  assign n23105 = n11208 | n23099 ;
  assign n23106 = n23103 | n23105 ;
  assign n23107 = ( n2816 & n23104 ) | ( n2816 & n23106 ) | ( n23104 & n23106 ) ;
  assign n23108 = x50 & n23106 ;
  assign n23109 = x50 & n23099 ;
  assign n23110 = ( x50 & n23103 ) | ( x50 & n23109 ) | ( n23103 & n23109 ) ;
  assign n23111 = ( n2816 & n23108 ) | ( n2816 & n23110 ) | ( n23108 & n23110 ) ;
  assign n23112 = x50 & ~n23110 ;
  assign n23113 = x50 & ~n23106 ;
  assign n23114 = ( ~n2816 & n23112 ) | ( ~n2816 & n23113 ) | ( n23112 & n23113 ) ;
  assign n23115 = ( n23107 & ~n23111 ) | ( n23107 & n23114 ) | ( ~n23111 & n23114 ) ;
  assign n23117 = ( ~n23098 & n23115 ) | ( ~n23098 & n23116 ) | ( n23115 & n23116 ) ;
  assign n23118 = ( n23098 & ~n23115 ) | ( n23098 & n23117 ) | ( ~n23115 & n23117 ) ;
  assign n23119 = ( ~n23116 & n23117 ) | ( ~n23116 & n23118 ) | ( n23117 & n23118 ) ;
  assign n23120 = ( n22444 & n22445 ) | ( n22444 & n22464 ) | ( n22445 & n22464 ) ;
  assign n23121 = n23119 & n23120 ;
  assign n23122 = n23119 | n23120 ;
  assign n23123 = ~n23121 & n23122 ;
  assign n23124 = x90 & n9933 ;
  assign n23125 = x89 & n9928 ;
  assign n23126 = x88 & ~n9927 ;
  assign n23127 = n10379 & n23126 ;
  assign n23128 = n23125 | n23127 ;
  assign n23129 = n23124 | n23128 ;
  assign n23130 = n9936 | n23124 ;
  assign n23131 = n23128 | n23130 ;
  assign n23132 = ( n3519 & n23129 ) | ( n3519 & n23131 ) | ( n23129 & n23131 ) ;
  assign n23133 = x47 & n23131 ;
  assign n23134 = x47 & n23124 ;
  assign n23135 = ( x47 & n23128 ) | ( x47 & n23134 ) | ( n23128 & n23134 ) ;
  assign n23136 = ( n3519 & n23133 ) | ( n3519 & n23135 ) | ( n23133 & n23135 ) ;
  assign n23137 = x47 & ~n23135 ;
  assign n23138 = x47 & ~n23131 ;
  assign n23139 = ( ~n3519 & n23137 ) | ( ~n3519 & n23138 ) | ( n23137 & n23138 ) ;
  assign n23140 = ( n23132 & ~n23136 ) | ( n23132 & n23139 ) | ( ~n23136 & n23139 ) ;
  assign n23141 = n23123 & ~n23140 ;
  assign n23142 = n23123 | n23140 ;
  assign n23143 = ( ~n23123 & n23141 ) | ( ~n23123 & n23142 ) | ( n23141 & n23142 ) ;
  assign n23144 = ( n22474 & n22475 ) | ( n22474 & n22497 ) | ( n22475 & n22497 ) ;
  assign n23145 = n23143 | n23144 ;
  assign n23146 = n23143 & n23144 ;
  assign n23147 = n23145 & ~n23146 ;
  assign n23148 = x93 & n8724 ;
  assign n23149 = x92 & n8719 ;
  assign n23150 = x91 & ~n8718 ;
  assign n23151 = n9149 & n23150 ;
  assign n23152 = n23149 | n23151 ;
  assign n23153 = n23148 | n23152 ;
  assign n23154 = n8727 | n23148 ;
  assign n23155 = n23152 | n23154 ;
  assign n23156 = ( n4305 & n23153 ) | ( n4305 & n23155 ) | ( n23153 & n23155 ) ;
  assign n23157 = x44 & n23155 ;
  assign n23158 = x44 & n23148 ;
  assign n23159 = ( x44 & n23152 ) | ( x44 & n23158 ) | ( n23152 & n23158 ) ;
  assign n23160 = ( n4305 & n23157 ) | ( n4305 & n23159 ) | ( n23157 & n23159 ) ;
  assign n23161 = x44 & ~n23159 ;
  assign n23162 = x44 & ~n23155 ;
  assign n23163 = ( ~n4305 & n23161 ) | ( ~n4305 & n23162 ) | ( n23161 & n23162 ) ;
  assign n23164 = ( n23156 & ~n23160 ) | ( n23156 & n23163 ) | ( ~n23160 & n23163 ) ;
  assign n23165 = ~n23147 & n23164 ;
  assign n23166 = n23143 | n23164 ;
  assign n23167 = ( n23144 & n23164 ) | ( n23144 & n23166 ) | ( n23164 & n23166 ) ;
  assign n23168 = n23145 & ~n23167 ;
  assign n23169 = n23165 | n23168 ;
  assign n23170 = n22500 | n22520 ;
  assign n23171 = ( n22500 & n22503 ) | ( n22500 & n23170 ) | ( n22503 & n23170 ) ;
  assign n23172 = n23169 | n23171 ;
  assign n23173 = n23169 & n23171 ;
  assign n23174 = n23172 & ~n23173 ;
  assign n23175 = x96 & n7566 ;
  assign n23176 = x95 & n7561 ;
  assign n23177 = x94 & ~n7560 ;
  assign n23178 = n7953 & n23177 ;
  assign n23179 = n23176 | n23178 ;
  assign n23180 = n23175 | n23179 ;
  assign n23181 = n7569 | n23175 ;
  assign n23182 = n23179 | n23181 ;
  assign n23183 = ( n5202 & n23180 ) | ( n5202 & n23182 ) | ( n23180 & n23182 ) ;
  assign n23184 = x41 & n23182 ;
  assign n23185 = x41 & n23175 ;
  assign n23186 = ( x41 & n23179 ) | ( x41 & n23185 ) | ( n23179 & n23185 ) ;
  assign n23187 = ( n5202 & n23184 ) | ( n5202 & n23186 ) | ( n23184 & n23186 ) ;
  assign n23188 = x41 & ~n23186 ;
  assign n23189 = x41 & ~n23182 ;
  assign n23190 = ( ~n5202 & n23188 ) | ( ~n5202 & n23189 ) | ( n23188 & n23189 ) ;
  assign n23191 = ( n23183 & ~n23187 ) | ( n23183 & n23190 ) | ( ~n23187 & n23190 ) ;
  assign n23192 = n23174 | n23191 ;
  assign n23193 = n23174 & n23191 ;
  assign n23194 = n23192 & ~n23193 ;
  assign n23195 = n22529 | n22547 ;
  assign n23196 = ( n22529 & n22530 ) | ( n22529 & n23195 ) | ( n22530 & n23195 ) ;
  assign n23197 = n23194 & n23196 ;
  assign n23198 = n23194 | n23196 ;
  assign n23199 = ~n23197 & n23198 ;
  assign n23200 = x99 & n6536 ;
  assign n23201 = x98 & n6531 ;
  assign n23202 = x97 & ~n6530 ;
  assign n23203 = n6871 & n23202 ;
  assign n23204 = n23201 | n23203 ;
  assign n23205 = n23200 | n23204 ;
  assign n23206 = n6539 | n23200 ;
  assign n23207 = n23204 | n23206 ;
  assign n23208 = ( n6164 & n23205 ) | ( n6164 & n23207 ) | ( n23205 & n23207 ) ;
  assign n23209 = x38 & n23207 ;
  assign n23210 = x38 & n23200 ;
  assign n23211 = ( x38 & n23204 ) | ( x38 & n23210 ) | ( n23204 & n23210 ) ;
  assign n23212 = ( n6164 & n23209 ) | ( n6164 & n23211 ) | ( n23209 & n23211 ) ;
  assign n23213 = x38 & ~n23211 ;
  assign n23214 = x38 & ~n23207 ;
  assign n23215 = ( ~n6164 & n23213 ) | ( ~n6164 & n23214 ) | ( n23213 & n23214 ) ;
  assign n23216 = ( n23208 & ~n23212 ) | ( n23208 & n23215 ) | ( ~n23212 & n23215 ) ;
  assign n23217 = n23199 & ~n23216 ;
  assign n23218 = n23199 | n23216 ;
  assign n23219 = ( ~n23199 & n23217 ) | ( ~n23199 & n23218 ) | ( n23217 & n23218 ) ;
  assign n23220 = n22550 | n22578 ;
  assign n23221 = ( n22552 & n22578 ) | ( n22552 & n23220 ) | ( n22578 & n23220 ) ;
  assign n23222 = ( n22553 & n22555 ) | ( n22553 & n23221 ) | ( n22555 & n23221 ) ;
  assign n23223 = n23219 | n23222 ;
  assign n23224 = n23219 & n23222 ;
  assign n23225 = n23223 & ~n23224 ;
  assign n23226 = ( n22963 & n22985 ) | ( n22963 & ~n23225 ) | ( n22985 & ~n23225 ) ;
  assign n23227 = ( ~n22985 & n23225 ) | ( ~n22985 & n23226 ) | ( n23225 & n23226 ) ;
  assign n23228 = ( ~n22963 & n23226 ) | ( ~n22963 & n23227 ) | ( n23226 & n23227 ) ;
  assign n23229 = ~n22609 & n22942 ;
  assign n23230 = ~n22330 & n22942 ;
  assign n23231 = ( ~n22331 & n23229 ) | ( ~n22331 & n23230 ) | ( n23229 & n23230 ) ;
  assign n23232 = n23228 & n23231 ;
  assign n23233 = ( n22946 & n23228 ) | ( n22946 & n23232 ) | ( n23228 & n23232 ) ;
  assign n23234 = n23228 | n23231 ;
  assign n23235 = n22946 | n23234 ;
  assign n23236 = ~n23233 & n23235 ;
  assign n23237 = n22916 & ~n22917 ;
  assign n23238 = ( ~n22630 & n22916 ) | ( ~n22630 & n23237 ) | ( n22916 & n23237 ) ;
  assign n23239 = ~n22895 & n23238 ;
  assign n23240 = ~n22611 & n23237 ;
  assign n23241 = ~n22611 & n22916 ;
  assign n23242 = ( ~n22630 & n23240 ) | ( ~n22630 & n23241 ) | ( n23240 & n23241 ) ;
  assign n23243 = ( ~n22892 & n23239 ) | ( ~n22892 & n23242 ) | ( n23239 & n23242 ) ;
  assign n23244 = n23236 & n23243 ;
  assign n23245 = ( n22924 & n23236 ) | ( n22924 & n23244 ) | ( n23236 & n23244 ) ;
  assign n23246 = n23236 | n23243 ;
  assign n23247 = n22924 | n23246 ;
  assign n23248 = ~n23245 & n23247 ;
  assign n23249 = n22890 | n23248 ;
  assign n23250 = n22890 & n23248 ;
  assign n23251 = n23249 & ~n23250 ;
  assign n23252 = n21841 & n22265 ;
  assign n23253 = n22265 & n22269 ;
  assign n23254 = n22265 & n22266 ;
  assign n23255 = ( n20962 & n23253 ) | ( n20962 & n23254 ) | ( n23253 & n23254 ) ;
  assign n23256 = ( n21591 & n23252 ) | ( n21591 & n23255 ) | ( n23252 & n23255 ) ;
  assign n23257 = ( n21563 & n23252 ) | ( n21563 & n23255 ) | ( n23252 & n23255 ) ;
  assign n23258 = ( n21586 & n23256 ) | ( n21586 & n23257 ) | ( n23256 & n23257 ) ;
  assign n23259 = ( n22265 & n22282 ) | ( n22265 & n23258 ) | ( n22282 & n23258 ) ;
  assign n23260 = n22283 & ~n23259 ;
  assign n23261 = n22265 & ~n23252 ;
  assign n23262 = n22265 & ~n23253 ;
  assign n23263 = n22265 & ~n23254 ;
  assign n23264 = ( ~n20962 & n23262 ) | ( ~n20962 & n23263 ) | ( n23262 & n23263 ) ;
  assign n23265 = ( ~n21591 & n23261 ) | ( ~n21591 & n23264 ) | ( n23261 & n23264 ) ;
  assign n23266 = ( ~n21563 & n23261 ) | ( ~n21563 & n23264 ) | ( n23261 & n23264 ) ;
  assign n23267 = ( ~n21586 & n23265 ) | ( ~n21586 & n23266 ) | ( n23265 & n23266 ) ;
  assign n23268 = n22636 & n23267 ;
  assign n23269 = ~n22282 & n23268 ;
  assign n23270 = n23259 | n23269 ;
  assign n23271 = n22636 | n23259 ;
  assign n23272 = ( n23260 & n23270 ) | ( n23260 & n23271 ) | ( n23270 & n23271 ) ;
  assign n23274 = x116 & n1854 ;
  assign n23275 = x115 & ~n1853 ;
  assign n23276 = n2037 & n23275 ;
  assign n23277 = n23274 | n23276 ;
  assign n23273 = x117 & n1859 ;
  assign n23279 = n1862 | n23273 ;
  assign n23280 = n23277 | n23279 ;
  assign n23278 = n23273 | n23277 ;
  assign n23281 = n23278 & n23280 ;
  assign n23282 = ( ~n13522 & n23280 ) | ( ~n13522 & n23281 ) | ( n23280 & n23281 ) ;
  assign n23283 = n23280 & n23281 ;
  assign n23284 = ( n13503 & n23282 ) | ( n13503 & n23283 ) | ( n23282 & n23283 ) ;
  assign n23285 = x20 & n23284 ;
  assign n23286 = x20 & ~n23284 ;
  assign n23287 = ( n23284 & ~n23285 ) | ( n23284 & n23286 ) | ( ~n23285 & n23286 ) ;
  assign n23288 = n23258 & n23287 ;
  assign n23289 = n22265 & n23287 ;
  assign n23290 = ( n22282 & n23288 ) | ( n22282 & n23289 ) | ( n23288 & n23289 ) ;
  assign n23291 = ( n23269 & n23287 ) | ( n23269 & n23290 ) | ( n23287 & n23290 ) ;
  assign n23292 = ( n22636 & n23287 ) | ( n22636 & n23290 ) | ( n23287 & n23290 ) ;
  assign n23293 = ( n23260 & n23291 ) | ( n23260 & n23292 ) | ( n23291 & n23292 ) ;
  assign n23294 = n23272 & ~n23293 ;
  assign n23295 = n23287 & ~n23289 ;
  assign n23296 = ~n23258 & n23287 ;
  assign n23297 = ( ~n22282 & n23295 ) | ( ~n22282 & n23296 ) | ( n23295 & n23296 ) ;
  assign n23298 = ~n23269 & n23297 ;
  assign n23299 = ~n22636 & n23297 ;
  assign n23300 = ( ~n23260 & n23298 ) | ( ~n23260 & n23299 ) | ( n23298 & n23299 ) ;
  assign n23301 = n23251 & n23300 ;
  assign n23302 = ( n23251 & n23294 ) | ( n23251 & n23301 ) | ( n23294 & n23301 ) ;
  assign n23303 = n23251 | n23300 ;
  assign n23304 = n23294 | n23303 ;
  assign n23305 = ~n23302 & n23304 ;
  assign n23306 = ~n22871 & n23305 ;
  assign n23307 = ( n22247 & n22251 ) | ( n22247 & n22648 ) | ( n22251 & n22648 ) ;
  assign n23308 = n22864 | n23305 ;
  assign n23309 = ( n23305 & n23307 ) | ( n23305 & n23308 ) | ( n23307 & n23308 ) ;
  assign n23310 = n22870 & ~n23309 ;
  assign n23311 = n23306 | n23310 ;
  assign n23312 = x123 & n962 ;
  assign n23313 = x122 & n957 ;
  assign n23314 = x121 & ~n956 ;
  assign n23315 = n1105 & n23314 ;
  assign n23316 = n23313 | n23315 ;
  assign n23317 = n23312 | n23316 ;
  assign n23318 = n965 | n23312 ;
  assign n23319 = n23316 | n23318 ;
  assign n23320 = ( n16086 & n23317 ) | ( n16086 & n23319 ) | ( n23317 & n23319 ) ;
  assign n23321 = x14 & n23319 ;
  assign n23322 = x14 & n23312 ;
  assign n23323 = ( x14 & n23316 ) | ( x14 & n23322 ) | ( n23316 & n23322 ) ;
  assign n23324 = ( n16086 & n23321 ) | ( n16086 & n23323 ) | ( n23321 & n23323 ) ;
  assign n23325 = x14 & ~n23323 ;
  assign n23326 = x14 & ~n23319 ;
  assign n23327 = ( ~n16086 & n23325 ) | ( ~n16086 & n23326 ) | ( n23325 & n23326 ) ;
  assign n23328 = ( n23320 & ~n23324 ) | ( n23320 & n23327 ) | ( ~n23324 & n23327 ) ;
  assign n23329 = n22650 | n22704 ;
  assign n23330 = ( n22704 & n22705 ) | ( n22704 & n23329 ) | ( n22705 & n23329 ) ;
  assign n23331 = ( n23311 & n23328 ) | ( n23311 & ~n23330 ) | ( n23328 & ~n23330 ) ;
  assign n23332 = ( ~n23328 & n23330 ) | ( ~n23328 & n23331 ) | ( n23330 & n23331 ) ;
  assign n23333 = ( ~n23311 & n23331 ) | ( ~n23311 & n23332 ) | ( n23331 & n23332 ) ;
  assign n23334 = n22843 | n23331 ;
  assign n23335 = ~n22843 & n23311 ;
  assign n23336 = ( n23332 & n23334 ) | ( n23332 & ~n23335 ) | ( n23334 & ~n23335 ) ;
  assign n23337 = ( ~n22825 & n23333 ) | ( ~n22825 & n23336 ) | ( n23333 & n23336 ) ;
  assign n23338 = ( ~n22672 & n23333 ) | ( ~n22672 & n23336 ) | ( n23333 & n23336 ) ;
  assign n23339 = ( ~n22678 & n23337 ) | ( ~n22678 & n23338 ) | ( n23337 & n23338 ) ;
  assign n23340 = n22847 | n23339 ;
  assign n23341 = n22843 & n23331 ;
  assign n23342 = n22843 & ~n23311 ;
  assign n23343 = ( n23332 & n23341 ) | ( n23332 & n23342 ) | ( n23341 & n23342 ) ;
  assign n23344 = ~n22825 & n23343 ;
  assign n23345 = ~n22672 & n23343 ;
  assign n23346 = ( ~n22678 & n23344 ) | ( ~n22678 & n23345 ) | ( n23344 & n23345 ) ;
  assign n23347 = ( n22847 & n23333 ) | ( n22847 & n23346 ) | ( n23333 & n23346 ) ;
  assign n23348 = n23340 & ~n23347 ;
  assign n23349 = n22815 & n23348 ;
  assign n23350 = ~n22817 & n23349 ;
  assign n23351 = ( n22819 & n23348 ) | ( n22819 & n23350 ) | ( n23348 & n23350 ) ;
  assign n23352 = n22815 | n23348 ;
  assign n23353 = ( ~n22817 & n23348 ) | ( ~n22817 & n23352 ) | ( n23348 & n23352 ) ;
  assign n23354 = n22819 | n23353 ;
  assign n23355 = ~n23351 & n23354 ;
  assign n23356 = n22783 | n22796 ;
  assign n23357 = n22708 & n22755 ;
  assign n23358 = n22708 | n22755 ;
  assign n23359 = ~n23357 & n23358 ;
  assign n23360 = n22723 | n23359 ;
  assign n23361 = ( n22725 & n23359 ) | ( n22725 & n23360 ) | ( n23359 & n23360 ) ;
  assign n23362 = ( n22726 & n22728 ) | ( n22726 & n23361 ) | ( n22728 & n23361 ) ;
  assign n23363 = ( n23355 & ~n23356 ) | ( n23355 & n23362 ) | ( ~n23356 & n23362 ) ;
  assign n23364 = ( n23356 & ~n23362 ) | ( n23356 & n23363 ) | ( ~n23362 & n23363 ) ;
  assign n23365 = ( ~n23355 & n23363 ) | ( ~n23355 & n23364 ) | ( n23363 & n23364 ) ;
  assign n23366 = x127 & n636 ;
  assign n23367 = x126 & n631 ;
  assign n23368 = x125 & ~n630 ;
  assign n23369 = n764 & n23368 ;
  assign n23370 = n23367 | n23369 ;
  assign n23371 = n23366 | n23370 ;
  assign n23372 = n639 | n23366 ;
  assign n23373 = n23370 | n23372 ;
  assign n23374 = ( n18763 & n23371 ) | ( n18763 & n23373 ) | ( n23371 & n23373 ) ;
  assign n23375 = x11 & n23373 ;
  assign n23376 = x11 & n23366 ;
  assign n23377 = ( x11 & n23370 ) | ( x11 & n23376 ) | ( n23370 & n23376 ) ;
  assign n23378 = ( n18763 & n23375 ) | ( n18763 & n23377 ) | ( n23375 & n23377 ) ;
  assign n23379 = x11 & ~n23377 ;
  assign n23380 = x11 & ~n23373 ;
  assign n23381 = ( ~n18763 & n23379 ) | ( ~n18763 & n23380 ) | ( n23379 & n23380 ) ;
  assign n23382 = ( n23374 & ~n23378 ) | ( n23374 & n23381 ) | ( ~n23378 & n23381 ) ;
  assign n23383 = n23293 | n23302 ;
  assign n23384 = x118 & n1859 ;
  assign n23385 = x117 & n1854 ;
  assign n23386 = x116 & ~n1853 ;
  assign n23387 = n2037 & n23386 ;
  assign n23388 = n23385 | n23387 ;
  assign n23389 = n23384 | n23388 ;
  assign n23390 = n1862 | n23384 ;
  assign n23391 = n23388 | n23390 ;
  assign n23392 = ( ~n14002 & n23389 ) | ( ~n14002 & n23391 ) | ( n23389 & n23391 ) ;
  assign n23393 = n23389 & n23391 ;
  assign n23394 = ( n13981 & n23392 ) | ( n13981 & n23393 ) | ( n23392 & n23393 ) ;
  assign n23395 = x20 & n23394 ;
  assign n23396 = x20 & ~n23394 ;
  assign n23397 = ( n23394 & ~n23395 ) | ( n23394 & n23396 ) | ( ~n23395 & n23396 ) ;
  assign n23398 = n23287 & n23397 ;
  assign n23399 = n23288 & n23397 ;
  assign n23400 = n23289 & n23397 ;
  assign n23401 = ( n22282 & n23399 ) | ( n22282 & n23400 ) | ( n23399 & n23400 ) ;
  assign n23402 = ( n23269 & n23398 ) | ( n23269 & n23401 ) | ( n23398 & n23401 ) ;
  assign n23403 = ( n22636 & n23398 ) | ( n22636 & n23401 ) | ( n23398 & n23401 ) ;
  assign n23404 = ( n23260 & n23402 ) | ( n23260 & n23403 ) | ( n23402 & n23403 ) ;
  assign n23405 = ( n23302 & n23397 ) | ( n23302 & n23404 ) | ( n23397 & n23404 ) ;
  assign n23406 = n23383 & ~n23405 ;
  assign n23407 = x115 & n2429 ;
  assign n23408 = x114 & n2424 ;
  assign n23409 = x113 & ~n2423 ;
  assign n23410 = n2631 & n23409 ;
  assign n23411 = n23408 | n23410 ;
  assign n23412 = n23407 | n23411 ;
  assign n23413 = n2432 | n23407 ;
  assign n23414 = n23411 | n23413 ;
  assign n23415 = ( ~n12550 & n23412 ) | ( ~n12550 & n23414 ) | ( n23412 & n23414 ) ;
  assign n23416 = n23412 & n23414 ;
  assign n23417 = ( n12532 & n23415 ) | ( n12532 & n23416 ) | ( n23415 & n23416 ) ;
  assign n23418 = x23 & n23417 ;
  assign n23419 = x23 & ~n23417 ;
  assign n23420 = ( n23417 & ~n23418 ) | ( n23417 & n23419 ) | ( ~n23418 & n23419 ) ;
  assign n23421 = n22885 | n23248 ;
  assign n23422 = ( n22887 & n23248 ) | ( n22887 & n23421 ) | ( n23248 & n23421 ) ;
  assign n23423 = n23420 & n23422 ;
  assign n23424 = n22889 & n23420 ;
  assign n23425 = ( n22890 & n23423 ) | ( n22890 & n23424 ) | ( n23423 & n23424 ) ;
  assign n23426 = n23420 | n23422 ;
  assign n23427 = n22889 | n23420 ;
  assign n23428 = ( n22890 & n23426 ) | ( n22890 & n23427 ) | ( n23426 & n23427 ) ;
  assign n23429 = ~n23425 & n23428 ;
  assign n23430 = x112 & n3085 ;
  assign n23431 = x111 & n3080 ;
  assign n23432 = x110 & ~n3079 ;
  assign n23433 = n3309 & n23432 ;
  assign n23434 = n23431 | n23433 ;
  assign n23435 = n23430 | n23434 ;
  assign n23436 = n3088 | n23430 ;
  assign n23437 = n23434 | n23436 ;
  assign n23438 = ( n11172 & n23435 ) | ( n11172 & n23437 ) | ( n23435 & n23437 ) ;
  assign n23439 = x26 & n23437 ;
  assign n23440 = x26 & n23430 ;
  assign n23441 = ( x26 & n23434 ) | ( x26 & n23440 ) | ( n23434 & n23440 ) ;
  assign n23442 = ( n11172 & n23439 ) | ( n11172 & n23441 ) | ( n23439 & n23441 ) ;
  assign n23443 = x26 & ~n23441 ;
  assign n23444 = x26 & ~n23437 ;
  assign n23445 = ( ~n11172 & n23443 ) | ( ~n11172 & n23444 ) | ( n23443 & n23444 ) ;
  assign n23446 = ( n23438 & ~n23442 ) | ( n23438 & n23445 ) | ( ~n23442 & n23445 ) ;
  assign n23447 = n22923 & n23446 ;
  assign n23448 = ( n23245 & n23446 ) | ( n23245 & n23447 ) | ( n23446 & n23447 ) ;
  assign n23449 = n22923 | n23446 ;
  assign n23450 = n23245 | n23449 ;
  assign n23451 = ~n23448 & n23450 ;
  assign n23452 = x109 & n3816 ;
  assign n23453 = x108 & n3811 ;
  assign n23454 = x107 & ~n3810 ;
  assign n23455 = n4067 & n23454 ;
  assign n23456 = n23453 | n23455 ;
  assign n23457 = n23452 | n23456 ;
  assign n23458 = n3819 | n23452 ;
  assign n23459 = n23456 | n23458 ;
  assign n23460 = ( n9878 & n23457 ) | ( n9878 & n23459 ) | ( n23457 & n23459 ) ;
  assign n23461 = x29 & n23459 ;
  assign n23462 = x29 & n23452 ;
  assign n23463 = ( x29 & n23456 ) | ( x29 & n23462 ) | ( n23456 & n23462 ) ;
  assign n23464 = ( n9878 & n23461 ) | ( n9878 & n23463 ) | ( n23461 & n23463 ) ;
  assign n23465 = x29 & ~n23463 ;
  assign n23466 = x29 & ~n23459 ;
  assign n23467 = ( ~n9878 & n23465 ) | ( ~n9878 & n23466 ) | ( n23465 & n23466 ) ;
  assign n23468 = ( n23460 & ~n23464 ) | ( n23460 & n23467 ) | ( ~n23464 & n23467 ) ;
  assign n23470 = n22963 & n23225 ;
  assign n23471 = n22963 | n23225 ;
  assign n23472 = ~n23470 & n23471 ;
  assign n23473 = n22980 | n23472 ;
  assign n23474 = ( n22982 & n23472 ) | ( n22982 & n23473 ) | ( n23472 & n23473 ) ;
  assign n23475 = ( n22984 & n22985 ) | ( n22984 & n23474 ) | ( n22985 & n23474 ) ;
  assign n23476 = x106 & n4631 ;
  assign n23477 = x105 & n4626 ;
  assign n23478 = x104 & ~n4625 ;
  assign n23479 = n4943 & n23478 ;
  assign n23480 = n23477 | n23479 ;
  assign n23481 = n23476 | n23480 ;
  assign n23482 = n4634 | n23476 ;
  assign n23483 = n23480 | n23482 ;
  assign n23484 = ( n8656 & n23481 ) | ( n8656 & n23483 ) | ( n23481 & n23483 ) ;
  assign n23485 = x32 & n23483 ;
  assign n23486 = x32 & n23476 ;
  assign n23487 = ( x32 & n23480 ) | ( x32 & n23486 ) | ( n23480 & n23486 ) ;
  assign n23488 = ( n8656 & n23485 ) | ( n8656 & n23487 ) | ( n23485 & n23487 ) ;
  assign n23489 = x32 & ~n23487 ;
  assign n23490 = x32 & ~n23483 ;
  assign n23491 = ( ~n8656 & n23489 ) | ( ~n8656 & n23490 ) | ( n23489 & n23490 ) ;
  assign n23492 = ( n23484 & ~n23488 ) | ( n23484 & n23491 ) | ( ~n23488 & n23491 ) ;
  assign n23493 = n23474 & n23492 ;
  assign n23494 = n22984 & n23492 ;
  assign n23495 = ( n22985 & n23493 ) | ( n22985 & n23494 ) | ( n23493 & n23494 ) ;
  assign n23496 = n23475 & ~n23495 ;
  assign n23691 = ( n23146 & n23147 ) | ( n23146 & n23167 ) | ( n23147 & n23167 ) ;
  assign n23497 = x73 & n18290 ;
  assign n23498 = x63 & x72 ;
  assign n23499 = ~n18290 & n23498 ;
  assign n23500 = n23497 | n23499 ;
  assign n23501 = x8 & n22989 ;
  assign n23502 = x8 | n22989 ;
  assign n23503 = ~n23501 & n23502 ;
  assign n23504 = n23500 & ~n23503 ;
  assign n23505 = ~n23500 & n23503 ;
  assign n23506 = n23504 | n23505 ;
  assign n23507 = n22991 & ~n23506 ;
  assign n23508 = ( n23000 & n23506 ) | ( n23000 & ~n23507 ) | ( n23506 & ~n23507 ) ;
  assign n23509 = ~n22991 & n23506 ;
  assign n23510 = n23000 & n23509 ;
  assign n23511 = n23508 & ~n23510 ;
  assign n23512 = x76 & n17146 ;
  assign n23513 = x75 & n17141 ;
  assign n23514 = x74 & ~n17140 ;
  assign n23515 = n17724 & n23514 ;
  assign n23516 = n23513 | n23515 ;
  assign n23517 = n23512 | n23516 ;
  assign n23518 = n17149 | n23512 ;
  assign n23519 = n23516 | n23518 ;
  assign n23520 = ( n923 & n23517 ) | ( n923 & n23519 ) | ( n23517 & n23519 ) ;
  assign n23521 = x62 & n23519 ;
  assign n23522 = x62 & n23512 ;
  assign n23523 = ( x62 & n23516 ) | ( x62 & n23522 ) | ( n23516 & n23522 ) ;
  assign n23524 = ( n923 & n23521 ) | ( n923 & n23523 ) | ( n23521 & n23523 ) ;
  assign n23525 = x62 & ~n23523 ;
  assign n23526 = x62 & ~n23519 ;
  assign n23527 = ( ~n923 & n23525 ) | ( ~n923 & n23526 ) | ( n23525 & n23526 ) ;
  assign n23528 = ( n23520 & ~n23524 ) | ( n23520 & n23527 ) | ( ~n23524 & n23527 ) ;
  assign n23529 = n23511 & ~n23528 ;
  assign n23530 = ~n23511 & n23528 ;
  assign n23531 = n23529 | n23530 ;
  assign n23532 = x79 & n15552 ;
  assign n23533 = x78 & n15547 ;
  assign n23534 = x77 & ~n15546 ;
  assign n23535 = n16123 & n23534 ;
  assign n23536 = n23533 | n23535 ;
  assign n23537 = n23532 | n23536 ;
  assign n23538 = n15555 | n23532 ;
  assign n23539 = n23536 | n23538 ;
  assign n23540 = ( n1332 & n23537 ) | ( n1332 & n23539 ) | ( n23537 & n23539 ) ;
  assign n23541 = x59 & n23539 ;
  assign n23542 = x59 & n23532 ;
  assign n23543 = ( x59 & n23536 ) | ( x59 & n23542 ) | ( n23536 & n23542 ) ;
  assign n23544 = ( n1332 & n23541 ) | ( n1332 & n23543 ) | ( n23541 & n23543 ) ;
  assign n23545 = x59 & ~n23543 ;
  assign n23546 = x59 & ~n23539 ;
  assign n23547 = ( ~n1332 & n23545 ) | ( ~n1332 & n23546 ) | ( n23545 & n23546 ) ;
  assign n23548 = ( n23540 & ~n23544 ) | ( n23540 & n23547 ) | ( ~n23544 & n23547 ) ;
  assign n23549 = n23531 & n23548 ;
  assign n23550 = n23531 | n23548 ;
  assign n23551 = ~n23549 & n23550 ;
  assign n23552 = ( n23003 & n23020 ) | ( n23003 & n23040 ) | ( n23020 & n23040 ) ;
  assign n23553 = n23551 | n23552 ;
  assign n23554 = n23551 & n23552 ;
  assign n23555 = n23553 & ~n23554 ;
  assign n23556 = x82 & n14045 ;
  assign n23557 = x81 & n14040 ;
  assign n23558 = x80 & ~n14039 ;
  assign n23559 = n14552 & n23558 ;
  assign n23560 = n23557 | n23559 ;
  assign n23561 = n23556 | n23560 ;
  assign n23562 = n14048 | n23556 ;
  assign n23563 = n23560 | n23562 ;
  assign n23564 = ( n1811 & n23561 ) | ( n1811 & n23563 ) | ( n23561 & n23563 ) ;
  assign n23565 = x56 & n23563 ;
  assign n23566 = x56 & n23556 ;
  assign n23567 = ( x56 & n23560 ) | ( x56 & n23566 ) | ( n23560 & n23566 ) ;
  assign n23568 = ( n1811 & n23565 ) | ( n1811 & n23567 ) | ( n23565 & n23567 ) ;
  assign n23569 = x56 & ~n23567 ;
  assign n23570 = x56 & ~n23563 ;
  assign n23571 = ( ~n1811 & n23569 ) | ( ~n1811 & n23570 ) | ( n23569 & n23570 ) ;
  assign n23572 = ( n23564 & ~n23568 ) | ( n23564 & n23571 ) | ( ~n23568 & n23571 ) ;
  assign n23573 = n23555 & n23572 ;
  assign n23574 = n23555 & ~n23573 ;
  assign n23576 = ( n23048 & n23049 ) | ( n23048 & n23071 ) | ( n23049 & n23071 ) ;
  assign n23575 = ~n23555 & n23572 ;
  assign n23577 = n23575 & n23576 ;
  assign n23578 = ( n23574 & n23576 ) | ( n23574 & n23577 ) | ( n23576 & n23577 ) ;
  assign n23579 = n23575 | n23576 ;
  assign n23580 = n23574 | n23579 ;
  assign n23581 = ~n23578 & n23580 ;
  assign n23582 = x85 & n12574 ;
  assign n23583 = x84 & n12569 ;
  assign n23584 = x83 & ~n12568 ;
  assign n23585 = n13076 & n23584 ;
  assign n23586 = n23583 | n23585 ;
  assign n23587 = n23582 | n23586 ;
  assign n23588 = n12577 | n23582 ;
  assign n23589 = n23586 | n23588 ;
  assign n23590 = ( n2381 & n23587 ) | ( n2381 & n23589 ) | ( n23587 & n23589 ) ;
  assign n23591 = x53 & n23589 ;
  assign n23592 = x53 & n23582 ;
  assign n23593 = ( x53 & n23586 ) | ( x53 & n23592 ) | ( n23586 & n23592 ) ;
  assign n23594 = ( n2381 & n23591 ) | ( n2381 & n23593 ) | ( n23591 & n23593 ) ;
  assign n23595 = x53 & ~n23593 ;
  assign n23596 = x53 & ~n23589 ;
  assign n23597 = ( ~n2381 & n23595 ) | ( ~n2381 & n23596 ) | ( n23595 & n23596 ) ;
  assign n23598 = ( n23590 & ~n23594 ) | ( n23590 & n23597 ) | ( ~n23594 & n23597 ) ;
  assign n23599 = n23581 & n23598 ;
  assign n23600 = n23581 & ~n23599 ;
  assign n23601 = n23075 | n23095 ;
  assign n23602 = ( n23073 & n23095 ) | ( n23073 & n23601 ) | ( n23095 & n23601 ) ;
  assign n23603 = ( n23077 & n23078 ) | ( n23077 & n23602 ) | ( n23078 & n23602 ) ;
  assign n23604 = ~n23581 & n23598 ;
  assign n23605 = n23603 & n23604 ;
  assign n23606 = ( n23600 & n23603 ) | ( n23600 & n23605 ) | ( n23603 & n23605 ) ;
  assign n23607 = n23603 | n23604 ;
  assign n23608 = n23600 | n23607 ;
  assign n23609 = ~n23606 & n23608 ;
  assign n23610 = x88 & n11205 ;
  assign n23611 = x87 & n11200 ;
  assign n23612 = x86 & ~n11199 ;
  assign n23613 = n11679 & n23612 ;
  assign n23614 = n23611 | n23613 ;
  assign n23615 = n23610 | n23614 ;
  assign n23616 = n11208 | n23610 ;
  assign n23617 = n23614 | n23616 ;
  assign n23618 = ( ~n3039 & n23615 ) | ( ~n3039 & n23617 ) | ( n23615 & n23617 ) ;
  assign n23619 = n23615 & n23617 ;
  assign n23620 = ( n3023 & n23618 ) | ( n3023 & n23619 ) | ( n23618 & n23619 ) ;
  assign n23621 = x50 & n23617 ;
  assign n23622 = x50 & n23610 ;
  assign n23623 = ( x50 & n23614 ) | ( x50 & n23622 ) | ( n23614 & n23622 ) ;
  assign n23624 = ( ~n3039 & n23621 ) | ( ~n3039 & n23623 ) | ( n23621 & n23623 ) ;
  assign n23625 = n23621 & n23623 ;
  assign n23626 = ( n3023 & n23624 ) | ( n3023 & n23625 ) | ( n23624 & n23625 ) ;
  assign n23627 = x50 & ~n23623 ;
  assign n23628 = x50 & ~n23617 ;
  assign n23629 = ( n3039 & n23627 ) | ( n3039 & n23628 ) | ( n23627 & n23628 ) ;
  assign n23630 = n23627 | n23628 ;
  assign n23631 = ( ~n3023 & n23629 ) | ( ~n3023 & n23630 ) | ( n23629 & n23630 ) ;
  assign n23632 = ( n23620 & ~n23626 ) | ( n23620 & n23631 ) | ( ~n23626 & n23631 ) ;
  assign n23633 = n23609 & n23632 ;
  assign n23634 = n23609 & ~n23633 ;
  assign n23635 = ~n23609 & n23632 ;
  assign n23636 = n23098 & n23116 ;
  assign n23637 = n23098 & ~n23636 ;
  assign n23638 = ~n23098 & n23116 ;
  assign n23639 = n23115 | n23116 ;
  assign n23640 = ( n23098 & n23115 ) | ( n23098 & n23639 ) | ( n23115 & n23639 ) ;
  assign n23641 = ( n23636 & n23638 ) | ( n23636 & n23640 ) | ( n23638 & n23640 ) ;
  assign n23642 = n23636 | n23640 ;
  assign n23643 = ( n23637 & n23641 ) | ( n23637 & n23642 ) | ( n23641 & n23642 ) ;
  assign n23644 = ~n23635 & n23643 ;
  assign n23645 = ~n23634 & n23644 ;
  assign n23646 = n23635 & ~n23643 ;
  assign n23647 = ( n23634 & ~n23643 ) | ( n23634 & n23646 ) | ( ~n23643 & n23646 ) ;
  assign n23648 = n23645 | n23647 ;
  assign n23649 = x91 & n9933 ;
  assign n23650 = x90 & n9928 ;
  assign n23651 = x89 & ~n9927 ;
  assign n23652 = n10379 & n23651 ;
  assign n23653 = n23650 | n23652 ;
  assign n23654 = n23649 | n23653 ;
  assign n23655 = n9936 | n23649 ;
  assign n23656 = n23653 | n23655 ;
  assign n23657 = ( n3768 & n23654 ) | ( n3768 & n23656 ) | ( n23654 & n23656 ) ;
  assign n23658 = x47 & n23656 ;
  assign n23659 = x47 & n23649 ;
  assign n23660 = ( x47 & n23653 ) | ( x47 & n23659 ) | ( n23653 & n23659 ) ;
  assign n23661 = ( n3768 & n23658 ) | ( n3768 & n23660 ) | ( n23658 & n23660 ) ;
  assign n23662 = x47 & ~n23660 ;
  assign n23663 = x47 & ~n23656 ;
  assign n23664 = ( ~n3768 & n23662 ) | ( ~n3768 & n23663 ) | ( n23662 & n23663 ) ;
  assign n23665 = ( n23657 & ~n23661 ) | ( n23657 & n23664 ) | ( ~n23661 & n23664 ) ;
  assign n23666 = n23648 & n23665 ;
  assign n23667 = n23648 | n23665 ;
  assign n23668 = ~n23666 & n23667 ;
  assign n23669 = n23121 | n23140 ;
  assign n23670 = ( n23121 & n23123 ) | ( n23121 & n23669 ) | ( n23123 & n23669 ) ;
  assign n23671 = n23668 | n23670 ;
  assign n23672 = n23668 & n23670 ;
  assign n23673 = n23671 & ~n23672 ;
  assign n23674 = x94 & n8724 ;
  assign n23675 = x93 & n8719 ;
  assign n23676 = x92 & ~n8718 ;
  assign n23677 = n9149 & n23676 ;
  assign n23678 = n23675 | n23677 ;
  assign n23679 = n23674 | n23678 ;
  assign n23680 = n8727 | n23674 ;
  assign n23681 = n23678 | n23680 ;
  assign n23682 = ( n4583 & n23679 ) | ( n4583 & n23681 ) | ( n23679 & n23681 ) ;
  assign n23683 = x44 & n23681 ;
  assign n23684 = x44 & n23674 ;
  assign n23685 = ( x44 & n23678 ) | ( x44 & n23684 ) | ( n23678 & n23684 ) ;
  assign n23686 = ( n4583 & n23683 ) | ( n4583 & n23685 ) | ( n23683 & n23685 ) ;
  assign n23687 = x44 & ~n23685 ;
  assign n23688 = x44 & ~n23681 ;
  assign n23689 = ( ~n4583 & n23687 ) | ( ~n4583 & n23688 ) | ( n23687 & n23688 ) ;
  assign n23690 = ( n23682 & ~n23686 ) | ( n23682 & n23689 ) | ( ~n23686 & n23689 ) ;
  assign n23692 = ( n23673 & ~n23690 ) | ( n23673 & n23691 ) | ( ~n23690 & n23691 ) ;
  assign n23693 = ( ~n23673 & n23690 ) | ( ~n23673 & n23691 ) | ( n23690 & n23691 ) ;
  assign n23694 = ( ~n23691 & n23692 ) | ( ~n23691 & n23693 ) | ( n23692 & n23693 ) ;
  assign n23695 = x97 & n7566 ;
  assign n23696 = x96 & n7561 ;
  assign n23697 = x95 & ~n7560 ;
  assign n23698 = n7953 & n23697 ;
  assign n23699 = n23696 | n23698 ;
  assign n23700 = n23695 | n23699 ;
  assign n23701 = n7569 | n23695 ;
  assign n23702 = n23699 | n23701 ;
  assign n23703 = ( n5505 & n23700 ) | ( n5505 & n23702 ) | ( n23700 & n23702 ) ;
  assign n23704 = x41 & n23702 ;
  assign n23705 = x41 & n23695 ;
  assign n23706 = ( x41 & n23699 ) | ( x41 & n23705 ) | ( n23699 & n23705 ) ;
  assign n23707 = ( n5505 & n23704 ) | ( n5505 & n23706 ) | ( n23704 & n23706 ) ;
  assign n23708 = x41 & ~n23706 ;
  assign n23709 = x41 & ~n23702 ;
  assign n23710 = ( ~n5505 & n23708 ) | ( ~n5505 & n23709 ) | ( n23708 & n23709 ) ;
  assign n23711 = ( n23703 & ~n23707 ) | ( n23703 & n23710 ) | ( ~n23707 & n23710 ) ;
  assign n23712 = n23694 & n23711 ;
  assign n23713 = n23694 & ~n23712 ;
  assign n23714 = ~n23694 & n23711 ;
  assign n23715 = n23713 | n23714 ;
  assign n23716 = n23171 | n23191 ;
  assign n23717 = ( n23169 & n23191 ) | ( n23169 & n23716 ) | ( n23191 & n23716 ) ;
  assign n23718 = ( n23173 & n23174 ) | ( n23173 & n23717 ) | ( n23174 & n23717 ) ;
  assign n23719 = ~n23715 & n23718 ;
  assign n23720 = n23715 & ~n23718 ;
  assign n23721 = n23719 | n23720 ;
  assign n23722 = x100 & n6536 ;
  assign n23723 = x99 & n6531 ;
  assign n23724 = x98 & ~n6530 ;
  assign n23725 = n6871 & n23724 ;
  assign n23726 = n23723 | n23725 ;
  assign n23727 = n23722 | n23726 ;
  assign n23728 = n6539 | n23722 ;
  assign n23729 = n23726 | n23728 ;
  assign n23730 = ( n6483 & n23727 ) | ( n6483 & n23729 ) | ( n23727 & n23729 ) ;
  assign n23731 = x38 & n23729 ;
  assign n23732 = x38 & n23722 ;
  assign n23733 = ( x38 & n23726 ) | ( x38 & n23732 ) | ( n23726 & n23732 ) ;
  assign n23734 = ( n6483 & n23731 ) | ( n6483 & n23733 ) | ( n23731 & n23733 ) ;
  assign n23735 = x38 & ~n23733 ;
  assign n23736 = x38 & ~n23729 ;
  assign n23737 = ( ~n6483 & n23735 ) | ( ~n6483 & n23736 ) | ( n23735 & n23736 ) ;
  assign n23738 = ( n23730 & ~n23734 ) | ( n23730 & n23737 ) | ( ~n23734 & n23737 ) ;
  assign n23739 = n23721 & n23738 ;
  assign n23740 = n23721 | n23738 ;
  assign n23741 = ~n23739 & n23740 ;
  assign n23742 = n23196 | n23216 ;
  assign n23743 = ( n23194 & n23216 ) | ( n23194 & n23742 ) | ( n23216 & n23742 ) ;
  assign n23744 = ( n23197 & n23199 ) | ( n23197 & n23743 ) | ( n23199 & n23743 ) ;
  assign n23745 = n23741 | n23744 ;
  assign n23746 = n23741 & n23744 ;
  assign n23747 = n23745 & ~n23746 ;
  assign n23748 = x103 & n5554 ;
  assign n23749 = x102 & n5549 ;
  assign n23750 = x101 & ~n5548 ;
  assign n23751 = n5893 & n23750 ;
  assign n23752 = n23749 | n23751 ;
  assign n23753 = n23748 | n23752 ;
  assign n23754 = n5557 | n23748 ;
  assign n23755 = n23752 | n23754 ;
  assign n23756 = ( n7529 & n23753 ) | ( n7529 & n23755 ) | ( n23753 & n23755 ) ;
  assign n23757 = x35 & n23755 ;
  assign n23758 = x35 & n23748 ;
  assign n23759 = ( x35 & n23752 ) | ( x35 & n23758 ) | ( n23752 & n23758 ) ;
  assign n23760 = ( n7529 & n23757 ) | ( n7529 & n23759 ) | ( n23757 & n23759 ) ;
  assign n23761 = x35 & ~n23759 ;
  assign n23762 = x35 & ~n23755 ;
  assign n23763 = ( ~n7529 & n23761 ) | ( ~n7529 & n23762 ) | ( n23761 & n23762 ) ;
  assign n23764 = ( n23756 & ~n23760 ) | ( n23756 & n23763 ) | ( ~n23760 & n23763 ) ;
  assign n23765 = n23747 & n23764 ;
  assign n23766 = n23747 & ~n23765 ;
  assign n23767 = ~n23747 & n23764 ;
  assign n23768 = n22963 | n23224 ;
  assign n23769 = ( n23224 & n23225 ) | ( n23224 & n23768 ) | ( n23225 & n23768 ) ;
  assign n23770 = ~n23767 & n23769 ;
  assign n23771 = ~n23766 & n23770 ;
  assign n23772 = n23767 & ~n23769 ;
  assign n23773 = ( n23766 & ~n23769 ) | ( n23766 & n23772 ) | ( ~n23769 & n23772 ) ;
  assign n23774 = n23771 | n23773 ;
  assign n23775 = ~n23474 & n23492 ;
  assign n23776 = ~n22984 & n23492 ;
  assign n23777 = ( ~n22985 & n23775 ) | ( ~n22985 & n23776 ) | ( n23775 & n23776 ) ;
  assign n23778 = n23774 & n23777 ;
  assign n23779 = ( n23496 & n23774 ) | ( n23496 & n23778 ) | ( n23774 & n23778 ) ;
  assign n23780 = n23774 | n23777 ;
  assign n23781 = n23496 | n23780 ;
  assign n23782 = ~n23779 & n23781 ;
  assign n23783 = ( ~n22945 & n23468 ) | ( ~n22945 & n23782 ) | ( n23468 & n23782 ) ;
  assign n23784 = n23468 & n23782 ;
  assign n23785 = ( ~n23233 & n23783 ) | ( ~n23233 & n23784 ) | ( n23783 & n23784 ) ;
  assign n23469 = n22945 | n23233 ;
  assign n23786 = ( n23469 & ~n23782 ) | ( n23469 & n23785 ) | ( ~n23782 & n23785 ) ;
  assign n23787 = ( ~n23468 & n23785 ) | ( ~n23468 & n23786 ) | ( n23785 & n23786 ) ;
  assign n23788 = n23451 & ~n23787 ;
  assign n23789 = n23451 | n23787 ;
  assign n23790 = ( ~n23451 & n23788 ) | ( ~n23451 & n23789 ) | ( n23788 & n23789 ) ;
  assign n23791 = n23429 & ~n23790 ;
  assign n23792 = n23429 | n23790 ;
  assign n23793 = ( ~n23429 & n23791 ) | ( ~n23429 & n23792 ) | ( n23791 & n23792 ) ;
  assign n23794 = ( n22636 & n23260 ) | ( n22636 & n23269 ) | ( n23260 & n23269 ) ;
  assign n23795 = n23397 & ~n23401 ;
  assign n23796 = n23397 & ~n23398 ;
  assign n23797 = ( ~n23794 & n23795 ) | ( ~n23794 & n23796 ) | ( n23795 & n23796 ) ;
  assign n23798 = n23793 & n23797 ;
  assign n23799 = ~n23302 & n23798 ;
  assign n23800 = ( n23406 & n23793 ) | ( n23406 & n23799 ) | ( n23793 & n23799 ) ;
  assign n23801 = n23793 | n23797 ;
  assign n23802 = ( ~n23302 & n23793 ) | ( ~n23302 & n23801 ) | ( n23793 & n23801 ) ;
  assign n23803 = n23406 | n23802 ;
  assign n23804 = ~n23800 & n23803 ;
  assign n23805 = x121 & n1383 ;
  assign n23806 = x120 & n1378 ;
  assign n23807 = x119 & ~n1377 ;
  assign n23808 = n1542 & n23807 ;
  assign n23809 = n23806 | n23808 ;
  assign n23810 = n23805 | n23809 ;
  assign n23811 = n1386 | n23805 ;
  assign n23812 = n23809 | n23811 ;
  assign n23813 = ( n15501 & n23810 ) | ( n15501 & n23812 ) | ( n23810 & n23812 ) ;
  assign n23814 = x17 & n23812 ;
  assign n23815 = x17 & n23805 ;
  assign n23816 = ( x17 & n23809 ) | ( x17 & n23815 ) | ( n23809 & n23815 ) ;
  assign n23817 = ( n15501 & n23814 ) | ( n15501 & n23816 ) | ( n23814 & n23816 ) ;
  assign n23818 = x17 & ~n23816 ;
  assign n23819 = x17 & ~n23812 ;
  assign n23820 = ( ~n15501 & n23818 ) | ( ~n15501 & n23819 ) | ( n23818 & n23819 ) ;
  assign n23821 = ( n23813 & ~n23817 ) | ( n23813 & n23820 ) | ( ~n23817 & n23820 ) ;
  assign n23822 = ( n22867 & n22871 ) | ( n22867 & n23309 ) | ( n22871 & n23309 ) ;
  assign n23823 = n23821 | n23822 ;
  assign n23824 = n23821 & n23822 ;
  assign n23825 = n23823 & ~n23824 ;
  assign n23826 = n23328 & n23330 ;
  assign n23827 = n23330 & ~n23826 ;
  assign n23828 = n23311 & n23328 ;
  assign n23829 = ~n23330 & n23828 ;
  assign n23830 = n23826 | n23829 ;
  assign n23831 = n23311 | n23826 ;
  assign n23832 = ( n23827 & n23830 ) | ( n23827 & n23831 ) | ( n23830 & n23831 ) ;
  assign n23833 = x124 & n962 ;
  assign n23834 = x123 & n957 ;
  assign n23835 = x122 & ~n956 ;
  assign n23836 = n1105 & n23835 ;
  assign n23837 = n23834 | n23836 ;
  assign n23838 = n23833 | n23837 ;
  assign n23839 = n965 | n23833 ;
  assign n23840 = n23837 | n23839 ;
  assign n23841 = ( n17084 & n23838 ) | ( n17084 & n23840 ) | ( n23838 & n23840 ) ;
  assign n23842 = x14 & n23840 ;
  assign n23843 = x14 & n23833 ;
  assign n23844 = ( x14 & n23837 ) | ( x14 & n23843 ) | ( n23837 & n23843 ) ;
  assign n23845 = ( n17084 & n23842 ) | ( n17084 & n23844 ) | ( n23842 & n23844 ) ;
  assign n23846 = x14 & ~n23844 ;
  assign n23847 = x14 & ~n23840 ;
  assign n23848 = ( ~n17084 & n23846 ) | ( ~n17084 & n23847 ) | ( n23846 & n23847 ) ;
  assign n23849 = ( n23841 & ~n23845 ) | ( n23841 & n23848 ) | ( ~n23845 & n23848 ) ;
  assign n23850 = n23328 | n23849 ;
  assign n23851 = ( n23330 & n23849 ) | ( n23330 & n23850 ) | ( n23849 & n23850 ) ;
  assign n23852 = n23829 | n23851 ;
  assign n23853 = n23311 | n23851 ;
  assign n23854 = ( n23827 & n23852 ) | ( n23827 & n23853 ) | ( n23852 & n23853 ) ;
  assign n23855 = ~n23849 & n23850 ;
  assign n23856 = n23330 & n23855 ;
  assign n23857 = ( n23829 & ~n23849 ) | ( n23829 & n23856 ) | ( ~n23849 & n23856 ) ;
  assign n23858 = ( n23311 & ~n23849 ) | ( n23311 & n23856 ) | ( ~n23849 & n23856 ) ;
  assign n23859 = ( n23827 & n23857 ) | ( n23827 & n23858 ) | ( n23857 & n23858 ) ;
  assign n23860 = ( ~n23832 & n23854 ) | ( ~n23832 & n23859 ) | ( n23854 & n23859 ) ;
  assign n23861 = ( n23804 & ~n23825 ) | ( n23804 & n23860 ) | ( ~n23825 & n23860 ) ;
  assign n23862 = ( n23825 & ~n23860 ) | ( n23825 & n23861 ) | ( ~n23860 & n23861 ) ;
  assign n23863 = ( ~n23804 & n23861 ) | ( ~n23804 & n23862 ) | ( n23861 & n23862 ) ;
  assign n23864 = n22846 | n23346 ;
  assign n23865 = n22846 | n23333 ;
  assign n23866 = ( n22847 & n23864 ) | ( n22847 & n23865 ) | ( n23864 & n23865 ) ;
  assign n23867 = ( n23382 & n23863 ) | ( n23382 & ~n23866 ) | ( n23863 & ~n23866 ) ;
  assign n23868 = ( ~n23863 & n23866 ) | ( ~n23863 & n23867 ) | ( n23866 & n23867 ) ;
  assign n23869 = ( ~n23382 & n23867 ) | ( ~n23382 & n23868 ) | ( n23867 & n23868 ) ;
  assign n23870 = n22818 & n23869 ;
  assign n23871 = ( n23351 & n23869 ) | ( n23351 & n23870 ) | ( n23869 & n23870 ) ;
  assign n23872 = n22818 | n23350 ;
  assign n23873 = n22818 | n23348 ;
  assign n23874 = ( n22819 & n23872 ) | ( n22819 & n23873 ) | ( n23872 & n23873 ) ;
  assign n23875 = ~n23871 & n23874 ;
  assign n23876 = n23355 & n23362 ;
  assign n23877 = n23362 & ~n23876 ;
  assign n23878 = n23355 & ~n23362 ;
  assign n23879 = n23877 | n23878 ;
  assign n23880 = n22783 & n23879 ;
  assign n23881 = n23876 | n23880 ;
  assign n23882 = n23876 | n23878 ;
  assign n23883 = n23877 | n23882 ;
  assign n23884 = ( n22796 & n23881 ) | ( n22796 & n23883 ) | ( n23881 & n23883 ) ;
  assign n23885 = n23869 & ~n23870 ;
  assign n23886 = ~n23351 & n23885 ;
  assign n23887 = n23884 | n23886 ;
  assign n23888 = n23875 | n23887 ;
  assign n23889 = n23875 | n23886 ;
  assign n23890 = n23883 & n23889 ;
  assign n23891 = n23876 & n23889 ;
  assign n23892 = ( n23880 & n23889 ) | ( n23880 & n23891 ) | ( n23889 & n23891 ) ;
  assign n23893 = ( n22796 & n23890 ) | ( n22796 & n23892 ) | ( n23890 & n23892 ) ;
  assign n23894 = n23888 & ~n23893 ;
  assign n23912 = n23328 & n23849 ;
  assign n23913 = n23330 & n23912 ;
  assign n23914 = ( n23829 & n23849 ) | ( n23829 & n23913 ) | ( n23849 & n23913 ) ;
  assign n23915 = ( n23311 & n23849 ) | ( n23311 & n23913 ) | ( n23849 & n23913 ) ;
  assign n23916 = ( n23827 & n23914 ) | ( n23827 & n23915 ) | ( n23914 & n23915 ) ;
  assign n23909 = n23804 & n23825 ;
  assign n23910 = n23804 | n23825 ;
  assign n23911 = ~n23909 & n23910 ;
  assign n23917 = n23911 | n23916 ;
  assign n23918 = ( n23860 & n23916 ) | ( n23860 & n23917 ) | ( n23916 & n23917 ) ;
  assign n23895 = x127 & n631 ;
  assign n23896 = x126 & ~n630 ;
  assign n23897 = n764 & n23896 ;
  assign n23898 = n23895 | n23897 ;
  assign n23899 = n639 | n23898 ;
  assign n23900 = ( n19328 & n23898 ) | ( n19328 & n23899 ) | ( n23898 & n23899 ) ;
  assign n23901 = x11 & n23898 ;
  assign n23902 = ( x11 & n1532 ) | ( x11 & n23898 ) | ( n1532 & n23898 ) ;
  assign n23903 = ( n19328 & n23901 ) | ( n19328 & n23902 ) | ( n23901 & n23902 ) ;
  assign n23904 = x11 & ~n1532 ;
  assign n23905 = ~n23898 & n23904 ;
  assign n23906 = x11 & ~n23898 ;
  assign n23907 = ( ~n19328 & n23905 ) | ( ~n19328 & n23906 ) | ( n23905 & n23906 ) ;
  assign n23908 = ( n23900 & ~n23903 ) | ( n23900 & n23907 ) | ( ~n23903 & n23907 ) ;
  assign n23919 = n23908 & n23918 ;
  assign n23920 = n23918 & ~n23919 ;
  assign n23938 = n23804 | n23824 ;
  assign n23939 = ( n23824 & n23825 ) | ( n23824 & n23938 ) | ( n23825 & n23938 ) ;
  assign n23921 = x125 & n962 ;
  assign n23922 = x124 & n957 ;
  assign n23923 = x123 & ~n956 ;
  assign n23924 = n1105 & n23923 ;
  assign n23925 = n23922 | n23924 ;
  assign n23926 = n23921 | n23925 ;
  assign n23927 = n965 | n23921 ;
  assign n23928 = n23925 | n23927 ;
  assign n23929 = ( n17670 & n23926 ) | ( n17670 & n23928 ) | ( n23926 & n23928 ) ;
  assign n23930 = x14 & n23928 ;
  assign n23931 = x14 & n23921 ;
  assign n23932 = ( x14 & n23925 ) | ( x14 & n23931 ) | ( n23925 & n23931 ) ;
  assign n23933 = ( n17670 & n23930 ) | ( n17670 & n23932 ) | ( n23930 & n23932 ) ;
  assign n23934 = x14 & ~n23932 ;
  assign n23935 = x14 & ~n23928 ;
  assign n23936 = ( ~n17670 & n23934 ) | ( ~n17670 & n23935 ) | ( n23934 & n23935 ) ;
  assign n23937 = ( n23929 & ~n23933 ) | ( n23929 & n23936 ) | ( ~n23933 & n23936 ) ;
  assign n23940 = n23937 & n23939 ;
  assign n23941 = n23939 & ~n23940 ;
  assign n23942 = n23405 | n23799 ;
  assign n23943 = n23405 | n23793 ;
  assign n23944 = ( n23406 & n23942 ) | ( n23406 & n23943 ) | ( n23942 & n23943 ) ;
  assign n23946 = x121 & n1378 ;
  assign n23947 = x120 & ~n1377 ;
  assign n23948 = n1542 & n23947 ;
  assign n23949 = n23946 | n23948 ;
  assign n23945 = x122 & n1383 ;
  assign n23951 = n1386 | n23945 ;
  assign n23952 = n23949 | n23951 ;
  assign n23950 = n23945 | n23949 ;
  assign n23953 = n23950 & n23952 ;
  assign n23954 = ( n16043 & n23952 ) | ( n16043 & n23953 ) | ( n23952 & n23953 ) ;
  assign n23955 = x17 & n23953 ;
  assign n23956 = x17 & n23952 ;
  assign n23957 = ( n16043 & n23955 ) | ( n16043 & n23956 ) | ( n23955 & n23956 ) ;
  assign n23958 = x17 & ~n23953 ;
  assign n23959 = x17 & ~n23952 ;
  assign n23960 = ( ~n16043 & n23958 ) | ( ~n16043 & n23959 ) | ( n23958 & n23959 ) ;
  assign n23961 = ( n23954 & ~n23957 ) | ( n23954 & n23960 ) | ( ~n23957 & n23960 ) ;
  assign n23962 = n23404 & n23961 ;
  assign n23963 = n23397 & n23961 ;
  assign n23964 = ( n23302 & n23962 ) | ( n23302 & n23963 ) | ( n23962 & n23963 ) ;
  assign n23965 = ( n23799 & n23961 ) | ( n23799 & n23964 ) | ( n23961 & n23964 ) ;
  assign n23966 = ( n23793 & n23961 ) | ( n23793 & n23964 ) | ( n23961 & n23964 ) ;
  assign n23967 = ( n23406 & n23965 ) | ( n23406 & n23966 ) | ( n23965 & n23966 ) ;
  assign n23968 = n23944 & ~n23967 ;
  assign n23969 = n22942 & n23468 ;
  assign n23970 = n22609 & n23969 ;
  assign n23971 = n22330 & n23969 ;
  assign n23972 = ( n22331 & n23970 ) | ( n22331 & n23971 ) | ( n23970 & n23971 ) ;
  assign n23973 = ( n23233 & n23468 ) | ( n23233 & n23972 ) | ( n23468 & n23972 ) ;
  assign n23974 = n23469 & ~n23973 ;
  assign n23975 = n23468 & ~n23969 ;
  assign n23976 = ( ~n22609 & n23468 ) | ( ~n22609 & n23975 ) | ( n23468 & n23975 ) ;
  assign n23977 = ( ~n22330 & n23468 ) | ( ~n22330 & n23975 ) | ( n23468 & n23975 ) ;
  assign n23978 = ( ~n22331 & n23976 ) | ( ~n22331 & n23977 ) | ( n23976 & n23977 ) ;
  assign n23979 = n23782 & n23978 ;
  assign n23980 = ~n23233 & n23979 ;
  assign n23981 = n23973 | n23980 ;
  assign n23982 = n23782 | n23973 ;
  assign n23983 = ( n23974 & n23981 ) | ( n23974 & n23982 ) | ( n23981 & n23982 ) ;
  assign n23984 = x113 & n3085 ;
  assign n23985 = x112 & n3080 ;
  assign n23986 = x111 & ~n3079 ;
  assign n23987 = n3309 & n23986 ;
  assign n23988 = n23985 | n23987 ;
  assign n23989 = n23984 | n23988 ;
  assign n23990 = n3088 | n23984 ;
  assign n23991 = n23988 | n23990 ;
  assign n23992 = ( ~n11642 & n23989 ) | ( ~n11642 & n23991 ) | ( n23989 & n23991 ) ;
  assign n23993 = n23989 & n23991 ;
  assign n23994 = ( n11626 & n23992 ) | ( n11626 & n23993 ) | ( n23992 & n23993 ) ;
  assign n23995 = x26 & n23994 ;
  assign n23996 = x26 & ~n23994 ;
  assign n23997 = ( n23994 & ~n23995 ) | ( n23994 & n23996 ) | ( ~n23995 & n23996 ) ;
  assign n23998 = n23972 & n23997 ;
  assign n23999 = n23468 & n23997 ;
  assign n24000 = ( n23233 & n23998 ) | ( n23233 & n23999 ) | ( n23998 & n23999 ) ;
  assign n24001 = ( n23980 & n23997 ) | ( n23980 & n24000 ) | ( n23997 & n24000 ) ;
  assign n24002 = ( n23782 & n23997 ) | ( n23782 & n24000 ) | ( n23997 & n24000 ) ;
  assign n24003 = ( n23974 & n24001 ) | ( n23974 & n24002 ) | ( n24001 & n24002 ) ;
  assign n24004 = n23983 & ~n24003 ;
  assign n24005 = n23766 | n23767 ;
  assign n24006 = x107 & n4631 ;
  assign n24007 = x106 & n4626 ;
  assign n24008 = x105 & ~n4625 ;
  assign n24009 = n4943 & n24008 ;
  assign n24010 = n24007 | n24009 ;
  assign n24011 = n24006 | n24010 ;
  assign n24012 = n4634 | n24006 ;
  assign n24013 = n24010 | n24012 ;
  assign n24014 = ( n9084 & n24011 ) | ( n9084 & n24013 ) | ( n24011 & n24013 ) ;
  assign n24015 = x32 & n24013 ;
  assign n24016 = x32 & n24006 ;
  assign n24017 = ( x32 & n24010 ) | ( x32 & n24016 ) | ( n24010 & n24016 ) ;
  assign n24018 = ( n9084 & n24015 ) | ( n9084 & n24017 ) | ( n24015 & n24017 ) ;
  assign n24019 = x32 & ~n24017 ;
  assign n24020 = x32 & ~n24013 ;
  assign n24021 = ( ~n9084 & n24019 ) | ( ~n9084 & n24020 ) | ( n24019 & n24020 ) ;
  assign n24022 = ( n24014 & ~n24018 ) | ( n24014 & n24021 ) | ( ~n24018 & n24021 ) ;
  assign n24023 = n23765 | n23769 ;
  assign n24024 = n24022 | n24023 ;
  assign n24025 = n23765 | n24022 ;
  assign n24026 = ( n24005 & n24024 ) | ( n24005 & n24025 ) | ( n24024 & n24025 ) ;
  assign n24027 = n24022 & n24023 ;
  assign n24028 = n23765 & n24022 ;
  assign n24029 = ( n24005 & n24027 ) | ( n24005 & n24028 ) | ( n24027 & n24028 ) ;
  assign n24030 = n24026 & ~n24029 ;
  assign n24279 = ( n23694 & n23711 ) | ( n23694 & n23717 ) | ( n23711 & n23717 ) ;
  assign n24280 = ( n23173 & n23694 ) | ( n23173 & n23711 ) | ( n23694 & n23711 ) ;
  assign n24281 = ( n23174 & n24279 ) | ( n23174 & n24280 ) | ( n24279 & n24280 ) ;
  assign n24031 = n23599 | n23606 ;
  assign n24032 = n23573 | n23578 ;
  assign n24033 = n23548 | n23552 ;
  assign n24034 = ( n23531 & n23552 ) | ( n23531 & n24033 ) | ( n23552 & n24033 ) ;
  assign n24035 = ( n23549 & n23551 ) | ( n23549 & n24034 ) | ( n23551 & n24034 ) ;
  assign n24036 = x76 & n17141 ;
  assign n24037 = x75 & ~n17140 ;
  assign n24038 = n17724 & n24037 ;
  assign n24039 = n24036 | n24038 ;
  assign n24040 = x77 & n17146 ;
  assign n24041 = n17149 | n24040 ;
  assign n24042 = n24039 | n24041 ;
  assign n24043 = ~x62 & n24042 ;
  assign n24044 = ~x62 & n24040 ;
  assign n24045 = ( ~x62 & n24039 ) | ( ~x62 & n24044 ) | ( n24039 & n24044 ) ;
  assign n24046 = ( n1059 & n24043 ) | ( n1059 & n24045 ) | ( n24043 & n24045 ) ;
  assign n24047 = x62 & ~n24042 ;
  assign n24048 = x62 & x77 ;
  assign n24049 = n17146 & n24048 ;
  assign n24050 = x62 & ~n24049 ;
  assign n24051 = ~n24039 & n24050 ;
  assign n24052 = ( ~n1059 & n24047 ) | ( ~n1059 & n24051 ) | ( n24047 & n24051 ) ;
  assign n24053 = n24046 | n24052 ;
  assign n24054 = ( ~x8 & n22989 ) | ( ~x8 & n23500 ) | ( n22989 & n23500 ) ;
  assign n24055 = x74 & n18290 ;
  assign n24056 = x63 & x73 ;
  assign n24057 = ~n18290 & n24056 ;
  assign n24058 = n24055 | n24057 ;
  assign n24059 = n24054 & ~n24058 ;
  assign n24060 = n24054 & ~n24059 ;
  assign n24061 = n24054 | n24058 ;
  assign n24062 = ~n24060 & n24061 ;
  assign n24063 = n24053 & ~n24062 ;
  assign n24064 = ~n24053 & n24062 ;
  assign n24065 = n24063 | n24064 ;
  assign n24066 = ( n22991 & ~n23506 ) | ( n22991 & n23528 ) | ( ~n23506 & n23528 ) ;
  assign n24067 = n23506 & ~n23528 ;
  assign n24068 = ( n23000 & ~n24066 ) | ( n23000 & n24067 ) | ( ~n24066 & n24067 ) ;
  assign n24069 = n24065 | n24068 ;
  assign n24070 = ~n24065 & n24069 ;
  assign n24071 = x80 & n15552 ;
  assign n24072 = x79 & n15547 ;
  assign n24073 = x78 & ~n15546 ;
  assign n24074 = n16123 & n24073 ;
  assign n24075 = n24072 | n24074 ;
  assign n24076 = n24071 | n24075 ;
  assign n24077 = n15555 | n24071 ;
  assign n24078 = n24075 | n24077 ;
  assign n24079 = ( n1499 & n24076 ) | ( n1499 & n24078 ) | ( n24076 & n24078 ) ;
  assign n24080 = x59 & n24078 ;
  assign n24081 = x59 & n24071 ;
  assign n24082 = ( x59 & n24075 ) | ( x59 & n24081 ) | ( n24075 & n24081 ) ;
  assign n24083 = ( n1499 & n24080 ) | ( n1499 & n24082 ) | ( n24080 & n24082 ) ;
  assign n24084 = x59 & ~n24082 ;
  assign n24085 = x59 & ~n24078 ;
  assign n24086 = ( ~n1499 & n24084 ) | ( ~n1499 & n24085 ) | ( n24084 & n24085 ) ;
  assign n24087 = ( n24079 & ~n24083 ) | ( n24079 & n24086 ) | ( ~n24083 & n24086 ) ;
  assign n24088 = n24068 | n24087 ;
  assign n24089 = n24065 & ~n24088 ;
  assign n24090 = ( n24070 & ~n24087 ) | ( n24070 & n24089 ) | ( ~n24087 & n24089 ) ;
  assign n24091 = n24068 & n24087 ;
  assign n24092 = ( ~n24065 & n24087 ) | ( ~n24065 & n24091 ) | ( n24087 & n24091 ) ;
  assign n24093 = ~n24070 & n24092 ;
  assign n24094 = n24034 & n24093 ;
  assign n24095 = n23549 & n24093 ;
  assign n24096 = ( n23551 & n24094 ) | ( n23551 & n24095 ) | ( n24094 & n24095 ) ;
  assign n24097 = ( n24035 & n24090 ) | ( n24035 & n24096 ) | ( n24090 & n24096 ) ;
  assign n24098 = n24090 | n24093 ;
  assign n24099 = n24035 | n24098 ;
  assign n24100 = ~n24097 & n24099 ;
  assign n24101 = x83 & n14045 ;
  assign n24102 = x82 & n14040 ;
  assign n24103 = x81 & ~n14039 ;
  assign n24104 = n14552 & n24103 ;
  assign n24105 = n24102 | n24104 ;
  assign n24106 = n24101 | n24105 ;
  assign n24107 = n14048 | n24101 ;
  assign n24108 = n24105 | n24107 ;
  assign n24109 = ( n2009 & n24106 ) | ( n2009 & n24108 ) | ( n24106 & n24108 ) ;
  assign n24110 = x56 & n24108 ;
  assign n24111 = x56 & n24101 ;
  assign n24112 = ( x56 & n24105 ) | ( x56 & n24111 ) | ( n24105 & n24111 ) ;
  assign n24113 = ( n2009 & n24110 ) | ( n2009 & n24112 ) | ( n24110 & n24112 ) ;
  assign n24114 = x56 & ~n24112 ;
  assign n24115 = x56 & ~n24108 ;
  assign n24116 = ( ~n2009 & n24114 ) | ( ~n2009 & n24115 ) | ( n24114 & n24115 ) ;
  assign n24117 = ( n24109 & ~n24113 ) | ( n24109 & n24116 ) | ( ~n24113 & n24116 ) ;
  assign n24118 = n24098 & ~n24117 ;
  assign n24119 = ( n24035 & ~n24117 ) | ( n24035 & n24118 ) | ( ~n24117 & n24118 ) ;
  assign n24120 = ~n24097 & n24119 ;
  assign n24121 = n24117 | n24120 ;
  assign n24122 = ( ~n24100 & n24120 ) | ( ~n24100 & n24121 ) | ( n24120 & n24121 ) ;
  assign n24123 = n24032 | n24122 ;
  assign n24124 = n24032 & n24122 ;
  assign n24125 = n24123 & ~n24124 ;
  assign n24126 = x86 & n12574 ;
  assign n24127 = x85 & n12569 ;
  assign n24128 = x84 & ~n12568 ;
  assign n24129 = n13076 & n24128 ;
  assign n24130 = n24127 | n24129 ;
  assign n24131 = n24126 | n24130 ;
  assign n24132 = n12577 | n24126 ;
  assign n24133 = n24130 | n24132 ;
  assign n24134 = ( n2606 & n24131 ) | ( n2606 & n24133 ) | ( n24131 & n24133 ) ;
  assign n24135 = x53 & n24133 ;
  assign n24136 = x53 & n24126 ;
  assign n24137 = ( x53 & n24130 ) | ( x53 & n24136 ) | ( n24130 & n24136 ) ;
  assign n24138 = ( n2606 & n24135 ) | ( n2606 & n24137 ) | ( n24135 & n24137 ) ;
  assign n24139 = x53 & ~n24137 ;
  assign n24140 = x53 & ~n24133 ;
  assign n24141 = ( ~n2606 & n24139 ) | ( ~n2606 & n24140 ) | ( n24139 & n24140 ) ;
  assign n24142 = ( n24134 & ~n24138 ) | ( n24134 & n24141 ) | ( ~n24138 & n24141 ) ;
  assign n24143 = ~n24125 & n24142 ;
  assign n24144 = n24031 & n24143 ;
  assign n24145 = n24122 | n24142 ;
  assign n24146 = ( n24032 & n24142 ) | ( n24032 & n24145 ) | ( n24142 & n24145 ) ;
  assign n24147 = n24123 & ~n24146 ;
  assign n24148 = ( n24031 & n24144 ) | ( n24031 & n24147 ) | ( n24144 & n24147 ) ;
  assign n24149 = n24143 | n24147 ;
  assign n24150 = n24031 | n24149 ;
  assign n24151 = ~n24148 & n24150 ;
  assign n24152 = x89 & n11205 ;
  assign n24153 = x88 & n11200 ;
  assign n24154 = x87 & ~n11199 ;
  assign n24155 = n11679 & n24154 ;
  assign n24156 = n24153 | n24155 ;
  assign n24157 = n24152 | n24156 ;
  assign n24158 = n11208 | n24152 ;
  assign n24159 = n24156 | n24158 ;
  assign n24160 = ( n3282 & n24157 ) | ( n3282 & n24159 ) | ( n24157 & n24159 ) ;
  assign n24161 = x50 & n24159 ;
  assign n24162 = x50 & n24152 ;
  assign n24163 = ( x50 & n24156 ) | ( x50 & n24162 ) | ( n24156 & n24162 ) ;
  assign n24164 = ( n3282 & n24161 ) | ( n3282 & n24163 ) | ( n24161 & n24163 ) ;
  assign n24165 = x50 & ~n24163 ;
  assign n24166 = x50 & ~n24159 ;
  assign n24167 = ( ~n3282 & n24165 ) | ( ~n3282 & n24166 ) | ( n24165 & n24166 ) ;
  assign n24168 = ( n24160 & ~n24164 ) | ( n24160 & n24167 ) | ( ~n24164 & n24167 ) ;
  assign n24169 = n24150 & ~n24168 ;
  assign n24170 = ~n24148 & n24169 ;
  assign n24171 = n24168 | n24170 ;
  assign n24172 = ( ~n24151 & n24170 ) | ( ~n24151 & n24171 ) | ( n24170 & n24171 ) ;
  assign n24173 = n23634 | n23635 ;
  assign n24174 = n23633 | n23643 ;
  assign n24175 = ( n23633 & n24173 ) | ( n23633 & n24174 ) | ( n24173 & n24174 ) ;
  assign n24176 = n24172 | n24175 ;
  assign n24177 = n24172 & n24175 ;
  assign n24178 = n24176 & ~n24177 ;
  assign n24179 = x92 & n9933 ;
  assign n24180 = x91 & n9928 ;
  assign n24181 = x90 & ~n9927 ;
  assign n24182 = n10379 & n24181 ;
  assign n24183 = n24180 | n24182 ;
  assign n24184 = n24179 | n24183 ;
  assign n24185 = n9936 | n24179 ;
  assign n24186 = n24183 | n24185 ;
  assign n24187 = ( n4040 & n24184 ) | ( n4040 & n24186 ) | ( n24184 & n24186 ) ;
  assign n24188 = x47 & n24186 ;
  assign n24189 = x47 & n24179 ;
  assign n24190 = ( x47 & n24183 ) | ( x47 & n24189 ) | ( n24183 & n24189 ) ;
  assign n24191 = ( n4040 & n24188 ) | ( n4040 & n24190 ) | ( n24188 & n24190 ) ;
  assign n24192 = x47 & ~n24190 ;
  assign n24193 = x47 & ~n24186 ;
  assign n24194 = ( ~n4040 & n24192 ) | ( ~n4040 & n24193 ) | ( n24192 & n24193 ) ;
  assign n24195 = ( n24187 & ~n24191 ) | ( n24187 & n24194 ) | ( ~n24191 & n24194 ) ;
  assign n24196 = ~n24178 & n24195 ;
  assign n24197 = n24174 | n24195 ;
  assign n24198 = n23633 | n24195 ;
  assign n24199 = ( n24173 & n24197 ) | ( n24173 & n24198 ) | ( n24197 & n24198 ) ;
  assign n24200 = ( n24172 & n24195 ) | ( n24172 & n24199 ) | ( n24195 & n24199 ) ;
  assign n24201 = n24176 & ~n24200 ;
  assign n24202 = n23666 | n23670 ;
  assign n24203 = ( n23666 & n23668 ) | ( n23666 & n24202 ) | ( n23668 & n24202 ) ;
  assign n24204 = n24201 | n24203 ;
  assign n24205 = n24196 | n24204 ;
  assign n24206 = n24201 & n24203 ;
  assign n24207 = ( n24196 & n24203 ) | ( n24196 & n24206 ) | ( n24203 & n24206 ) ;
  assign n24208 = n24205 & ~n24207 ;
  assign n24209 = x95 & n8724 ;
  assign n24210 = x94 & n8719 ;
  assign n24211 = x93 & ~n8718 ;
  assign n24212 = n9149 & n24211 ;
  assign n24213 = n24210 | n24212 ;
  assign n24214 = n24209 | n24213 ;
  assign n24215 = n8727 | n24209 ;
  assign n24216 = n24213 | n24215 ;
  assign n24217 = ( n4897 & n24214 ) | ( n4897 & n24216 ) | ( n24214 & n24216 ) ;
  assign n24218 = x44 & n24216 ;
  assign n24219 = x44 & n24209 ;
  assign n24220 = ( x44 & n24213 ) | ( x44 & n24219 ) | ( n24213 & n24219 ) ;
  assign n24221 = ( n4897 & n24218 ) | ( n4897 & n24220 ) | ( n24218 & n24220 ) ;
  assign n24222 = x44 & ~n24220 ;
  assign n24223 = x44 & ~n24216 ;
  assign n24224 = ( ~n4897 & n24222 ) | ( ~n4897 & n24223 ) | ( n24222 & n24223 ) ;
  assign n24225 = ( n24217 & ~n24221 ) | ( n24217 & n24224 ) | ( ~n24221 & n24224 ) ;
  assign n24226 = n24208 | n24225 ;
  assign n24227 = n24208 & n24225 ;
  assign n24228 = n24226 & ~n24227 ;
  assign n24229 = n23673 | n23690 ;
  assign n24230 = n23691 & n24229 ;
  assign n24231 = n23673 & n23690 ;
  assign n24232 = n24230 | n24231 ;
  assign n24233 = n24228 & n24232 ;
  assign n24234 = n24228 | n24232 ;
  assign n24235 = ~n24233 & n24234 ;
  assign n24236 = x98 & n7566 ;
  assign n24237 = x97 & n7561 ;
  assign n24238 = x96 & ~n7560 ;
  assign n24239 = n7953 & n24238 ;
  assign n24240 = n24237 | n24239 ;
  assign n24241 = n24236 | n24240 ;
  assign n24242 = n7569 | n24236 ;
  assign n24243 = n24240 | n24242 ;
  assign n24244 = ( ~n5850 & n24241 ) | ( ~n5850 & n24243 ) | ( n24241 & n24243 ) ;
  assign n24245 = n24241 & n24243 ;
  assign n24246 = ( n5834 & n24244 ) | ( n5834 & n24245 ) | ( n24244 & n24245 ) ;
  assign n24247 = x41 & n24243 ;
  assign n24248 = x41 & n24236 ;
  assign n24249 = ( x41 & n24240 ) | ( x41 & n24248 ) | ( n24240 & n24248 ) ;
  assign n24250 = ( ~n5850 & n24247 ) | ( ~n5850 & n24249 ) | ( n24247 & n24249 ) ;
  assign n24251 = n24247 & n24249 ;
  assign n24252 = ( n5834 & n24250 ) | ( n5834 & n24251 ) | ( n24250 & n24251 ) ;
  assign n24253 = x41 & ~n24249 ;
  assign n24254 = x41 & ~n24243 ;
  assign n24255 = ( n5850 & n24253 ) | ( n5850 & n24254 ) | ( n24253 & n24254 ) ;
  assign n24256 = n24253 | n24254 ;
  assign n24257 = ( ~n5834 & n24255 ) | ( ~n5834 & n24256 ) | ( n24255 & n24256 ) ;
  assign n24258 = ( n24246 & ~n24252 ) | ( n24246 & n24257 ) | ( ~n24252 & n24257 ) ;
  assign n24259 = n24235 & n24258 ;
  assign n24260 = n24235 | n24258 ;
  assign n24261 = ~n24259 & n24260 ;
  assign n24262 = x101 & n6536 ;
  assign n24263 = x100 & n6531 ;
  assign n24264 = x99 & ~n6530 ;
  assign n24265 = n6871 & n24264 ;
  assign n24266 = n24263 | n24265 ;
  assign n24267 = n24262 | n24266 ;
  assign n24268 = n6539 | n24262 ;
  assign n24269 = n24266 | n24268 ;
  assign n24270 = ( n6844 & n24267 ) | ( n6844 & n24269 ) | ( n24267 & n24269 ) ;
  assign n24271 = x38 & n24269 ;
  assign n24272 = x38 & n24262 ;
  assign n24273 = ( x38 & n24266 ) | ( x38 & n24272 ) | ( n24266 & n24272 ) ;
  assign n24274 = ( n6844 & n24271 ) | ( n6844 & n24273 ) | ( n24271 & n24273 ) ;
  assign n24275 = x38 & ~n24273 ;
  assign n24276 = x38 & ~n24269 ;
  assign n24277 = ( ~n6844 & n24275 ) | ( ~n6844 & n24276 ) | ( n24275 & n24276 ) ;
  assign n24278 = ( n24270 & ~n24274 ) | ( n24270 & n24277 ) | ( ~n24274 & n24277 ) ;
  assign n24282 = ( ~n24261 & n24278 ) | ( ~n24261 & n24281 ) | ( n24278 & n24281 ) ;
  assign n24283 = ( n24261 & ~n24278 ) | ( n24261 & n24282 ) | ( ~n24278 & n24282 ) ;
  assign n24284 = ( ~n24281 & n24282 ) | ( ~n24281 & n24283 ) | ( n24282 & n24283 ) ;
  assign n24285 = n23739 | n23744 ;
  assign n24286 = ( n23739 & n23741 ) | ( n23739 & n24285 ) | ( n23741 & n24285 ) ;
  assign n24287 = n24284 & n24286 ;
  assign n24288 = n24284 & ~n24287 ;
  assign n24289 = x104 & n5554 ;
  assign n24290 = x103 & n5549 ;
  assign n24291 = x102 & ~n5548 ;
  assign n24292 = n5893 & n24291 ;
  assign n24293 = n24290 | n24292 ;
  assign n24294 = n24289 | n24293 ;
  assign n24295 = n5557 | n24289 ;
  assign n24296 = n24293 | n24295 ;
  assign n24297 = ( n7911 & n24294 ) | ( n7911 & n24296 ) | ( n24294 & n24296 ) ;
  assign n24298 = x35 & n24296 ;
  assign n24299 = x35 & n24289 ;
  assign n24300 = ( x35 & n24293 ) | ( x35 & n24299 ) | ( n24293 & n24299 ) ;
  assign n24301 = ( n7911 & n24298 ) | ( n7911 & n24300 ) | ( n24298 & n24300 ) ;
  assign n24302 = x35 & ~n24300 ;
  assign n24303 = x35 & ~n24296 ;
  assign n24304 = ( ~n7911 & n24302 ) | ( ~n7911 & n24303 ) | ( n24302 & n24303 ) ;
  assign n24305 = ( n24297 & ~n24301 ) | ( n24297 & n24304 ) | ( ~n24301 & n24304 ) ;
  assign n24306 = ~n24284 & n24286 ;
  assign n24307 = n24305 & n24306 ;
  assign n24308 = ( n24288 & n24305 ) | ( n24288 & n24307 ) | ( n24305 & n24307 ) ;
  assign n24309 = n24305 | n24306 ;
  assign n24310 = n24288 | n24309 ;
  assign n24311 = ~n24308 & n24310 ;
  assign n24312 = ~n24030 & n24311 ;
  assign n24313 = ( n23765 & n24005 ) | ( n23765 & n24023 ) | ( n24005 & n24023 ) ;
  assign n24314 = n24022 | n24311 ;
  assign n24315 = ( n24311 & n24313 ) | ( n24311 & n24314 ) | ( n24313 & n24314 ) ;
  assign n24316 = n24026 & ~n24315 ;
  assign n24317 = n24312 | n24316 ;
  assign n24318 = n23495 | n23779 ;
  assign n24320 = x109 & n3811 ;
  assign n24321 = x108 & ~n3810 ;
  assign n24322 = n4067 & n24321 ;
  assign n24323 = n24320 | n24322 ;
  assign n24319 = x110 & n3816 ;
  assign n24325 = n3819 | n24319 ;
  assign n24326 = n24323 | n24325 ;
  assign n24324 = n24319 | n24323 ;
  assign n24327 = n24324 & n24326 ;
  assign n24328 = ( n10330 & n24326 ) | ( n10330 & n24327 ) | ( n24326 & n24327 ) ;
  assign n24329 = x29 & n24327 ;
  assign n24330 = x29 & n24326 ;
  assign n24331 = ( n10330 & n24329 ) | ( n10330 & n24330 ) | ( n24329 & n24330 ) ;
  assign n24332 = x29 & ~n24327 ;
  assign n24333 = x29 & ~n24326 ;
  assign n24334 = ( ~n10330 & n24332 ) | ( ~n10330 & n24333 ) | ( n24332 & n24333 ) ;
  assign n24335 = ( n24328 & ~n24331 ) | ( n24328 & n24334 ) | ( ~n24331 & n24334 ) ;
  assign n24336 = n23492 & n24335 ;
  assign n24337 = n23474 & n24336 ;
  assign n24338 = n22984 & n24336 ;
  assign n24339 = ( n22985 & n24337 ) | ( n22985 & n24338 ) | ( n24337 & n24338 ) ;
  assign n24340 = ( n23779 & n24335 ) | ( n23779 & n24339 ) | ( n24335 & n24339 ) ;
  assign n24341 = n24318 & ~n24340 ;
  assign n24342 = n24335 & ~n24336 ;
  assign n24343 = ( ~n23474 & n24335 ) | ( ~n23474 & n24342 ) | ( n24335 & n24342 ) ;
  assign n24344 = ( ~n22984 & n24335 ) | ( ~n22984 & n24342 ) | ( n24335 & n24342 ) ;
  assign n24345 = ( ~n22985 & n24343 ) | ( ~n22985 & n24344 ) | ( n24343 & n24344 ) ;
  assign n24346 = n24317 & n24345 ;
  assign n24347 = ~n23779 & n24346 ;
  assign n24348 = ( n24317 & n24341 ) | ( n24317 & n24347 ) | ( n24341 & n24347 ) ;
  assign n24349 = n24317 | n24345 ;
  assign n24350 = ( ~n23779 & n24317 ) | ( ~n23779 & n24349 ) | ( n24317 & n24349 ) ;
  assign n24351 = n24341 | n24350 ;
  assign n24352 = ~n24348 & n24351 ;
  assign n24353 = n23997 & ~n23999 ;
  assign n24354 = ~n23972 & n23997 ;
  assign n24355 = ( ~n23233 & n24353 ) | ( ~n23233 & n24354 ) | ( n24353 & n24354 ) ;
  assign n24356 = ~n23980 & n24355 ;
  assign n24357 = ~n23782 & n24355 ;
  assign n24358 = ( ~n23974 & n24356 ) | ( ~n23974 & n24357 ) | ( n24356 & n24357 ) ;
  assign n24359 = n24352 & n24358 ;
  assign n24360 = ( n24004 & n24352 ) | ( n24004 & n24359 ) | ( n24352 & n24359 ) ;
  assign n24361 = n24352 | n24358 ;
  assign n24362 = n24004 | n24361 ;
  assign n24363 = ~n24360 & n24362 ;
  assign n24364 = x119 & n1859 ;
  assign n24365 = x118 & n1854 ;
  assign n24366 = x117 & ~n1853 ;
  assign n24367 = n2037 & n24366 ;
  assign n24368 = n24365 | n24367 ;
  assign n24369 = n24364 | n24368 ;
  assign n24370 = n1862 | n24364 ;
  assign n24371 = n24368 | n24370 ;
  assign n24372 = ( n14496 & n24369 ) | ( n14496 & n24371 ) | ( n24369 & n24371 ) ;
  assign n24373 = x20 & n24371 ;
  assign n24374 = x20 & n24364 ;
  assign n24375 = ( x20 & n24368 ) | ( x20 & n24374 ) | ( n24368 & n24374 ) ;
  assign n24376 = ( n14496 & n24373 ) | ( n14496 & n24375 ) | ( n24373 & n24375 ) ;
  assign n24377 = x20 & ~n24375 ;
  assign n24378 = x20 & ~n24371 ;
  assign n24379 = ( ~n14496 & n24377 ) | ( ~n14496 & n24378 ) | ( n24377 & n24378 ) ;
  assign n24380 = ( n24372 & ~n24376 ) | ( n24372 & n24379 ) | ( ~n24376 & n24379 ) ;
  assign n24381 = n23425 | n23790 ;
  assign n24382 = ( n23425 & n23429 ) | ( n23425 & n24381 ) | ( n23429 & n24381 ) ;
  assign n24383 = n24380 | n24382 ;
  assign n24384 = n24380 & n24382 ;
  assign n24385 = n24383 & ~n24384 ;
  assign n24386 = x116 & n2429 ;
  assign n24387 = x115 & n2424 ;
  assign n24388 = x114 & ~n2423 ;
  assign n24389 = n2631 & n24388 ;
  assign n24390 = n24387 | n24389 ;
  assign n24391 = n24386 | n24390 ;
  assign n24392 = n2432 | n24386 ;
  assign n24393 = n24390 | n24392 ;
  assign n24394 = ( ~n13040 & n24391 ) | ( ~n13040 & n24393 ) | ( n24391 & n24393 ) ;
  assign n24395 = n24391 & n24393 ;
  assign n24396 = ( n13022 & n24394 ) | ( n13022 & n24395 ) | ( n24394 & n24395 ) ;
  assign n24397 = x23 & n24396 ;
  assign n24398 = x23 & ~n24396 ;
  assign n24399 = ( n24396 & ~n24397 ) | ( n24396 & n24398 ) | ( ~n24397 & n24398 ) ;
  assign n24400 = n23447 | n23787 ;
  assign n24401 = n23446 | n23787 ;
  assign n24402 = ( n23245 & n24400 ) | ( n23245 & n24401 ) | ( n24400 & n24401 ) ;
  assign n24403 = n24399 & n24402 ;
  assign n24404 = n23448 & n24399 ;
  assign n24405 = ( n23451 & n24403 ) | ( n23451 & n24404 ) | ( n24403 & n24404 ) ;
  assign n24406 = n24399 | n24402 ;
  assign n24407 = n23448 | n24399 ;
  assign n24408 = ( n23451 & n24406 ) | ( n23451 & n24407 ) | ( n24406 & n24407 ) ;
  assign n24409 = ~n24405 & n24408 ;
  assign n24410 = ( n24363 & n24385 ) | ( n24363 & ~n24409 ) | ( n24385 & ~n24409 ) ;
  assign n24411 = ( ~n24385 & n24409 ) | ( ~n24385 & n24410 ) | ( n24409 & n24410 ) ;
  assign n24412 = ( ~n24363 & n24410 ) | ( ~n24363 & n24411 ) | ( n24410 & n24411 ) ;
  assign n24413 = n23961 & ~n23963 ;
  assign n24414 = ~n23404 & n23961 ;
  assign n24415 = ( ~n23302 & n24413 ) | ( ~n23302 & n24414 ) | ( n24413 & n24414 ) ;
  assign n24416 = ~n23799 & n24415 ;
  assign n24417 = ~n23793 & n24415 ;
  assign n24418 = ( ~n23406 & n24416 ) | ( ~n23406 & n24417 ) | ( n24416 & n24417 ) ;
  assign n24419 = n24412 & n24418 ;
  assign n24420 = ( n23968 & n24412 ) | ( n23968 & n24419 ) | ( n24412 & n24419 ) ;
  assign n24421 = n24412 | n24418 ;
  assign n24422 = n23968 | n24421 ;
  assign n24423 = ~n24420 & n24422 ;
  assign n24424 = n23937 & n24423 ;
  assign n24425 = ~n23939 & n24424 ;
  assign n24426 = ( n23941 & n24423 ) | ( n23941 & n24425 ) | ( n24423 & n24425 ) ;
  assign n24427 = n23937 | n24423 ;
  assign n24428 = ( ~n23939 & n24423 ) | ( ~n23939 & n24427 ) | ( n24423 & n24427 ) ;
  assign n24429 = n23941 | n24428 ;
  assign n24430 = ~n24426 & n24429 ;
  assign n24431 = n23908 | n24430 ;
  assign n24432 = ( ~n23918 & n24430 ) | ( ~n23918 & n24431 ) | ( n24430 & n24431 ) ;
  assign n24433 = n23920 | n24432 ;
  assign n24434 = n23908 & n24430 ;
  assign n24435 = ~n23918 & n24434 ;
  assign n24436 = ( n23920 & n24430 ) | ( n23920 & n24435 ) | ( n24430 & n24435 ) ;
  assign n24437 = n24433 & ~n24436 ;
  assign n24438 = n22843 & n23382 ;
  assign n24439 = n22825 & n24438 ;
  assign n24440 = n22672 & n24438 ;
  assign n24441 = ( n22678 & n24439 ) | ( n22678 & n24440 ) | ( n24439 & n24440 ) ;
  assign n24442 = ( n23346 & n23382 ) | ( n23346 & n24441 ) | ( n23382 & n24441 ) ;
  assign n24443 = ( n23333 & n23382 ) | ( n23333 & n24441 ) | ( n23382 & n24441 ) ;
  assign n24444 = ( n22847 & n24442 ) | ( n22847 & n24443 ) | ( n24442 & n24443 ) ;
  assign n24445 = n23866 & ~n24444 ;
  assign n24446 = n23382 & ~n24438 ;
  assign n24447 = ( ~n22825 & n23382 ) | ( ~n22825 & n24446 ) | ( n23382 & n24446 ) ;
  assign n24448 = ( ~n22672 & n23382 ) | ( ~n22672 & n24446 ) | ( n23382 & n24446 ) ;
  assign n24449 = ( ~n22678 & n24447 ) | ( ~n22678 & n24448 ) | ( n24447 & n24448 ) ;
  assign n24450 = ~n23346 & n24449 ;
  assign n24451 = ~n23333 & n24449 ;
  assign n24452 = ( ~n22847 & n24450 ) | ( ~n22847 & n24451 ) | ( n24450 & n24451 ) ;
  assign n24453 = n23863 & ~n24452 ;
  assign n24454 = ~n24445 & n24453 ;
  assign n24455 = ( n23863 & n24444 ) | ( n23863 & ~n24454 ) | ( n24444 & ~n24454 ) ;
  assign n24456 = n24437 & ~n24455 ;
  assign n24457 = n24437 & n24455 ;
  assign n24458 = n24455 & ~n24457 ;
  assign n24459 = n24456 | n24458 ;
  assign n24460 = n23871 | n23886 ;
  assign n24461 = n23875 | n24460 ;
  assign n24462 = n24459 & n24461 ;
  assign n24463 = n23871 & n24459 ;
  assign n24464 = ( n23883 & n24462 ) | ( n23883 & n24463 ) | ( n24462 & n24463 ) ;
  assign n24465 = ( n23891 & n24459 ) | ( n23891 & n24463 ) | ( n24459 & n24463 ) ;
  assign n24466 = ( n23879 & n24462 ) | ( n23879 & n24465 ) | ( n24462 & n24465 ) ;
  assign n24467 = n24462 & n24465 ;
  assign n24468 = ( n22783 & n24466 ) | ( n22783 & n24467 ) | ( n24466 & n24467 ) ;
  assign n24469 = ( n22796 & n24464 ) | ( n22796 & n24468 ) | ( n24464 & n24468 ) ;
  assign n24470 = n23871 | n23891 ;
  assign n24471 = ( n23880 & n24461 ) | ( n23880 & n24470 ) | ( n24461 & n24470 ) ;
  assign n24472 = ( n23871 & n23883 ) | ( n23871 & n24461 ) | ( n23883 & n24461 ) ;
  assign n24473 = ( n22796 & n24471 ) | ( n22796 & n24472 ) | ( n24471 & n24472 ) ;
  assign n24474 = ( ~n24437 & n24455 ) | ( ~n24437 & n24473 ) | ( n24455 & n24473 ) ;
  assign n24475 = ( n24456 & ~n24469 ) | ( n24456 & n24474 ) | ( ~n24469 & n24474 ) ;
  assign n24476 = x127 & ~n630 ;
  assign n24477 = n764 & n24476 ;
  assign n24478 = n639 & n19877 ;
  assign n24479 = n24477 | n24478 ;
  assign n24480 = n639 & n19880 ;
  assign n24481 = n24477 | n24480 ;
  assign n24482 = ( n18202 & n24479 ) | ( n18202 & n24481 ) | ( n24479 & n24481 ) ;
  assign n24483 = n24479 & n24481 ;
  assign n24484 = ( n18212 & n24482 ) | ( n18212 & n24483 ) | ( n24482 & n24483 ) ;
  assign n24485 = ( n18214 & n24482 ) | ( n18214 & n24483 ) | ( n24482 & n24483 ) ;
  assign n24486 = ( n14002 & n24484 ) | ( n14002 & n24485 ) | ( n24484 & n24485 ) ;
  assign n24487 = x11 & n24484 ;
  assign n24488 = x11 & n24485 ;
  assign n24489 = ( n14002 & n24487 ) | ( n14002 & n24488 ) | ( n24487 & n24488 ) ;
  assign n24490 = x11 & ~n24488 ;
  assign n24491 = x11 & ~n24487 ;
  assign n24492 = ( ~n14002 & n24490 ) | ( ~n14002 & n24491 ) | ( n24490 & n24491 ) ;
  assign n24493 = ( n24486 & ~n24489 ) | ( n24486 & n24492 ) | ( ~n24489 & n24492 ) ;
  assign n24911 = x125 & n957 ;
  assign n24912 = x124 & ~n956 ;
  assign n24913 = n1105 & n24912 ;
  assign n24914 = n24911 | n24913 ;
  assign n24910 = x126 & n962 ;
  assign n24916 = n965 | n24910 ;
  assign n24917 = n24914 | n24916 ;
  assign n24915 = n24910 | n24914 ;
  assign n24918 = n24915 & n24917 ;
  assign n24919 = ( n18220 & n24917 ) | ( n18220 & n24918 ) | ( n24917 & n24918 ) ;
  assign n24920 = x14 & n24918 ;
  assign n24921 = x14 & n24917 ;
  assign n24922 = ( n18220 & n24920 ) | ( n18220 & n24921 ) | ( n24920 & n24921 ) ;
  assign n24923 = x14 & ~n24918 ;
  assign n24924 = x14 & ~n24917 ;
  assign n24925 = ( ~n18220 & n24923 ) | ( ~n18220 & n24924 ) | ( n24923 & n24924 ) ;
  assign n24926 = ( n24919 & ~n24922 ) | ( n24919 & n24925 ) | ( ~n24922 & n24925 ) ;
  assign n24927 = n23961 & n24926 ;
  assign n24928 = n23962 & n24926 ;
  assign n24929 = n23963 & n24926 ;
  assign n24930 = ( n23302 & n24928 ) | ( n23302 & n24929 ) | ( n24928 & n24929 ) ;
  assign n24931 = ( n23799 & n24927 ) | ( n23799 & n24930 ) | ( n24927 & n24930 ) ;
  assign n24932 = ( n23793 & n24927 ) | ( n23793 & n24930 ) | ( n24927 & n24930 ) ;
  assign n24933 = ( n23406 & n24931 ) | ( n23406 & n24932 ) | ( n24931 & n24932 ) ;
  assign n24934 = ( n24420 & n24926 ) | ( n24420 & n24933 ) | ( n24926 & n24933 ) ;
  assign n24935 = n23961 | n24926 ;
  assign n24936 = n23962 | n24926 ;
  assign n24937 = n23963 | n24926 ;
  assign n24938 = ( n23302 & n24936 ) | ( n23302 & n24937 ) | ( n24936 & n24937 ) ;
  assign n24939 = ( n23799 & n24935 ) | ( n23799 & n24938 ) | ( n24935 & n24938 ) ;
  assign n24940 = ( n23793 & n24935 ) | ( n23793 & n24938 ) | ( n24935 & n24938 ) ;
  assign n24941 = ( n23406 & n24939 ) | ( n23406 & n24940 ) | ( n24939 & n24940 ) ;
  assign n24942 = n24420 | n24941 ;
  assign n24943 = ~n24934 & n24942 ;
  assign n24944 = x123 & n1383 ;
  assign n24945 = x122 & n1378 ;
  assign n24946 = x121 & ~n1377 ;
  assign n24947 = n1542 & n24946 ;
  assign n24948 = n24945 | n24947 ;
  assign n24949 = n24944 | n24948 ;
  assign n24950 = n1386 | n24944 ;
  assign n24951 = n24948 | n24950 ;
  assign n24952 = ( n16086 & n24949 ) | ( n16086 & n24951 ) | ( n24949 & n24951 ) ;
  assign n24953 = x17 & n24951 ;
  assign n24954 = x17 & n24944 ;
  assign n24955 = ( x17 & n24948 ) | ( x17 & n24954 ) | ( n24948 & n24954 ) ;
  assign n24956 = ( n16086 & n24953 ) | ( n16086 & n24955 ) | ( n24953 & n24955 ) ;
  assign n24957 = x17 & ~n24955 ;
  assign n24958 = x17 & ~n24951 ;
  assign n24959 = ( ~n16086 & n24957 ) | ( ~n16086 & n24958 ) | ( n24957 & n24958 ) ;
  assign n24960 = ( n24952 & ~n24956 ) | ( n24952 & n24959 ) | ( ~n24956 & n24959 ) ;
  assign n24961 = n24363 & n24409 ;
  assign n24962 = n24363 | n24409 ;
  assign n24963 = ~n24961 & n24962 ;
  assign n24964 = n24380 | n24963 ;
  assign n24965 = ( n24382 & n24963 ) | ( n24382 & n24964 ) | ( n24963 & n24964 ) ;
  assign n24966 = n24960 | n24965 ;
  assign n24967 = n24384 | n24960 ;
  assign n24968 = ( n24385 & n24966 ) | ( n24385 & n24967 ) | ( n24966 & n24967 ) ;
  assign n24969 = n24960 & n24965 ;
  assign n24970 = n24384 & n24960 ;
  assign n24971 = ( n24385 & n24969 ) | ( n24385 & n24970 ) | ( n24969 & n24970 ) ;
  assign n24972 = n24968 & ~n24971 ;
  assign n24511 = n24363 | n24405 ;
  assign n24512 = ( n24405 & n24409 ) | ( n24405 & n24511 ) | ( n24409 & n24511 ) ;
  assign n24494 = x120 & n1859 ;
  assign n24495 = x119 & n1854 ;
  assign n24496 = x118 & ~n1853 ;
  assign n24497 = n2037 & n24496 ;
  assign n24498 = n24495 | n24497 ;
  assign n24499 = n24494 | n24498 ;
  assign n24500 = n1862 | n24494 ;
  assign n24501 = n24498 | n24500 ;
  assign n24502 = ( n14991 & n24499 ) | ( n14991 & n24501 ) | ( n24499 & n24501 ) ;
  assign n24503 = x20 & n24501 ;
  assign n24504 = x20 & n24494 ;
  assign n24505 = ( x20 & n24498 ) | ( x20 & n24504 ) | ( n24498 & n24504 ) ;
  assign n24506 = ( n14991 & n24503 ) | ( n14991 & n24505 ) | ( n24503 & n24505 ) ;
  assign n24507 = x20 & ~n24505 ;
  assign n24508 = x20 & ~n24501 ;
  assign n24509 = ( ~n14991 & n24507 ) | ( ~n14991 & n24508 ) | ( n24507 & n24508 ) ;
  assign n24510 = ( n24502 & ~n24506 ) | ( n24502 & n24509 ) | ( ~n24506 & n24509 ) ;
  assign n24513 = n24510 & n24512 ;
  assign n24514 = n24512 & ~n24513 ;
  assign n24515 = n24003 | n24360 ;
  assign n24517 = x116 & n2424 ;
  assign n24518 = x115 & ~n2423 ;
  assign n24519 = n2631 & n24518 ;
  assign n24520 = n24517 | n24519 ;
  assign n24516 = x117 & n2429 ;
  assign n24522 = n2432 | n24516 ;
  assign n24523 = n24520 | n24522 ;
  assign n24521 = n24516 | n24520 ;
  assign n24524 = n24521 & n24523 ;
  assign n24525 = ( ~n13522 & n24523 ) | ( ~n13522 & n24524 ) | ( n24523 & n24524 ) ;
  assign n24526 = n24523 & n24524 ;
  assign n24527 = ( n13503 & n24525 ) | ( n13503 & n24526 ) | ( n24525 & n24526 ) ;
  assign n24528 = x23 & n24527 ;
  assign n24529 = x23 & ~n24527 ;
  assign n24530 = ( n24527 & ~n24528 ) | ( n24527 & n24529 ) | ( ~n24528 & n24529 ) ;
  assign n24531 = n23997 & n24530 ;
  assign n24532 = n23998 & n24530 ;
  assign n24533 = n23999 & n24530 ;
  assign n24534 = ( n23233 & n24532 ) | ( n23233 & n24533 ) | ( n24532 & n24533 ) ;
  assign n24535 = ( n23980 & n24531 ) | ( n23980 & n24534 ) | ( n24531 & n24534 ) ;
  assign n24536 = ( n23782 & n24531 ) | ( n23782 & n24534 ) | ( n24531 & n24534 ) ;
  assign n24537 = ( n23974 & n24535 ) | ( n23974 & n24536 ) | ( n24535 & n24536 ) ;
  assign n24538 = ( n24360 & n24530 ) | ( n24360 & n24537 ) | ( n24530 & n24537 ) ;
  assign n24539 = n24515 & ~n24538 ;
  assign n24541 = x107 & n4626 ;
  assign n24542 = x106 & ~n4625 ;
  assign n24543 = n4943 & n24542 ;
  assign n24544 = n24541 | n24543 ;
  assign n24540 = x108 & n4631 ;
  assign n24546 = n4634 | n24540 ;
  assign n24547 = n24544 | n24546 ;
  assign n24545 = n24540 | n24544 ;
  assign n24548 = n24545 & n24547 ;
  assign n24549 = ( n9479 & n24547 ) | ( n9479 & n24548 ) | ( n24547 & n24548 ) ;
  assign n24550 = x32 & n24548 ;
  assign n24551 = x32 & n24547 ;
  assign n24552 = ( n9479 & n24550 ) | ( n9479 & n24551 ) | ( n24550 & n24551 ) ;
  assign n24553 = x32 & ~n24548 ;
  assign n24554 = x32 & ~n24547 ;
  assign n24555 = ( ~n9479 & n24553 ) | ( ~n9479 & n24554 ) | ( n24553 & n24554 ) ;
  assign n24556 = ( n24549 & ~n24552 ) | ( n24549 & n24555 ) | ( ~n24552 & n24555 ) ;
  assign n24557 = n24287 & n24556 ;
  assign n24558 = ( n24308 & n24556 ) | ( n24308 & n24557 ) | ( n24556 & n24557 ) ;
  assign n24559 = n24287 | n24556 ;
  assign n24560 = n24308 | n24559 ;
  assign n24561 = ~n24558 & n24560 ;
  assign n24562 = x75 & n18290 ;
  assign n24563 = x63 & x74 ;
  assign n24564 = ~n18290 & n24563 ;
  assign n24565 = n24562 | n24564 ;
  assign n24566 = ~n24058 & n24565 ;
  assign n24567 = n24058 | n24566 ;
  assign n24568 = n24565 & ~n24566 ;
  assign n24569 = n24567 & ~n24568 ;
  assign n24570 = n24059 & ~n24569 ;
  assign n24571 = n24569 | n24570 ;
  assign n24572 = n24062 & ~n24571 ;
  assign n24573 = ( n24053 & n24571 ) | ( n24053 & ~n24572 ) | ( n24571 & ~n24572 ) ;
  assign n24574 = ~n24059 & n24061 ;
  assign n24575 = ~n24060 & n24574 ;
  assign n24576 = n24569 & ~n24575 ;
  assign n24577 = n24059 & n24569 ;
  assign n24578 = ( n24053 & n24576 ) | ( n24053 & n24577 ) | ( n24576 & n24577 ) ;
  assign n24579 = n24573 & ~n24578 ;
  assign n24580 = x78 & n17146 ;
  assign n24581 = x77 & n17141 ;
  assign n24582 = x76 & ~n17140 ;
  assign n24583 = n17724 & n24582 ;
  assign n24584 = n24581 | n24583 ;
  assign n24585 = n24580 | n24584 ;
  assign n24586 = n17149 | n24580 ;
  assign n24587 = n24584 | n24586 ;
  assign n24588 = ( n1192 & n24585 ) | ( n1192 & n24587 ) | ( n24585 & n24587 ) ;
  assign n24589 = x62 & n24587 ;
  assign n24590 = x62 & n24580 ;
  assign n24591 = ( x62 & n24584 ) | ( x62 & n24590 ) | ( n24584 & n24590 ) ;
  assign n24592 = ( n1192 & n24589 ) | ( n1192 & n24591 ) | ( n24589 & n24591 ) ;
  assign n24593 = x62 & ~n24591 ;
  assign n24594 = x62 & ~n24587 ;
  assign n24595 = ( ~n1192 & n24593 ) | ( ~n1192 & n24594 ) | ( n24593 & n24594 ) ;
  assign n24596 = ( n24588 & ~n24592 ) | ( n24588 & n24595 ) | ( ~n24592 & n24595 ) ;
  assign n24597 = ~n24579 & n24596 ;
  assign n24598 = n24579 & ~n24596 ;
  assign n24599 = n24597 | n24598 ;
  assign n24600 = x81 & n15552 ;
  assign n24601 = x80 & n15547 ;
  assign n24602 = x79 & ~n15546 ;
  assign n24603 = n16123 & n24602 ;
  assign n24604 = n24601 | n24603 ;
  assign n24605 = n24600 | n24604 ;
  assign n24606 = n15555 | n24600 ;
  assign n24607 = n24604 | n24606 ;
  assign n24608 = ( n1651 & n24605 ) | ( n1651 & n24607 ) | ( n24605 & n24607 ) ;
  assign n24609 = x59 & n24607 ;
  assign n24610 = x59 & n24600 ;
  assign n24611 = ( x59 & n24604 ) | ( x59 & n24610 ) | ( n24604 & n24610 ) ;
  assign n24612 = ( n1651 & n24609 ) | ( n1651 & n24611 ) | ( n24609 & n24611 ) ;
  assign n24613 = x59 & ~n24611 ;
  assign n24614 = x59 & ~n24607 ;
  assign n24615 = ( ~n1651 & n24613 ) | ( ~n1651 & n24614 ) | ( n24613 & n24614 ) ;
  assign n24616 = ( n24608 & ~n24612 ) | ( n24608 & n24615 ) | ( ~n24612 & n24615 ) ;
  assign n24617 = ~n24599 & n24616 ;
  assign n24618 = n24599 | n24617 ;
  assign n24620 = ~n24068 & n24087 ;
  assign n24621 = n24065 & n24620 ;
  assign n24622 = n24069 & ~n24621 ;
  assign n24623 = n24069 & ~n24087 ;
  assign n24624 = ( ~n24070 & n24622 ) | ( ~n24070 & n24623 ) | ( n24622 & n24623 ) ;
  assign n24619 = n24599 & n24616 ;
  assign n24625 = n24619 & ~n24624 ;
  assign n24626 = ( n24618 & n24624 ) | ( n24618 & ~n24625 ) | ( n24624 & ~n24625 ) ;
  assign n24627 = ~n24619 & n24624 ;
  assign n24628 = n24618 & n24627 ;
  assign n24629 = n24626 & ~n24628 ;
  assign n24630 = x84 & n14045 ;
  assign n24631 = x83 & n14040 ;
  assign n24632 = x82 & ~n14039 ;
  assign n24633 = n14552 & n24632 ;
  assign n24634 = n24631 | n24633 ;
  assign n24635 = n24630 | n24634 ;
  assign n24636 = n14048 | n24630 ;
  assign n24637 = n24634 | n24636 ;
  assign n24638 = ( n2194 & n24635 ) | ( n2194 & n24637 ) | ( n24635 & n24637 ) ;
  assign n24639 = x56 & n24637 ;
  assign n24640 = x56 & n24630 ;
  assign n24641 = ( x56 & n24634 ) | ( x56 & n24640 ) | ( n24634 & n24640 ) ;
  assign n24642 = ( n2194 & n24639 ) | ( n2194 & n24641 ) | ( n24639 & n24641 ) ;
  assign n24643 = x56 & ~n24641 ;
  assign n24644 = x56 & ~n24637 ;
  assign n24645 = ( ~n2194 & n24643 ) | ( ~n2194 & n24644 ) | ( n24643 & n24644 ) ;
  assign n24646 = ( n24638 & ~n24642 ) | ( n24638 & n24645 ) | ( ~n24642 & n24645 ) ;
  assign n24647 = n24629 | n24646 ;
  assign n24648 = n24629 & n24646 ;
  assign n24649 = n24647 & ~n24648 ;
  assign n24650 = n24098 & n24117 ;
  assign n24651 = ( n24035 & n24117 ) | ( n24035 & n24650 ) | ( n24117 & n24650 ) ;
  assign n24652 = ~n24097 & n24651 ;
  assign n24653 = n24097 | n24652 ;
  assign n24654 = ~n24649 & n24653 ;
  assign n24655 = n24649 & n24653 ;
  assign n24656 = x87 & n12574 ;
  assign n24657 = x86 & n12569 ;
  assign n24658 = x85 & ~n12568 ;
  assign n24659 = n13076 & n24658 ;
  assign n24660 = n24657 | n24659 ;
  assign n24661 = n24656 | n24660 ;
  assign n24662 = n12577 | n24656 ;
  assign n24663 = n24660 | n24662 ;
  assign n24664 = ( n2816 & n24661 ) | ( n2816 & n24663 ) | ( n24661 & n24663 ) ;
  assign n24665 = x53 & n24663 ;
  assign n24666 = x53 & n24656 ;
  assign n24667 = ( x53 & n24660 ) | ( x53 & n24666 ) | ( n24660 & n24666 ) ;
  assign n24668 = ( n2816 & n24665 ) | ( n2816 & n24667 ) | ( n24665 & n24667 ) ;
  assign n24669 = x53 & ~n24667 ;
  assign n24670 = x53 & ~n24663 ;
  assign n24671 = ( ~n2816 & n24669 ) | ( ~n2816 & n24670 ) | ( n24669 & n24670 ) ;
  assign n24672 = ( n24664 & ~n24668 ) | ( n24664 & n24671 ) | ( ~n24668 & n24671 ) ;
  assign n24673 = n24649 | n24672 ;
  assign n24674 = ( ~n24655 & n24672 ) | ( ~n24655 & n24673 ) | ( n24672 & n24673 ) ;
  assign n24675 = n24654 | n24674 ;
  assign n24676 = n24649 & ~n24655 ;
  assign n24677 = n24654 & n24672 ;
  assign n24678 = ( n24672 & n24676 ) | ( n24672 & n24677 ) | ( n24676 & n24677 ) ;
  assign n24679 = n24675 & ~n24678 ;
  assign n24680 = ( n24124 & n24125 ) | ( n24124 & n24146 ) | ( n24125 & n24146 ) ;
  assign n24681 = n24679 & n24680 ;
  assign n24682 = n24679 | n24680 ;
  assign n24683 = ~n24681 & n24682 ;
  assign n24684 = x90 & n11205 ;
  assign n24685 = x89 & n11200 ;
  assign n24686 = x88 & ~n11199 ;
  assign n24687 = n11679 & n24686 ;
  assign n24688 = n24685 | n24687 ;
  assign n24689 = n24684 | n24688 ;
  assign n24690 = n11208 | n24684 ;
  assign n24691 = n24688 | n24690 ;
  assign n24692 = ( n3519 & n24689 ) | ( n3519 & n24691 ) | ( n24689 & n24691 ) ;
  assign n24693 = x50 & n24691 ;
  assign n24694 = x50 & n24684 ;
  assign n24695 = ( x50 & n24688 ) | ( x50 & n24694 ) | ( n24688 & n24694 ) ;
  assign n24696 = ( n3519 & n24693 ) | ( n3519 & n24695 ) | ( n24693 & n24695 ) ;
  assign n24697 = x50 & ~n24695 ;
  assign n24698 = x50 & ~n24691 ;
  assign n24699 = ( ~n3519 & n24697 ) | ( ~n3519 & n24698 ) | ( n24697 & n24698 ) ;
  assign n24700 = ( n24692 & ~n24696 ) | ( n24692 & n24699 ) | ( ~n24696 & n24699 ) ;
  assign n24701 = n24683 & n24700 ;
  assign n24702 = n24683 | n24700 ;
  assign n24703 = ~n24701 & n24702 ;
  assign n24704 = n24150 & n24168 ;
  assign n24705 = ~n24148 & n24704 ;
  assign n24706 = n24148 | n24705 ;
  assign n24707 = n24703 & n24706 ;
  assign n24708 = n24703 | n24706 ;
  assign n24709 = ~n24707 & n24708 ;
  assign n24710 = x93 & n9933 ;
  assign n24711 = x92 & n9928 ;
  assign n24712 = x91 & ~n9927 ;
  assign n24713 = n10379 & n24712 ;
  assign n24714 = n24711 | n24713 ;
  assign n24715 = n24710 | n24714 ;
  assign n24716 = n9936 | n24710 ;
  assign n24717 = n24714 | n24716 ;
  assign n24718 = ( n4305 & n24715 ) | ( n4305 & n24717 ) | ( n24715 & n24717 ) ;
  assign n24719 = x47 & n24717 ;
  assign n24720 = x47 & n24710 ;
  assign n24721 = ( x47 & n24714 ) | ( x47 & n24720 ) | ( n24714 & n24720 ) ;
  assign n24722 = ( n4305 & n24719 ) | ( n4305 & n24721 ) | ( n24719 & n24721 ) ;
  assign n24723 = x47 & ~n24721 ;
  assign n24724 = x47 & ~n24717 ;
  assign n24725 = ( ~n4305 & n24723 ) | ( ~n4305 & n24724 ) | ( n24723 & n24724 ) ;
  assign n24726 = ( n24718 & ~n24722 ) | ( n24718 & n24725 ) | ( ~n24722 & n24725 ) ;
  assign n24727 = n24709 & ~n24726 ;
  assign n24728 = n24709 | n24726 ;
  assign n24729 = ( ~n24709 & n24727 ) | ( ~n24709 & n24728 ) | ( n24727 & n24728 ) ;
  assign n24730 = n24175 | n24195 ;
  assign n24731 = ( n24172 & n24195 ) | ( n24172 & n24730 ) | ( n24195 & n24730 ) ;
  assign n24732 = ( n24177 & n24178 ) | ( n24177 & n24731 ) | ( n24178 & n24731 ) ;
  assign n24733 = n24729 | n24732 ;
  assign n24734 = n24729 & n24732 ;
  assign n24735 = n24733 & ~n24734 ;
  assign n24736 = x96 & n8724 ;
  assign n24737 = x95 & n8719 ;
  assign n24738 = x94 & ~n8718 ;
  assign n24739 = n9149 & n24738 ;
  assign n24740 = n24737 | n24739 ;
  assign n24741 = n24736 | n24740 ;
  assign n24742 = n8727 | n24736 ;
  assign n24743 = n24740 | n24742 ;
  assign n24744 = ( n5202 & n24741 ) | ( n5202 & n24743 ) | ( n24741 & n24743 ) ;
  assign n24745 = x44 & n24743 ;
  assign n24746 = x44 & n24736 ;
  assign n24747 = ( x44 & n24740 ) | ( x44 & n24746 ) | ( n24740 & n24746 ) ;
  assign n24748 = ( n5202 & n24745 ) | ( n5202 & n24747 ) | ( n24745 & n24747 ) ;
  assign n24749 = x44 & ~n24747 ;
  assign n24750 = x44 & ~n24743 ;
  assign n24751 = ( ~n5202 & n24749 ) | ( ~n5202 & n24750 ) | ( n24749 & n24750 ) ;
  assign n24752 = ( n24744 & ~n24748 ) | ( n24744 & n24751 ) | ( ~n24748 & n24751 ) ;
  assign n24753 = n24735 | n24752 ;
  assign n24754 = n24735 & n24752 ;
  assign n24755 = n24753 & ~n24754 ;
  assign n24756 = n24207 | n24225 ;
  assign n24757 = ( n24207 & n24208 ) | ( n24207 & n24756 ) | ( n24208 & n24756 ) ;
  assign n24758 = n24755 & n24757 ;
  assign n24759 = n24755 | n24757 ;
  assign n24760 = ~n24758 & n24759 ;
  assign n24761 = x99 & n7566 ;
  assign n24762 = x98 & n7561 ;
  assign n24763 = x97 & ~n7560 ;
  assign n24764 = n7953 & n24763 ;
  assign n24765 = n24762 | n24764 ;
  assign n24766 = n24761 | n24765 ;
  assign n24767 = n7569 | n24761 ;
  assign n24768 = n24765 | n24767 ;
  assign n24769 = ( n6164 & n24766 ) | ( n6164 & n24768 ) | ( n24766 & n24768 ) ;
  assign n24770 = x41 & n24768 ;
  assign n24771 = x41 & n24761 ;
  assign n24772 = ( x41 & n24765 ) | ( x41 & n24771 ) | ( n24765 & n24771 ) ;
  assign n24773 = ( n6164 & n24770 ) | ( n6164 & n24772 ) | ( n24770 & n24772 ) ;
  assign n24774 = x41 & ~n24772 ;
  assign n24775 = x41 & ~n24768 ;
  assign n24776 = ( ~n6164 & n24774 ) | ( ~n6164 & n24775 ) | ( n24774 & n24775 ) ;
  assign n24777 = ( n24769 & ~n24773 ) | ( n24769 & n24776 ) | ( ~n24773 & n24776 ) ;
  assign n24778 = n24760 & ~n24777 ;
  assign n24779 = n24760 | n24777 ;
  assign n24780 = ( ~n24760 & n24778 ) | ( ~n24760 & n24779 ) | ( n24778 & n24779 ) ;
  assign n24781 = n24232 | n24258 ;
  assign n24782 = ( n24228 & n24258 ) | ( n24228 & n24781 ) | ( n24258 & n24781 ) ;
  assign n24783 = ( n24233 & n24235 ) | ( n24233 & n24782 ) | ( n24235 & n24782 ) ;
  assign n24784 = n24780 | n24783 ;
  assign n24785 = n24780 & n24783 ;
  assign n24786 = n24784 & ~n24785 ;
  assign n24787 = x102 & n6536 ;
  assign n24788 = x101 & n6531 ;
  assign n24789 = x100 & ~n6530 ;
  assign n24790 = n6871 & n24789 ;
  assign n24791 = n24788 | n24790 ;
  assign n24792 = n24787 | n24791 ;
  assign n24793 = n6539 | n24787 ;
  assign n24794 = n24791 | n24793 ;
  assign n24795 = ( n7178 & n24792 ) | ( n7178 & n24794 ) | ( n24792 & n24794 ) ;
  assign n24796 = x38 & n24794 ;
  assign n24797 = x38 & n24787 ;
  assign n24798 = ( x38 & n24791 ) | ( x38 & n24797 ) | ( n24791 & n24797 ) ;
  assign n24799 = ( n7178 & n24796 ) | ( n7178 & n24798 ) | ( n24796 & n24798 ) ;
  assign n24800 = x38 & ~n24798 ;
  assign n24801 = x38 & ~n24794 ;
  assign n24802 = ( ~n7178 & n24800 ) | ( ~n7178 & n24801 ) | ( n24800 & n24801 ) ;
  assign n24803 = ( n24795 & ~n24799 ) | ( n24795 & n24802 ) | ( ~n24799 & n24802 ) ;
  assign n24804 = n24786 | n24803 ;
  assign n24805 = n24786 & n24803 ;
  assign n24806 = n24804 & ~n24805 ;
  assign n24807 = n24261 & n24281 ;
  assign n24808 = n24261 & ~n24807 ;
  assign n24809 = n24278 & n24281 ;
  assign n24810 = ~n24261 & n24809 ;
  assign n24811 = n24807 | n24810 ;
  assign n24812 = n24278 | n24807 ;
  assign n24813 = ( n24808 & n24811 ) | ( n24808 & n24812 ) | ( n24811 & n24812 ) ;
  assign n24814 = n24806 & n24813 ;
  assign n24815 = n24806 | n24813 ;
  assign n24816 = ~n24814 & n24815 ;
  assign n24817 = x105 & n5554 ;
  assign n24818 = x104 & n5549 ;
  assign n24819 = x103 & ~n5548 ;
  assign n24820 = n5893 & n24819 ;
  assign n24821 = n24818 | n24820 ;
  assign n24822 = n24817 | n24821 ;
  assign n24823 = n5557 | n24817 ;
  assign n24824 = n24821 | n24823 ;
  assign n24825 = ( n8273 & n24822 ) | ( n8273 & n24824 ) | ( n24822 & n24824 ) ;
  assign n24826 = x35 & n24824 ;
  assign n24827 = x35 & n24817 ;
  assign n24828 = ( x35 & n24821 ) | ( x35 & n24827 ) | ( n24821 & n24827 ) ;
  assign n24829 = ( n8273 & n24826 ) | ( n8273 & n24828 ) | ( n24826 & n24828 ) ;
  assign n24830 = x35 & ~n24828 ;
  assign n24831 = x35 & ~n24824 ;
  assign n24832 = ( ~n8273 & n24830 ) | ( ~n8273 & n24831 ) | ( n24830 & n24831 ) ;
  assign n24833 = ( n24825 & ~n24829 ) | ( n24825 & n24832 ) | ( ~n24829 & n24832 ) ;
  assign n24834 = n24816 & ~n24833 ;
  assign n24835 = n24816 | n24833 ;
  assign n24836 = ( ~n24816 & n24834 ) | ( ~n24816 & n24835 ) | ( n24834 & n24835 ) ;
  assign n24837 = n24561 & ~n24836 ;
  assign n24838 = n24836 | n24837 ;
  assign n24839 = ( ~n24561 & n24837 ) | ( ~n24561 & n24838 ) | ( n24837 & n24838 ) ;
  assign n24841 = x113 & n3080 ;
  assign n24842 = x112 & ~n3079 ;
  assign n24843 = n3309 & n24842 ;
  assign n24844 = n24841 | n24843 ;
  assign n24840 = x114 & n3085 ;
  assign n24846 = n3088 | n24840 ;
  assign n24847 = n24844 | n24846 ;
  assign n24845 = n24840 | n24844 ;
  assign n24848 = n24845 & n24847 ;
  assign n24849 = ( ~n12095 & n24847 ) | ( ~n12095 & n24848 ) | ( n24847 & n24848 ) ;
  assign n24850 = n24847 & n24848 ;
  assign n24851 = ( n12079 & n24849 ) | ( n12079 & n24850 ) | ( n24849 & n24850 ) ;
  assign n24852 = x26 & n24851 ;
  assign n24853 = x26 & ~n24851 ;
  assign n24854 = ( n24851 & ~n24852 ) | ( n24851 & n24853 ) | ( ~n24852 & n24853 ) ;
  assign n24855 = n24339 & n24854 ;
  assign n24856 = n24335 & n24854 ;
  assign n24857 = ( n23779 & n24855 ) | ( n23779 & n24856 ) | ( n24855 & n24856 ) ;
  assign n24858 = ( n24347 & n24854 ) | ( n24347 & n24857 ) | ( n24854 & n24857 ) ;
  assign n24859 = ( n24317 & n24854 ) | ( n24317 & n24857 ) | ( n24854 & n24857 ) ;
  assign n24860 = ( n24341 & n24858 ) | ( n24341 & n24859 ) | ( n24858 & n24859 ) ;
  assign n24861 = n24339 | n24854 ;
  assign n24862 = n24335 | n24854 ;
  assign n24863 = ( n23779 & n24861 ) | ( n23779 & n24862 ) | ( n24861 & n24862 ) ;
  assign n24864 = n24347 | n24863 ;
  assign n24865 = n24317 | n24863 ;
  assign n24866 = ( n24341 & n24864 ) | ( n24341 & n24865 ) | ( n24864 & n24865 ) ;
  assign n24867 = ~n24860 & n24866 ;
  assign n24868 = x111 & n3816 ;
  assign n24869 = x110 & n3811 ;
  assign n24870 = x109 & ~n3810 ;
  assign n24871 = n4067 & n24870 ;
  assign n24872 = n24869 | n24871 ;
  assign n24873 = n24868 | n24872 ;
  assign n24874 = n3819 | n24868 ;
  assign n24875 = n24872 | n24874 ;
  assign n24876 = ( n10749 & n24873 ) | ( n10749 & n24875 ) | ( n24873 & n24875 ) ;
  assign n24877 = x29 & n24875 ;
  assign n24878 = x29 & n24868 ;
  assign n24879 = ( x29 & n24872 ) | ( x29 & n24878 ) | ( n24872 & n24878 ) ;
  assign n24880 = ( n10749 & n24877 ) | ( n10749 & n24879 ) | ( n24877 & n24879 ) ;
  assign n24881 = x29 & ~n24879 ;
  assign n24882 = x29 & ~n24875 ;
  assign n24883 = ( ~n10749 & n24881 ) | ( ~n10749 & n24882 ) | ( n24881 & n24882 ) ;
  assign n24884 = ( n24876 & ~n24880 ) | ( n24876 & n24883 ) | ( ~n24880 & n24883 ) ;
  assign n24885 = n24029 | n24311 ;
  assign n24886 = ( n24029 & n24030 ) | ( n24029 & n24885 ) | ( n24030 & n24885 ) ;
  assign n24887 = n24884 | n24886 ;
  assign n24888 = n24884 & n24886 ;
  assign n24889 = n24887 & ~n24888 ;
  assign n24890 = ( n24839 & n24867 ) | ( n24839 & ~n24889 ) | ( n24867 & ~n24889 ) ;
  assign n24891 = ( ~n24867 & n24889 ) | ( ~n24867 & n24890 ) | ( n24889 & n24890 ) ;
  assign n24892 = ( ~n24839 & n24890 ) | ( ~n24839 & n24891 ) | ( n24890 & n24891 ) ;
  assign n24893 = ( n23782 & n23974 ) | ( n23782 & n23980 ) | ( n23974 & n23980 ) ;
  assign n24894 = n24530 & ~n24534 ;
  assign n24895 = n24530 & ~n24531 ;
  assign n24896 = ( ~n24893 & n24894 ) | ( ~n24893 & n24895 ) | ( n24894 & n24895 ) ;
  assign n24897 = ~n24360 & n24896 ;
  assign n24898 = n24892 & n24897 ;
  assign n24899 = ( n24539 & n24892 ) | ( n24539 & n24898 ) | ( n24892 & n24898 ) ;
  assign n24900 = n24892 | n24897 ;
  assign n24901 = n24539 | n24900 ;
  assign n24902 = ~n24899 & n24901 ;
  assign n24903 = n24510 & n24902 ;
  assign n24904 = ~n24512 & n24903 ;
  assign n24905 = ( n24514 & n24902 ) | ( n24514 & n24904 ) | ( n24902 & n24904 ) ;
  assign n24906 = n24510 | n24902 ;
  assign n24907 = ( ~n24512 & n24902 ) | ( ~n24512 & n24906 ) | ( n24902 & n24906 ) ;
  assign n24908 = n24514 | n24907 ;
  assign n24909 = ~n24905 & n24908 ;
  assign n24973 = ( n24909 & n24943 ) | ( n24909 & ~n24972 ) | ( n24943 & ~n24972 ) ;
  assign n24974 = ( ~n24943 & n24972 ) | ( ~n24943 & n24973 ) | ( n24972 & n24973 ) ;
  assign n24976 = ( ~n23940 & n24493 ) | ( ~n23940 & n24973 ) | ( n24493 & n24973 ) ;
  assign n24977 = ( n23940 & ~n24493 ) | ( n23940 & n24909 ) | ( ~n24493 & n24909 ) ;
  assign n24978 = ( n24974 & n24976 ) | ( n24974 & ~n24977 ) | ( n24976 & ~n24977 ) ;
  assign n24979 = n24493 & n24973 ;
  assign n24980 = n24493 & ~n24909 ;
  assign n24981 = ( n24974 & n24979 ) | ( n24974 & n24980 ) | ( n24979 & n24980 ) ;
  assign n24982 = ( ~n24426 & n24978 ) | ( ~n24426 & n24981 ) | ( n24978 & n24981 ) ;
  assign n24975 = ( ~n24909 & n24973 ) | ( ~n24909 & n24974 ) | ( n24973 & n24974 ) ;
  assign n24983 = n23940 | n24425 ;
  assign n24984 = n23940 | n24423 ;
  assign n24985 = ( n23941 & n24983 ) | ( n23941 & n24984 ) | ( n24983 & n24984 ) ;
  assign n24986 = ( ~n24975 & n24982 ) | ( ~n24975 & n24985 ) | ( n24982 & n24985 ) ;
  assign n24987 = ( ~n24493 & n24982 ) | ( ~n24493 & n24986 ) | ( n24982 & n24986 ) ;
  assign n24988 = n23919 & n24987 ;
  assign n24989 = ( n24436 & n24987 ) | ( n24436 & n24988 ) | ( n24987 & n24988 ) ;
  assign n24990 = n23919 | n24435 ;
  assign n24991 = n23919 | n24430 ;
  assign n24992 = ( n23920 & n24990 ) | ( n23920 & n24991 ) | ( n24990 & n24991 ) ;
  assign n24993 = ~n24989 & n24992 ;
  assign n24994 = n24987 & ~n24988 ;
  assign n24995 = ~n24436 & n24994 ;
  assign n24996 = n24993 | n24995 ;
  assign n24997 = n24457 | n24463 ;
  assign n24998 = n24457 | n24459 ;
  assign n24999 = ( n24457 & n24461 ) | ( n24457 & n24998 ) | ( n24461 & n24998 ) ;
  assign n25000 = ( n23883 & n24997 ) | ( n23883 & n24999 ) | ( n24997 & n24999 ) ;
  assign n25001 = n24996 & n25000 ;
  assign n25002 = n24457 & n24996 ;
  assign n25003 = ( n24468 & n24996 ) | ( n24468 & n25002 ) | ( n24996 & n25002 ) ;
  assign n25004 = ( n22796 & n25001 ) | ( n22796 & n25003 ) | ( n25001 & n25003 ) ;
  assign n25005 = n24457 | n24468 ;
  assign n25006 = ( n22796 & n25000 ) | ( n22796 & n25005 ) | ( n25000 & n25005 ) ;
  assign n25007 = ~n25004 & n25006 ;
  assign n25008 = ( n24996 & ~n25004 ) | ( n24996 & n25007 ) | ( ~n25004 & n25007 ) ;
  assign n25009 = n23937 & n24493 ;
  assign n25010 = n23939 & n25009 ;
  assign n25011 = ( n24425 & n24493 ) | ( n24425 & n25010 ) | ( n24493 & n25010 ) ;
  assign n25012 = ( n24423 & n24493 ) | ( n24423 & n25010 ) | ( n24493 & n25010 ) ;
  assign n25013 = ( n23941 & n25011 ) | ( n23941 & n25012 ) | ( n25011 & n25012 ) ;
  assign n25014 = n24985 & ~n25013 ;
  assign n25015 = ~n23937 & n24493 ;
  assign n25016 = ( ~n23939 & n24493 ) | ( ~n23939 & n25015 ) | ( n24493 & n25015 ) ;
  assign n25017 = n24973 & n25016 ;
  assign n25018 = ~n24909 & n25016 ;
  assign n25019 = ( n24974 & n25017 ) | ( n24974 & n25018 ) | ( n25017 & n25018 ) ;
  assign n25020 = ~n24426 & n25019 ;
  assign n25021 = ( n24975 & n25014 ) | ( n24975 & n25020 ) | ( n25014 & n25020 ) ;
  assign n25022 = x115 & n3085 ;
  assign n25023 = x114 & n3080 ;
  assign n25024 = x113 & ~n3079 ;
  assign n25025 = n3309 & n25024 ;
  assign n25026 = n25023 | n25025 ;
  assign n25027 = n25022 | n25026 ;
  assign n25028 = n3088 | n25022 ;
  assign n25029 = n25026 | n25028 ;
  assign n25030 = ( ~n12550 & n25027 ) | ( ~n12550 & n25029 ) | ( n25027 & n25029 ) ;
  assign n25031 = n25027 & n25029 ;
  assign n25032 = ( n12532 & n25030 ) | ( n12532 & n25031 ) | ( n25030 & n25031 ) ;
  assign n25033 = x26 & n25032 ;
  assign n25034 = x26 & ~n25032 ;
  assign n25035 = ( n25032 & ~n25033 ) | ( n25032 & n25034 ) | ( ~n25033 & n25034 ) ;
  assign n25036 = n24839 & n24889 ;
  assign n25037 = n24839 | n24889 ;
  assign n25038 = ~n25036 & n25037 ;
  assign n25039 = n24860 | n25038 ;
  assign n25040 = ( n24860 & n24867 ) | ( n24860 & n25039 ) | ( n24867 & n25039 ) ;
  assign n25041 = n25035 | n25040 ;
  assign n25042 = n25035 & n25040 ;
  assign n25043 = n25041 & ~n25042 ;
  assign n25044 = n24538 | n24899 ;
  assign n25045 = x118 & n2429 ;
  assign n25046 = x117 & n2424 ;
  assign n25047 = x116 & ~n2423 ;
  assign n25048 = n2631 & n25047 ;
  assign n25049 = n25046 | n25048 ;
  assign n25050 = n25045 | n25049 ;
  assign n25051 = n2432 | n25045 ;
  assign n25052 = n25049 | n25051 ;
  assign n25053 = ( ~n14002 & n25050 ) | ( ~n14002 & n25052 ) | ( n25050 & n25052 ) ;
  assign n25054 = n25050 & n25052 ;
  assign n25055 = ( n13981 & n25053 ) | ( n13981 & n25054 ) | ( n25053 & n25054 ) ;
  assign n25056 = x23 & n25055 ;
  assign n25057 = x23 & ~n25055 ;
  assign n25058 = ( n25055 & ~n25056 ) | ( n25055 & n25057 ) | ( ~n25056 & n25057 ) ;
  assign n25059 = n24537 & n25058 ;
  assign n25060 = n24530 & n25058 ;
  assign n25061 = ( n24360 & n25059 ) | ( n24360 & n25060 ) | ( n25059 & n25060 ) ;
  assign n25062 = ( n24899 & n25058 ) | ( n24899 & n25061 ) | ( n25058 & n25061 ) ;
  assign n25063 = n25044 & ~n25062 ;
  assign n25266 = n24734 | n24752 ;
  assign n25267 = ( n24734 & n24735 ) | ( n24734 & n25266 ) | ( n24735 & n25266 ) ;
  assign n25069 = x78 & n17141 ;
  assign n25070 = x77 & ~n17140 ;
  assign n25071 = n17724 & n25070 ;
  assign n25072 = n25069 | n25071 ;
  assign n25073 = x79 & n17146 ;
  assign n25074 = n17149 | n25073 ;
  assign n25075 = n25072 | n25074 ;
  assign n25076 = ~x62 & n25075 ;
  assign n25077 = ~x62 & n25073 ;
  assign n25078 = ( ~x62 & n25072 ) | ( ~x62 & n25077 ) | ( n25072 & n25077 ) ;
  assign n25079 = ( n1332 & n25076 ) | ( n1332 & n25078 ) | ( n25076 & n25078 ) ;
  assign n25080 = x62 & ~n25075 ;
  assign n25081 = x62 & x79 ;
  assign n25082 = n17146 & n25081 ;
  assign n25083 = x62 & ~n25082 ;
  assign n25084 = ~n25072 & n25083 ;
  assign n25085 = ( ~n1332 & n25080 ) | ( ~n1332 & n25084 ) | ( n25080 & n25084 ) ;
  assign n25086 = n25079 | n25085 ;
  assign n25087 = x76 & n18290 ;
  assign n25088 = x63 & x75 ;
  assign n25089 = ~n18290 & n25088 ;
  assign n25090 = n25087 | n25089 ;
  assign n25091 = x11 & n24058 ;
  assign n25092 = x11 | n24058 ;
  assign n25093 = ~n25091 & n25092 ;
  assign n25094 = n25090 & ~n25093 ;
  assign n25095 = ~n25090 & n25093 ;
  assign n25096 = n25094 | n25095 ;
  assign n25097 = n25086 & ~n25096 ;
  assign n25098 = ~n25086 & n25096 ;
  assign n25099 = n25097 | n25098 ;
  assign n25100 = ( n24062 & n24569 ) | ( n24062 & ~n24570 ) | ( n24569 & ~n24570 ) ;
  assign n25101 = ~n24566 & n25100 ;
  assign n25102 = ~n24566 & n24569 ;
  assign n25103 = ( n24566 & n24570 ) | ( n24566 & ~n25102 ) | ( n24570 & ~n25102 ) ;
  assign n25104 = ( n24053 & ~n25101 ) | ( n24053 & n25103 ) | ( ~n25101 & n25103 ) ;
  assign n25105 = ~n25099 & n25104 ;
  assign n25106 = n25099 | n25105 ;
  assign n25107 = x82 & n15552 ;
  assign n25108 = x81 & n15547 ;
  assign n25109 = x80 & ~n15546 ;
  assign n25110 = n16123 & n25109 ;
  assign n25111 = n25108 | n25110 ;
  assign n25112 = n25107 | n25111 ;
  assign n25113 = n15555 | n25107 ;
  assign n25114 = n25111 | n25113 ;
  assign n25115 = ( n1811 & n25112 ) | ( n1811 & n25114 ) | ( n25112 & n25114 ) ;
  assign n25116 = x59 & n25114 ;
  assign n25117 = x59 & n25107 ;
  assign n25118 = ( x59 & n25111 ) | ( x59 & n25117 ) | ( n25111 & n25117 ) ;
  assign n25119 = ( n1811 & n25116 ) | ( n1811 & n25118 ) | ( n25116 & n25118 ) ;
  assign n25120 = x59 & ~n25118 ;
  assign n25121 = x59 & ~n25114 ;
  assign n25122 = ( ~n1811 & n25120 ) | ( ~n1811 & n25121 ) | ( n25120 & n25121 ) ;
  assign n25123 = ( n25115 & ~n25119 ) | ( n25115 & n25122 ) | ( ~n25119 & n25122 ) ;
  assign n25124 = n25104 & n25123 ;
  assign n25125 = n25099 & n25124 ;
  assign n25126 = ( ~n25106 & n25123 ) | ( ~n25106 & n25125 ) | ( n25123 & n25125 ) ;
  assign n25127 = n25104 | n25123 ;
  assign n25128 = ( n25099 & n25123 ) | ( n25099 & n25127 ) | ( n25123 & n25127 ) ;
  assign n25129 = n25106 & ~n25128 ;
  assign n25130 = n25126 | n25129 ;
  assign n25131 = n24596 | n24616 ;
  assign n25132 = ( ~n24579 & n24616 ) | ( ~n24579 & n25131 ) | ( n24616 & n25131 ) ;
  assign n25133 = ( n24597 & ~n24599 ) | ( n24597 & n25132 ) | ( ~n24599 & n25132 ) ;
  assign n25134 = n25130 & ~n25133 ;
  assign n25135 = ~n25130 & n25133 ;
  assign n25136 = n25134 | n25135 ;
  assign n25137 = x85 & n14045 ;
  assign n25138 = x84 & n14040 ;
  assign n25139 = x83 & ~n14039 ;
  assign n25140 = n14552 & n25139 ;
  assign n25141 = n25138 | n25140 ;
  assign n25142 = n25137 | n25141 ;
  assign n25143 = n14048 | n25137 ;
  assign n25144 = n25141 | n25143 ;
  assign n25145 = ( n2381 & n25142 ) | ( n2381 & n25144 ) | ( n25142 & n25144 ) ;
  assign n25146 = x56 & n25144 ;
  assign n25147 = x56 & n25137 ;
  assign n25148 = ( x56 & n25141 ) | ( x56 & n25147 ) | ( n25141 & n25147 ) ;
  assign n25149 = ( n2381 & n25146 ) | ( n2381 & n25148 ) | ( n25146 & n25148 ) ;
  assign n25150 = x56 & ~n25148 ;
  assign n25151 = x56 & ~n25144 ;
  assign n25152 = ( ~n2381 & n25150 ) | ( ~n2381 & n25151 ) | ( n25150 & n25151 ) ;
  assign n25153 = ( n25145 & ~n25149 ) | ( n25145 & n25152 ) | ( ~n25149 & n25152 ) ;
  assign n25154 = ~n25136 & n25153 ;
  assign n25155 = n25136 | n25154 ;
  assign n25157 = n24626 & ~n24646 ;
  assign n25158 = ( n24626 & ~n24629 ) | ( n24626 & n25157 ) | ( ~n24629 & n25157 ) ;
  assign n25156 = n25136 & n25153 ;
  assign n25159 = n25156 & ~n25158 ;
  assign n25160 = ( n25155 & n25158 ) | ( n25155 & ~n25159 ) | ( n25158 & ~n25159 ) ;
  assign n25161 = ~n25156 & n25158 ;
  assign n25162 = n25155 & n25161 ;
  assign n25163 = n25160 & ~n25162 ;
  assign n25164 = x88 & n12574 ;
  assign n25165 = x87 & n12569 ;
  assign n25166 = x86 & ~n12568 ;
  assign n25167 = n13076 & n25166 ;
  assign n25168 = n25165 | n25167 ;
  assign n25169 = n25164 | n25168 ;
  assign n25170 = n12577 | n25164 ;
  assign n25171 = n25168 | n25170 ;
  assign n25172 = ( ~n3039 & n25169 ) | ( ~n3039 & n25171 ) | ( n25169 & n25171 ) ;
  assign n25173 = n25169 & n25171 ;
  assign n25174 = ( n3023 & n25172 ) | ( n3023 & n25173 ) | ( n25172 & n25173 ) ;
  assign n25175 = x53 & n25171 ;
  assign n25176 = x53 & n25164 ;
  assign n25177 = ( x53 & n25168 ) | ( x53 & n25176 ) | ( n25168 & n25176 ) ;
  assign n25178 = ( ~n3039 & n25175 ) | ( ~n3039 & n25177 ) | ( n25175 & n25177 ) ;
  assign n25179 = n25175 & n25177 ;
  assign n25180 = ( n3023 & n25178 ) | ( n3023 & n25179 ) | ( n25178 & n25179 ) ;
  assign n25181 = x53 & ~n25177 ;
  assign n25182 = x53 & ~n25171 ;
  assign n25183 = ( n3039 & n25181 ) | ( n3039 & n25182 ) | ( n25181 & n25182 ) ;
  assign n25184 = n25181 | n25182 ;
  assign n25185 = ( ~n3023 & n25183 ) | ( ~n3023 & n25184 ) | ( n25183 & n25184 ) ;
  assign n25186 = ( n25174 & ~n25180 ) | ( n25174 & n25185 ) | ( ~n25180 & n25185 ) ;
  assign n25187 = n25163 & n25186 ;
  assign n25188 = n25163 & ~n25187 ;
  assign n25189 = ~n25163 & n25186 ;
  assign n25190 = n25188 | n25189 ;
  assign n25191 = n24655 | n24678 ;
  assign n25192 = ~n25190 & n25191 ;
  assign n25193 = n25190 & ~n25191 ;
  assign n25194 = n25192 | n25193 ;
  assign n25195 = x91 & n11205 ;
  assign n25196 = x90 & n11200 ;
  assign n25197 = x89 & ~n11199 ;
  assign n25198 = n11679 & n25197 ;
  assign n25199 = n25196 | n25198 ;
  assign n25200 = n25195 | n25199 ;
  assign n25201 = n11208 | n25195 ;
  assign n25202 = n25199 | n25201 ;
  assign n25203 = ( n3768 & n25200 ) | ( n3768 & n25202 ) | ( n25200 & n25202 ) ;
  assign n25204 = x50 & n25202 ;
  assign n25205 = x50 & n25195 ;
  assign n25206 = ( x50 & n25199 ) | ( x50 & n25205 ) | ( n25199 & n25205 ) ;
  assign n25207 = ( n3768 & n25204 ) | ( n3768 & n25206 ) | ( n25204 & n25206 ) ;
  assign n25208 = x50 & ~n25206 ;
  assign n25209 = x50 & ~n25202 ;
  assign n25210 = ( ~n3768 & n25208 ) | ( ~n3768 & n25209 ) | ( n25208 & n25209 ) ;
  assign n25211 = ( n25203 & ~n25207 ) | ( n25203 & n25210 ) | ( ~n25207 & n25210 ) ;
  assign n25212 = n25194 & n25211 ;
  assign n25213 = n25194 | n25211 ;
  assign n25214 = ~n25212 & n25213 ;
  assign n25215 = n24679 | n24700 ;
  assign n25216 = ( n24680 & n24700 ) | ( n24680 & n25215 ) | ( n24700 & n25215 ) ;
  assign n25217 = ( n24681 & n24683 ) | ( n24681 & n25216 ) | ( n24683 & n25216 ) ;
  assign n25218 = n25214 | n25217 ;
  assign n25219 = n25214 & n25217 ;
  assign n25220 = n25218 & ~n25219 ;
  assign n25221 = x94 & n9933 ;
  assign n25222 = x93 & n9928 ;
  assign n25223 = x92 & ~n9927 ;
  assign n25224 = n10379 & n25223 ;
  assign n25225 = n25222 | n25224 ;
  assign n25226 = n25221 | n25225 ;
  assign n25227 = n9936 | n25221 ;
  assign n25228 = n25225 | n25227 ;
  assign n25229 = ( n4583 & n25226 ) | ( n4583 & n25228 ) | ( n25226 & n25228 ) ;
  assign n25230 = x47 & n25228 ;
  assign n25231 = x47 & n25221 ;
  assign n25232 = ( x47 & n25225 ) | ( x47 & n25231 ) | ( n25225 & n25231 ) ;
  assign n25233 = ( n4583 & n25230 ) | ( n4583 & n25232 ) | ( n25230 & n25232 ) ;
  assign n25234 = x47 & ~n25232 ;
  assign n25235 = x47 & ~n25228 ;
  assign n25236 = ( ~n4583 & n25234 ) | ( ~n4583 & n25235 ) | ( n25234 & n25235 ) ;
  assign n25237 = ( n25229 & ~n25233 ) | ( n25229 & n25236 ) | ( ~n25233 & n25236 ) ;
  assign n25238 = n25220 & n25237 ;
  assign n25240 = n24703 | n24726 ;
  assign n25241 = ( n24706 & n24726 ) | ( n24706 & n25240 ) | ( n24726 & n25240 ) ;
  assign n25242 = ( n24707 & n24709 ) | ( n24707 & n25241 ) | ( n24709 & n25241 ) ;
  assign n25239 = n25220 | n25237 ;
  assign n25243 = n25239 & n25242 ;
  assign n25244 = n25238 & n25242 ;
  assign n25245 = ( n25242 & ~n25243 ) | ( n25242 & n25244 ) | ( ~n25243 & n25244 ) ;
  assign n25246 = ( n25220 & n25237 ) | ( n25220 & ~n25239 ) | ( n25237 & ~n25239 ) ;
  assign n25247 = ( n25239 & ~n25242 ) | ( n25239 & n25246 ) | ( ~n25242 & n25246 ) ;
  assign n25248 = ( ~n25238 & n25245 ) | ( ~n25238 & n25247 ) | ( n25245 & n25247 ) ;
  assign n25249 = x97 & n8724 ;
  assign n25250 = x96 & n8719 ;
  assign n25251 = x95 & ~n8718 ;
  assign n25252 = n9149 & n25251 ;
  assign n25253 = n25250 | n25252 ;
  assign n25254 = n25249 | n25253 ;
  assign n25255 = n8727 | n25249 ;
  assign n25256 = n25253 | n25255 ;
  assign n25257 = ( n5505 & n25254 ) | ( n5505 & n25256 ) | ( n25254 & n25256 ) ;
  assign n25258 = x44 & n25256 ;
  assign n25259 = x44 & n25249 ;
  assign n25260 = ( x44 & n25253 ) | ( x44 & n25259 ) | ( n25253 & n25259 ) ;
  assign n25261 = ( n5505 & n25258 ) | ( n5505 & n25260 ) | ( n25258 & n25260 ) ;
  assign n25262 = x44 & ~n25260 ;
  assign n25263 = x44 & ~n25256 ;
  assign n25264 = ( ~n5505 & n25262 ) | ( ~n5505 & n25263 ) | ( n25262 & n25263 ) ;
  assign n25265 = ( n25257 & ~n25261 ) | ( n25257 & n25264 ) | ( ~n25261 & n25264 ) ;
  assign n25268 = ( n25248 & ~n25265 ) | ( n25248 & n25267 ) | ( ~n25265 & n25267 ) ;
  assign n25269 = ( ~n25248 & n25265 ) | ( ~n25248 & n25267 ) | ( n25265 & n25267 ) ;
  assign n25270 = ( ~n25267 & n25268 ) | ( ~n25267 & n25269 ) | ( n25268 & n25269 ) ;
  assign n25271 = x100 & n7566 ;
  assign n25272 = x99 & n7561 ;
  assign n25273 = x98 & ~n7560 ;
  assign n25274 = n7953 & n25273 ;
  assign n25275 = n25272 | n25274 ;
  assign n25276 = n25271 | n25275 ;
  assign n25277 = n7569 | n25271 ;
  assign n25278 = n25275 | n25277 ;
  assign n25279 = ( n6483 & n25276 ) | ( n6483 & n25278 ) | ( n25276 & n25278 ) ;
  assign n25280 = x41 & n25278 ;
  assign n25281 = x41 & n25271 ;
  assign n25282 = ( x41 & n25275 ) | ( x41 & n25281 ) | ( n25275 & n25281 ) ;
  assign n25283 = ( n6483 & n25280 ) | ( n6483 & n25282 ) | ( n25280 & n25282 ) ;
  assign n25284 = x41 & ~n25282 ;
  assign n25285 = x41 & ~n25278 ;
  assign n25286 = ( ~n6483 & n25284 ) | ( ~n6483 & n25285 ) | ( n25284 & n25285 ) ;
  assign n25287 = ( n25279 & ~n25283 ) | ( n25279 & n25286 ) | ( ~n25283 & n25286 ) ;
  assign n25288 = n25270 & n25287 ;
  assign n25289 = n25270 | n25287 ;
  assign n25290 = ~n25288 & n25289 ;
  assign n25291 = n24757 | n24777 ;
  assign n25292 = ( n24755 & n24777 ) | ( n24755 & n25291 ) | ( n24777 & n25291 ) ;
  assign n25293 = ( n24758 & n24760 ) | ( n24758 & n25292 ) | ( n24760 & n25292 ) ;
  assign n25294 = n25290 | n25293 ;
  assign n25295 = n25290 & n25293 ;
  assign n25296 = n25294 & ~n25295 ;
  assign n25297 = x103 & n6536 ;
  assign n25298 = x102 & n6531 ;
  assign n25299 = x101 & ~n6530 ;
  assign n25300 = n6871 & n25299 ;
  assign n25301 = n25298 | n25300 ;
  assign n25302 = n25297 | n25301 ;
  assign n25303 = n6539 | n25297 ;
  assign n25304 = n25301 | n25303 ;
  assign n25305 = ( n7529 & n25302 ) | ( n7529 & n25304 ) | ( n25302 & n25304 ) ;
  assign n25306 = x38 & n25304 ;
  assign n25307 = x38 & n25297 ;
  assign n25308 = ( x38 & n25301 ) | ( x38 & n25307 ) | ( n25301 & n25307 ) ;
  assign n25309 = ( n7529 & n25306 ) | ( n7529 & n25308 ) | ( n25306 & n25308 ) ;
  assign n25310 = x38 & ~n25308 ;
  assign n25311 = x38 & ~n25304 ;
  assign n25312 = ( ~n7529 & n25310 ) | ( ~n7529 & n25311 ) | ( n25310 & n25311 ) ;
  assign n25313 = ( n25305 & ~n25309 ) | ( n25305 & n25312 ) | ( ~n25309 & n25312 ) ;
  assign n25314 = n25296 & n25313 ;
  assign n25315 = n25296 & ~n25314 ;
  assign n25316 = ~n25296 & n25313 ;
  assign n25317 = n25315 | n25316 ;
  assign n25318 = n24783 | n24803 ;
  assign n25319 = ( n24780 & n24803 ) | ( n24780 & n25318 ) | ( n24803 & n25318 ) ;
  assign n25320 = ( n24785 & n24786 ) | ( n24785 & n25319 ) | ( n24786 & n25319 ) ;
  assign n25321 = ~n25317 & n25320 ;
  assign n25322 = n25317 & ~n25320 ;
  assign n25323 = n25321 | n25322 ;
  assign n25324 = x106 & n5554 ;
  assign n25325 = x105 & n5549 ;
  assign n25326 = x104 & ~n5548 ;
  assign n25327 = n5893 & n25326 ;
  assign n25328 = n25325 | n25327 ;
  assign n25329 = n25324 | n25328 ;
  assign n25330 = n5557 | n25324 ;
  assign n25331 = n25328 | n25330 ;
  assign n25332 = ( n8656 & n25329 ) | ( n8656 & n25331 ) | ( n25329 & n25331 ) ;
  assign n25333 = x35 & n25331 ;
  assign n25334 = x35 & n25324 ;
  assign n25335 = ( x35 & n25328 ) | ( x35 & n25334 ) | ( n25328 & n25334 ) ;
  assign n25336 = ( n8656 & n25333 ) | ( n8656 & n25335 ) | ( n25333 & n25335 ) ;
  assign n25337 = x35 & ~n25335 ;
  assign n25338 = x35 & ~n25331 ;
  assign n25339 = ( ~n8656 & n25337 ) | ( ~n8656 & n25338 ) | ( n25337 & n25338 ) ;
  assign n25340 = ( n25332 & ~n25336 ) | ( n25332 & n25339 ) | ( ~n25336 & n25339 ) ;
  assign n25341 = n25323 & n25340 ;
  assign n25342 = n25323 | n25340 ;
  assign n25343 = ~n25341 & n25342 ;
  assign n25344 = n24813 | n24833 ;
  assign n25345 = ( n24806 & n24833 ) | ( n24806 & n25344 ) | ( n24833 & n25344 ) ;
  assign n25346 = ( n24814 & n24816 ) | ( n24814 & n25345 ) | ( n24816 & n25345 ) ;
  assign n25347 = n25343 | n25346 ;
  assign n25348 = n25343 & n25346 ;
  assign n25349 = n25347 & ~n25348 ;
  assign n25350 = n24561 & n24836 ;
  assign n25351 = n24558 | n25350 ;
  assign n25352 = x109 & n4631 ;
  assign n25353 = x108 & n4626 ;
  assign n25354 = x107 & ~n4625 ;
  assign n25355 = n4943 & n25354 ;
  assign n25356 = n25353 | n25355 ;
  assign n25357 = n25352 | n25356 ;
  assign n25358 = n4634 | n25352 ;
  assign n25359 = n25356 | n25358 ;
  assign n25360 = ( n9878 & n25357 ) | ( n9878 & n25359 ) | ( n25357 & n25359 ) ;
  assign n25361 = x32 & n25359 ;
  assign n25362 = x32 & n25352 ;
  assign n25363 = ( x32 & n25356 ) | ( x32 & n25362 ) | ( n25356 & n25362 ) ;
  assign n25364 = ( n9878 & n25361 ) | ( n9878 & n25363 ) | ( n25361 & n25363 ) ;
  assign n25365 = x32 & ~n25363 ;
  assign n25366 = x32 & ~n25359 ;
  assign n25367 = ( ~n9878 & n25365 ) | ( ~n9878 & n25366 ) | ( n25365 & n25366 ) ;
  assign n25368 = ( n25360 & ~n25364 ) | ( n25360 & n25367 ) | ( ~n25364 & n25367 ) ;
  assign n25369 = n24557 & n25368 ;
  assign n25370 = n24556 & n25368 ;
  assign n25371 = ( n24308 & n25369 ) | ( n24308 & n25370 ) | ( n25369 & n25370 ) ;
  assign n25372 = ( n25350 & n25368 ) | ( n25350 & n25371 ) | ( n25368 & n25371 ) ;
  assign n25373 = n25351 & ~n25372 ;
  assign n25374 = ~n24557 & n25368 ;
  assign n25375 = ~n24556 & n25368 ;
  assign n25376 = ( ~n24308 & n25374 ) | ( ~n24308 & n25375 ) | ( n25374 & n25375 ) ;
  assign n25377 = ~n25350 & n25376 ;
  assign n25378 = n25349 & n25377 ;
  assign n25379 = ( n25349 & n25373 ) | ( n25349 & n25378 ) | ( n25373 & n25378 ) ;
  assign n25380 = n25349 | n25377 ;
  assign n25381 = n25373 | n25380 ;
  assign n25382 = ~n25379 & n25381 ;
  assign n25383 = x112 & n3816 ;
  assign n25384 = x111 & n3811 ;
  assign n25385 = x110 & ~n3810 ;
  assign n25386 = n4067 & n25385 ;
  assign n25387 = n25384 | n25386 ;
  assign n25388 = n25383 | n25387 ;
  assign n25389 = n3819 | n25383 ;
  assign n25390 = n25387 | n25389 ;
  assign n25391 = ( n11172 & n25388 ) | ( n11172 & n25390 ) | ( n25388 & n25390 ) ;
  assign n25392 = x29 & n25390 ;
  assign n25393 = x29 & n25383 ;
  assign n25394 = ( x29 & n25387 ) | ( x29 & n25393 ) | ( n25387 & n25393 ) ;
  assign n25395 = ( n11172 & n25392 ) | ( n11172 & n25394 ) | ( n25392 & n25394 ) ;
  assign n25396 = x29 & ~n25394 ;
  assign n25397 = x29 & ~n25390 ;
  assign n25398 = ( ~n11172 & n25396 ) | ( ~n11172 & n25397 ) | ( n25396 & n25397 ) ;
  assign n25399 = ( n25391 & ~n25395 ) | ( n25391 & n25398 ) | ( ~n25395 & n25398 ) ;
  assign n25400 = n24839 | n24888 ;
  assign n25401 = ( n24888 & n24889 ) | ( n24888 & n25400 ) | ( n24889 & n25400 ) ;
  assign n25402 = ~n25399 & n25401 ;
  assign n25403 = n25399 & ~n25401 ;
  assign n25404 = n25402 | n25403 ;
  assign n25405 = n25382 & n25404 ;
  assign n25406 = n25404 & ~n25405 ;
  assign n25407 = ( n25382 & ~n25405 ) | ( n25382 & n25406 ) | ( ~n25405 & n25406 ) ;
  assign n25408 = n25043 & n25407 ;
  assign n25409 = n25043 | n25407 ;
  assign n25064 = n25058 & ~n25060 ;
  assign n25065 = ~n24537 & n25058 ;
  assign n25066 = ( ~n24360 & n25064 ) | ( ~n24360 & n25065 ) | ( n25064 & n25065 ) ;
  assign n25410 = ( n25043 & ~n25066 ) | ( n25043 & n25407 ) | ( ~n25066 & n25407 ) ;
  assign n25411 = ( n24899 & n25409 ) | ( n24899 & n25410 ) | ( n25409 & n25410 ) ;
  assign n25412 = ( ~n25063 & n25408 ) | ( ~n25063 & n25411 ) | ( n25408 & n25411 ) ;
  assign n25067 = ~n24899 & n25066 ;
  assign n25068 = n25063 | n25067 ;
  assign n25413 = ( n25068 & ~n25407 ) | ( n25068 & n25412 ) | ( ~n25407 & n25412 ) ;
  assign n25414 = ( ~n25043 & n25412 ) | ( ~n25043 & n25413 ) | ( n25412 & n25413 ) ;
  assign n25415 = x124 & n1383 ;
  assign n25416 = x123 & n1378 ;
  assign n25417 = x122 & ~n1377 ;
  assign n25418 = n1542 & n25417 ;
  assign n25419 = n25416 | n25418 ;
  assign n25420 = n25415 | n25419 ;
  assign n25421 = n1386 | n25415 ;
  assign n25422 = n25419 | n25421 ;
  assign n25423 = ( n17084 & n25420 ) | ( n17084 & n25422 ) | ( n25420 & n25422 ) ;
  assign n25424 = x17 & n25422 ;
  assign n25425 = x17 & n25415 ;
  assign n25426 = ( x17 & n25419 ) | ( x17 & n25425 ) | ( n25419 & n25425 ) ;
  assign n25427 = ( n17084 & n25424 ) | ( n17084 & n25426 ) | ( n25424 & n25426 ) ;
  assign n25428 = x17 & ~n25426 ;
  assign n25429 = x17 & ~n25422 ;
  assign n25430 = ( ~n17084 & n25428 ) | ( ~n17084 & n25429 ) | ( n25428 & n25429 ) ;
  assign n25431 = ( n25423 & ~n25427 ) | ( n25423 & n25430 ) | ( ~n25427 & n25430 ) ;
  assign n25432 = n24909 | n24971 ;
  assign n25433 = ( n24971 & n24972 ) | ( n24971 & n25432 ) | ( n24972 & n25432 ) ;
  assign n25434 = ~n25431 & n25433 ;
  assign n25435 = n25431 & ~n25433 ;
  assign n25436 = n25434 | n25435 ;
  assign n25437 = x121 & n1859 ;
  assign n25438 = x120 & n1854 ;
  assign n25439 = x119 & ~n1853 ;
  assign n25440 = n2037 & n25439 ;
  assign n25441 = n25438 | n25440 ;
  assign n25442 = n25437 | n25441 ;
  assign n25443 = n1862 | n25437 ;
  assign n25444 = n25441 | n25443 ;
  assign n25445 = ( n15501 & n25442 ) | ( n15501 & n25444 ) | ( n25442 & n25444 ) ;
  assign n25446 = x20 & n25444 ;
  assign n25447 = x20 & n25437 ;
  assign n25448 = ( x20 & n25441 ) | ( x20 & n25447 ) | ( n25441 & n25447 ) ;
  assign n25449 = ( n15501 & n25446 ) | ( n15501 & n25448 ) | ( n25446 & n25448 ) ;
  assign n25450 = x20 & ~n25448 ;
  assign n25451 = x20 & ~n25444 ;
  assign n25452 = ( ~n15501 & n25450 ) | ( ~n15501 & n25451 ) | ( n25450 & n25451 ) ;
  assign n25453 = ( n25445 & ~n25449 ) | ( n25445 & n25452 ) | ( ~n25449 & n25452 ) ;
  assign n25454 = n24510 & n25453 ;
  assign n25455 = n24512 & n25454 ;
  assign n25456 = ( n24904 & n25453 ) | ( n24904 & n25455 ) | ( n25453 & n25455 ) ;
  assign n25457 = ( n24902 & n25453 ) | ( n24902 & n25455 ) | ( n25453 & n25455 ) ;
  assign n25458 = ( n24514 & n25456 ) | ( n24514 & n25457 ) | ( n25456 & n25457 ) ;
  assign n25459 = n24510 | n25453 ;
  assign n25460 = ( n24512 & n25453 ) | ( n24512 & n25459 ) | ( n25453 & n25459 ) ;
  assign n25461 = n24904 | n25460 ;
  assign n25462 = n24902 | n25460 ;
  assign n25463 = ( n24514 & n25461 ) | ( n24514 & n25462 ) | ( n25461 & n25462 ) ;
  assign n25464 = ~n25458 & n25463 ;
  assign n25465 = ( n25414 & n25436 ) | ( n25414 & ~n25464 ) | ( n25436 & ~n25464 ) ;
  assign n25466 = ( ~n25436 & n25464 ) | ( ~n25436 & n25465 ) | ( n25464 & n25465 ) ;
  assign n25467 = ( ~n25414 & n25465 ) | ( ~n25414 & n25466 ) | ( n25465 & n25466 ) ;
  assign n25468 = x127 & n962 ;
  assign n25469 = x126 & n957 ;
  assign n25470 = x125 & ~n956 ;
  assign n25471 = n1105 & n25470 ;
  assign n25472 = n25469 | n25471 ;
  assign n25473 = n25468 | n25472 ;
  assign n25474 = n965 | n25468 ;
  assign n25475 = n25472 | n25474 ;
  assign n25476 = ( n18763 & n25473 ) | ( n18763 & n25475 ) | ( n25473 & n25475 ) ;
  assign n25477 = x14 & n25475 ;
  assign n25478 = x14 & n25468 ;
  assign n25479 = ( x14 & n25472 ) | ( x14 & n25478 ) | ( n25472 & n25478 ) ;
  assign n25480 = ( n18763 & n25477 ) | ( n18763 & n25479 ) | ( n25477 & n25479 ) ;
  assign n25481 = x14 & ~n25479 ;
  assign n25482 = x14 & ~n25475 ;
  assign n25483 = ( ~n18763 & n25481 ) | ( ~n18763 & n25482 ) | ( n25481 & n25482 ) ;
  assign n25484 = ( n25476 & ~n25480 ) | ( n25476 & n25483 ) | ( ~n25480 & n25483 ) ;
  assign n25485 = n24909 & n24972 ;
  assign n25486 = n24909 | n24972 ;
  assign n25487 = ~n25485 & n25486 ;
  assign n25488 = n24933 | n25487 ;
  assign n25489 = n24926 | n25487 ;
  assign n25490 = ( n24420 & n25488 ) | ( n24420 & n25489 ) | ( n25488 & n25489 ) ;
  assign n25491 = ( n24934 & n24943 ) | ( n24934 & n25490 ) | ( n24943 & n25490 ) ;
  assign n25492 = ( n25467 & n25484 ) | ( n25467 & ~n25491 ) | ( n25484 & ~n25491 ) ;
  assign n25493 = ( n25467 & ~n25484 ) | ( n25467 & n25491 ) | ( ~n25484 & n25491 ) ;
  assign n25494 = ( ~n25467 & n25492 ) | ( ~n25467 & n25493 ) | ( n25492 & n25493 ) ;
  assign n25495 = n25013 & n25494 ;
  assign n25496 = ( n25021 & n25494 ) | ( n25021 & n25495 ) | ( n25494 & n25495 ) ;
  assign n25497 = n25013 | n25020 ;
  assign n25498 = n24975 | n25013 ;
  assign n25499 = ( n25014 & n25497 ) | ( n25014 & n25498 ) | ( n25497 & n25498 ) ;
  assign n25500 = ~n25496 & n25499 ;
  assign n25501 = n24989 | n25002 ;
  assign n25502 = n24989 | n24995 ;
  assign n25503 = n24993 | n25502 ;
  assign n25504 = ( n24468 & n25501 ) | ( n24468 & n25503 ) | ( n25501 & n25503 ) ;
  assign n25505 = ( n24989 & n25000 ) | ( n24989 & n25503 ) | ( n25000 & n25503 ) ;
  assign n25506 = ( n22796 & n25504 ) | ( n22796 & n25505 ) | ( n25504 & n25505 ) ;
  assign n25507 = ~n25013 & n25494 ;
  assign n25508 = ~n25021 & n25507 ;
  assign n25509 = n25506 | n25508 ;
  assign n25510 = n25500 | n25509 ;
  assign n25511 = n25500 | n25508 ;
  assign n25512 = n25503 & n25511 ;
  assign n25513 = n24989 & n25511 ;
  assign n25514 = ( n25002 & n25511 ) | ( n25002 & n25513 ) | ( n25511 & n25513 ) ;
  assign n25515 = ( n24468 & n25512 ) | ( n24468 & n25514 ) | ( n25512 & n25514 ) ;
  assign n25516 = ( n24999 & n25512 ) | ( n24999 & n25513 ) | ( n25512 & n25513 ) ;
  assign n25517 = ( n24997 & n25512 ) | ( n24997 & n25513 ) | ( n25512 & n25513 ) ;
  assign n25518 = ( n23883 & n25516 ) | ( n23883 & n25517 ) | ( n25516 & n25517 ) ;
  assign n25519 = ( n22786 & n25515 ) | ( n22786 & n25518 ) | ( n25515 & n25518 ) ;
  assign n25520 = n25514 & n25518 ;
  assign n25521 = n25512 & n25518 ;
  assign n25522 = ( n24468 & n25520 ) | ( n24468 & n25521 ) | ( n25520 & n25521 ) ;
  assign n25523 = ( n22794 & n25519 ) | ( n22794 & n25522 ) | ( n25519 & n25522 ) ;
  assign n25524 = n25510 & ~n25523 ;
  assign n25525 = n25484 & n25490 ;
  assign n25526 = n24934 & n25484 ;
  assign n25527 = ( n24943 & n25525 ) | ( n24943 & n25526 ) | ( n25525 & n25526 ) ;
  assign n25528 = n25491 & ~n25527 ;
  assign n25529 = n25484 & ~n25490 ;
  assign n25530 = ~n24934 & n25484 ;
  assign n25531 = ( ~n24943 & n25529 ) | ( ~n24943 & n25530 ) | ( n25529 & n25530 ) ;
  assign n25532 = n25467 & ~n25531 ;
  assign n25533 = ~n25528 & n25532 ;
  assign n25534 = ( n25467 & n25527 ) | ( n25467 & ~n25533 ) | ( n25527 & ~n25533 ) ;
  assign n25535 = n25431 & n25433 ;
  assign n25536 = n25414 & n25464 ;
  assign n25537 = n25414 | n25464 ;
  assign n25538 = ~n25536 & n25537 ;
  assign n25539 = n25431 | n25538 ;
  assign n25540 = ( n25433 & n25538 ) | ( n25433 & n25539 ) | ( n25538 & n25539 ) ;
  assign n25541 = ( n25436 & n25535 ) | ( n25436 & n25540 ) | ( n25535 & n25540 ) ;
  assign n25542 = x127 & n957 ;
  assign n25543 = x126 & ~n956 ;
  assign n25544 = n1105 & n25543 ;
  assign n25545 = n25542 | n25544 ;
  assign n25546 = n965 | n25545 ;
  assign n25547 = ( n19328 & n25545 ) | ( n19328 & n25546 ) | ( n25545 & n25546 ) ;
  assign n25548 = x14 & n25545 ;
  assign n25549 = ( x14 & n2082 ) | ( x14 & n25545 ) | ( n2082 & n25545 ) ;
  assign n25550 = ( n19328 & n25548 ) | ( n19328 & n25549 ) | ( n25548 & n25549 ) ;
  assign n25551 = x14 & ~n2082 ;
  assign n25552 = ~n25545 & n25551 ;
  assign n25553 = x14 & ~n25545 ;
  assign n25554 = ( ~n19328 & n25552 ) | ( ~n19328 & n25553 ) | ( n25552 & n25553 ) ;
  assign n25555 = ( n25547 & ~n25550 ) | ( n25547 & n25554 ) | ( ~n25550 & n25554 ) ;
  assign n25556 = n25540 & n25555 ;
  assign n25557 = n25535 & n25555 ;
  assign n25558 = ( n25436 & n25556 ) | ( n25436 & n25557 ) | ( n25556 & n25557 ) ;
  assign n25559 = n25541 & ~n25558 ;
  assign n25577 = n25414 | n25458 ;
  assign n25578 = ( n25458 & n25464 ) | ( n25458 & n25577 ) | ( n25464 & n25577 ) ;
  assign n25560 = x125 & n1383 ;
  assign n25561 = x124 & n1378 ;
  assign n25562 = x123 & ~n1377 ;
  assign n25563 = n1542 & n25562 ;
  assign n25564 = n25561 | n25563 ;
  assign n25565 = n25560 | n25564 ;
  assign n25566 = n1386 | n25560 ;
  assign n25567 = n25564 | n25566 ;
  assign n25568 = ( n17670 & n25565 ) | ( n17670 & n25567 ) | ( n25565 & n25567 ) ;
  assign n25569 = x17 & n25567 ;
  assign n25570 = x17 & n25560 ;
  assign n25571 = ( x17 & n25564 ) | ( x17 & n25570 ) | ( n25564 & n25570 ) ;
  assign n25572 = ( n17670 & n25569 ) | ( n17670 & n25571 ) | ( n25569 & n25571 ) ;
  assign n25573 = x17 & ~n25571 ;
  assign n25574 = x17 & ~n25567 ;
  assign n25575 = ( ~n17670 & n25573 ) | ( ~n17670 & n25574 ) | ( n25573 & n25574 ) ;
  assign n25576 = ( n25568 & ~n25572 ) | ( n25568 & n25575 ) | ( ~n25572 & n25575 ) ;
  assign n25579 = n25576 & n25578 ;
  assign n25580 = n25578 & ~n25579 ;
  assign n25582 = x121 & n1854 ;
  assign n25583 = x120 & ~n1853 ;
  assign n25584 = n2037 & n25583 ;
  assign n25585 = n25582 | n25584 ;
  assign n25581 = x122 & n1859 ;
  assign n25587 = n1862 | n25581 ;
  assign n25588 = n25585 | n25587 ;
  assign n25586 = n25581 | n25585 ;
  assign n25589 = n25586 & n25588 ;
  assign n25590 = ( n16043 & n25588 ) | ( n16043 & n25589 ) | ( n25588 & n25589 ) ;
  assign n25591 = x20 & n25589 ;
  assign n25592 = x20 & n25588 ;
  assign n25593 = ( n16043 & n25591 ) | ( n16043 & n25592 ) | ( n25591 & n25592 ) ;
  assign n25594 = x20 & ~n25589 ;
  assign n25595 = x20 & ~n25588 ;
  assign n25596 = ( ~n16043 & n25594 ) | ( ~n16043 & n25595 ) | ( n25594 & n25595 ) ;
  assign n25597 = ( n25590 & ~n25593 ) | ( n25590 & n25596 ) | ( ~n25593 & n25596 ) ;
  assign n25598 = n25066 & n25409 ;
  assign n25599 = ~n24899 & n25598 ;
  assign n25600 = ~n25061 & n25408 ;
  assign n25601 = ~n25058 & n25407 ;
  assign n25602 = n25043 & n25601 ;
  assign n25603 = ( ~n24899 & n25600 ) | ( ~n24899 & n25602 ) | ( n25600 & n25602 ) ;
  assign n25604 = ( n25062 & n25599 ) | ( n25062 & ~n25603 ) | ( n25599 & ~n25603 ) ;
  assign n25605 = ( n25062 & n25409 ) | ( n25062 & ~n25603 ) | ( n25409 & ~n25603 ) ;
  assign n25606 = ( n25063 & n25604 ) | ( n25063 & n25605 ) | ( n25604 & n25605 ) ;
  assign n25607 = n25597 & n25606 ;
  assign n25608 = n25597 | n25606 ;
  assign n25609 = ~n25607 & n25608 ;
  assign n25627 = n25042 | n25407 ;
  assign n25628 = ( n25042 & n25043 ) | ( n25042 & n25627 ) | ( n25043 & n25627 ) ;
  assign n25610 = x119 & n2429 ;
  assign n25611 = x118 & n2424 ;
  assign n25612 = x117 & ~n2423 ;
  assign n25613 = n2631 & n25612 ;
  assign n25614 = n25611 | n25613 ;
  assign n25615 = n25610 | n25614 ;
  assign n25616 = n2432 | n25610 ;
  assign n25617 = n25614 | n25616 ;
  assign n25618 = ( n14496 & n25615 ) | ( n14496 & n25617 ) | ( n25615 & n25617 ) ;
  assign n25619 = x23 & n25617 ;
  assign n25620 = x23 & n25610 ;
  assign n25621 = ( x23 & n25614 ) | ( x23 & n25620 ) | ( n25614 & n25620 ) ;
  assign n25622 = ( n14496 & n25619 ) | ( n14496 & n25621 ) | ( n25619 & n25621 ) ;
  assign n25623 = x23 & ~n25621 ;
  assign n25624 = x23 & ~n25617 ;
  assign n25625 = ( ~n14496 & n25623 ) | ( ~n14496 & n25624 ) | ( n25623 & n25624 ) ;
  assign n25626 = ( n25618 & ~n25622 ) | ( n25618 & n25625 ) | ( ~n25622 & n25625 ) ;
  assign n25629 = n25626 & n25628 ;
  assign n25630 = n25628 & ~n25629 ;
  assign n25632 = x115 & n3080 ;
  assign n25633 = x114 & ~n3079 ;
  assign n25634 = n3309 & n25633 ;
  assign n25635 = n25632 | n25634 ;
  assign n25631 = x116 & n3085 ;
  assign n25637 = n3088 | n25631 ;
  assign n25638 = n25635 | n25637 ;
  assign n25636 = n25631 | n25635 ;
  assign n25639 = n25636 & n25638 ;
  assign n25640 = ( ~n13040 & n25638 ) | ( ~n13040 & n25639 ) | ( n25638 & n25639 ) ;
  assign n25641 = n25638 & n25639 ;
  assign n25642 = ( n13022 & n25640 ) | ( n13022 & n25641 ) | ( n25640 & n25641 ) ;
  assign n25643 = x26 & n25642 ;
  assign n25644 = x26 & ~n25642 ;
  assign n25645 = ( n25642 & ~n25643 ) | ( n25642 & n25644 ) | ( ~n25643 & n25644 ) ;
  assign n25646 = n25399 & n25401 ;
  assign n25647 = n25382 | n25646 ;
  assign n25648 = ( n25404 & n25646 ) | ( n25404 & n25647 ) | ( n25646 & n25647 ) ;
  assign n25649 = n25645 & n25648 ;
  assign n25650 = n25645 | n25648 ;
  assign n25651 = ~n25649 & n25650 ;
  assign n25652 = n25372 | n25379 ;
  assign n25653 = x113 & n3816 ;
  assign n25654 = x112 & n3811 ;
  assign n25655 = x111 & ~n3810 ;
  assign n25656 = n4067 & n25655 ;
  assign n25657 = n25654 | n25656 ;
  assign n25658 = n25653 | n25657 ;
  assign n25659 = n3819 | n25653 ;
  assign n25660 = n25657 | n25659 ;
  assign n25661 = ( ~n11642 & n25658 ) | ( ~n11642 & n25660 ) | ( n25658 & n25660 ) ;
  assign n25662 = n25658 & n25660 ;
  assign n25663 = ( n11626 & n25661 ) | ( n11626 & n25662 ) | ( n25661 & n25662 ) ;
  assign n25664 = x29 & n25663 ;
  assign n25665 = x29 & ~n25663 ;
  assign n25666 = ( n25663 & ~n25664 ) | ( n25663 & n25665 ) | ( ~n25664 & n25665 ) ;
  assign n25667 = n25371 & n25666 ;
  assign n25668 = n25368 & n25666 ;
  assign n25669 = ( n25350 & n25667 ) | ( n25350 & n25668 ) | ( n25667 & n25668 ) ;
  assign n25670 = ( n25379 & n25666 ) | ( n25379 & n25669 ) | ( n25666 & n25669 ) ;
  assign n25671 = n25652 & ~n25670 ;
  assign n25672 = n25341 | n25346 ;
  assign n25673 = ( n25341 & n25343 ) | ( n25341 & n25672 ) | ( n25343 & n25672 ) ;
  assign n25675 = x109 & n4626 ;
  assign n25676 = x108 & ~n4625 ;
  assign n25677 = n4943 & n25676 ;
  assign n25678 = n25675 | n25677 ;
  assign n25674 = x110 & n4631 ;
  assign n25680 = n4634 | n25674 ;
  assign n25681 = n25678 | n25680 ;
  assign n25679 = n25674 | n25678 ;
  assign n25682 = n25679 & n25681 ;
  assign n25683 = ( n10330 & n25681 ) | ( n10330 & n25682 ) | ( n25681 & n25682 ) ;
  assign n25684 = x32 & n25682 ;
  assign n25685 = x32 & n25681 ;
  assign n25686 = ( n10330 & n25684 ) | ( n10330 & n25685 ) | ( n25684 & n25685 ) ;
  assign n25687 = x32 & ~n25682 ;
  assign n25688 = x32 & ~n25681 ;
  assign n25689 = ( ~n10330 & n25687 ) | ( ~n10330 & n25688 ) | ( n25687 & n25688 ) ;
  assign n25690 = ( n25683 & ~n25686 ) | ( n25683 & n25689 ) | ( ~n25686 & n25689 ) ;
  assign n25691 = n25340 & n25690 ;
  assign n25692 = n25323 & n25691 ;
  assign n25693 = ( n25346 & n25690 ) | ( n25346 & n25692 ) | ( n25690 & n25692 ) ;
  assign n25694 = n25690 & n25692 ;
  assign n25695 = ( n25343 & n25693 ) | ( n25343 & n25694 ) | ( n25693 & n25694 ) ;
  assign n25696 = n25673 & ~n25695 ;
  assign n25886 = ~n25247 & n25265 ;
  assign n25887 = n25238 & n25265 ;
  assign n25888 = ( ~n25245 & n25886 ) | ( ~n25245 & n25887 ) | ( n25886 & n25887 ) ;
  assign n25889 = n25267 & ~n25888 ;
  assign n25890 = n25247 & n25265 ;
  assign n25891 = ~n25238 & n25265 ;
  assign n25892 = ( n25245 & n25890 ) | ( n25245 & n25891 ) | ( n25890 & n25891 ) ;
  assign n25893 = n25248 & ~n25892 ;
  assign n25894 = ( n25267 & n25892 ) | ( n25267 & n25893 ) | ( n25892 & n25893 ) ;
  assign n25895 = n25267 | n25892 ;
  assign n25896 = ( ~n25889 & n25894 ) | ( ~n25889 & n25895 ) | ( n25894 & n25895 ) ;
  assign n25850 = n25212 | n25217 ;
  assign n25851 = ( n25212 & n25214 ) | ( n25212 & n25850 ) | ( n25214 & n25850 ) ;
  assign n25697 = x79 & n17141 ;
  assign n25698 = x78 & ~n17140 ;
  assign n25699 = n17724 & n25698 ;
  assign n25700 = n25697 | n25699 ;
  assign n25701 = x80 & n17146 ;
  assign n25702 = n17149 | n25701 ;
  assign n25703 = n25700 | n25702 ;
  assign n25704 = ~x62 & n25703 ;
  assign n25705 = ~x62 & n25701 ;
  assign n25706 = ( ~x62 & n25700 ) | ( ~x62 & n25705 ) | ( n25700 & n25705 ) ;
  assign n25707 = ( n1499 & n25704 ) | ( n1499 & n25706 ) | ( n25704 & n25706 ) ;
  assign n25708 = x62 & ~n25703 ;
  assign n25709 = x62 & x80 ;
  assign n25710 = n17146 & n25709 ;
  assign n25711 = x62 & ~n25710 ;
  assign n25712 = ~n25700 & n25711 ;
  assign n25713 = ( ~n1499 & n25708 ) | ( ~n1499 & n25712 ) | ( n25708 & n25712 ) ;
  assign n25714 = n25707 | n25713 ;
  assign n25715 = ( ~x11 & n24058 ) | ( ~x11 & n25090 ) | ( n24058 & n25090 ) ;
  assign n25716 = x77 & n18290 ;
  assign n25717 = x63 & x76 ;
  assign n25718 = ~n18290 & n25717 ;
  assign n25719 = n25716 | n25718 ;
  assign n25720 = n25715 & ~n25719 ;
  assign n25721 = n25715 & ~n25720 ;
  assign n25722 = n25715 | n25719 ;
  assign n25723 = ~n25721 & n25722 ;
  assign n25724 = n25714 | n25723 ;
  assign n25725 = n25714 & ~n25723 ;
  assign n25726 = ( ~n25714 & n25724 ) | ( ~n25714 & n25725 ) | ( n25724 & n25725 ) ;
  assign n25727 = n25097 | n25104 ;
  assign n25728 = ( n25097 & ~n25099 ) | ( n25097 & n25727 ) | ( ~n25099 & n25727 ) ;
  assign n25729 = n25726 & ~n25728 ;
  assign n25730 = ~n25726 & n25728 ;
  assign n25731 = n25729 | n25730 ;
  assign n25732 = x83 & n15552 ;
  assign n25733 = x82 & n15547 ;
  assign n25734 = x81 & ~n15546 ;
  assign n25735 = n16123 & n25734 ;
  assign n25736 = n25733 | n25735 ;
  assign n25737 = n25732 | n25736 ;
  assign n25738 = n15555 | n25732 ;
  assign n25739 = n25736 | n25738 ;
  assign n25740 = ( n2009 & n25737 ) | ( n2009 & n25739 ) | ( n25737 & n25739 ) ;
  assign n25741 = x59 & n25739 ;
  assign n25742 = x59 & n25732 ;
  assign n25743 = ( x59 & n25736 ) | ( x59 & n25742 ) | ( n25736 & n25742 ) ;
  assign n25744 = ( n2009 & n25741 ) | ( n2009 & n25743 ) | ( n25741 & n25743 ) ;
  assign n25745 = x59 & ~n25743 ;
  assign n25746 = x59 & ~n25739 ;
  assign n25747 = ( ~n2009 & n25745 ) | ( ~n2009 & n25746 ) | ( n25745 & n25746 ) ;
  assign n25748 = ( n25740 & ~n25744 ) | ( n25740 & n25747 ) | ( ~n25744 & n25747 ) ;
  assign n25749 = n25731 & n25748 ;
  assign n25750 = n25726 & ~n25748 ;
  assign n25751 = ( n25728 & n25748 ) | ( n25728 & ~n25750 ) | ( n25748 & ~n25750 ) ;
  assign n25752 = n25729 | n25751 ;
  assign n25753 = ~n25749 & n25752 ;
  assign n25754 = n25126 | n25133 ;
  assign n25755 = ( n25126 & ~n25130 ) | ( n25126 & n25754 ) | ( ~n25130 & n25754 ) ;
  assign n25756 = n25753 & ~n25755 ;
  assign n25757 = ~n25753 & n25755 ;
  assign n25758 = n25756 | n25757 ;
  assign n25759 = x86 & n14045 ;
  assign n25760 = x85 & n14040 ;
  assign n25761 = x84 & ~n14039 ;
  assign n25762 = n14552 & n25761 ;
  assign n25763 = n25760 | n25762 ;
  assign n25764 = n25759 | n25763 ;
  assign n25765 = n14048 | n25759 ;
  assign n25766 = n25763 | n25765 ;
  assign n25767 = ( n2606 & n25764 ) | ( n2606 & n25766 ) | ( n25764 & n25766 ) ;
  assign n25768 = x56 & n25766 ;
  assign n25769 = x56 & n25759 ;
  assign n25770 = ( x56 & n25763 ) | ( x56 & n25769 ) | ( n25763 & n25769 ) ;
  assign n25771 = ( n2606 & n25768 ) | ( n2606 & n25770 ) | ( n25768 & n25770 ) ;
  assign n25772 = x56 & ~n25770 ;
  assign n25773 = x56 & ~n25766 ;
  assign n25774 = ( ~n2606 & n25772 ) | ( ~n2606 & n25773 ) | ( n25772 & n25773 ) ;
  assign n25775 = ( n25767 & ~n25771 ) | ( n25767 & n25774 ) | ( ~n25771 & n25774 ) ;
  assign n25776 = n25758 & n25775 ;
  assign n25777 = n25757 | n25775 ;
  assign n25778 = n25756 | n25777 ;
  assign n25779 = ~n25776 & n25778 ;
  assign n25780 = ~n25154 & n25158 ;
  assign n25781 = ~n25154 & n25155 ;
  assign n25782 = ( ~n25159 & n25780 ) | ( ~n25159 & n25781 ) | ( n25780 & n25781 ) ;
  assign n25783 = n25779 & n25782 ;
  assign n25784 = n25779 | n25782 ;
  assign n25785 = ~n25783 & n25784 ;
  assign n25786 = x89 & n12574 ;
  assign n25787 = x88 & n12569 ;
  assign n25788 = x87 & ~n12568 ;
  assign n25789 = n13076 & n25788 ;
  assign n25790 = n25787 | n25789 ;
  assign n25791 = n25786 | n25790 ;
  assign n25792 = n12577 | n25786 ;
  assign n25793 = n25790 | n25792 ;
  assign n25794 = ( n3282 & n25791 ) | ( n3282 & n25793 ) | ( n25791 & n25793 ) ;
  assign n25795 = x53 & n25793 ;
  assign n25796 = x53 & n25786 ;
  assign n25797 = ( x53 & n25790 ) | ( x53 & n25796 ) | ( n25790 & n25796 ) ;
  assign n25798 = ( n3282 & n25795 ) | ( n3282 & n25797 ) | ( n25795 & n25797 ) ;
  assign n25799 = x53 & ~n25797 ;
  assign n25800 = x53 & ~n25793 ;
  assign n25801 = ( ~n3282 & n25799 ) | ( ~n3282 & n25800 ) | ( n25799 & n25800 ) ;
  assign n25802 = ( n25794 & ~n25798 ) | ( n25794 & n25801 ) | ( ~n25798 & n25801 ) ;
  assign n25803 = ~n25785 & n25802 ;
  assign n25804 = n25779 & ~n25802 ;
  assign n25805 = ( n25782 & ~n25802 ) | ( n25782 & n25804 ) | ( ~n25802 & n25804 ) ;
  assign n25806 = ~n25783 & n25805 ;
  assign n25807 = n25803 | n25806 ;
  assign n25808 = n25187 | n25191 ;
  assign n25809 = ( n25187 & n25190 ) | ( n25187 & n25808 ) | ( n25190 & n25808 ) ;
  assign n25810 = n25807 | n25809 ;
  assign n25811 = n25807 & n25809 ;
  assign n25812 = n25810 & ~n25811 ;
  assign n25813 = x92 & n11205 ;
  assign n25814 = x91 & n11200 ;
  assign n25815 = x90 & ~n11199 ;
  assign n25816 = n11679 & n25815 ;
  assign n25817 = n25814 | n25816 ;
  assign n25818 = n25813 | n25817 ;
  assign n25819 = n11208 | n25813 ;
  assign n25820 = n25817 | n25819 ;
  assign n25821 = ( n4040 & n25818 ) | ( n4040 & n25820 ) | ( n25818 & n25820 ) ;
  assign n25822 = x50 & n25820 ;
  assign n25823 = x50 & n25813 ;
  assign n25824 = ( x50 & n25817 ) | ( x50 & n25823 ) | ( n25817 & n25823 ) ;
  assign n25825 = ( n4040 & n25822 ) | ( n4040 & n25824 ) | ( n25822 & n25824 ) ;
  assign n25826 = x50 & ~n25824 ;
  assign n25827 = x50 & ~n25820 ;
  assign n25828 = ( ~n4040 & n25826 ) | ( ~n4040 & n25827 ) | ( n25826 & n25827 ) ;
  assign n25829 = ( n25821 & ~n25825 ) | ( n25821 & n25828 ) | ( ~n25825 & n25828 ) ;
  assign n25830 = n25812 | n25829 ;
  assign n25831 = n25812 & n25829 ;
  assign n25832 = n25830 & ~n25831 ;
  assign n25833 = x95 & n9933 ;
  assign n25834 = x94 & n9928 ;
  assign n25835 = x93 & ~n9927 ;
  assign n25836 = n10379 & n25835 ;
  assign n25837 = n25834 | n25836 ;
  assign n25838 = n25833 | n25837 ;
  assign n25839 = n9936 | n25833 ;
  assign n25840 = n25837 | n25839 ;
  assign n25841 = ( n4897 & n25838 ) | ( n4897 & n25840 ) | ( n25838 & n25840 ) ;
  assign n25842 = x47 & n25840 ;
  assign n25843 = x47 & n25833 ;
  assign n25844 = ( x47 & n25837 ) | ( x47 & n25843 ) | ( n25837 & n25843 ) ;
  assign n25845 = ( n4897 & n25842 ) | ( n4897 & n25844 ) | ( n25842 & n25844 ) ;
  assign n25846 = x47 & ~n25844 ;
  assign n25847 = x47 & ~n25840 ;
  assign n25848 = ( ~n4897 & n25846 ) | ( ~n4897 & n25847 ) | ( n25846 & n25847 ) ;
  assign n25849 = ( n25841 & ~n25845 ) | ( n25841 & n25848 ) | ( ~n25845 & n25848 ) ;
  assign n25852 = ( ~n25832 & n25849 ) | ( ~n25832 & n25851 ) | ( n25849 & n25851 ) ;
  assign n25853 = ( n25832 & ~n25849 ) | ( n25832 & n25852 ) | ( ~n25849 & n25852 ) ;
  assign n25854 = ( ~n25851 & n25852 ) | ( ~n25851 & n25853 ) | ( n25852 & n25853 ) ;
  assign n25855 = n25238 | n25239 ;
  assign n25856 = ( n25238 & n25242 ) | ( n25238 & n25855 ) | ( n25242 & n25855 ) ;
  assign n25857 = n25854 & n25856 ;
  assign n25858 = n25854 | n25856 ;
  assign n25859 = ~n25857 & n25858 ;
  assign n25860 = x98 & n8724 ;
  assign n25861 = x97 & n8719 ;
  assign n25862 = x96 & ~n8718 ;
  assign n25863 = n9149 & n25862 ;
  assign n25864 = n25861 | n25863 ;
  assign n25865 = n25860 | n25864 ;
  assign n25866 = n8727 | n25860 ;
  assign n25867 = n25864 | n25866 ;
  assign n25868 = ( ~n5850 & n25865 ) | ( ~n5850 & n25867 ) | ( n25865 & n25867 ) ;
  assign n25869 = n25865 & n25867 ;
  assign n25870 = ( n5834 & n25868 ) | ( n5834 & n25869 ) | ( n25868 & n25869 ) ;
  assign n25871 = x44 & n25867 ;
  assign n25872 = x44 & n25860 ;
  assign n25873 = ( x44 & n25864 ) | ( x44 & n25872 ) | ( n25864 & n25872 ) ;
  assign n25874 = ( ~n5850 & n25871 ) | ( ~n5850 & n25873 ) | ( n25871 & n25873 ) ;
  assign n25875 = n25871 & n25873 ;
  assign n25876 = ( n5834 & n25874 ) | ( n5834 & n25875 ) | ( n25874 & n25875 ) ;
  assign n25877 = x44 & ~n25873 ;
  assign n25878 = x44 & ~n25867 ;
  assign n25879 = ( n5850 & n25877 ) | ( n5850 & n25878 ) | ( n25877 & n25878 ) ;
  assign n25880 = n25877 | n25878 ;
  assign n25881 = ( ~n5834 & n25879 ) | ( ~n5834 & n25880 ) | ( n25879 & n25880 ) ;
  assign n25882 = ( n25870 & ~n25876 ) | ( n25870 & n25881 ) | ( ~n25876 & n25881 ) ;
  assign n25883 = n25859 & n25882 ;
  assign n25884 = n25859 | n25882 ;
  assign n25885 = ~n25883 & n25884 ;
  assign n25897 = n25885 & n25896 ;
  assign n25898 = n25896 & ~n25897 ;
  assign n25899 = x101 & n7566 ;
  assign n25900 = x100 & n7561 ;
  assign n25901 = x99 & ~n7560 ;
  assign n25902 = n7953 & n25901 ;
  assign n25903 = n25900 | n25902 ;
  assign n25904 = n25899 | n25903 ;
  assign n25905 = n7569 | n25899 ;
  assign n25906 = n25903 | n25905 ;
  assign n25907 = ( n6844 & n25904 ) | ( n6844 & n25906 ) | ( n25904 & n25906 ) ;
  assign n25908 = x41 & n25906 ;
  assign n25909 = x41 & n25899 ;
  assign n25910 = ( x41 & n25903 ) | ( x41 & n25909 ) | ( n25903 & n25909 ) ;
  assign n25911 = ( n6844 & n25908 ) | ( n6844 & n25910 ) | ( n25908 & n25910 ) ;
  assign n25912 = x41 & ~n25910 ;
  assign n25913 = x41 & ~n25906 ;
  assign n25914 = ( ~n6844 & n25912 ) | ( ~n6844 & n25913 ) | ( n25912 & n25913 ) ;
  assign n25915 = ( n25907 & ~n25911 ) | ( n25907 & n25914 ) | ( ~n25911 & n25914 ) ;
  assign n25916 = n25885 | n25915 ;
  assign n25917 = ( ~n25896 & n25915 ) | ( ~n25896 & n25916 ) | ( n25915 & n25916 ) ;
  assign n25918 = n25898 | n25917 ;
  assign n25919 = n25885 & n25915 ;
  assign n25920 = ~n25885 & n25915 ;
  assign n25921 = ( ~n25896 & n25915 ) | ( ~n25896 & n25920 ) | ( n25915 & n25920 ) ;
  assign n25922 = ( n25898 & n25919 ) | ( n25898 & n25921 ) | ( n25919 & n25921 ) ;
  assign n25923 = n25918 & ~n25922 ;
  assign n25924 = n25288 | n25295 ;
  assign n25925 = n25923 & n25924 ;
  assign n25926 = n25923 & ~n25925 ;
  assign n25927 = x104 & n6536 ;
  assign n25928 = x103 & n6531 ;
  assign n25929 = x102 & ~n6530 ;
  assign n25930 = n6871 & n25929 ;
  assign n25931 = n25928 | n25930 ;
  assign n25932 = n25927 | n25931 ;
  assign n25933 = n6539 | n25927 ;
  assign n25934 = n25931 | n25933 ;
  assign n25935 = ( n7911 & n25932 ) | ( n7911 & n25934 ) | ( n25932 & n25934 ) ;
  assign n25936 = x38 & n25934 ;
  assign n25937 = x38 & n25927 ;
  assign n25938 = ( x38 & n25931 ) | ( x38 & n25937 ) | ( n25931 & n25937 ) ;
  assign n25939 = ( n7911 & n25936 ) | ( n7911 & n25938 ) | ( n25936 & n25938 ) ;
  assign n25940 = x38 & ~n25938 ;
  assign n25941 = x38 & ~n25934 ;
  assign n25942 = ( ~n7911 & n25940 ) | ( ~n7911 & n25941 ) | ( n25940 & n25941 ) ;
  assign n25943 = ( n25935 & ~n25939 ) | ( n25935 & n25942 ) | ( ~n25939 & n25942 ) ;
  assign n25944 = ~n25923 & n25924 ;
  assign n25945 = n25943 & n25944 ;
  assign n25946 = ( n25926 & n25943 ) | ( n25926 & n25945 ) | ( n25943 & n25945 ) ;
  assign n25947 = n25943 | n25944 ;
  assign n25948 = n25926 | n25947 ;
  assign n25949 = ~n25946 & n25948 ;
  assign n25950 = ( n25296 & n25313 ) | ( n25296 & n25319 ) | ( n25313 & n25319 ) ;
  assign n25951 = ( n24785 & n25296 ) | ( n24785 & n25313 ) | ( n25296 & n25313 ) ;
  assign n25952 = ( n24786 & n25950 ) | ( n24786 & n25951 ) | ( n25950 & n25951 ) ;
  assign n25953 = n25949 | n25952 ;
  assign n25954 = n25949 & n25952 ;
  assign n25955 = n25953 & ~n25954 ;
  assign n25956 = x107 & n5554 ;
  assign n25957 = x106 & n5549 ;
  assign n25958 = x105 & ~n5548 ;
  assign n25959 = n5893 & n25958 ;
  assign n25960 = n25957 | n25959 ;
  assign n25961 = n25956 | n25960 ;
  assign n25962 = n5557 | n25956 ;
  assign n25963 = n25960 | n25962 ;
  assign n25964 = ( n9084 & n25961 ) | ( n9084 & n25963 ) | ( n25961 & n25963 ) ;
  assign n25965 = x35 & n25963 ;
  assign n25966 = x35 & n25956 ;
  assign n25967 = ( x35 & n25960 ) | ( x35 & n25966 ) | ( n25960 & n25966 ) ;
  assign n25968 = ( n9084 & n25965 ) | ( n9084 & n25967 ) | ( n25965 & n25967 ) ;
  assign n25969 = x35 & ~n25967 ;
  assign n25970 = x35 & ~n25963 ;
  assign n25971 = ( ~n9084 & n25969 ) | ( ~n9084 & n25970 ) | ( n25969 & n25970 ) ;
  assign n25972 = ( n25964 & ~n25968 ) | ( n25964 & n25971 ) | ( ~n25968 & n25971 ) ;
  assign n25973 = n25955 & ~n25972 ;
  assign n25974 = n25955 | n25972 ;
  assign n25975 = ( ~n25955 & n25973 ) | ( ~n25955 & n25974 ) | ( n25973 & n25974 ) ;
  assign n25976 = ~n25340 & n25690 ;
  assign n25977 = ( ~n25323 & n25690 ) | ( ~n25323 & n25976 ) | ( n25690 & n25976 ) ;
  assign n25978 = ~n25346 & n25977 ;
  assign n25979 = ( ~n25343 & n25977 ) | ( ~n25343 & n25978 ) | ( n25977 & n25978 ) ;
  assign n25980 = n25975 & ~n25979 ;
  assign n25981 = ~n25696 & n25980 ;
  assign n25982 = ~n25975 & n25979 ;
  assign n25983 = ( n25696 & ~n25975 ) | ( n25696 & n25982 ) | ( ~n25975 & n25982 ) ;
  assign n25984 = n25981 | n25983 ;
  assign n25985 = n25666 & ~n25667 ;
  assign n25986 = n25666 & ~n25668 ;
  assign n25987 = ( ~n25350 & n25985 ) | ( ~n25350 & n25986 ) | ( n25985 & n25986 ) ;
  assign n25988 = ~n25379 & n25987 ;
  assign n25989 = n25984 & n25988 ;
  assign n25990 = ( n25671 & n25984 ) | ( n25671 & n25989 ) | ( n25984 & n25989 ) ;
  assign n25991 = n25984 | n25988 ;
  assign n25992 = n25671 | n25991 ;
  assign n25993 = ~n25990 & n25992 ;
  assign n25994 = n25651 & ~n25993 ;
  assign n25995 = n25651 | n25993 ;
  assign n25996 = ( ~n25651 & n25994 ) | ( ~n25651 & n25995 ) | ( n25994 & n25995 ) ;
  assign n25997 = n25626 & ~n25628 ;
  assign n25998 = n25996 & n25997 ;
  assign n25999 = ( n25630 & n25996 ) | ( n25630 & n25998 ) | ( n25996 & n25998 ) ;
  assign n26000 = n25996 | n25997 ;
  assign n26001 = n25630 | n26000 ;
  assign n26002 = ~n25999 & n26001 ;
  assign n26003 = n25609 & n26002 ;
  assign n26004 = n25609 & ~n26003 ;
  assign n26005 = ~n25609 & n26002 ;
  assign n26006 = n26004 | n26005 ;
  assign n26007 = n25576 & ~n25578 ;
  assign n26008 = n26006 & n26007 ;
  assign n26009 = ( n25580 & n26006 ) | ( n25580 & n26008 ) | ( n26006 & n26008 ) ;
  assign n26010 = n26006 | n26007 ;
  assign n26011 = n25580 | n26010 ;
  assign n26012 = ~n26009 & n26011 ;
  assign n26013 = n25555 | n26012 ;
  assign n26014 = ( ~n25541 & n26012 ) | ( ~n25541 & n26013 ) | ( n26012 & n26013 ) ;
  assign n26015 = n25559 | n26014 ;
  assign n26016 = n25555 & n26012 ;
  assign n26017 = ~n25541 & n26016 ;
  assign n26018 = ( n25559 & n26012 ) | ( n25559 & n26017 ) | ( n26012 & n26017 ) ;
  assign n26019 = n26015 & ~n26018 ;
  assign n26020 = n25527 & n26019 ;
  assign n26021 = n25467 & n26019 ;
  assign n26022 = ( ~n25533 & n26020 ) | ( ~n25533 & n26021 ) | ( n26020 & n26021 ) ;
  assign n26023 = n25534 & ~n26022 ;
  assign n26024 = ~n25527 & n26019 ;
  assign n26025 = ~n25467 & n26019 ;
  assign n26026 = ( n25533 & n26024 ) | ( n25533 & n26025 ) | ( n26024 & n26025 ) ;
  assign n26027 = n26023 | n26026 ;
  assign n26028 = n25496 | n25522 ;
  assign n26029 = n25496 | n25519 ;
  assign n26030 = ( n22794 & n26028 ) | ( n22794 & n26029 ) | ( n26028 & n26029 ) ;
  assign n26031 = n26027 | n26030 ;
  assign n26032 = ~n26030 & n26031 ;
  assign n26033 = ( ~n26027 & n26031 ) | ( ~n26027 & n26032 ) | ( n26031 & n26032 ) ;
  assign n26034 = n25579 | n26009 ;
  assign n26035 = x127 & ~n956 ;
  assign n26036 = n1105 & n26035 ;
  assign n26037 = n965 & n19877 ;
  assign n26038 = n26036 | n26037 ;
  assign n26039 = n965 & n19880 ;
  assign n26040 = n26036 | n26039 ;
  assign n26041 = ( n18202 & n26038 ) | ( n18202 & n26040 ) | ( n26038 & n26040 ) ;
  assign n26042 = n26038 & n26040 ;
  assign n26043 = ( n18212 & n26041 ) | ( n18212 & n26042 ) | ( n26041 & n26042 ) ;
  assign n26044 = ( n18214 & n26041 ) | ( n18214 & n26042 ) | ( n26041 & n26042 ) ;
  assign n26045 = ( n14002 & n26043 ) | ( n14002 & n26044 ) | ( n26043 & n26044 ) ;
  assign n26046 = x14 & n26043 ;
  assign n26047 = x14 & n26044 ;
  assign n26048 = ( n14002 & n26046 ) | ( n14002 & n26047 ) | ( n26046 & n26047 ) ;
  assign n26049 = x14 & ~n26047 ;
  assign n26050 = x14 & ~n26046 ;
  assign n26051 = ( ~n14002 & n26049 ) | ( ~n14002 & n26050 ) | ( n26049 & n26050 ) ;
  assign n26052 = ( n26045 & ~n26048 ) | ( n26045 & n26051 ) | ( ~n26048 & n26051 ) ;
  assign n26053 = n25576 & n26052 ;
  assign n26054 = n25578 & n26053 ;
  assign n26055 = ( n26009 & n26052 ) | ( n26009 & n26054 ) | ( n26052 & n26054 ) ;
  assign n26056 = n26034 & ~n26055 ;
  assign n26057 = n25597 | n26002 ;
  assign n26058 = ( n25606 & n26002 ) | ( n25606 & n26057 ) | ( n26002 & n26057 ) ;
  assign n26059 = ( n25607 & n25609 ) | ( n25607 & n26058 ) | ( n25609 & n26058 ) ;
  assign n26061 = x125 & n1378 ;
  assign n26062 = x124 & ~n1377 ;
  assign n26063 = n1542 & n26062 ;
  assign n26064 = n26061 | n26063 ;
  assign n26060 = x126 & n1383 ;
  assign n26066 = n1386 | n26060 ;
  assign n26067 = n26064 | n26066 ;
  assign n26065 = n26060 | n26064 ;
  assign n26068 = n26065 & n26067 ;
  assign n26069 = ( n18220 & n26067 ) | ( n18220 & n26068 ) | ( n26067 & n26068 ) ;
  assign n26070 = x17 & n26068 ;
  assign n26071 = x17 & n26067 ;
  assign n26072 = ( n18220 & n26070 ) | ( n18220 & n26071 ) | ( n26070 & n26071 ) ;
  assign n26073 = x17 & ~n26068 ;
  assign n26074 = x17 & ~n26067 ;
  assign n26075 = ( ~n18220 & n26073 ) | ( ~n18220 & n26074 ) | ( n26073 & n26074 ) ;
  assign n26076 = ( n26069 & ~n26072 ) | ( n26069 & n26075 ) | ( ~n26072 & n26075 ) ;
  assign n26077 = n26058 & n26076 ;
  assign n26078 = n25607 & n26076 ;
  assign n26079 = ( n25609 & n26077 ) | ( n25609 & n26078 ) | ( n26077 & n26078 ) ;
  assign n26080 = n26059 & ~n26079 ;
  assign n26081 = x117 & n3085 ;
  assign n26082 = x116 & n3080 ;
  assign n26083 = x115 & ~n3079 ;
  assign n26084 = n3309 & n26083 ;
  assign n26085 = n26082 | n26084 ;
  assign n26086 = n26081 | n26085 ;
  assign n26087 = n3088 | n26081 ;
  assign n26088 = n26085 | n26087 ;
  assign n26089 = ( ~n13522 & n26086 ) | ( ~n13522 & n26088 ) | ( n26086 & n26088 ) ;
  assign n26090 = n26086 & n26088 ;
  assign n26091 = ( n13503 & n26089 ) | ( n13503 & n26090 ) | ( n26089 & n26090 ) ;
  assign n26092 = x26 & n26091 ;
  assign n26093 = x26 & ~n26091 ;
  assign n26094 = ( n26091 & ~n26092 ) | ( n26091 & n26093 ) | ( ~n26092 & n26093 ) ;
  assign n26095 = n25666 & n26094 ;
  assign n26096 = n25667 & n26094 ;
  assign n26097 = n25668 & n26094 ;
  assign n26098 = ( n25350 & n26096 ) | ( n25350 & n26097 ) | ( n26096 & n26097 ) ;
  assign n26099 = ( n25379 & n26095 ) | ( n25379 & n26098 ) | ( n26095 & n26098 ) ;
  assign n26100 = ( n25990 & n26094 ) | ( n25990 & n26099 ) | ( n26094 & n26099 ) ;
  assign n26101 = n25666 | n26094 ;
  assign n26102 = n25667 | n26094 ;
  assign n26103 = n25668 | n26094 ;
  assign n26104 = ( n25350 & n26102 ) | ( n25350 & n26103 ) | ( n26102 & n26103 ) ;
  assign n26105 = ( n25379 & n26101 ) | ( n25379 & n26104 ) | ( n26101 & n26104 ) ;
  assign n26106 = n25990 | n26105 ;
  assign n26107 = ~n26100 & n26106 ;
  assign n26109 = x113 & n3811 ;
  assign n26110 = x112 & ~n3810 ;
  assign n26111 = n4067 & n26110 ;
  assign n26112 = n26109 | n26111 ;
  assign n26108 = x114 & n3816 ;
  assign n26114 = n3819 | n26108 ;
  assign n26115 = n26112 | n26114 ;
  assign n26113 = n26108 | n26112 ;
  assign n26116 = n26113 & n26115 ;
  assign n26117 = ( ~n12095 & n26115 ) | ( ~n12095 & n26116 ) | ( n26115 & n26116 ) ;
  assign n26118 = n26115 & n26116 ;
  assign n26119 = ( n12079 & n26117 ) | ( n12079 & n26118 ) | ( n26117 & n26118 ) ;
  assign n26120 = x29 & n26119 ;
  assign n26121 = x29 & ~n26119 ;
  assign n26122 = ( n26119 & ~n26120 ) | ( n26119 & n26121 ) | ( ~n26120 & n26121 ) ;
  assign n26123 = n25975 & n25979 ;
  assign n26124 = ( n25696 & n25975 ) | ( n25696 & n26123 ) | ( n25975 & n26123 ) ;
  assign n26125 = n25695 & n26122 ;
  assign n26126 = ( n26122 & n26124 ) | ( n26122 & n26125 ) | ( n26124 & n26125 ) ;
  assign n26127 = n25695 | n26122 ;
  assign n26128 = n26124 | n26127 ;
  assign n26129 = ~n26126 & n26128 ;
  assign n26131 = x110 & n4626 ;
  assign n26132 = x109 & ~n4625 ;
  assign n26133 = n4943 & n26132 ;
  assign n26134 = n26131 | n26133 ;
  assign n26130 = x111 & n4631 ;
  assign n26136 = n4634 | n26130 ;
  assign n26137 = n26134 | n26136 ;
  assign n26135 = n26130 | n26134 ;
  assign n26138 = n26135 & n26137 ;
  assign n26139 = ( n10749 & n26137 ) | ( n10749 & n26138 ) | ( n26137 & n26138 ) ;
  assign n26140 = x32 & n26138 ;
  assign n26141 = x32 & n26137 ;
  assign n26142 = ( n10749 & n26140 ) | ( n10749 & n26141 ) | ( n26140 & n26141 ) ;
  assign n26143 = x32 & ~n26138 ;
  assign n26144 = x32 & ~n26137 ;
  assign n26145 = ( ~n10749 & n26143 ) | ( ~n10749 & n26144 ) | ( n26143 & n26144 ) ;
  assign n26146 = ( n26139 & ~n26142 ) | ( n26139 & n26145 ) | ( ~n26142 & n26145 ) ;
  assign n26147 = n25952 | n25972 ;
  assign n26148 = ( n25949 & n25972 ) | ( n25949 & n26147 ) | ( n25972 & n26147 ) ;
  assign n26149 = n26146 & n26148 ;
  assign n26150 = n25954 & n26146 ;
  assign n26151 = ( n25955 & n26149 ) | ( n25955 & n26150 ) | ( n26149 & n26150 ) ;
  assign n26152 = n26146 | n26148 ;
  assign n26153 = n25954 | n26146 ;
  assign n26154 = ( n25955 & n26152 ) | ( n25955 & n26153 ) | ( n26152 & n26153 ) ;
  assign n26155 = ~n26151 & n26154 ;
  assign n26279 = n25811 | n25829 ;
  assign n26280 = ( n25811 & n25812 ) | ( n25811 & n26279 ) | ( n25812 & n26279 ) ;
  assign n26156 = x78 & n18290 ;
  assign n26157 = x63 & x77 ;
  assign n26158 = ~n18290 & n26157 ;
  assign n26159 = n26156 | n26158 ;
  assign n26160 = ~n25719 & n26159 ;
  assign n26161 = n25719 & ~n26159 ;
  assign n26162 = n26160 | n26161 ;
  assign n26164 = x80 & n17141 ;
  assign n26165 = x79 & ~n17140 ;
  assign n26166 = n17724 & n26165 ;
  assign n26167 = n26164 | n26166 ;
  assign n26163 = x81 & n17146 ;
  assign n26169 = n17149 | n26163 ;
  assign n26170 = n26167 | n26169 ;
  assign n26168 = n26163 | n26167 ;
  assign n26171 = n26168 & n26170 ;
  assign n26172 = ( n1651 & n26170 ) | ( n1651 & n26171 ) | ( n26170 & n26171 ) ;
  assign n26173 = x62 & n26171 ;
  assign n26174 = x62 & n26170 ;
  assign n26175 = ( n1651 & n26173 ) | ( n1651 & n26174 ) | ( n26173 & n26174 ) ;
  assign n26176 = x62 & ~n26171 ;
  assign n26177 = x62 & ~n26170 ;
  assign n26178 = ( ~n1651 & n26176 ) | ( ~n1651 & n26177 ) | ( n26176 & n26177 ) ;
  assign n26179 = ( n26172 & ~n26175 ) | ( n26172 & n26178 ) | ( ~n26175 & n26178 ) ;
  assign n26180 = ~n26162 & n26179 ;
  assign n26181 = n26162 & ~n26179 ;
  assign n26182 = n26180 | n26181 ;
  assign n26183 = ( n25714 & n25715 ) | ( n25714 & ~n25719 ) | ( n25715 & ~n25719 ) ;
  assign n26184 = ~n26182 & n26183 ;
  assign n26185 = n26182 & ~n26183 ;
  assign n26186 = n26184 | n26185 ;
  assign n26187 = x84 & n15552 ;
  assign n26188 = x83 & n15547 ;
  assign n26189 = x82 & ~n15546 ;
  assign n26190 = n16123 & n26189 ;
  assign n26191 = n26188 | n26190 ;
  assign n26192 = n26187 | n26191 ;
  assign n26193 = n15555 | n26187 ;
  assign n26194 = n26191 | n26193 ;
  assign n26195 = ( n2194 & n26192 ) | ( n2194 & n26194 ) | ( n26192 & n26194 ) ;
  assign n26196 = x59 & n26194 ;
  assign n26197 = x59 & n26187 ;
  assign n26198 = ( x59 & n26191 ) | ( x59 & n26197 ) | ( n26191 & n26197 ) ;
  assign n26199 = ( n2194 & n26196 ) | ( n2194 & n26198 ) | ( n26196 & n26198 ) ;
  assign n26200 = x59 & ~n26198 ;
  assign n26201 = x59 & ~n26194 ;
  assign n26202 = ( ~n2194 & n26200 ) | ( ~n2194 & n26201 ) | ( n26200 & n26201 ) ;
  assign n26203 = ( n26195 & ~n26199 ) | ( n26195 & n26202 ) | ( ~n26199 & n26202 ) ;
  assign n26204 = n26186 | n26203 ;
  assign n26205 = n26186 & ~n26203 ;
  assign n26206 = ( ~n26186 & n26204 ) | ( ~n26186 & n26205 ) | ( n26204 & n26205 ) ;
  assign n26207 = ( n25730 & ~n25731 ) | ( n25730 & n25751 ) | ( ~n25731 & n25751 ) ;
  assign n26208 = n26206 & ~n26207 ;
  assign n26209 = ~n26206 & n26207 ;
  assign n26210 = n26208 | n26209 ;
  assign n26211 = x87 & n14045 ;
  assign n26212 = x86 & n14040 ;
  assign n26213 = x85 & ~n14039 ;
  assign n26214 = n14552 & n26213 ;
  assign n26215 = n26212 | n26214 ;
  assign n26216 = n26211 | n26215 ;
  assign n26217 = n14048 | n26211 ;
  assign n26218 = n26215 | n26217 ;
  assign n26219 = ( n2816 & n26216 ) | ( n2816 & n26218 ) | ( n26216 & n26218 ) ;
  assign n26220 = x56 & n26218 ;
  assign n26221 = x56 & n26211 ;
  assign n26222 = ( x56 & n26215 ) | ( x56 & n26221 ) | ( n26215 & n26221 ) ;
  assign n26223 = ( n2816 & n26220 ) | ( n2816 & n26222 ) | ( n26220 & n26222 ) ;
  assign n26224 = x56 & ~n26222 ;
  assign n26225 = x56 & ~n26218 ;
  assign n26226 = ( ~n2816 & n26224 ) | ( ~n2816 & n26225 ) | ( n26224 & n26225 ) ;
  assign n26227 = ( n26219 & ~n26223 ) | ( n26219 & n26226 ) | ( ~n26223 & n26226 ) ;
  assign n26228 = n26210 & ~n26227 ;
  assign n26229 = ~n26210 & n26227 ;
  assign n26230 = n26228 | n26229 ;
  assign n26231 = ( n25757 & ~n25758 ) | ( n25757 & n25777 ) | ( ~n25758 & n25777 ) ;
  assign n26232 = ~n26230 & n26231 ;
  assign n26233 = n26230 & ~n26231 ;
  assign n26234 = n26232 | n26233 ;
  assign n26235 = x90 & n12574 ;
  assign n26236 = x89 & n12569 ;
  assign n26237 = x88 & ~n12568 ;
  assign n26238 = n13076 & n26237 ;
  assign n26239 = n26236 | n26238 ;
  assign n26240 = n26235 | n26239 ;
  assign n26241 = n12577 | n26235 ;
  assign n26242 = n26239 | n26241 ;
  assign n26243 = ( n3519 & n26240 ) | ( n3519 & n26242 ) | ( n26240 & n26242 ) ;
  assign n26244 = x53 & n26242 ;
  assign n26245 = x53 & n26235 ;
  assign n26246 = ( x53 & n26239 ) | ( x53 & n26245 ) | ( n26239 & n26245 ) ;
  assign n26247 = ( n3519 & n26244 ) | ( n3519 & n26246 ) | ( n26244 & n26246 ) ;
  assign n26248 = x53 & ~n26246 ;
  assign n26249 = x53 & ~n26242 ;
  assign n26250 = ( ~n3519 & n26248 ) | ( ~n3519 & n26249 ) | ( n26248 & n26249 ) ;
  assign n26251 = ( n26243 & ~n26247 ) | ( n26243 & n26250 ) | ( ~n26247 & n26250 ) ;
  assign n26252 = ~n26234 & n26251 ;
  assign n26253 = n26234 & ~n26251 ;
  assign n26254 = n26252 | n26253 ;
  assign n26255 = ( n25784 & ~n25785 ) | ( n25784 & n25805 ) | ( ~n25785 & n25805 ) ;
  assign n26256 = n26254 | n26255 ;
  assign n26257 = n26254 & n26255 ;
  assign n26258 = n26256 & ~n26257 ;
  assign n26259 = x93 & n11205 ;
  assign n26260 = x92 & n11200 ;
  assign n26261 = x91 & ~n11199 ;
  assign n26262 = n11679 & n26261 ;
  assign n26263 = n26260 | n26262 ;
  assign n26264 = n26259 | n26263 ;
  assign n26265 = n11208 | n26259 ;
  assign n26266 = n26263 | n26265 ;
  assign n26267 = ( n4305 & n26264 ) | ( n4305 & n26266 ) | ( n26264 & n26266 ) ;
  assign n26268 = x50 & n26266 ;
  assign n26269 = x50 & n26259 ;
  assign n26270 = ( x50 & n26263 ) | ( x50 & n26269 ) | ( n26263 & n26269 ) ;
  assign n26271 = ( n4305 & n26268 ) | ( n4305 & n26270 ) | ( n26268 & n26270 ) ;
  assign n26272 = x50 & ~n26270 ;
  assign n26273 = x50 & ~n26266 ;
  assign n26274 = ( ~n4305 & n26272 ) | ( ~n4305 & n26273 ) | ( n26272 & n26273 ) ;
  assign n26275 = ( n26267 & ~n26271 ) | ( n26267 & n26274 ) | ( ~n26271 & n26274 ) ;
  assign n26276 = n26258 & ~n26275 ;
  assign n26277 = n26258 | n26275 ;
  assign n26278 = ( ~n26258 & n26276 ) | ( ~n26258 & n26277 ) | ( n26276 & n26277 ) ;
  assign n26281 = n26278 & n26280 ;
  assign n26282 = n26280 & ~n26281 ;
  assign n26283 = x96 & n9933 ;
  assign n26284 = x95 & n9928 ;
  assign n26285 = x94 & ~n9927 ;
  assign n26286 = n10379 & n26285 ;
  assign n26287 = n26284 | n26286 ;
  assign n26288 = n26283 | n26287 ;
  assign n26289 = n9936 | n26283 ;
  assign n26290 = n26287 | n26289 ;
  assign n26291 = ( n5202 & n26288 ) | ( n5202 & n26290 ) | ( n26288 & n26290 ) ;
  assign n26292 = x47 & n26290 ;
  assign n26293 = x47 & n26283 ;
  assign n26294 = ( x47 & n26287 ) | ( x47 & n26293 ) | ( n26287 & n26293 ) ;
  assign n26295 = ( n5202 & n26292 ) | ( n5202 & n26294 ) | ( n26292 & n26294 ) ;
  assign n26296 = x47 & ~n26294 ;
  assign n26297 = x47 & ~n26290 ;
  assign n26298 = ( ~n5202 & n26296 ) | ( ~n5202 & n26297 ) | ( n26296 & n26297 ) ;
  assign n26299 = ( n26291 & ~n26295 ) | ( n26291 & n26298 ) | ( ~n26295 & n26298 ) ;
  assign n26300 = n26278 & ~n26280 ;
  assign n26301 = ~n26299 & n26300 ;
  assign n26302 = ( n26282 & ~n26299 ) | ( n26282 & n26301 ) | ( ~n26299 & n26301 ) ;
  assign n26303 = n26299 & ~n26300 ;
  assign n26304 = ~n26282 & n26303 ;
  assign n26305 = n26302 | n26304 ;
  assign n26306 = n25832 & n25851 ;
  assign n26307 = n25851 & ~n26306 ;
  assign n26308 = n25832 & ~n26306 ;
  assign n26309 = n26307 | n26308 ;
  assign n26310 = n25849 | n26306 ;
  assign n26311 = ( n26306 & n26309 ) | ( n26306 & n26310 ) | ( n26309 & n26310 ) ;
  assign n26312 = n26305 | n26311 ;
  assign n26313 = n26305 & n26311 ;
  assign n26314 = n26312 & ~n26313 ;
  assign n26315 = x99 & n8724 ;
  assign n26316 = x98 & n8719 ;
  assign n26317 = x97 & ~n8718 ;
  assign n26318 = n9149 & n26317 ;
  assign n26319 = n26316 | n26318 ;
  assign n26320 = n26315 | n26319 ;
  assign n26321 = n8727 | n26315 ;
  assign n26322 = n26319 | n26321 ;
  assign n26323 = ( n6164 & n26320 ) | ( n6164 & n26322 ) | ( n26320 & n26322 ) ;
  assign n26324 = x44 & n26322 ;
  assign n26325 = x44 & n26315 ;
  assign n26326 = ( x44 & n26319 ) | ( x44 & n26325 ) | ( n26319 & n26325 ) ;
  assign n26327 = ( n6164 & n26324 ) | ( n6164 & n26326 ) | ( n26324 & n26326 ) ;
  assign n26328 = x44 & ~n26326 ;
  assign n26329 = x44 & ~n26322 ;
  assign n26330 = ( ~n6164 & n26328 ) | ( ~n6164 & n26329 ) | ( n26328 & n26329 ) ;
  assign n26331 = ( n26323 & ~n26327 ) | ( n26323 & n26330 ) | ( ~n26327 & n26330 ) ;
  assign n26332 = ~n26314 & n26331 ;
  assign n26333 = n26305 | n26331 ;
  assign n26334 = ( n26311 & n26331 ) | ( n26311 & n26333 ) | ( n26331 & n26333 ) ;
  assign n26335 = n26312 & ~n26334 ;
  assign n26336 = n26332 | n26335 ;
  assign n26337 = n25854 | n25882 ;
  assign n26338 = ( n25856 & n25882 ) | ( n25856 & n26337 ) | ( n25882 & n26337 ) ;
  assign n26339 = ( n25857 & n25859 ) | ( n25857 & n26338 ) | ( n25859 & n26338 ) ;
  assign n26340 = n26336 | n26339 ;
  assign n26341 = n26336 & n26339 ;
  assign n26342 = n26340 & ~n26341 ;
  assign n26343 = x102 & n7566 ;
  assign n26344 = x101 & n7561 ;
  assign n26345 = x100 & ~n7560 ;
  assign n26346 = n7953 & n26345 ;
  assign n26347 = n26344 | n26346 ;
  assign n26348 = n26343 | n26347 ;
  assign n26349 = n7569 | n26343 ;
  assign n26350 = n26347 | n26349 ;
  assign n26351 = ( n7178 & n26348 ) | ( n7178 & n26350 ) | ( n26348 & n26350 ) ;
  assign n26352 = x41 & n26350 ;
  assign n26353 = x41 & n26343 ;
  assign n26354 = ( x41 & n26347 ) | ( x41 & n26353 ) | ( n26347 & n26353 ) ;
  assign n26355 = ( n7178 & n26352 ) | ( n7178 & n26354 ) | ( n26352 & n26354 ) ;
  assign n26356 = x41 & ~n26354 ;
  assign n26357 = x41 & ~n26350 ;
  assign n26358 = ( ~n7178 & n26356 ) | ( ~n7178 & n26357 ) | ( n26356 & n26357 ) ;
  assign n26359 = ( n26351 & ~n26355 ) | ( n26351 & n26358 ) | ( ~n26355 & n26358 ) ;
  assign n26360 = n26342 | n26359 ;
  assign n26361 = n26342 & n26359 ;
  assign n26362 = n26360 & ~n26361 ;
  assign n26363 = n25897 | n25921 ;
  assign n26364 = n25897 | n25919 ;
  assign n26365 = ( n25898 & n26363 ) | ( n25898 & n26364 ) | ( n26363 & n26364 ) ;
  assign n26366 = n26362 & n26365 ;
  assign n26367 = n26362 | n26365 ;
  assign n26368 = ~n26366 & n26367 ;
  assign n26369 = x105 & n6536 ;
  assign n26370 = x104 & n6531 ;
  assign n26371 = x103 & ~n6530 ;
  assign n26372 = n6871 & n26371 ;
  assign n26373 = n26370 | n26372 ;
  assign n26374 = n26369 | n26373 ;
  assign n26375 = n6539 | n26369 ;
  assign n26376 = n26373 | n26375 ;
  assign n26377 = ( n8273 & n26374 ) | ( n8273 & n26376 ) | ( n26374 & n26376 ) ;
  assign n26378 = x38 & n26376 ;
  assign n26379 = x38 & n26369 ;
  assign n26380 = ( x38 & n26373 ) | ( x38 & n26379 ) | ( n26373 & n26379 ) ;
  assign n26381 = ( n8273 & n26378 ) | ( n8273 & n26380 ) | ( n26378 & n26380 ) ;
  assign n26382 = x38 & ~n26380 ;
  assign n26383 = x38 & ~n26376 ;
  assign n26384 = ( ~n8273 & n26382 ) | ( ~n8273 & n26383 ) | ( n26382 & n26383 ) ;
  assign n26385 = ( n26377 & ~n26381 ) | ( n26377 & n26384 ) | ( ~n26381 & n26384 ) ;
  assign n26386 = n26368 & n26385 ;
  assign n26387 = n26368 | n26385 ;
  assign n26388 = ~n26386 & n26387 ;
  assign n26389 = n25925 | n25946 ;
  assign n26390 = n26388 & n26389 ;
  assign n26391 = n26388 | n26389 ;
  assign n26392 = ~n26390 & n26391 ;
  assign n26393 = x108 & n5554 ;
  assign n26394 = x107 & n5549 ;
  assign n26395 = x106 & ~n5548 ;
  assign n26396 = n5893 & n26395 ;
  assign n26397 = n26394 | n26396 ;
  assign n26398 = n26393 | n26397 ;
  assign n26399 = n5557 | n26393 ;
  assign n26400 = n26397 | n26399 ;
  assign n26401 = ( n9479 & n26398 ) | ( n9479 & n26400 ) | ( n26398 & n26400 ) ;
  assign n26402 = x35 & n26400 ;
  assign n26403 = x35 & n26393 ;
  assign n26404 = ( x35 & n26397 ) | ( x35 & n26403 ) | ( n26397 & n26403 ) ;
  assign n26405 = ( n9479 & n26402 ) | ( n9479 & n26404 ) | ( n26402 & n26404 ) ;
  assign n26406 = x35 & ~n26404 ;
  assign n26407 = x35 & ~n26400 ;
  assign n26408 = ( ~n9479 & n26406 ) | ( ~n9479 & n26407 ) | ( n26406 & n26407 ) ;
  assign n26409 = ( n26401 & ~n26405 ) | ( n26401 & n26408 ) | ( ~n26405 & n26408 ) ;
  assign n26410 = n26392 & n26409 ;
  assign n26411 = n26392 & ~n26410 ;
  assign n26412 = ~n26392 & n26409 ;
  assign n26413 = n26411 | n26412 ;
  assign n26414 = ~n26155 & n26413 ;
  assign n26415 = n26155 & ~n26413 ;
  assign n26416 = n26414 | n26415 ;
  assign n26417 = n26129 & ~n26416 ;
  assign n26418 = n26129 | n26416 ;
  assign n26419 = ( ~n26129 & n26417 ) | ( ~n26129 & n26418 ) | ( n26417 & n26418 ) ;
  assign n26420 = n26107 & ~n26419 ;
  assign n26421 = n26107 | n26419 ;
  assign n26422 = ( ~n26107 & n26420 ) | ( ~n26107 & n26421 ) | ( n26420 & n26421 ) ;
  assign n26423 = x123 & n1859 ;
  assign n26424 = x122 & n1854 ;
  assign n26425 = x121 & ~n1853 ;
  assign n26426 = n2037 & n26425 ;
  assign n26427 = n26424 | n26426 ;
  assign n26428 = n26423 | n26427 ;
  assign n26429 = n1862 | n26423 ;
  assign n26430 = n26427 | n26429 ;
  assign n26431 = ( n16086 & n26428 ) | ( n16086 & n26430 ) | ( n26428 & n26430 ) ;
  assign n26432 = x20 & n26430 ;
  assign n26433 = x20 & n26423 ;
  assign n26434 = ( x20 & n26427 ) | ( x20 & n26433 ) | ( n26427 & n26433 ) ;
  assign n26435 = ( n16086 & n26432 ) | ( n16086 & n26434 ) | ( n26432 & n26434 ) ;
  assign n26436 = x20 & ~n26434 ;
  assign n26437 = x20 & ~n26430 ;
  assign n26438 = ( ~n16086 & n26436 ) | ( ~n16086 & n26437 ) | ( n26436 & n26437 ) ;
  assign n26439 = ( n26431 & ~n26435 ) | ( n26431 & n26438 ) | ( ~n26435 & n26438 ) ;
  assign n26440 = n25626 & n26439 ;
  assign n26441 = n25628 & n26440 ;
  assign n26442 = ( n25999 & n26439 ) | ( n25999 & n26441 ) | ( n26439 & n26441 ) ;
  assign n26443 = n25626 | n26439 ;
  assign n26444 = ( n25628 & n26439 ) | ( n25628 & n26443 ) | ( n26439 & n26443 ) ;
  assign n26445 = n25999 | n26444 ;
  assign n26446 = ~n26442 & n26445 ;
  assign n26447 = x120 & n2429 ;
  assign n26448 = x119 & n2424 ;
  assign n26449 = x118 & ~n2423 ;
  assign n26450 = n2631 & n26449 ;
  assign n26451 = n26448 | n26450 ;
  assign n26452 = n26447 | n26451 ;
  assign n26453 = n2432 | n26447 ;
  assign n26454 = n26451 | n26453 ;
  assign n26455 = ( n14991 & n26452 ) | ( n14991 & n26454 ) | ( n26452 & n26454 ) ;
  assign n26456 = x23 & n26454 ;
  assign n26457 = x23 & n26447 ;
  assign n26458 = ( x23 & n26451 ) | ( x23 & n26457 ) | ( n26451 & n26457 ) ;
  assign n26459 = ( n14991 & n26456 ) | ( n14991 & n26458 ) | ( n26456 & n26458 ) ;
  assign n26460 = x23 & ~n26458 ;
  assign n26461 = x23 & ~n26454 ;
  assign n26462 = ( ~n14991 & n26460 ) | ( ~n14991 & n26461 ) | ( n26460 & n26461 ) ;
  assign n26463 = ( n26455 & ~n26459 ) | ( n26455 & n26462 ) | ( ~n26459 & n26462 ) ;
  assign n26464 = n25649 | n25993 ;
  assign n26465 = ( n25649 & n25651 ) | ( n25649 & n26464 ) | ( n25651 & n26464 ) ;
  assign n26466 = n26463 | n26465 ;
  assign n26467 = n26463 & n26465 ;
  assign n26468 = n26466 & ~n26467 ;
  assign n26469 = ( n26422 & n26446 ) | ( n26422 & ~n26468 ) | ( n26446 & ~n26468 ) ;
  assign n26470 = ( ~n26446 & n26468 ) | ( ~n26446 & n26469 ) | ( n26468 & n26469 ) ;
  assign n26471 = ( ~n26422 & n26469 ) | ( ~n26422 & n26470 ) | ( n26469 & n26470 ) ;
  assign n26472 = ~n26058 & n26076 ;
  assign n26473 = ~n25607 & n26076 ;
  assign n26474 = ( ~n25609 & n26472 ) | ( ~n25609 & n26473 ) | ( n26472 & n26473 ) ;
  assign n26475 = n26471 | n26474 ;
  assign n26476 = n26080 | n26475 ;
  assign n26477 = n26471 & n26474 ;
  assign n26478 = ( n26080 & n26471 ) | ( n26080 & n26477 ) | ( n26471 & n26477 ) ;
  assign n26479 = n26476 & ~n26478 ;
  assign n26480 = ~n25576 & n26052 ;
  assign n26481 = ( ~n25578 & n26052 ) | ( ~n25578 & n26480 ) | ( n26052 & n26480 ) ;
  assign n26482 = n26479 & n26481 ;
  assign n26483 = ~n26009 & n26482 ;
  assign n26484 = ( n26056 & n26479 ) | ( n26056 & n26483 ) | ( n26479 & n26483 ) ;
  assign n26485 = n26479 | n26481 ;
  assign n26486 = ( ~n26009 & n26479 ) | ( ~n26009 & n26485 ) | ( n26479 & n26485 ) ;
  assign n26487 = n26056 | n26486 ;
  assign n26488 = ~n26484 & n26487 ;
  assign n26489 = n25558 & n26488 ;
  assign n26490 = ( n26018 & n26488 ) | ( n26018 & n26489 ) | ( n26488 & n26489 ) ;
  assign n26491 = n25558 | n26488 ;
  assign n26492 = n26018 | n26491 ;
  assign n26493 = ~n26490 & n26492 ;
  assign n26494 = n26022 | n26026 ;
  assign n26495 = n26023 | n26494 ;
  assign n26496 = ( n26022 & n26030 ) | ( n26022 & n26495 ) | ( n26030 & n26495 ) ;
  assign n26497 = n26493 | n26496 ;
  assign n26498 = n26493 & n26495 ;
  assign n26499 = n26022 & n26493 ;
  assign n26500 = ( n26030 & n26498 ) | ( n26030 & n26499 ) | ( n26498 & n26499 ) ;
  assign n26501 = n26497 & ~n26500 ;
  assign n26591 = n26209 | n26227 ;
  assign n26592 = ( n26209 & ~n26210 ) | ( n26209 & n26591 ) | ( ~n26210 & n26591 ) ;
  assign n26502 = x81 & n17141 ;
  assign n26503 = x80 & ~n17140 ;
  assign n26504 = n17724 & n26503 ;
  assign n26505 = n26502 | n26504 ;
  assign n26506 = x82 & n17146 ;
  assign n26507 = n17149 | n26506 ;
  assign n26508 = n26505 | n26507 ;
  assign n26509 = ~x62 & n26508 ;
  assign n26510 = ~x62 & n26506 ;
  assign n26511 = ( ~x62 & n26505 ) | ( ~x62 & n26510 ) | ( n26505 & n26510 ) ;
  assign n26512 = ( n1811 & n26509 ) | ( n1811 & n26511 ) | ( n26509 & n26511 ) ;
  assign n26513 = x62 & ~n26508 ;
  assign n26514 = x62 & x82 ;
  assign n26515 = n17146 & n26514 ;
  assign n26516 = x62 & ~n26515 ;
  assign n26517 = ~n26505 & n26516 ;
  assign n26518 = ( ~n1811 & n26513 ) | ( ~n1811 & n26517 ) | ( n26513 & n26517 ) ;
  assign n26519 = n26512 | n26518 ;
  assign n26520 = x79 & n18290 ;
  assign n26521 = x63 & x78 ;
  assign n26522 = ~n18290 & n26521 ;
  assign n26523 = n26520 | n26522 ;
  assign n26524 = ~x14 & n26523 ;
  assign n26525 = n26523 & ~n26524 ;
  assign n26526 = x14 | n26523 ;
  assign n26527 = n25719 & ~n26526 ;
  assign n26528 = ( n25719 & n26525 ) | ( n25719 & n26527 ) | ( n26525 & n26527 ) ;
  assign n26529 = ~n25719 & n26526 ;
  assign n26530 = ~n26525 & n26529 ;
  assign n26531 = n26528 | n26530 ;
  assign n26532 = n26519 & ~n26531 ;
  assign n26533 = ~n26519 & n26531 ;
  assign n26534 = n26532 | n26533 ;
  assign n26535 = ~n26160 & n26162 ;
  assign n26536 = ( n26160 & n26179 ) | ( n26160 & ~n26535 ) | ( n26179 & ~n26535 ) ;
  assign n26537 = n26534 & ~n26536 ;
  assign n26538 = ~n26534 & n26536 ;
  assign n26539 = n26537 | n26538 ;
  assign n26540 = x85 & n15552 ;
  assign n26541 = x84 & n15547 ;
  assign n26542 = x83 & ~n15546 ;
  assign n26543 = n16123 & n26542 ;
  assign n26544 = n26541 | n26543 ;
  assign n26545 = n26540 | n26544 ;
  assign n26546 = n15555 | n26540 ;
  assign n26547 = n26544 | n26546 ;
  assign n26548 = ( n2381 & n26545 ) | ( n2381 & n26547 ) | ( n26545 & n26547 ) ;
  assign n26549 = x59 & n26547 ;
  assign n26550 = x59 & n26540 ;
  assign n26551 = ( x59 & n26544 ) | ( x59 & n26550 ) | ( n26544 & n26550 ) ;
  assign n26552 = ( n2381 & n26549 ) | ( n2381 & n26551 ) | ( n26549 & n26551 ) ;
  assign n26553 = x59 & ~n26551 ;
  assign n26554 = x59 & ~n26547 ;
  assign n26555 = ( ~n2381 & n26553 ) | ( ~n2381 & n26554 ) | ( n26553 & n26554 ) ;
  assign n26556 = ( n26548 & ~n26552 ) | ( n26548 & n26555 ) | ( ~n26552 & n26555 ) ;
  assign n26557 = ~n26539 & n26556 ;
  assign n26558 = n26539 | n26557 ;
  assign n26560 = n26183 | n26203 ;
  assign n26561 = ( ~n26182 & n26203 ) | ( ~n26182 & n26560 ) | ( n26203 & n26560 ) ;
  assign n26562 = ( n26184 & ~n26186 ) | ( n26184 & n26561 ) | ( ~n26186 & n26561 ) ;
  assign n26559 = n26539 & n26556 ;
  assign n26563 = n26559 & n26562 ;
  assign n26564 = ( ~n26558 & n26562 ) | ( ~n26558 & n26563 ) | ( n26562 & n26563 ) ;
  assign n26565 = n26559 | n26562 ;
  assign n26566 = n26558 & ~n26565 ;
  assign n26567 = n26564 | n26566 ;
  assign n26568 = x88 & n14045 ;
  assign n26569 = x87 & n14040 ;
  assign n26570 = x86 & ~n14039 ;
  assign n26571 = n14552 & n26570 ;
  assign n26572 = n26569 | n26571 ;
  assign n26573 = n26568 | n26572 ;
  assign n26574 = n14048 | n26568 ;
  assign n26575 = n26572 | n26574 ;
  assign n26576 = ( ~n3039 & n26573 ) | ( ~n3039 & n26575 ) | ( n26573 & n26575 ) ;
  assign n26577 = n26573 & n26575 ;
  assign n26578 = ( n3023 & n26576 ) | ( n3023 & n26577 ) | ( n26576 & n26577 ) ;
  assign n26579 = x56 & n26575 ;
  assign n26580 = x56 & n26568 ;
  assign n26581 = ( x56 & n26572 ) | ( x56 & n26580 ) | ( n26572 & n26580 ) ;
  assign n26582 = ( ~n3039 & n26579 ) | ( ~n3039 & n26581 ) | ( n26579 & n26581 ) ;
  assign n26583 = n26579 & n26581 ;
  assign n26584 = ( n3023 & n26582 ) | ( n3023 & n26583 ) | ( n26582 & n26583 ) ;
  assign n26585 = x56 & ~n26581 ;
  assign n26586 = x56 & ~n26575 ;
  assign n26587 = ( n3039 & n26585 ) | ( n3039 & n26586 ) | ( n26585 & n26586 ) ;
  assign n26588 = n26585 | n26586 ;
  assign n26589 = ( ~n3023 & n26587 ) | ( ~n3023 & n26588 ) | ( n26587 & n26588 ) ;
  assign n26590 = ( n26578 & ~n26584 ) | ( n26578 & n26589 ) | ( ~n26584 & n26589 ) ;
  assign n26593 = ( n26567 & ~n26590 ) | ( n26567 & n26592 ) | ( ~n26590 & n26592 ) ;
  assign n26594 = ( ~n26567 & n26590 ) | ( ~n26567 & n26592 ) | ( n26590 & n26592 ) ;
  assign n26595 = ( ~n26592 & n26593 ) | ( ~n26592 & n26594 ) | ( n26593 & n26594 ) ;
  assign n26596 = x91 & n12574 ;
  assign n26597 = x90 & n12569 ;
  assign n26598 = x89 & ~n12568 ;
  assign n26599 = n13076 & n26598 ;
  assign n26600 = n26597 | n26599 ;
  assign n26601 = n26596 | n26600 ;
  assign n26602 = n12577 | n26596 ;
  assign n26603 = n26600 | n26602 ;
  assign n26604 = ( n3768 & n26601 ) | ( n3768 & n26603 ) | ( n26601 & n26603 ) ;
  assign n26605 = x53 & n26603 ;
  assign n26606 = x53 & n26596 ;
  assign n26607 = ( x53 & n26600 ) | ( x53 & n26606 ) | ( n26600 & n26606 ) ;
  assign n26608 = ( n3768 & n26605 ) | ( n3768 & n26607 ) | ( n26605 & n26607 ) ;
  assign n26609 = x53 & ~n26607 ;
  assign n26610 = x53 & ~n26603 ;
  assign n26611 = ( ~n3768 & n26609 ) | ( ~n3768 & n26610 ) | ( n26609 & n26610 ) ;
  assign n26612 = ( n26604 & ~n26608 ) | ( n26604 & n26611 ) | ( ~n26608 & n26611 ) ;
  assign n26613 = ~n26595 & n26612 ;
  assign n26614 = n26595 | n26613 ;
  assign n26616 = n26232 | n26251 ;
  assign n26617 = ( n26232 & ~n26234 ) | ( n26232 & n26616 ) | ( ~n26234 & n26616 ) ;
  assign n26615 = n26595 & n26612 ;
  assign n26618 = n26615 & n26617 ;
  assign n26619 = ( ~n26614 & n26617 ) | ( ~n26614 & n26618 ) | ( n26617 & n26618 ) ;
  assign n26620 = n26615 | n26617 ;
  assign n26621 = n26614 & ~n26620 ;
  assign n26622 = n26619 | n26621 ;
  assign n26623 = x94 & n11205 ;
  assign n26624 = x93 & n11200 ;
  assign n26625 = x92 & ~n11199 ;
  assign n26626 = n11679 & n26625 ;
  assign n26627 = n26624 | n26626 ;
  assign n26628 = n26623 | n26627 ;
  assign n26629 = n11208 | n26623 ;
  assign n26630 = n26627 | n26629 ;
  assign n26631 = ( n4583 & n26628 ) | ( n4583 & n26630 ) | ( n26628 & n26630 ) ;
  assign n26632 = x50 & n26630 ;
  assign n26633 = x50 & n26623 ;
  assign n26634 = ( x50 & n26627 ) | ( x50 & n26633 ) | ( n26627 & n26633 ) ;
  assign n26635 = ( n4583 & n26632 ) | ( n4583 & n26634 ) | ( n26632 & n26634 ) ;
  assign n26636 = x50 & ~n26634 ;
  assign n26637 = x50 & ~n26630 ;
  assign n26638 = ( ~n4583 & n26636 ) | ( ~n4583 & n26637 ) | ( n26636 & n26637 ) ;
  assign n26639 = ( n26631 & ~n26635 ) | ( n26631 & n26638 ) | ( ~n26635 & n26638 ) ;
  assign n26640 = ~n26622 & n26639 ;
  assign n26641 = n26622 | n26640 ;
  assign n26642 = n26254 & ~n26275 ;
  assign n26643 = ( n26255 & ~n26275 ) | ( n26255 & n26642 ) | ( ~n26275 & n26642 ) ;
  assign n26644 = ( n26256 & ~n26258 ) | ( n26256 & n26643 ) | ( ~n26258 & n26643 ) ;
  assign n26645 = n26622 & n26639 ;
  assign n26646 = ~n26644 & n26645 ;
  assign n26647 = ( n26641 & n26644 ) | ( n26641 & ~n26646 ) | ( n26644 & ~n26646 ) ;
  assign n26648 = n26644 & ~n26645 ;
  assign n26649 = n26641 & n26648 ;
  assign n26650 = n26647 & ~n26649 ;
  assign n26651 = x97 & n9933 ;
  assign n26652 = x96 & n9928 ;
  assign n26653 = x95 & ~n9927 ;
  assign n26654 = n10379 & n26653 ;
  assign n26655 = n26652 | n26654 ;
  assign n26656 = n26651 | n26655 ;
  assign n26657 = n9936 | n26651 ;
  assign n26658 = n26655 | n26657 ;
  assign n26659 = ( n5505 & n26656 ) | ( n5505 & n26658 ) | ( n26656 & n26658 ) ;
  assign n26660 = x47 & n26658 ;
  assign n26661 = x47 & n26651 ;
  assign n26662 = ( x47 & n26655 ) | ( x47 & n26661 ) | ( n26655 & n26661 ) ;
  assign n26663 = ( n5505 & n26660 ) | ( n5505 & n26662 ) | ( n26660 & n26662 ) ;
  assign n26664 = x47 & ~n26662 ;
  assign n26665 = x47 & ~n26658 ;
  assign n26666 = ( ~n5505 & n26664 ) | ( ~n5505 & n26665 ) | ( n26664 & n26665 ) ;
  assign n26667 = ( n26659 & ~n26663 ) | ( n26659 & n26666 ) | ( ~n26663 & n26666 ) ;
  assign n26668 = n26650 & n26667 ;
  assign n26669 = n26650 & ~n26668 ;
  assign n26670 = ~n26650 & n26667 ;
  assign n26671 = n26669 | n26670 ;
  assign n26672 = n26278 | n26299 ;
  assign n26673 = ( n26280 & n26299 ) | ( n26280 & n26672 ) | ( n26299 & n26672 ) ;
  assign n26674 = ( n26281 & n26300 ) | ( n26281 & n26673 ) | ( n26300 & n26673 ) ;
  assign n26675 = n26281 | n26673 ;
  assign n26676 = ( n26282 & n26674 ) | ( n26282 & n26675 ) | ( n26674 & n26675 ) ;
  assign n26677 = n26671 & n26676 ;
  assign n26678 = n26671 & ~n26677 ;
  assign n26679 = x100 & n8724 ;
  assign n26680 = x99 & n8719 ;
  assign n26681 = x98 & ~n8718 ;
  assign n26682 = n9149 & n26681 ;
  assign n26683 = n26680 | n26682 ;
  assign n26684 = n26679 | n26683 ;
  assign n26685 = n8727 | n26679 ;
  assign n26686 = n26683 | n26685 ;
  assign n26687 = ( n6483 & n26684 ) | ( n6483 & n26686 ) | ( n26684 & n26686 ) ;
  assign n26688 = x44 & n26686 ;
  assign n26689 = x44 & n26679 ;
  assign n26690 = ( x44 & n26683 ) | ( x44 & n26689 ) | ( n26683 & n26689 ) ;
  assign n26691 = ( n6483 & n26688 ) | ( n6483 & n26690 ) | ( n26688 & n26690 ) ;
  assign n26692 = x44 & ~n26690 ;
  assign n26693 = x44 & ~n26686 ;
  assign n26694 = ( ~n6483 & n26692 ) | ( ~n6483 & n26693 ) | ( n26692 & n26693 ) ;
  assign n26695 = ( n26687 & ~n26691 ) | ( n26687 & n26694 ) | ( ~n26691 & n26694 ) ;
  assign n26696 = n26676 & n26695 ;
  assign n26697 = ~n26676 & n26695 ;
  assign n26698 = ( ~n26671 & n26695 ) | ( ~n26671 & n26697 ) | ( n26695 & n26697 ) ;
  assign n26699 = ( n26678 & n26696 ) | ( n26678 & n26698 ) | ( n26696 & n26698 ) ;
  assign n26700 = n26676 | n26695 ;
  assign n26701 = n26676 & ~n26695 ;
  assign n26702 = n26671 & n26701 ;
  assign n26703 = ( n26678 & n26700 ) | ( n26678 & ~n26702 ) | ( n26700 & ~n26702 ) ;
  assign n26704 = ~n26699 & n26703 ;
  assign n26705 = ( n26313 & n26314 ) | ( n26313 & n26334 ) | ( n26314 & n26334 ) ;
  assign n26706 = n26704 | n26705 ;
  assign n26707 = n26704 & n26705 ;
  assign n26708 = n26706 & ~n26707 ;
  assign n26709 = x103 & n7566 ;
  assign n26710 = x102 & n7561 ;
  assign n26711 = x101 & ~n7560 ;
  assign n26712 = n7953 & n26711 ;
  assign n26713 = n26710 | n26712 ;
  assign n26714 = n26709 | n26713 ;
  assign n26715 = n7569 | n26709 ;
  assign n26716 = n26713 | n26715 ;
  assign n26717 = ( n7529 & n26714 ) | ( n7529 & n26716 ) | ( n26714 & n26716 ) ;
  assign n26718 = x41 & n26716 ;
  assign n26719 = x41 & n26709 ;
  assign n26720 = ( x41 & n26713 ) | ( x41 & n26719 ) | ( n26713 & n26719 ) ;
  assign n26721 = ( n7529 & n26718 ) | ( n7529 & n26720 ) | ( n26718 & n26720 ) ;
  assign n26722 = x41 & ~n26720 ;
  assign n26723 = x41 & ~n26716 ;
  assign n26724 = ( ~n7529 & n26722 ) | ( ~n7529 & n26723 ) | ( n26722 & n26723 ) ;
  assign n26725 = ( n26717 & ~n26721 ) | ( n26717 & n26724 ) | ( ~n26721 & n26724 ) ;
  assign n26726 = n26708 & n26725 ;
  assign n26727 = n26708 & ~n26726 ;
  assign n26728 = ~n26708 & n26725 ;
  assign n26729 = n26339 | n26359 ;
  assign n26730 = ( n26336 & n26359 ) | ( n26336 & n26729 ) | ( n26359 & n26729 ) ;
  assign n26731 = ( n26341 & n26342 ) | ( n26341 & n26730 ) | ( n26342 & n26730 ) ;
  assign n26732 = ~n26728 & n26731 ;
  assign n26733 = ~n26727 & n26732 ;
  assign n26734 = n26728 & ~n26731 ;
  assign n26735 = ( n26727 & ~n26731 ) | ( n26727 & n26734 ) | ( ~n26731 & n26734 ) ;
  assign n26736 = n26733 | n26735 ;
  assign n26737 = x106 & n6536 ;
  assign n26738 = x105 & n6531 ;
  assign n26739 = x104 & ~n6530 ;
  assign n26740 = n6871 & n26739 ;
  assign n26741 = n26738 | n26740 ;
  assign n26742 = n26737 | n26741 ;
  assign n26743 = n6539 | n26737 ;
  assign n26744 = n26741 | n26743 ;
  assign n26745 = ( n8656 & n26742 ) | ( n8656 & n26744 ) | ( n26742 & n26744 ) ;
  assign n26746 = x38 & n26744 ;
  assign n26747 = x38 & n26737 ;
  assign n26748 = ( x38 & n26741 ) | ( x38 & n26747 ) | ( n26741 & n26747 ) ;
  assign n26749 = ( n8656 & n26746 ) | ( n8656 & n26748 ) | ( n26746 & n26748 ) ;
  assign n26750 = x38 & ~n26748 ;
  assign n26751 = x38 & ~n26744 ;
  assign n26752 = ( ~n8656 & n26750 ) | ( ~n8656 & n26751 ) | ( n26750 & n26751 ) ;
  assign n26753 = ( n26745 & ~n26749 ) | ( n26745 & n26752 ) | ( ~n26749 & n26752 ) ;
  assign n26754 = n26736 & n26753 ;
  assign n26755 = n26736 | n26753 ;
  assign n26756 = ~n26754 & n26755 ;
  assign n26757 = n26366 | n26385 ;
  assign n26758 = ( n26366 & n26368 ) | ( n26366 & n26757 ) | ( n26368 & n26757 ) ;
  assign n26759 = n26756 | n26758 ;
  assign n26760 = n26756 & n26758 ;
  assign n26761 = n26759 & ~n26760 ;
  assign n26762 = x109 & n5554 ;
  assign n26763 = x108 & n5549 ;
  assign n26764 = x107 & ~n5548 ;
  assign n26765 = n5893 & n26764 ;
  assign n26766 = n26763 | n26765 ;
  assign n26767 = n26762 | n26766 ;
  assign n26768 = n5557 | n26762 ;
  assign n26769 = n26766 | n26768 ;
  assign n26770 = ( n9878 & n26767 ) | ( n9878 & n26769 ) | ( n26767 & n26769 ) ;
  assign n26771 = x35 & n26769 ;
  assign n26772 = x35 & n26762 ;
  assign n26773 = ( x35 & n26766 ) | ( x35 & n26772 ) | ( n26766 & n26772 ) ;
  assign n26774 = ( n9878 & n26771 ) | ( n9878 & n26773 ) | ( n26771 & n26773 ) ;
  assign n26775 = x35 & ~n26773 ;
  assign n26776 = x35 & ~n26769 ;
  assign n26777 = ( ~n9878 & n26775 ) | ( ~n9878 & n26776 ) | ( n26775 & n26776 ) ;
  assign n26778 = ( n26770 & ~n26774 ) | ( n26770 & n26777 ) | ( ~n26774 & n26777 ) ;
  assign n26779 = n26761 & n26778 ;
  assign n26780 = n26761 & ~n26779 ;
  assign n26781 = ~n26761 & n26778 ;
  assign n26782 = n26780 | n26781 ;
  assign n26783 = n26388 | n26409 ;
  assign n26784 = ( n26389 & n26409 ) | ( n26389 & n26783 ) | ( n26409 & n26783 ) ;
  assign n26785 = ( n26390 & n26392 ) | ( n26390 & n26784 ) | ( n26392 & n26784 ) ;
  assign n26786 = n26782 | n26785 ;
  assign n26787 = n26782 & n26785 ;
  assign n26788 = n26786 & ~n26787 ;
  assign n26789 = n26151 | n26155 ;
  assign n26790 = ( n26151 & n26413 ) | ( n26151 & n26789 ) | ( n26413 & n26789 ) ;
  assign n26791 = x112 & n4631 ;
  assign n26792 = x111 & n4626 ;
  assign n26793 = x110 & ~n4625 ;
  assign n26794 = n4943 & n26793 ;
  assign n26795 = n26792 | n26794 ;
  assign n26796 = n26791 | n26795 ;
  assign n26797 = n4634 | n26791 ;
  assign n26798 = n26795 | n26797 ;
  assign n26799 = ( n11172 & n26796 ) | ( n11172 & n26798 ) | ( n26796 & n26798 ) ;
  assign n26800 = x32 & n26798 ;
  assign n26801 = x32 & n26791 ;
  assign n26802 = ( x32 & n26795 ) | ( x32 & n26801 ) | ( n26795 & n26801 ) ;
  assign n26803 = ( n11172 & n26800 ) | ( n11172 & n26802 ) | ( n26800 & n26802 ) ;
  assign n26804 = x32 & ~n26802 ;
  assign n26805 = x32 & ~n26798 ;
  assign n26806 = ( ~n11172 & n26804 ) | ( ~n11172 & n26805 ) | ( n26804 & n26805 ) ;
  assign n26807 = ( n26799 & ~n26803 ) | ( n26799 & n26806 ) | ( ~n26803 & n26806 ) ;
  assign n26808 = n26151 & n26807 ;
  assign n26809 = ( n26155 & n26807 ) | ( n26155 & n26808 ) | ( n26807 & n26808 ) ;
  assign n26810 = n26807 & n26808 ;
  assign n26811 = ( n26413 & n26809 ) | ( n26413 & n26810 ) | ( n26809 & n26810 ) ;
  assign n26812 = n26790 & ~n26811 ;
  assign n26813 = ~n26151 & n26807 ;
  assign n26814 = ~n26155 & n26813 ;
  assign n26815 = ( ~n26413 & n26813 ) | ( ~n26413 & n26814 ) | ( n26813 & n26814 ) ;
  assign n26816 = n26788 & n26815 ;
  assign n26817 = ( n26788 & n26812 ) | ( n26788 & n26816 ) | ( n26812 & n26816 ) ;
  assign n26818 = n26788 | n26815 ;
  assign n26819 = n26812 | n26818 ;
  assign n26820 = ~n26817 & n26819 ;
  assign n26821 = x115 & n3816 ;
  assign n26822 = x114 & n3811 ;
  assign n26823 = x113 & ~n3810 ;
  assign n26824 = n4067 & n26823 ;
  assign n26825 = n26822 | n26824 ;
  assign n26826 = n26821 | n26825 ;
  assign n26827 = n3819 | n26821 ;
  assign n26828 = n26825 | n26827 ;
  assign n26829 = ( ~n12550 & n26826 ) | ( ~n12550 & n26828 ) | ( n26826 & n26828 ) ;
  assign n26830 = n26826 & n26828 ;
  assign n26831 = ( n12532 & n26829 ) | ( n12532 & n26830 ) | ( n26829 & n26830 ) ;
  assign n26832 = x29 & n26831 ;
  assign n26833 = x29 & ~n26831 ;
  assign n26834 = ( n26831 & ~n26832 ) | ( n26831 & n26833 ) | ( ~n26832 & n26833 ) ;
  assign n26835 = n26126 | n26416 ;
  assign n26836 = ( n26126 & n26129 ) | ( n26126 & n26835 ) | ( n26129 & n26835 ) ;
  assign n26837 = n26834 | n26836 ;
  assign n26838 = n26834 & n26836 ;
  assign n26839 = n26837 & ~n26838 ;
  assign n26840 = n26820 & n26839 ;
  assign n26841 = n26839 & ~n26840 ;
  assign n26842 = ( n26820 & ~n26840 ) | ( n26820 & n26841 ) | ( ~n26840 & n26841 ) ;
  assign n26843 = x121 & n2429 ;
  assign n26844 = x120 & n2424 ;
  assign n26845 = x119 & ~n2423 ;
  assign n26846 = n2631 & n26845 ;
  assign n26847 = n26844 | n26846 ;
  assign n26848 = n26843 | n26847 ;
  assign n26849 = n2432 | n26843 ;
  assign n26850 = n26847 | n26849 ;
  assign n26851 = ( n15501 & n26848 ) | ( n15501 & n26850 ) | ( n26848 & n26850 ) ;
  assign n26852 = x23 & n26850 ;
  assign n26853 = x23 & n26843 ;
  assign n26854 = ( x23 & n26847 ) | ( x23 & n26853 ) | ( n26847 & n26853 ) ;
  assign n26855 = ( n15501 & n26852 ) | ( n15501 & n26854 ) | ( n26852 & n26854 ) ;
  assign n26856 = x23 & ~n26854 ;
  assign n26857 = x23 & ~n26850 ;
  assign n26858 = ( ~n15501 & n26856 ) | ( ~n15501 & n26857 ) | ( n26856 & n26857 ) ;
  assign n26859 = ( n26851 & ~n26855 ) | ( n26851 & n26858 ) | ( ~n26855 & n26858 ) ;
  assign n26860 = n26422 | n26467 ;
  assign n26861 = ( n26467 & n26468 ) | ( n26467 & n26860 ) | ( n26468 & n26860 ) ;
  assign n26862 = ~n26859 & n26861 ;
  assign n26863 = n26859 & ~n26861 ;
  assign n26864 = n26862 | n26863 ;
  assign n26865 = x118 & n3085 ;
  assign n26866 = x117 & n3080 ;
  assign n26867 = x116 & ~n3079 ;
  assign n26868 = n3309 & n26867 ;
  assign n26869 = n26866 | n26868 ;
  assign n26870 = n26865 | n26869 ;
  assign n26871 = n3088 | n26865 ;
  assign n26872 = n26869 | n26871 ;
  assign n26873 = ( ~n14002 & n26870 ) | ( ~n14002 & n26872 ) | ( n26870 & n26872 ) ;
  assign n26874 = n26870 & n26872 ;
  assign n26875 = ( n13981 & n26873 ) | ( n13981 & n26874 ) | ( n26873 & n26874 ) ;
  assign n26876 = x26 & n26875 ;
  assign n26877 = x26 & ~n26875 ;
  assign n26878 = ( n26875 & ~n26876 ) | ( n26875 & n26877 ) | ( ~n26876 & n26877 ) ;
  assign n26879 = n26100 | n26419 ;
  assign n26880 = ( n26100 & n26107 ) | ( n26100 & n26879 ) | ( n26107 & n26879 ) ;
  assign n26881 = n26878 | n26880 ;
  assign n26882 = n26878 & n26880 ;
  assign n26883 = n26881 & ~n26882 ;
  assign n26884 = ( n26842 & n26864 ) | ( n26842 & ~n26883 ) | ( n26864 & ~n26883 ) ;
  assign n26885 = ( ~n26864 & n26883 ) | ( ~n26864 & n26884 ) | ( n26883 & n26884 ) ;
  assign n26886 = ( ~n26842 & n26884 ) | ( ~n26842 & n26885 ) | ( n26884 & n26885 ) ;
  assign n26887 = x124 & n1859 ;
  assign n26888 = x123 & n1854 ;
  assign n26889 = x122 & ~n1853 ;
  assign n26890 = n2037 & n26889 ;
  assign n26891 = n26888 | n26890 ;
  assign n26892 = n26887 | n26891 ;
  assign n26893 = n1862 | n26887 ;
  assign n26894 = n26891 | n26893 ;
  assign n26895 = ( n17084 & n26892 ) | ( n17084 & n26894 ) | ( n26892 & n26894 ) ;
  assign n26896 = x20 & n26894 ;
  assign n26897 = x20 & n26887 ;
  assign n26898 = ( x20 & n26891 ) | ( x20 & n26897 ) | ( n26891 & n26897 ) ;
  assign n26899 = ( n17084 & n26896 ) | ( n17084 & n26898 ) | ( n26896 & n26898 ) ;
  assign n26900 = x20 & ~n26898 ;
  assign n26901 = x20 & ~n26894 ;
  assign n26902 = ( ~n17084 & n26900 ) | ( ~n17084 & n26901 ) | ( n26900 & n26901 ) ;
  assign n26903 = ( n26895 & ~n26899 ) | ( n26895 & n26902 ) | ( ~n26899 & n26902 ) ;
  assign n26904 = n26422 & n26468 ;
  assign n26905 = n26422 | n26468 ;
  assign n26906 = ~n26904 & n26905 ;
  assign n26907 = n26442 | n26906 ;
  assign n26908 = ( n26442 & n26446 ) | ( n26442 & n26907 ) | ( n26446 & n26907 ) ;
  assign n26909 = n26903 | n26908 ;
  assign n26910 = n26903 & n26908 ;
  assign n26911 = n26909 & ~n26910 ;
  assign n26912 = n26080 | n26474 ;
  assign n26913 = n26079 | n26471 ;
  assign n26914 = x127 & n1383 ;
  assign n26915 = x126 & n1378 ;
  assign n26916 = x125 & ~n1377 ;
  assign n26917 = n1542 & n26916 ;
  assign n26918 = n26915 | n26917 ;
  assign n26919 = n26914 | n26918 ;
  assign n26920 = n1386 | n26914 ;
  assign n26921 = n26918 | n26920 ;
  assign n26922 = ( n18763 & n26919 ) | ( n18763 & n26921 ) | ( n26919 & n26921 ) ;
  assign n26923 = x17 & n26921 ;
  assign n26924 = x17 & n26914 ;
  assign n26925 = ( x17 & n26918 ) | ( x17 & n26924 ) | ( n26918 & n26924 ) ;
  assign n26926 = ( n18763 & n26923 ) | ( n18763 & n26925 ) | ( n26923 & n26925 ) ;
  assign n26927 = x17 & ~n26925 ;
  assign n26928 = x17 & ~n26921 ;
  assign n26929 = ( ~n18763 & n26927 ) | ( ~n18763 & n26928 ) | ( n26927 & n26928 ) ;
  assign n26930 = ( n26922 & ~n26926 ) | ( n26922 & n26929 ) | ( ~n26926 & n26929 ) ;
  assign n26931 = n26913 & n26930 ;
  assign n26932 = n26079 & n26930 ;
  assign n26933 = ( n26912 & n26931 ) | ( n26912 & n26932 ) | ( n26931 & n26932 ) ;
  assign n26934 = n26913 | n26930 ;
  assign n26935 = n26079 | n26930 ;
  assign n26936 = ( n26912 & n26934 ) | ( n26912 & n26935 ) | ( n26934 & n26935 ) ;
  assign n26937 = ~n26933 & n26936 ;
  assign n26938 = ( n26886 & ~n26911 ) | ( n26886 & n26937 ) | ( ~n26911 & n26937 ) ;
  assign n26939 = ( n26911 & ~n26937 ) | ( n26911 & n26938 ) | ( ~n26937 & n26938 ) ;
  assign n26940 = ( ~n26886 & n26938 ) | ( ~n26886 & n26939 ) | ( n26938 & n26939 ) ;
  assign n26941 = n26055 | n26483 ;
  assign n26942 = n26054 | n26479 ;
  assign n26943 = n26052 | n26479 ;
  assign n26944 = ( n26009 & n26942 ) | ( n26009 & n26943 ) | ( n26942 & n26943 ) ;
  assign n26945 = ( n26056 & n26941 ) | ( n26056 & n26944 ) | ( n26941 & n26944 ) ;
  assign n26946 = n26940 | n26945 ;
  assign n26947 = n26940 & n26945 ;
  assign n26948 = n26946 & ~n26947 ;
  assign n26949 = n26490 | n26493 ;
  assign n26950 = ( n26490 & n26495 ) | ( n26490 & n26949 ) | ( n26495 & n26949 ) ;
  assign n26951 = ( n26022 & n26490 ) | ( n26022 & n26949 ) | ( n26490 & n26949 ) ;
  assign n26952 = ( n26030 & n26950 ) | ( n26030 & n26951 ) | ( n26950 & n26951 ) ;
  assign n26953 = n26948 | n26952 ;
  assign n26954 = n26948 & n26951 ;
  assign n26955 = n26490 & n26948 ;
  assign n26956 = ( n26493 & n26948 ) | ( n26493 & n26955 ) | ( n26948 & n26955 ) ;
  assign n26957 = ( n26495 & n26955 ) | ( n26495 & n26956 ) | ( n26955 & n26956 ) ;
  assign n26958 = ( n26030 & n26954 ) | ( n26030 & n26957 ) | ( n26954 & n26957 ) ;
  assign n26959 = n26953 & ~n26958 ;
  assign n26960 = x113 & n4631 ;
  assign n26961 = x112 & n4626 ;
  assign n26962 = x111 & ~n4625 ;
  assign n26963 = n4943 & n26962 ;
  assign n26964 = n26961 | n26963 ;
  assign n26965 = n26960 | n26964 ;
  assign n26966 = n4634 | n26960 ;
  assign n26967 = n26964 | n26966 ;
  assign n26968 = ( ~n11642 & n26965 ) | ( ~n11642 & n26967 ) | ( n26965 & n26967 ) ;
  assign n26969 = n26965 & n26967 ;
  assign n26970 = ( n11626 & n26968 ) | ( n11626 & n26969 ) | ( n26968 & n26969 ) ;
  assign n26971 = x32 & n26970 ;
  assign n26972 = x32 & ~n26970 ;
  assign n26973 = ( n26970 & ~n26971 ) | ( n26970 & n26972 ) | ( ~n26971 & n26972 ) ;
  assign n26974 = n26779 | n26785 ;
  assign n26975 = ( n26779 & n26782 ) | ( n26779 & n26974 ) | ( n26782 & n26974 ) ;
  assign n26976 = n26973 | n26975 ;
  assign n26977 = n26973 & n26975 ;
  assign n26978 = n26976 & ~n26977 ;
  assign n26979 = n26811 | n26817 ;
  assign n26980 = x116 & n3816 ;
  assign n26981 = x115 & n3811 ;
  assign n26982 = x114 & ~n3810 ;
  assign n26983 = n4067 & n26982 ;
  assign n26984 = n26981 | n26983 ;
  assign n26985 = n26980 | n26984 ;
  assign n26986 = n3819 | n26980 ;
  assign n26987 = n26984 | n26986 ;
  assign n26988 = ( ~n13040 & n26985 ) | ( ~n13040 & n26987 ) | ( n26985 & n26987 ) ;
  assign n26989 = n26985 & n26987 ;
  assign n26990 = ( n13022 & n26988 ) | ( n13022 & n26989 ) | ( n26988 & n26989 ) ;
  assign n26991 = x29 & n26990 ;
  assign n26992 = x29 & ~n26990 ;
  assign n26993 = ( n26990 & ~n26991 ) | ( n26990 & n26992 ) | ( ~n26991 & n26992 ) ;
  assign n26994 = n26807 & n26993 ;
  assign n26995 = n26151 & n26994 ;
  assign n26996 = ( n26155 & n26994 ) | ( n26155 & n26995 ) | ( n26994 & n26995 ) ;
  assign n26997 = n26994 & n26995 ;
  assign n26998 = ( n26413 & n26996 ) | ( n26413 & n26997 ) | ( n26996 & n26997 ) ;
  assign n26999 = ( n26817 & n26993 ) | ( n26817 & n26998 ) | ( n26993 & n26998 ) ;
  assign n27000 = n26979 & ~n26999 ;
  assign n27004 = ( n26708 & n26725 ) | ( n26708 & n26731 ) | ( n26725 & n26731 ) ;
  assign n27171 = n26668 | n26676 ;
  assign n27172 = ( n26668 & n26671 ) | ( n26668 & n27171 ) | ( n26671 & n27171 ) ;
  assign n27005 = n26567 & ~n26590 ;
  assign n27006 = n26592 & ~n27005 ;
  assign n27007 = ~n26567 & n26590 ;
  assign n27008 = n27006 | n27007 ;
  assign n27009 = n26557 | n26564 ;
  assign n27010 = x80 & n18290 ;
  assign n27011 = x63 & x79 ;
  assign n27012 = ~n18290 & n27011 ;
  assign n27013 = n27010 | n27012 ;
  assign n27014 = n26524 & ~n27013 ;
  assign n27015 = ( n26528 & ~n27013 ) | ( n26528 & n27014 ) | ( ~n27013 & n27014 ) ;
  assign n27016 = ~n26524 & n27013 ;
  assign n27017 = ~n26528 & n27016 ;
  assign n27018 = n27015 | n27017 ;
  assign n27020 = x82 & n17141 ;
  assign n27021 = x81 & ~n17140 ;
  assign n27022 = n17724 & n27021 ;
  assign n27023 = n27020 | n27022 ;
  assign n27019 = x83 & n17146 ;
  assign n27025 = n17149 | n27019 ;
  assign n27026 = n27023 | n27025 ;
  assign n27024 = n27019 | n27023 ;
  assign n27027 = n27024 & n27026 ;
  assign n27028 = ( n2009 & n27026 ) | ( n2009 & n27027 ) | ( n27026 & n27027 ) ;
  assign n27029 = x62 & n27027 ;
  assign n27030 = x62 & n27026 ;
  assign n27031 = ( n2009 & n27029 ) | ( n2009 & n27030 ) | ( n27029 & n27030 ) ;
  assign n27032 = x62 & ~n27027 ;
  assign n27033 = x62 & ~n27026 ;
  assign n27034 = ( ~n2009 & n27032 ) | ( ~n2009 & n27033 ) | ( n27032 & n27033 ) ;
  assign n27035 = ( n27028 & ~n27031 ) | ( n27028 & n27034 ) | ( ~n27031 & n27034 ) ;
  assign n27036 = ~n27018 & n27035 ;
  assign n27037 = n27018 & ~n27035 ;
  assign n27038 = n27036 | n27037 ;
  assign n27039 = n26532 | n26536 ;
  assign n27040 = ( n26532 & ~n26534 ) | ( n26532 & n27039 ) | ( ~n26534 & n27039 ) ;
  assign n27041 = ~n27038 & n27040 ;
  assign n27042 = n27038 & ~n27040 ;
  assign n27043 = n27041 | n27042 ;
  assign n27044 = x86 & n15552 ;
  assign n27045 = x85 & n15547 ;
  assign n27046 = x84 & ~n15546 ;
  assign n27047 = n16123 & n27046 ;
  assign n27048 = n27045 | n27047 ;
  assign n27049 = n27044 | n27048 ;
  assign n27050 = n15555 | n27044 ;
  assign n27051 = n27048 | n27050 ;
  assign n27052 = ( n2606 & n27049 ) | ( n2606 & n27051 ) | ( n27049 & n27051 ) ;
  assign n27053 = x59 & n27051 ;
  assign n27054 = x59 & n27044 ;
  assign n27055 = ( x59 & n27048 ) | ( x59 & n27054 ) | ( n27048 & n27054 ) ;
  assign n27056 = ( n2606 & n27053 ) | ( n2606 & n27055 ) | ( n27053 & n27055 ) ;
  assign n27057 = x59 & ~n27055 ;
  assign n27058 = x59 & ~n27051 ;
  assign n27059 = ( ~n2606 & n27057 ) | ( ~n2606 & n27058 ) | ( n27057 & n27058 ) ;
  assign n27060 = ( n27052 & ~n27056 ) | ( n27052 & n27059 ) | ( ~n27056 & n27059 ) ;
  assign n27061 = n27043 | n27060 ;
  assign n27062 = n27043 & ~n27060 ;
  assign n27063 = ( ~n27043 & n27061 ) | ( ~n27043 & n27062 ) | ( n27061 & n27062 ) ;
  assign n27064 = ~n27009 & n27063 ;
  assign n27065 = n27009 & ~n27063 ;
  assign n27066 = n27064 | n27065 ;
  assign n27067 = x89 & n14045 ;
  assign n27068 = x88 & n14040 ;
  assign n27069 = x87 & ~n14039 ;
  assign n27070 = n14552 & n27069 ;
  assign n27071 = n27068 | n27070 ;
  assign n27072 = n27067 | n27071 ;
  assign n27073 = n14048 | n27067 ;
  assign n27074 = n27071 | n27073 ;
  assign n27075 = ( n3282 & n27072 ) | ( n3282 & n27074 ) | ( n27072 & n27074 ) ;
  assign n27076 = x56 & n27074 ;
  assign n27077 = x56 & n27067 ;
  assign n27078 = ( x56 & n27071 ) | ( x56 & n27077 ) | ( n27071 & n27077 ) ;
  assign n27079 = ( n3282 & n27076 ) | ( n3282 & n27078 ) | ( n27076 & n27078 ) ;
  assign n27080 = x56 & ~n27078 ;
  assign n27081 = x56 & ~n27074 ;
  assign n27082 = ( ~n3282 & n27080 ) | ( ~n3282 & n27081 ) | ( n27080 & n27081 ) ;
  assign n27083 = ( n27075 & ~n27079 ) | ( n27075 & n27082 ) | ( ~n27079 & n27082 ) ;
  assign n27084 = n27066 & n27083 ;
  assign n27085 = n27008 & ~n27084 ;
  assign n27086 = n27063 & ~n27083 ;
  assign n27087 = ( n27009 & n27083 ) | ( n27009 & ~n27086 ) | ( n27083 & ~n27086 ) ;
  assign n27088 = n27064 | n27087 ;
  assign n27089 = n27085 & n27088 ;
  assign n27090 = ~n27008 & n27084 ;
  assign n27091 = ( n27008 & n27088 ) | ( n27008 & ~n27090 ) | ( n27088 & ~n27090 ) ;
  assign n27092 = ~n27089 & n27091 ;
  assign n27093 = x92 & n12574 ;
  assign n27094 = x91 & n12569 ;
  assign n27095 = x90 & ~n12568 ;
  assign n27096 = n13076 & n27095 ;
  assign n27097 = n27094 | n27096 ;
  assign n27098 = n27093 | n27097 ;
  assign n27099 = n12577 | n27093 ;
  assign n27100 = n27097 | n27099 ;
  assign n27101 = ( n4040 & n27098 ) | ( n4040 & n27100 ) | ( n27098 & n27100 ) ;
  assign n27102 = x53 & n27100 ;
  assign n27103 = x53 & n27093 ;
  assign n27104 = ( x53 & n27097 ) | ( x53 & n27103 ) | ( n27097 & n27103 ) ;
  assign n27105 = ( n4040 & n27102 ) | ( n4040 & n27104 ) | ( n27102 & n27104 ) ;
  assign n27106 = x53 & ~n27104 ;
  assign n27107 = x53 & ~n27100 ;
  assign n27108 = ( ~n4040 & n27106 ) | ( ~n4040 & n27107 ) | ( n27106 & n27107 ) ;
  assign n27109 = ( n27101 & ~n27105 ) | ( n27101 & n27108 ) | ( ~n27105 & n27108 ) ;
  assign n27110 = n27092 & ~n27109 ;
  assign n27111 = ~n27092 & n27109 ;
  assign n27112 = n27110 | n27111 ;
  assign n27113 = n26613 | n26617 ;
  assign n27114 = ~n26613 & n26614 ;
  assign n27115 = ( n26618 & n27113 ) | ( n26618 & ~n27114 ) | ( n27113 & ~n27114 ) ;
  assign n27116 = ~n27112 & n27115 ;
  assign n27117 = n27112 & ~n27115 ;
  assign n27118 = n27116 | n27117 ;
  assign n27119 = x95 & n11205 ;
  assign n27120 = x94 & n11200 ;
  assign n27121 = x93 & ~n11199 ;
  assign n27122 = n11679 & n27121 ;
  assign n27123 = n27120 | n27122 ;
  assign n27124 = n27119 | n27123 ;
  assign n27125 = n11208 | n27119 ;
  assign n27126 = n27123 | n27125 ;
  assign n27127 = ( n4897 & n27124 ) | ( n4897 & n27126 ) | ( n27124 & n27126 ) ;
  assign n27128 = x50 & n27126 ;
  assign n27129 = x50 & n27119 ;
  assign n27130 = ( x50 & n27123 ) | ( x50 & n27129 ) | ( n27123 & n27129 ) ;
  assign n27131 = ( n4897 & n27128 ) | ( n4897 & n27130 ) | ( n27128 & n27130 ) ;
  assign n27132 = x50 & ~n27130 ;
  assign n27133 = x50 & ~n27126 ;
  assign n27134 = ( ~n4897 & n27132 ) | ( ~n4897 & n27133 ) | ( n27132 & n27133 ) ;
  assign n27135 = ( n27127 & ~n27131 ) | ( n27127 & n27134 ) | ( ~n27131 & n27134 ) ;
  assign n27136 = n27118 | n27135 ;
  assign n27137 = n27118 & ~n27135 ;
  assign n27138 = ( ~n27118 & n27136 ) | ( ~n27118 & n27137 ) | ( n27136 & n27137 ) ;
  assign n27139 = ~n26640 & n26644 ;
  assign n27140 = ~n26640 & n26641 ;
  assign n27141 = ( ~n26646 & n27139 ) | ( ~n26646 & n27140 ) | ( n27139 & n27140 ) ;
  assign n27142 = n27138 & n27141 ;
  assign n27143 = n27138 | n27141 ;
  assign n27144 = ~n27142 & n27143 ;
  assign n27145 = x98 & n9933 ;
  assign n27146 = x97 & n9928 ;
  assign n27147 = x96 & ~n9927 ;
  assign n27148 = n10379 & n27147 ;
  assign n27149 = n27146 | n27148 ;
  assign n27150 = n27145 | n27149 ;
  assign n27151 = n9936 | n27145 ;
  assign n27152 = n27149 | n27151 ;
  assign n27153 = ( ~n5850 & n27150 ) | ( ~n5850 & n27152 ) | ( n27150 & n27152 ) ;
  assign n27154 = n27150 & n27152 ;
  assign n27155 = ( n5834 & n27153 ) | ( n5834 & n27154 ) | ( n27153 & n27154 ) ;
  assign n27156 = x47 & n27152 ;
  assign n27157 = x47 & n27145 ;
  assign n27158 = ( x47 & n27149 ) | ( x47 & n27157 ) | ( n27149 & n27157 ) ;
  assign n27159 = ( ~n5850 & n27156 ) | ( ~n5850 & n27158 ) | ( n27156 & n27158 ) ;
  assign n27160 = n27156 & n27158 ;
  assign n27161 = ( n5834 & n27159 ) | ( n5834 & n27160 ) | ( n27159 & n27160 ) ;
  assign n27162 = x47 & ~n27158 ;
  assign n27163 = x47 & ~n27152 ;
  assign n27164 = ( n5850 & n27162 ) | ( n5850 & n27163 ) | ( n27162 & n27163 ) ;
  assign n27165 = n27162 | n27163 ;
  assign n27166 = ( ~n5834 & n27164 ) | ( ~n5834 & n27165 ) | ( n27164 & n27165 ) ;
  assign n27167 = ( n27155 & ~n27161 ) | ( n27155 & n27166 ) | ( ~n27161 & n27166 ) ;
  assign n27168 = n27144 | n27167 ;
  assign n27169 = n27144 & n27167 ;
  assign n27170 = n27168 & ~n27169 ;
  assign n27173 = n27170 & n27172 ;
  assign n27174 = n27172 & ~n27173 ;
  assign n27175 = x101 & n8724 ;
  assign n27176 = x100 & n8719 ;
  assign n27177 = x99 & ~n8718 ;
  assign n27178 = n9149 & n27177 ;
  assign n27179 = n27176 | n27178 ;
  assign n27180 = n27175 | n27179 ;
  assign n27181 = n8727 | n27175 ;
  assign n27182 = n27179 | n27181 ;
  assign n27183 = ( n6844 & n27180 ) | ( n6844 & n27182 ) | ( n27180 & n27182 ) ;
  assign n27184 = x44 & n27182 ;
  assign n27185 = x44 & n27175 ;
  assign n27186 = ( x44 & n27179 ) | ( x44 & n27185 ) | ( n27179 & n27185 ) ;
  assign n27187 = ( n6844 & n27184 ) | ( n6844 & n27186 ) | ( n27184 & n27186 ) ;
  assign n27188 = x44 & ~n27186 ;
  assign n27189 = x44 & ~n27182 ;
  assign n27190 = ( ~n6844 & n27188 ) | ( ~n6844 & n27189 ) | ( n27188 & n27189 ) ;
  assign n27191 = ( n27183 & ~n27187 ) | ( n27183 & n27190 ) | ( ~n27187 & n27190 ) ;
  assign n27192 = n27170 | n27191 ;
  assign n27193 = ( ~n27172 & n27191 ) | ( ~n27172 & n27192 ) | ( n27191 & n27192 ) ;
  assign n27194 = n27174 | n27193 ;
  assign n27195 = ( n27170 & n27172 ) | ( n27170 & n27191 ) | ( n27172 & n27191 ) ;
  assign n27196 = ~n27173 & n27195 ;
  assign n27197 = n27194 & ~n27196 ;
  assign n27198 = x104 & n7566 ;
  assign n27199 = x103 & n7561 ;
  assign n27200 = x102 & ~n7560 ;
  assign n27201 = n7953 & n27200 ;
  assign n27202 = n27199 | n27201 ;
  assign n27203 = n27198 | n27202 ;
  assign n27204 = n7569 | n27198 ;
  assign n27205 = n27202 | n27204 ;
  assign n27206 = ( n7911 & n27203 ) | ( n7911 & n27205 ) | ( n27203 & n27205 ) ;
  assign n27207 = x41 & n27205 ;
  assign n27208 = x41 & n27198 ;
  assign n27209 = ( x41 & n27202 ) | ( x41 & n27208 ) | ( n27202 & n27208 ) ;
  assign n27210 = ( n7911 & n27207 ) | ( n7911 & n27209 ) | ( n27207 & n27209 ) ;
  assign n27211 = x41 & ~n27209 ;
  assign n27212 = x41 & ~n27205 ;
  assign n27213 = ( ~n7911 & n27211 ) | ( ~n7911 & n27212 ) | ( n27211 & n27212 ) ;
  assign n27214 = ( n27206 & ~n27210 ) | ( n27206 & n27213 ) | ( ~n27210 & n27213 ) ;
  assign n27215 = n26699 | n26705 ;
  assign n27216 = ( n26699 & n26704 ) | ( n26699 & n27215 ) | ( n26704 & n27215 ) ;
  assign n27217 = ( n27197 & n27214 ) | ( n27197 & ~n27216 ) | ( n27214 & ~n27216 ) ;
  assign n27218 = ( ~n27214 & n27216 ) | ( ~n27214 & n27217 ) | ( n27216 & n27217 ) ;
  assign n27219 = ( ~n27197 & n27217 ) | ( ~n27197 & n27218 ) | ( n27217 & n27218 ) ;
  assign n27220 = n27004 | n27219 ;
  assign n27221 = n27004 & n27219 ;
  assign n27222 = n27220 & ~n27221 ;
  assign n27223 = x107 & n6536 ;
  assign n27224 = x106 & n6531 ;
  assign n27225 = x105 & ~n6530 ;
  assign n27226 = n6871 & n27225 ;
  assign n27227 = n27224 | n27226 ;
  assign n27228 = n27223 | n27227 ;
  assign n27229 = n6539 | n27223 ;
  assign n27230 = n27227 | n27229 ;
  assign n27231 = ( n9084 & n27228 ) | ( n9084 & n27230 ) | ( n27228 & n27230 ) ;
  assign n27232 = x38 & n27230 ;
  assign n27233 = x38 & n27223 ;
  assign n27234 = ( x38 & n27227 ) | ( x38 & n27233 ) | ( n27227 & n27233 ) ;
  assign n27235 = ( n9084 & n27232 ) | ( n9084 & n27234 ) | ( n27232 & n27234 ) ;
  assign n27236 = x38 & ~n27234 ;
  assign n27237 = x38 & ~n27230 ;
  assign n27238 = ( ~n9084 & n27236 ) | ( ~n9084 & n27237 ) | ( n27236 & n27237 ) ;
  assign n27239 = ( n27231 & ~n27235 ) | ( n27231 & n27238 ) | ( ~n27235 & n27238 ) ;
  assign n27240 = n27222 & ~n27239 ;
  assign n27241 = n27222 | n27239 ;
  assign n27242 = ( ~n27222 & n27240 ) | ( ~n27222 & n27241 ) | ( n27240 & n27241 ) ;
  assign n27243 = n26754 & n27242 ;
  assign n27244 = ( n26760 & n27242 ) | ( n26760 & n27243 ) | ( n27242 & n27243 ) ;
  assign n27245 = n26754 | n27242 ;
  assign n27246 = n26760 | n27245 ;
  assign n27247 = ~n27244 & n27246 ;
  assign n27248 = x110 & n5554 ;
  assign n27249 = x109 & n5549 ;
  assign n27250 = x108 & ~n5548 ;
  assign n27251 = n5893 & n27250 ;
  assign n27252 = n27249 | n27251 ;
  assign n27253 = n27248 | n27252 ;
  assign n27254 = n5557 | n27248 ;
  assign n27255 = n27252 | n27254 ;
  assign n27256 = ( n10330 & n27253 ) | ( n10330 & n27255 ) | ( n27253 & n27255 ) ;
  assign n27257 = x35 & n27255 ;
  assign n27258 = x35 & n27248 ;
  assign n27259 = ( x35 & n27252 ) | ( x35 & n27258 ) | ( n27252 & n27258 ) ;
  assign n27260 = ( n10330 & n27257 ) | ( n10330 & n27259 ) | ( n27257 & n27259 ) ;
  assign n27261 = x35 & ~n27259 ;
  assign n27262 = x35 & ~n27255 ;
  assign n27263 = ( ~n10330 & n27261 ) | ( ~n10330 & n27262 ) | ( n27261 & n27262 ) ;
  assign n27264 = ( n27256 & ~n27260 ) | ( n27256 & n27263 ) | ( ~n27260 & n27263 ) ;
  assign n27265 = ~n27247 & n27264 ;
  assign n27266 = n27244 | n27264 ;
  assign n27267 = n27246 & ~n27266 ;
  assign n27268 = n27265 | n27267 ;
  assign n27269 = n26978 & n27268 ;
  assign n27270 = n26978 | n27268 ;
  assign n27001 = n26993 & ~n26998 ;
  assign n27271 = ( n26978 & ~n27001 ) | ( n26978 & n27268 ) | ( ~n27001 & n27268 ) ;
  assign n27272 = ( n26817 & n27270 ) | ( n26817 & n27271 ) | ( n27270 & n27271 ) ;
  assign n27273 = ( ~n27000 & n27269 ) | ( ~n27000 & n27272 ) | ( n27269 & n27272 ) ;
  assign n27002 = ~n26817 & n27001 ;
  assign n27003 = n27000 | n27002 ;
  assign n27274 = ( n27003 & ~n27268 ) | ( n27003 & n27273 ) | ( ~n27268 & n27273 ) ;
  assign n27275 = ( ~n26978 & n27273 ) | ( ~n26978 & n27274 ) | ( n27273 & n27274 ) ;
  assign n27277 = x121 & n2424 ;
  assign n27278 = x120 & ~n2423 ;
  assign n27279 = n2631 & n27278 ;
  assign n27280 = n27277 | n27279 ;
  assign n27276 = x122 & n2429 ;
  assign n27282 = n2432 | n27276 ;
  assign n27283 = n27280 | n27282 ;
  assign n27281 = n27276 | n27280 ;
  assign n27284 = n27281 & n27283 ;
  assign n27285 = ( n16043 & n27283 ) | ( n16043 & n27284 ) | ( n27283 & n27284 ) ;
  assign n27286 = x23 & n27284 ;
  assign n27287 = x23 & n27283 ;
  assign n27288 = ( n16043 & n27286 ) | ( n16043 & n27287 ) | ( n27286 & n27287 ) ;
  assign n27289 = x23 & ~n27284 ;
  assign n27290 = x23 & ~n27283 ;
  assign n27291 = ( ~n16043 & n27289 ) | ( ~n16043 & n27290 ) | ( n27289 & n27290 ) ;
  assign n27292 = ( n27285 & ~n27288 ) | ( n27285 & n27291 ) | ( ~n27288 & n27291 ) ;
  assign n27293 = n26842 | n26882 ;
  assign n27294 = ( n26882 & n26883 ) | ( n26882 & n27293 ) | ( n26883 & n27293 ) ;
  assign n27295 = n27292 & n27294 ;
  assign n27296 = n27292 | n27294 ;
  assign n27297 = ~n27295 & n27296 ;
  assign n27298 = x119 & n3085 ;
  assign n27299 = x118 & n3080 ;
  assign n27300 = x117 & ~n3079 ;
  assign n27301 = n3309 & n27300 ;
  assign n27302 = n27299 | n27301 ;
  assign n27303 = n27298 | n27302 ;
  assign n27304 = n3088 | n27298 ;
  assign n27305 = n27302 | n27304 ;
  assign n27306 = ( n14496 & n27303 ) | ( n14496 & n27305 ) | ( n27303 & n27305 ) ;
  assign n27307 = x26 & n27305 ;
  assign n27308 = x26 & n27298 ;
  assign n27309 = ( x26 & n27302 ) | ( x26 & n27308 ) | ( n27302 & n27308 ) ;
  assign n27310 = ( n14496 & n27307 ) | ( n14496 & n27309 ) | ( n27307 & n27309 ) ;
  assign n27311 = x26 & ~n27309 ;
  assign n27312 = x26 & ~n27305 ;
  assign n27313 = ( ~n14496 & n27311 ) | ( ~n14496 & n27312 ) | ( n27311 & n27312 ) ;
  assign n27314 = ( n27306 & ~n27310 ) | ( n27306 & n27313 ) | ( ~n27310 & n27313 ) ;
  assign n27315 = n26820 | n26838 ;
  assign n27316 = ( n26838 & n26839 ) | ( n26838 & n27315 ) | ( n26839 & n27315 ) ;
  assign n27317 = n27314 | n27316 ;
  assign n27318 = n27314 & n27316 ;
  assign n27319 = n27317 & ~n27318 ;
  assign n27320 = ( n27275 & n27297 ) | ( n27275 & ~n27319 ) | ( n27297 & ~n27319 ) ;
  assign n27321 = ( ~n27297 & n27319 ) | ( ~n27297 & n27320 ) | ( n27319 & n27320 ) ;
  assign n27322 = ( ~n27275 & n27320 ) | ( ~n27275 & n27321 ) | ( n27320 & n27321 ) ;
  assign n27323 = x127 & n1378 ;
  assign n27324 = x126 & ~n1377 ;
  assign n27325 = n1542 & n27324 ;
  assign n27326 = n27323 | n27325 ;
  assign n27327 = n1386 | n27326 ;
  assign n27328 = ( n19328 & n27326 ) | ( n19328 & n27327 ) | ( n27326 & n27327 ) ;
  assign n27329 = x17 & n27326 ;
  assign n27330 = ( x17 & n2676 ) | ( x17 & n27326 ) | ( n2676 & n27326 ) ;
  assign n27331 = ( n19328 & n27329 ) | ( n19328 & n27330 ) | ( n27329 & n27330 ) ;
  assign n27332 = x17 & ~n2676 ;
  assign n27333 = ~n27326 & n27332 ;
  assign n27334 = x17 & ~n27326 ;
  assign n27335 = ( ~n19328 & n27333 ) | ( ~n19328 & n27334 ) | ( n27333 & n27334 ) ;
  assign n27336 = ( n27328 & ~n27331 ) | ( n27328 & n27335 ) | ( ~n27331 & n27335 ) ;
  assign n27337 = n26886 | n26910 ;
  assign n27338 = ( n26910 & n26911 ) | ( n26910 & n27337 ) | ( n26911 & n27337 ) ;
  assign n27339 = n27336 & n27338 ;
  assign n27340 = n27336 | n27338 ;
  assign n27341 = ~n27339 & n27340 ;
  assign n27342 = x125 & n1859 ;
  assign n27343 = x124 & n1854 ;
  assign n27344 = x123 & ~n1853 ;
  assign n27345 = n2037 & n27344 ;
  assign n27346 = n27343 | n27345 ;
  assign n27347 = n27342 | n27346 ;
  assign n27348 = n1862 | n27342 ;
  assign n27349 = n27346 | n27348 ;
  assign n27350 = ( n17670 & n27347 ) | ( n17670 & n27349 ) | ( n27347 & n27349 ) ;
  assign n27351 = x20 & n27349 ;
  assign n27352 = x20 & n27342 ;
  assign n27353 = ( x20 & n27346 ) | ( x20 & n27352 ) | ( n27346 & n27352 ) ;
  assign n27354 = ( n17670 & n27351 ) | ( n17670 & n27353 ) | ( n27351 & n27353 ) ;
  assign n27355 = x20 & ~n27353 ;
  assign n27356 = x20 & ~n27349 ;
  assign n27357 = ( ~n17670 & n27355 ) | ( ~n17670 & n27356 ) | ( n27355 & n27356 ) ;
  assign n27358 = ( n27350 & ~n27354 ) | ( n27350 & n27357 ) | ( ~n27354 & n27357 ) ;
  assign n27359 = n26842 & n26883 ;
  assign n27360 = n26842 | n26883 ;
  assign n27361 = ~n27359 & n27360 ;
  assign n27362 = n27358 & n27361 ;
  assign n27363 = n26859 & n27358 ;
  assign n27364 = ( n26861 & n27362 ) | ( n26861 & n27363 ) | ( n27362 & n27363 ) ;
  assign n27365 = n27358 | n27361 ;
  assign n27366 = n26859 | n27358 ;
  assign n27367 = ( n26861 & n27365 ) | ( n26861 & n27366 ) | ( n27365 & n27366 ) ;
  assign n27368 = ~n27364 & n27367 ;
  assign n27369 = ( n27322 & n27341 ) | ( n27322 & ~n27368 ) | ( n27341 & ~n27368 ) ;
  assign n27370 = ( ~n27341 & n27368 ) | ( ~n27341 & n27369 ) | ( n27368 & n27369 ) ;
  assign n27371 = ( ~n27322 & n27369 ) | ( ~n27322 & n27370 ) | ( n27369 & n27370 ) ;
  assign n27372 = n26886 & n26911 ;
  assign n27373 = n26886 | n26911 ;
  assign n27374 = ~n27372 & n27373 ;
  assign n27375 = n26933 | n27374 ;
  assign n27376 = ( n26933 & n26937 ) | ( n26933 & n27375 ) | ( n26937 & n27375 ) ;
  assign n27377 = n27371 | n27376 ;
  assign n27378 = n27371 & n27376 ;
  assign n27379 = n27377 & ~n27378 ;
  assign n27380 = n26947 | n26956 ;
  assign n27381 = n26947 | n26948 ;
  assign n27382 = ( n26490 & n26947 ) | ( n26490 & n27381 ) | ( n26947 & n27381 ) ;
  assign n27383 = ( n26495 & n27380 ) | ( n26495 & n27382 ) | ( n27380 & n27382 ) ;
  assign n27384 = ( n26947 & n26951 ) | ( n26947 & n27381 ) | ( n26951 & n27381 ) ;
  assign n27385 = ( n26030 & n27383 ) | ( n26030 & n27384 ) | ( n27383 & n27384 ) ;
  assign n27386 = n27379 | n27385 ;
  assign n27387 = n27379 & n27383 ;
  assign n27388 = n26947 & n27379 ;
  assign n27389 = ( n26948 & n27379 ) | ( n26948 & n27388 ) | ( n27379 & n27388 ) ;
  assign n27390 = ( n26951 & n27388 ) | ( n26951 & n27389 ) | ( n27388 & n27389 ) ;
  assign n27391 = ( n26030 & n27387 ) | ( n26030 & n27390 ) | ( n27387 & n27390 ) ;
  assign n27392 = n27386 & ~n27391 ;
  assign n27833 = n27322 & n27368 ;
  assign n27834 = n27322 | n27368 ;
  assign n27835 = ~n27833 & n27834 ;
  assign n27836 = n27336 | n27835 ;
  assign n27837 = ( n27338 & n27835 ) | ( n27338 & n27836 ) | ( n27835 & n27836 ) ;
  assign n27838 = ( n27339 & n27341 ) | ( n27339 & n27837 ) | ( n27341 & n27837 ) ;
  assign n27411 = n27364 | n27368 ;
  assign n27412 = ( n27322 & n27364 ) | ( n27322 & n27411 ) | ( n27364 & n27411 ) ;
  assign n27393 = x127 & ~n1377 ;
  assign n27394 = n1542 & n27393 ;
  assign n27395 = n1386 & n19877 ;
  assign n27396 = n27394 | n27395 ;
  assign n27397 = n1386 & n19880 ;
  assign n27398 = n27394 | n27397 ;
  assign n27399 = ( n18202 & n27396 ) | ( n18202 & n27398 ) | ( n27396 & n27398 ) ;
  assign n27400 = n27396 & n27398 ;
  assign n27401 = ( n18212 & n27399 ) | ( n18212 & n27400 ) | ( n27399 & n27400 ) ;
  assign n27402 = ( n18214 & n27399 ) | ( n18214 & n27400 ) | ( n27399 & n27400 ) ;
  assign n27403 = ( n14002 & n27401 ) | ( n14002 & n27402 ) | ( n27401 & n27402 ) ;
  assign n27404 = x17 & n27401 ;
  assign n27405 = x17 & n27402 ;
  assign n27406 = ( n14002 & n27404 ) | ( n14002 & n27405 ) | ( n27404 & n27405 ) ;
  assign n27407 = x17 & ~n27405 ;
  assign n27408 = x17 & ~n27404 ;
  assign n27409 = ( ~n14002 & n27407 ) | ( ~n14002 & n27408 ) | ( n27407 & n27408 ) ;
  assign n27410 = ( n27403 & ~n27406 ) | ( n27403 & n27409 ) | ( ~n27406 & n27409 ) ;
  assign n27413 = n27410 & n27412 ;
  assign n27414 = n27412 & ~n27413 ;
  assign n27415 = x126 & n1859 ;
  assign n27416 = x125 & n1854 ;
  assign n27417 = x124 & ~n1853 ;
  assign n27418 = n2037 & n27417 ;
  assign n27419 = n27416 | n27418 ;
  assign n27420 = n27415 | n27419 ;
  assign n27421 = n1862 | n27415 ;
  assign n27422 = n27419 | n27421 ;
  assign n27423 = ( n18220 & n27420 ) | ( n18220 & n27422 ) | ( n27420 & n27422 ) ;
  assign n27424 = x20 & n27422 ;
  assign n27425 = x20 & n27415 ;
  assign n27426 = ( x20 & n27419 ) | ( x20 & n27425 ) | ( n27419 & n27425 ) ;
  assign n27427 = ( n18220 & n27424 ) | ( n18220 & n27426 ) | ( n27424 & n27426 ) ;
  assign n27428 = x20 & ~n27426 ;
  assign n27429 = x20 & ~n27422 ;
  assign n27430 = ( ~n18220 & n27428 ) | ( ~n18220 & n27429 ) | ( n27428 & n27429 ) ;
  assign n27431 = ( n27423 & ~n27427 ) | ( n27423 & n27430 ) | ( ~n27427 & n27430 ) ;
  assign n27432 = n27275 & n27319 ;
  assign n27433 = n27275 | n27319 ;
  assign n27434 = ~n27432 & n27433 ;
  assign n27435 = n27295 | n27434 ;
  assign n27436 = ( n27295 & n27297 ) | ( n27295 & n27435 ) | ( n27297 & n27435 ) ;
  assign n27437 = n27431 | n27436 ;
  assign n27438 = n27431 & n27436 ;
  assign n27439 = n27437 & ~n27438 ;
  assign n27440 = n27001 & n27270 ;
  assign n27441 = ~n26817 & n27440 ;
  assign n27442 = ~n26998 & n27268 ;
  assign n27443 = n26978 & n27442 ;
  assign n27444 = ~n26993 & n27268 ;
  assign n27445 = n26978 & n27444 ;
  assign n27446 = ( ~n26817 & n27443 ) | ( ~n26817 & n27445 ) | ( n27443 & n27445 ) ;
  assign n27447 = ( n26999 & n27441 ) | ( n26999 & ~n27446 ) | ( n27441 & ~n27446 ) ;
  assign n27448 = x120 & n3085 ;
  assign n27449 = x119 & n3080 ;
  assign n27450 = x118 & ~n3079 ;
  assign n27451 = n3309 & n27450 ;
  assign n27452 = n27449 | n27451 ;
  assign n27453 = n27448 | n27452 ;
  assign n27454 = n3088 | n27448 ;
  assign n27455 = n27452 | n27454 ;
  assign n27456 = ( n14991 & n27453 ) | ( n14991 & n27455 ) | ( n27453 & n27455 ) ;
  assign n27457 = x26 & n27455 ;
  assign n27458 = x26 & n27448 ;
  assign n27459 = ( x26 & n27452 ) | ( x26 & n27458 ) | ( n27452 & n27458 ) ;
  assign n27460 = ( n14991 & n27457 ) | ( n14991 & n27459 ) | ( n27457 & n27459 ) ;
  assign n27461 = x26 & ~n27459 ;
  assign n27462 = x26 & ~n27455 ;
  assign n27463 = ( ~n14991 & n27461 ) | ( ~n14991 & n27462 ) | ( n27461 & n27462 ) ;
  assign n27464 = ( n27456 & ~n27460 ) | ( n27456 & n27463 ) | ( ~n27460 & n27463 ) ;
  assign n27465 = ( n26999 & n27270 ) | ( n26999 & ~n27446 ) | ( n27270 & ~n27446 ) ;
  assign n27466 = n27464 & n27465 ;
  assign n27467 = n27000 & n27464 ;
  assign n27468 = ( n27447 & n27466 ) | ( n27447 & n27467 ) | ( n27466 & n27467 ) ;
  assign n27469 = n27464 | n27465 ;
  assign n27470 = n27000 | n27464 ;
  assign n27471 = ( n27447 & n27469 ) | ( n27447 & n27470 ) | ( n27469 & n27470 ) ;
  assign n27472 = ~n27468 & n27471 ;
  assign n27473 = n27275 | n27318 ;
  assign n27474 = ( n27318 & n27319 ) | ( n27318 & n27473 ) | ( n27319 & n27473 ) ;
  assign n27475 = x123 & n2429 ;
  assign n27476 = x122 & n2424 ;
  assign n27477 = x121 & ~n2423 ;
  assign n27478 = n2631 & n27477 ;
  assign n27479 = n27476 | n27478 ;
  assign n27480 = n27475 | n27479 ;
  assign n27481 = n2432 | n27475 ;
  assign n27482 = n27479 | n27481 ;
  assign n27483 = ( n16086 & n27480 ) | ( n16086 & n27482 ) | ( n27480 & n27482 ) ;
  assign n27484 = x23 & n27482 ;
  assign n27485 = x23 & n27475 ;
  assign n27486 = ( x23 & n27479 ) | ( x23 & n27485 ) | ( n27479 & n27485 ) ;
  assign n27487 = ( n16086 & n27484 ) | ( n16086 & n27486 ) | ( n27484 & n27486 ) ;
  assign n27488 = x23 & ~n27486 ;
  assign n27489 = x23 & ~n27482 ;
  assign n27490 = ( ~n16086 & n27488 ) | ( ~n16086 & n27489 ) | ( n27488 & n27489 ) ;
  assign n27491 = ( n27483 & ~n27487 ) | ( n27483 & n27490 ) | ( ~n27487 & n27490 ) ;
  assign n27492 = n27314 & n27491 ;
  assign n27493 = n27316 & n27492 ;
  assign n27494 = ( n27275 & n27491 ) | ( n27275 & n27493 ) | ( n27491 & n27493 ) ;
  assign n27495 = n27491 & n27493 ;
  assign n27496 = ( n27319 & n27494 ) | ( n27319 & n27495 ) | ( n27494 & n27495 ) ;
  assign n27497 = n27474 & ~n27496 ;
  assign n27503 = x114 & n4631 ;
  assign n27504 = x113 & n4626 ;
  assign n27505 = x112 & ~n4625 ;
  assign n27506 = n4943 & n27505 ;
  assign n27507 = n27504 | n27506 ;
  assign n27508 = n27503 | n27507 ;
  assign n27509 = n4634 | n27503 ;
  assign n27510 = n27507 | n27509 ;
  assign n27511 = ( ~n12095 & n27508 ) | ( ~n12095 & n27510 ) | ( n27508 & n27510 ) ;
  assign n27512 = n27508 & n27510 ;
  assign n27513 = ( n12079 & n27511 ) | ( n12079 & n27512 ) | ( n27511 & n27512 ) ;
  assign n27514 = x32 & n27513 ;
  assign n27515 = x32 & ~n27513 ;
  assign n27516 = ( n27513 & ~n27514 ) | ( n27513 & n27515 ) | ( ~n27514 & n27515 ) ;
  assign n27517 = ( n27244 & n27247 ) | ( n27244 & n27266 ) | ( n27247 & n27266 ) ;
  assign n27518 = n27516 | n27517 ;
  assign n27519 = n27516 & n27517 ;
  assign n27520 = n27518 & ~n27519 ;
  assign n27521 = x117 & n3816 ;
  assign n27522 = x116 & n3811 ;
  assign n27523 = x115 & ~n3810 ;
  assign n27524 = n4067 & n27523 ;
  assign n27525 = n27522 | n27524 ;
  assign n27526 = n27521 | n27525 ;
  assign n27527 = n3819 | n27521 ;
  assign n27528 = n27525 | n27527 ;
  assign n27529 = ( ~n13522 & n27526 ) | ( ~n13522 & n27528 ) | ( n27526 & n27528 ) ;
  assign n27530 = n27526 & n27528 ;
  assign n27531 = ( n13503 & n27529 ) | ( n13503 & n27530 ) | ( n27529 & n27530 ) ;
  assign n27532 = x29 & n27531 ;
  assign n27533 = x29 & ~n27531 ;
  assign n27534 = ( n27531 & ~n27532 ) | ( n27531 & n27533 ) | ( ~n27532 & n27533 ) ;
  assign n27535 = n26973 & n27534 ;
  assign n27536 = ( n27268 & n27534 ) | ( n27268 & n27535 ) | ( n27534 & n27535 ) ;
  assign n27537 = n27268 & n27534 ;
  assign n27538 = ( n26975 & n27536 ) | ( n26975 & n27537 ) | ( n27536 & n27537 ) ;
  assign n27539 = n27534 & n27535 ;
  assign n27540 = n26975 & n27539 ;
  assign n27541 = ( n26978 & n27538 ) | ( n26978 & n27540 ) | ( n27538 & n27540 ) ;
  assign n27542 = n26973 | n27268 ;
  assign n27543 = ( n26975 & n27268 ) | ( n26975 & n27542 ) | ( n27268 & n27542 ) ;
  assign n27544 = ( n26977 & n26978 ) | ( n26977 & n27543 ) | ( n26978 & n27543 ) ;
  assign n27545 = ~n27541 & n27544 ;
  assign n27553 = x102 & n8724 ;
  assign n27554 = x101 & n8719 ;
  assign n27555 = x100 & ~n8718 ;
  assign n27556 = n9149 & n27555 ;
  assign n27557 = n27554 | n27556 ;
  assign n27558 = n27553 | n27557 ;
  assign n27559 = n8727 | n27553 ;
  assign n27560 = n27557 | n27559 ;
  assign n27561 = ( n7178 & n27558 ) | ( n7178 & n27560 ) | ( n27558 & n27560 ) ;
  assign n27562 = x44 & n27560 ;
  assign n27563 = x44 & n27553 ;
  assign n27564 = ( x44 & n27557 ) | ( x44 & n27563 ) | ( n27557 & n27563 ) ;
  assign n27565 = ( n7178 & n27562 ) | ( n7178 & n27564 ) | ( n27562 & n27564 ) ;
  assign n27566 = x44 & ~n27564 ;
  assign n27567 = x44 & ~n27560 ;
  assign n27568 = ( ~n7178 & n27566 ) | ( ~n7178 & n27567 ) | ( n27566 & n27567 ) ;
  assign n27569 = ( n27561 & ~n27565 ) | ( n27561 & n27568 ) | ( ~n27565 & n27568 ) ;
  assign n27570 = x96 & n11205 ;
  assign n27571 = x95 & n11200 ;
  assign n27572 = x94 & ~n11199 ;
  assign n27573 = n11679 & n27572 ;
  assign n27574 = n27571 | n27573 ;
  assign n27575 = n27570 | n27574 ;
  assign n27576 = n11208 | n27570 ;
  assign n27577 = n27574 | n27576 ;
  assign n27578 = ( n5202 & n27575 ) | ( n5202 & n27577 ) | ( n27575 & n27577 ) ;
  assign n27579 = x50 & n27577 ;
  assign n27580 = x50 & n27570 ;
  assign n27581 = ( x50 & n27574 ) | ( x50 & n27580 ) | ( n27574 & n27580 ) ;
  assign n27582 = ( n5202 & n27579 ) | ( n5202 & n27581 ) | ( n27579 & n27581 ) ;
  assign n27583 = x50 & ~n27581 ;
  assign n27584 = x50 & ~n27577 ;
  assign n27585 = ( ~n5202 & n27583 ) | ( ~n5202 & n27584 ) | ( n27583 & n27584 ) ;
  assign n27586 = ( n27578 & ~n27582 ) | ( n27578 & n27585 ) | ( ~n27582 & n27585 ) ;
  assign n27587 = x83 & n17141 ;
  assign n27588 = x82 & ~n17140 ;
  assign n27589 = n17724 & n27588 ;
  assign n27590 = n27587 | n27589 ;
  assign n27591 = x84 & n17146 ;
  assign n27592 = n17149 | n27591 ;
  assign n27593 = n27590 | n27592 ;
  assign n27594 = ~x62 & n27593 ;
  assign n27595 = ~x62 & n27591 ;
  assign n27596 = ( ~x62 & n27590 ) | ( ~x62 & n27595 ) | ( n27590 & n27595 ) ;
  assign n27597 = ( n2194 & n27594 ) | ( n2194 & n27596 ) | ( n27594 & n27596 ) ;
  assign n27598 = x62 & ~n27593 ;
  assign n27599 = x62 & x84 ;
  assign n27600 = n17146 & n27599 ;
  assign n27601 = x62 & ~n27600 ;
  assign n27602 = ~n27590 & n27601 ;
  assign n27603 = ( ~n2194 & n27598 ) | ( ~n2194 & n27602 ) | ( n27598 & n27602 ) ;
  assign n27604 = n27597 | n27603 ;
  assign n27605 = x81 & n18290 ;
  assign n27606 = x63 & x80 ;
  assign n27607 = ~n18290 & n27606 ;
  assign n27608 = n27605 | n27607 ;
  assign n27609 = ~n27013 & n27608 ;
  assign n27610 = n27013 & ~n27608 ;
  assign n27611 = n27609 | n27610 ;
  assign n27612 = n27604 & ~n27611 ;
  assign n27613 = n27604 & ~n27612 ;
  assign n27614 = ~n27015 & n27018 ;
  assign n27615 = ( n27015 & n27035 ) | ( n27015 & ~n27614 ) | ( n27035 & ~n27614 ) ;
  assign n27616 = n27604 | n27611 ;
  assign n27617 = n27615 & ~n27616 ;
  assign n27618 = ( n27613 & n27615 ) | ( n27613 & n27617 ) | ( n27615 & n27617 ) ;
  assign n27619 = ~n27615 & n27616 ;
  assign n27620 = ~n27613 & n27619 ;
  assign n27621 = n27618 | n27620 ;
  assign n27622 = x87 & n15552 ;
  assign n27623 = x86 & n15547 ;
  assign n27624 = x85 & ~n15546 ;
  assign n27625 = n16123 & n27624 ;
  assign n27626 = n27623 | n27625 ;
  assign n27627 = n27622 | n27626 ;
  assign n27628 = n15555 | n27622 ;
  assign n27629 = n27626 | n27628 ;
  assign n27630 = ( n2816 & n27627 ) | ( n2816 & n27629 ) | ( n27627 & n27629 ) ;
  assign n27631 = x59 & n27629 ;
  assign n27632 = x59 & n27622 ;
  assign n27633 = ( x59 & n27626 ) | ( x59 & n27632 ) | ( n27626 & n27632 ) ;
  assign n27634 = ( n2816 & n27631 ) | ( n2816 & n27633 ) | ( n27631 & n27633 ) ;
  assign n27635 = x59 & ~n27633 ;
  assign n27636 = x59 & ~n27629 ;
  assign n27637 = ( ~n2816 & n27635 ) | ( ~n2816 & n27636 ) | ( n27635 & n27636 ) ;
  assign n27638 = ( n27630 & ~n27634 ) | ( n27630 & n27637 ) | ( ~n27634 & n27637 ) ;
  assign n27639 = n27621 & ~n27638 ;
  assign n27640 = ~n27621 & n27638 ;
  assign n27641 = n27639 | n27640 ;
  assign n27642 = n27038 & ~n27060 ;
  assign n27643 = ( n27040 & n27060 ) | ( n27040 & ~n27642 ) | ( n27060 & ~n27642 ) ;
  assign n27644 = ( n27041 & ~n27043 ) | ( n27041 & n27643 ) | ( ~n27043 & n27643 ) ;
  assign n27645 = ~n27641 & n27644 ;
  assign n27646 = n27641 & ~n27644 ;
  assign n27647 = n27645 | n27646 ;
  assign n27648 = x90 & n14045 ;
  assign n27649 = x89 & n14040 ;
  assign n27650 = x88 & ~n14039 ;
  assign n27651 = n14552 & n27650 ;
  assign n27652 = n27649 | n27651 ;
  assign n27653 = n27648 | n27652 ;
  assign n27654 = n14048 | n27648 ;
  assign n27655 = n27652 | n27654 ;
  assign n27656 = ( n3519 & n27653 ) | ( n3519 & n27655 ) | ( n27653 & n27655 ) ;
  assign n27657 = x56 & n27655 ;
  assign n27658 = x56 & n27648 ;
  assign n27659 = ( x56 & n27652 ) | ( x56 & n27658 ) | ( n27652 & n27658 ) ;
  assign n27660 = ( n3519 & n27657 ) | ( n3519 & n27659 ) | ( n27657 & n27659 ) ;
  assign n27661 = x56 & ~n27659 ;
  assign n27662 = x56 & ~n27655 ;
  assign n27663 = ( ~n3519 & n27661 ) | ( ~n3519 & n27662 ) | ( n27661 & n27662 ) ;
  assign n27664 = ( n27656 & ~n27660 ) | ( n27656 & n27663 ) | ( ~n27660 & n27663 ) ;
  assign n27665 = ~n27647 & n27664 ;
  assign n27666 = n27647 & ~n27664 ;
  assign n27667 = n27665 | n27666 ;
  assign n27668 = ( n27065 & ~n27066 ) | ( n27065 & n27087 ) | ( ~n27066 & n27087 ) ;
  assign n27669 = ~n27667 & n27668 ;
  assign n27670 = n27667 & ~n27668 ;
  assign n27671 = n27669 | n27670 ;
  assign n27672 = x93 & n12574 ;
  assign n27673 = x92 & n12569 ;
  assign n27674 = x91 & ~n12568 ;
  assign n27675 = n13076 & n27674 ;
  assign n27676 = n27673 | n27675 ;
  assign n27677 = n27672 | n27676 ;
  assign n27678 = n12577 | n27672 ;
  assign n27679 = n27676 | n27678 ;
  assign n27680 = ( n4305 & n27677 ) | ( n4305 & n27679 ) | ( n27677 & n27679 ) ;
  assign n27681 = x53 & n27679 ;
  assign n27682 = x53 & n27672 ;
  assign n27683 = ( x53 & n27676 ) | ( x53 & n27682 ) | ( n27676 & n27682 ) ;
  assign n27684 = ( n4305 & n27681 ) | ( n4305 & n27683 ) | ( n27681 & n27683 ) ;
  assign n27685 = x53 & ~n27683 ;
  assign n27686 = x53 & ~n27679 ;
  assign n27687 = ( ~n4305 & n27685 ) | ( ~n4305 & n27686 ) | ( n27685 & n27686 ) ;
  assign n27688 = ( n27680 & ~n27684 ) | ( n27680 & n27687 ) | ( ~n27684 & n27687 ) ;
  assign n27689 = n27671 | n27688 ;
  assign n27690 = n27671 & ~n27688 ;
  assign n27691 = ( ~n27671 & n27689 ) | ( ~n27671 & n27690 ) | ( n27689 & n27690 ) ;
  assign n27692 = ~n27084 & n27088 ;
  assign n27693 = ( n27008 & n27109 ) | ( n27008 & ~n27692 ) | ( n27109 & ~n27692 ) ;
  assign n27694 = ( n27586 & n27691 ) | ( n27586 & ~n27693 ) | ( n27691 & ~n27693 ) ;
  assign n27695 = ( ~n27691 & n27693 ) | ( ~n27691 & n27694 ) | ( n27693 & n27694 ) ;
  assign n27696 = ( ~n27586 & n27694 ) | ( ~n27586 & n27695 ) | ( n27694 & n27695 ) ;
  assign n27697 = n27115 | n27135 ;
  assign n27698 = ( ~n27112 & n27135 ) | ( ~n27112 & n27697 ) | ( n27135 & n27697 ) ;
  assign n27699 = ( n27116 & ~n27118 ) | ( n27116 & n27698 ) | ( ~n27118 & n27698 ) ;
  assign n27700 = n27696 & ~n27699 ;
  assign n27701 = ~n27696 & n27699 ;
  assign n27702 = n27700 | n27701 ;
  assign n27703 = x99 & n9933 ;
  assign n27704 = x98 & n9928 ;
  assign n27705 = x97 & ~n9927 ;
  assign n27706 = n10379 & n27705 ;
  assign n27707 = n27704 | n27706 ;
  assign n27708 = n27703 | n27707 ;
  assign n27709 = n9936 | n27703 ;
  assign n27710 = n27707 | n27709 ;
  assign n27711 = ( n6164 & n27708 ) | ( n6164 & n27710 ) | ( n27708 & n27710 ) ;
  assign n27712 = x47 & n27710 ;
  assign n27713 = x47 & n27703 ;
  assign n27714 = ( x47 & n27707 ) | ( x47 & n27713 ) | ( n27707 & n27713 ) ;
  assign n27715 = ( n6164 & n27712 ) | ( n6164 & n27714 ) | ( n27712 & n27714 ) ;
  assign n27716 = x47 & ~n27714 ;
  assign n27717 = x47 & ~n27710 ;
  assign n27718 = ( ~n6164 & n27716 ) | ( ~n6164 & n27717 ) | ( n27716 & n27717 ) ;
  assign n27719 = ( n27711 & ~n27715 ) | ( n27711 & n27718 ) | ( ~n27715 & n27718 ) ;
  assign n27720 = n27702 & n27719 ;
  assign n27721 = n27694 & ~n27719 ;
  assign n27722 = n27586 | n27719 ;
  assign n27723 = ( n27695 & n27721 ) | ( n27695 & ~n27722 ) | ( n27721 & ~n27722 ) ;
  assign n27724 = ( n27699 & n27719 ) | ( n27699 & ~n27723 ) | ( n27719 & ~n27723 ) ;
  assign n27725 = n27700 | n27724 ;
  assign n27726 = ~n27720 & n27725 ;
  assign n27727 = n27143 & ~n27167 ;
  assign n27728 = ( n27143 & ~n27144 ) | ( n27143 & n27727 ) | ( ~n27144 & n27727 ) ;
  assign n27729 = ( n27569 & n27726 ) | ( n27569 & ~n27728 ) | ( n27726 & ~n27728 ) ;
  assign n27730 = ( ~n27726 & n27728 ) | ( ~n27726 & n27729 ) | ( n27728 & n27729 ) ;
  assign n27731 = ( ~n27569 & n27729 ) | ( ~n27569 & n27730 ) | ( n27729 & n27730 ) ;
  assign n27732 = n27173 & n27731 ;
  assign n27733 = ( n27196 & n27731 ) | ( n27196 & n27732 ) | ( n27731 & n27732 ) ;
  assign n27734 = n27173 | n27731 ;
  assign n27735 = n27196 | n27734 ;
  assign n27736 = ~n27733 & n27735 ;
  assign n27737 = x105 & n7566 ;
  assign n27738 = x104 & n7561 ;
  assign n27739 = x103 & ~n7560 ;
  assign n27740 = n7953 & n27739 ;
  assign n27741 = n27738 | n27740 ;
  assign n27742 = n27737 | n27741 ;
  assign n27743 = n7569 | n27737 ;
  assign n27744 = n27741 | n27743 ;
  assign n27745 = ( n8273 & n27742 ) | ( n8273 & n27744 ) | ( n27742 & n27744 ) ;
  assign n27746 = x41 & n27744 ;
  assign n27747 = x41 & n27737 ;
  assign n27748 = ( x41 & n27741 ) | ( x41 & n27747 ) | ( n27741 & n27747 ) ;
  assign n27749 = ( n8273 & n27746 ) | ( n8273 & n27748 ) | ( n27746 & n27748 ) ;
  assign n27750 = x41 & ~n27748 ;
  assign n27751 = x41 & ~n27744 ;
  assign n27752 = ( ~n8273 & n27750 ) | ( ~n8273 & n27751 ) | ( n27750 & n27751 ) ;
  assign n27753 = ( n27745 & ~n27749 ) | ( n27745 & n27752 ) | ( ~n27749 & n27752 ) ;
  assign n27754 = n27736 & n27753 ;
  assign n27755 = n27736 | n27753 ;
  assign n27756 = ~n27754 & n27755 ;
  assign n27757 = n27197 & n27216 ;
  assign n27758 = n27216 & ~n27757 ;
  assign n27759 = n27197 & ~n27216 ;
  assign n27760 = n27214 & n27759 ;
  assign n27761 = ( n27214 & n27758 ) | ( n27214 & n27760 ) | ( n27758 & n27760 ) ;
  assign n27762 = n27756 & n27757 ;
  assign n27763 = ( n27756 & n27761 ) | ( n27756 & n27762 ) | ( n27761 & n27762 ) ;
  assign n27764 = n27756 | n27757 ;
  assign n27765 = n27761 | n27764 ;
  assign n27766 = ~n27763 & n27765 ;
  assign n27767 = x108 & n6536 ;
  assign n27768 = x107 & n6531 ;
  assign n27769 = x106 & ~n6530 ;
  assign n27770 = n6871 & n27769 ;
  assign n27771 = n27768 | n27770 ;
  assign n27772 = n27767 | n27771 ;
  assign n27773 = n6539 | n27767 ;
  assign n27774 = n27771 | n27773 ;
  assign n27775 = ( n9479 & n27772 ) | ( n9479 & n27774 ) | ( n27772 & n27774 ) ;
  assign n27776 = x38 & n27774 ;
  assign n27777 = x38 & n27767 ;
  assign n27778 = ( x38 & n27771 ) | ( x38 & n27777 ) | ( n27771 & n27777 ) ;
  assign n27779 = ( n9479 & n27776 ) | ( n9479 & n27778 ) | ( n27776 & n27778 ) ;
  assign n27780 = x38 & ~n27778 ;
  assign n27781 = x38 & ~n27774 ;
  assign n27782 = ( ~n9479 & n27780 ) | ( ~n9479 & n27781 ) | ( n27780 & n27781 ) ;
  assign n27783 = ( n27775 & ~n27779 ) | ( n27775 & n27782 ) | ( ~n27779 & n27782 ) ;
  assign n27784 = n27766 & n27783 ;
  assign n27785 = n27766 | n27783 ;
  assign n27786 = ~n27784 & n27785 ;
  assign n27787 = n27221 | n27239 ;
  assign n27788 = ( n27221 & n27222 ) | ( n27221 & n27787 ) | ( n27222 & n27787 ) ;
  assign n27789 = n27786 & n27788 ;
  assign n27790 = n27786 | n27788 ;
  assign n27791 = ~n27789 & n27790 ;
  assign n27792 = x111 & n5554 ;
  assign n27793 = x110 & n5549 ;
  assign n27794 = x109 & ~n5548 ;
  assign n27795 = n5893 & n27794 ;
  assign n27796 = n27793 | n27795 ;
  assign n27797 = n27792 | n27796 ;
  assign n27798 = n5557 | n27792 ;
  assign n27799 = n27796 | n27798 ;
  assign n27800 = ( n10749 & n27797 ) | ( n10749 & n27799 ) | ( n27797 & n27799 ) ;
  assign n27801 = x35 & n27799 ;
  assign n27802 = x35 & n27792 ;
  assign n27803 = ( x35 & n27796 ) | ( x35 & n27802 ) | ( n27796 & n27802 ) ;
  assign n27804 = ( n10749 & n27801 ) | ( n10749 & n27803 ) | ( n27801 & n27803 ) ;
  assign n27805 = x35 & ~n27803 ;
  assign n27806 = x35 & ~n27799 ;
  assign n27807 = ( ~n10749 & n27805 ) | ( ~n10749 & n27806 ) | ( n27805 & n27806 ) ;
  assign n27808 = ( n27800 & ~n27804 ) | ( n27800 & n27807 ) | ( ~n27804 & n27807 ) ;
  assign n27809 = n27791 & ~n27808 ;
  assign n27810 = n27791 | n27808 ;
  assign n27811 = ( ~n27791 & n27809 ) | ( ~n27791 & n27810 ) | ( n27809 & n27810 ) ;
  assign n27812 = n27520 & n27811 ;
  assign n27546 = n27534 & ~n27535 ;
  assign n27548 = ~n27268 & n27546 ;
  assign n27549 = ~n27268 & n27534 ;
  assign n27550 = ( ~n26975 & n27548 ) | ( ~n26975 & n27549 ) | ( n27548 & n27549 ) ;
  assign n27813 = ( n27520 & ~n27550 ) | ( n27520 & n27811 ) | ( ~n27550 & n27811 ) ;
  assign n27547 = ( ~n26975 & n27534 ) | ( ~n26975 & n27546 ) | ( n27534 & n27546 ) ;
  assign n27814 = ( n27520 & ~n27547 ) | ( n27520 & n27811 ) | ( ~n27547 & n27811 ) ;
  assign n27815 = ( n26978 & n27813 ) | ( n26978 & n27814 ) | ( n27813 & n27814 ) ;
  assign n27816 = ( ~n27545 & n27812 ) | ( ~n27545 & n27815 ) | ( n27812 & n27815 ) ;
  assign n27551 = ( ~n26978 & n27547 ) | ( ~n26978 & n27550 ) | ( n27547 & n27550 ) ;
  assign n27552 = n27545 | n27551 ;
  assign n27817 = ( n27552 & ~n27811 ) | ( n27552 & n27816 ) | ( ~n27811 & n27816 ) ;
  assign n27818 = ( ~n27520 & n27816 ) | ( ~n27520 & n27817 ) | ( n27816 & n27817 ) ;
  assign n27819 = n27472 & n27818 ;
  assign n27498 = n27491 & ~n27492 ;
  assign n27499 = ( ~n27316 & n27491 ) | ( ~n27316 & n27498 ) | ( n27491 & n27498 ) ;
  assign n27500 = ~n27275 & n27499 ;
  assign n27501 = ( ~n27319 & n27499 ) | ( ~n27319 & n27500 ) | ( n27499 & n27500 ) ;
  assign n27820 = ( n27472 & ~n27501 ) | ( n27472 & n27818 ) | ( ~n27501 & n27818 ) ;
  assign n27821 = ( ~n27497 & n27819 ) | ( ~n27497 & n27820 ) | ( n27819 & n27820 ) ;
  assign n27502 = n27497 | n27501 ;
  assign n27822 = ( n27502 & ~n27818 ) | ( n27502 & n27821 ) | ( ~n27818 & n27821 ) ;
  assign n27823 = ( ~n27472 & n27821 ) | ( ~n27472 & n27822 ) | ( n27821 & n27822 ) ;
  assign n27824 = n27439 | n27823 ;
  assign n27825 = n27439 & n27823 ;
  assign n27826 = n27824 & ~n27825 ;
  assign n27827 = n27410 & ~n27412 ;
  assign n27828 = n27826 & n27827 ;
  assign n27829 = ( n27414 & n27826 ) | ( n27414 & n27828 ) | ( n27826 & n27828 ) ;
  assign n27830 = n27826 | n27827 ;
  assign n27831 = n27414 | n27830 ;
  assign n27832 = ~n27829 & n27831 ;
  assign n27839 = n27832 & n27838 ;
  assign n27840 = n27838 & ~n27839 ;
  assign n27841 = n27378 | n27379 ;
  assign n27842 = ( n27378 & n27383 ) | ( n27378 & n27841 ) | ( n27383 & n27841 ) ;
  assign n27843 = n27378 | n27389 ;
  assign n27844 = ( n26947 & n27378 ) | ( n26947 & n27841 ) | ( n27378 & n27841 ) ;
  assign n27845 = ( n26951 & n27843 ) | ( n26951 & n27844 ) | ( n27843 & n27844 ) ;
  assign n27846 = ( n26030 & n27842 ) | ( n26030 & n27845 ) | ( n27842 & n27845 ) ;
  assign n27847 = n27832 & ~n27838 ;
  assign n27848 = n27846 | n27847 ;
  assign n27849 = n27840 | n27848 ;
  assign n27850 = n27840 | n27847 ;
  assign n27851 = n27378 & n27850 ;
  assign n27852 = ( n27379 & n27850 ) | ( n27379 & n27851 ) | ( n27850 & n27851 ) ;
  assign n27853 = ( n27383 & n27851 ) | ( n27383 & n27852 ) | ( n27851 & n27852 ) ;
  assign n27854 = n27844 & n27850 ;
  assign n27855 = ( n27389 & n27850 ) | ( n27389 & n27851 ) | ( n27850 & n27851 ) ;
  assign n27856 = ( n26951 & n27854 ) | ( n26951 & n27855 ) | ( n27854 & n27855 ) ;
  assign n27857 = ( n26030 & n27853 ) | ( n26030 & n27856 ) | ( n27853 & n27856 ) ;
  assign n27858 = n27849 & ~n27857 ;
  assign n27859 = n27413 | n27829 ;
  assign n27860 = x127 & n1859 ;
  assign n27861 = x126 & n1854 ;
  assign n27862 = x125 & ~n1853 ;
  assign n27863 = n2037 & n27862 ;
  assign n27864 = n27861 | n27863 ;
  assign n27865 = n27860 | n27864 ;
  assign n27866 = n1862 | n27860 ;
  assign n27867 = n27864 | n27866 ;
  assign n27868 = ( n18763 & n27865 ) | ( n18763 & n27867 ) | ( n27865 & n27867 ) ;
  assign n27869 = x20 & n27867 ;
  assign n27870 = x20 & n27860 ;
  assign n27871 = ( x20 & n27864 ) | ( x20 & n27870 ) | ( n27864 & n27870 ) ;
  assign n27872 = ( n18763 & n27869 ) | ( n18763 & n27871 ) | ( n27869 & n27871 ) ;
  assign n27873 = x20 & ~n27871 ;
  assign n27874 = x20 & ~n27867 ;
  assign n27875 = ( ~n18763 & n27873 ) | ( ~n18763 & n27874 ) | ( n27873 & n27874 ) ;
  assign n27876 = ( n27868 & ~n27872 ) | ( n27868 & n27875 ) | ( ~n27872 & n27875 ) ;
  assign n27877 = n27472 | n27818 ;
  assign n27878 = n27501 & n27877 ;
  assign n27879 = ( n27497 & n27877 ) | ( n27497 & n27878 ) | ( n27877 & n27878 ) ;
  assign n27880 = x124 & n2429 ;
  assign n27881 = x123 & n2424 ;
  assign n27882 = x122 & ~n2423 ;
  assign n27883 = n2631 & n27882 ;
  assign n27884 = n27881 | n27883 ;
  assign n27885 = n27880 | n27884 ;
  assign n27886 = n2432 | n27880 ;
  assign n27887 = n27884 | n27886 ;
  assign n27888 = ( n17084 & n27885 ) | ( n17084 & n27887 ) | ( n27885 & n27887 ) ;
  assign n27889 = x23 & n27887 ;
  assign n27890 = x23 & n27880 ;
  assign n27891 = ( x23 & n27884 ) | ( x23 & n27890 ) | ( n27884 & n27890 ) ;
  assign n27892 = ( n17084 & n27889 ) | ( n17084 & n27891 ) | ( n27889 & n27891 ) ;
  assign n27893 = x23 & ~n27891 ;
  assign n27894 = x23 & ~n27887 ;
  assign n27895 = ( ~n17084 & n27893 ) | ( ~n17084 & n27894 ) | ( n27893 & n27894 ) ;
  assign n27896 = ( n27888 & ~n27892 ) | ( n27888 & n27895 ) | ( ~n27892 & n27895 ) ;
  assign n27897 = n27496 & n27896 ;
  assign n27898 = ~n27819 & n27896 ;
  assign n27899 = ( n27496 & n27896 ) | ( n27496 & n27898 ) | ( n27896 & n27898 ) ;
  assign n27900 = ( n27879 & n27897 ) | ( n27879 & n27899 ) | ( n27897 & n27899 ) ;
  assign n27901 = n27496 | n27896 ;
  assign n27902 = n27819 & ~n27896 ;
  assign n27903 = ~n27496 & n27902 ;
  assign n27904 = ( n27879 & n27901 ) | ( n27879 & ~n27903 ) | ( n27901 & ~n27903 ) ;
  assign n27905 = ~n27900 & n27904 ;
  assign n27906 = x121 & n3085 ;
  assign n27907 = x120 & n3080 ;
  assign n27908 = x119 & ~n3079 ;
  assign n27909 = n3309 & n27908 ;
  assign n27910 = n27907 | n27909 ;
  assign n27911 = n27906 | n27910 ;
  assign n27912 = n3088 | n27906 ;
  assign n27913 = n27910 | n27912 ;
  assign n27914 = ( n15501 & n27911 ) | ( n15501 & n27913 ) | ( n27911 & n27913 ) ;
  assign n27915 = x26 & n27913 ;
  assign n27916 = x26 & n27906 ;
  assign n27917 = ( x26 & n27910 ) | ( x26 & n27916 ) | ( n27910 & n27916 ) ;
  assign n27918 = ( n15501 & n27915 ) | ( n15501 & n27917 ) | ( n27915 & n27917 ) ;
  assign n27919 = x26 & ~n27917 ;
  assign n27920 = x26 & ~n27913 ;
  assign n27921 = ( ~n15501 & n27919 ) | ( ~n15501 & n27920 ) | ( n27919 & n27920 ) ;
  assign n27922 = ( n27914 & ~n27918 ) | ( n27914 & n27921 ) | ( ~n27918 & n27921 ) ;
  assign n27923 = n27468 | n27818 ;
  assign n27924 = ( n27468 & n27472 ) | ( n27468 & n27923 ) | ( n27472 & n27923 ) ;
  assign n27925 = n27922 & n27924 ;
  assign n27926 = n27922 | n27924 ;
  assign n27927 = ~n27925 & n27926 ;
  assign n27928 = n27520 | n27811 ;
  assign n27929 = n27550 & n27928 ;
  assign n27930 = n27547 & n27928 ;
  assign n27931 = ( ~n26978 & n27929 ) | ( ~n26978 & n27930 ) | ( n27929 & n27930 ) ;
  assign n27932 = ( n27545 & n27928 ) | ( n27545 & n27931 ) | ( n27928 & n27931 ) ;
  assign n27933 = x118 & n3816 ;
  assign n27934 = x117 & n3811 ;
  assign n27935 = x116 & ~n3810 ;
  assign n27936 = n4067 & n27935 ;
  assign n27937 = n27934 | n27936 ;
  assign n27938 = n27933 | n27937 ;
  assign n27939 = n3819 | n27933 ;
  assign n27940 = n27937 | n27939 ;
  assign n27941 = ( ~n14002 & n27938 ) | ( ~n14002 & n27940 ) | ( n27938 & n27940 ) ;
  assign n27942 = n27938 & n27940 ;
  assign n27943 = ( n13981 & n27941 ) | ( n13981 & n27942 ) | ( n27941 & n27942 ) ;
  assign n27944 = x29 & n27943 ;
  assign n27945 = x29 & ~n27943 ;
  assign n27946 = ( n27943 & ~n27944 ) | ( n27943 & n27945 ) | ( ~n27944 & n27945 ) ;
  assign n27947 = ~n27540 & n27812 ;
  assign n27948 = ~n27538 & n27812 ;
  assign n27949 = ( ~n26978 & n27947 ) | ( ~n26978 & n27948 ) | ( n27947 & n27948 ) ;
  assign n27950 = n27946 & ~n27949 ;
  assign n27951 = n27540 & n27946 ;
  assign n27952 = n27538 & n27946 ;
  assign n27953 = ( n26978 & n27951 ) | ( n26978 & n27952 ) | ( n27951 & n27952 ) ;
  assign n27954 = ( n27932 & n27950 ) | ( n27932 & n27953 ) | ( n27950 & n27953 ) ;
  assign n27955 = ~n27946 & n27949 ;
  assign n27956 = n27540 | n27946 ;
  assign n27957 = n27538 | n27946 ;
  assign n27958 = ( n26978 & n27956 ) | ( n26978 & n27957 ) | ( n27956 & n27957 ) ;
  assign n27959 = ( n27932 & ~n27955 ) | ( n27932 & n27958 ) | ( ~n27955 & n27958 ) ;
  assign n27960 = ~n27954 & n27959 ;
  assign n27961 = x115 & n4631 ;
  assign n27962 = x114 & n4626 ;
  assign n27963 = x113 & ~n4625 ;
  assign n27964 = n4943 & n27963 ;
  assign n27965 = n27962 | n27964 ;
  assign n27966 = n27961 | n27965 ;
  assign n27967 = n4634 | n27961 ;
  assign n27968 = n27965 | n27967 ;
  assign n27969 = ( ~n12550 & n27966 ) | ( ~n12550 & n27968 ) | ( n27966 & n27968 ) ;
  assign n27970 = n27966 & n27968 ;
  assign n27971 = ( n12532 & n27969 ) | ( n12532 & n27970 ) | ( n27969 & n27970 ) ;
  assign n27972 = x32 & n27971 ;
  assign n27973 = x32 & ~n27971 ;
  assign n27974 = ( n27971 & ~n27972 ) | ( n27971 & n27973 ) | ( ~n27972 & n27973 ) ;
  assign n27975 = n27519 | n27811 ;
  assign n27976 = ( n27519 & n27520 ) | ( n27519 & n27975 ) | ( n27520 & n27975 ) ;
  assign n27977 = n27974 & n27976 ;
  assign n27978 = n27974 | n27976 ;
  assign n27979 = ~n27977 & n27978 ;
  assign n27980 = x88 & n15552 ;
  assign n27981 = x87 & n15547 ;
  assign n27982 = x86 & ~n15546 ;
  assign n27983 = n16123 & n27982 ;
  assign n27984 = n27981 | n27983 ;
  assign n27985 = n27980 | n27984 ;
  assign n27986 = n15555 | n27980 ;
  assign n27987 = n27984 | n27986 ;
  assign n27988 = ( ~n3039 & n27985 ) | ( ~n3039 & n27987 ) | ( n27985 & n27987 ) ;
  assign n27989 = n27985 & n27987 ;
  assign n27990 = ( n3023 & n27988 ) | ( n3023 & n27989 ) | ( n27988 & n27989 ) ;
  assign n27991 = x59 & n27987 ;
  assign n27992 = x59 & n27980 ;
  assign n27993 = ( x59 & n27984 ) | ( x59 & n27992 ) | ( n27984 & n27992 ) ;
  assign n27994 = ( ~n3039 & n27991 ) | ( ~n3039 & n27993 ) | ( n27991 & n27993 ) ;
  assign n27995 = n27991 & n27993 ;
  assign n27996 = ( n3023 & n27994 ) | ( n3023 & n27995 ) | ( n27994 & n27995 ) ;
  assign n27997 = x59 & ~n27993 ;
  assign n27998 = x59 & ~n27987 ;
  assign n27999 = ( n3039 & n27997 ) | ( n3039 & n27998 ) | ( n27997 & n27998 ) ;
  assign n28000 = n27997 | n27998 ;
  assign n28001 = ( ~n3023 & n27999 ) | ( ~n3023 & n28000 ) | ( n27999 & n28000 ) ;
  assign n28002 = ( n27990 & ~n27996 ) | ( n27990 & n28001 ) | ( ~n27996 & n28001 ) ;
  assign n28003 = x84 & n17141 ;
  assign n28004 = x83 & ~n17140 ;
  assign n28005 = n17724 & n28004 ;
  assign n28006 = n28003 | n28005 ;
  assign n28007 = x85 & n17146 ;
  assign n28008 = n17149 | n28007 ;
  assign n28009 = n28006 | n28008 ;
  assign n28010 = ~x62 & n28009 ;
  assign n28011 = ~x62 & n28007 ;
  assign n28012 = ( ~x62 & n28006 ) | ( ~x62 & n28011 ) | ( n28006 & n28011 ) ;
  assign n28013 = ( n2381 & n28010 ) | ( n2381 & n28012 ) | ( n28010 & n28012 ) ;
  assign n28014 = x62 & ~n28009 ;
  assign n28015 = x62 & x85 ;
  assign n28016 = n17146 & n28015 ;
  assign n28017 = x62 & ~n28016 ;
  assign n28018 = ~n28006 & n28017 ;
  assign n28019 = ( ~n2381 & n28014 ) | ( ~n2381 & n28018 ) | ( n28014 & n28018 ) ;
  assign n28020 = n28013 | n28019 ;
  assign n28021 = x82 & n18290 ;
  assign n28022 = x63 & x81 ;
  assign n28023 = ~n18290 & n28022 ;
  assign n28024 = n28021 | n28023 ;
  assign n28025 = ~x17 & n28024 ;
  assign n28026 = x17 & ~n28024 ;
  assign n28027 = n28025 | n28026 ;
  assign n28028 = n27608 & ~n28027 ;
  assign n28029 = ~n27608 & n28027 ;
  assign n28030 = n28028 | n28029 ;
  assign n28031 = n28020 & ~n28030 ;
  assign n28032 = ~n28020 & n28030 ;
  assign n28033 = n28031 | n28032 ;
  assign n28034 = n27609 & ~n27610 ;
  assign n28035 = n27610 & ~n28034 ;
  assign n28036 = ( n27604 & ~n28034 ) | ( n27604 & n28035 ) | ( ~n28034 & n28035 ) ;
  assign n28037 = n28033 | n28036 ;
  assign n28038 = n28002 & n28036 ;
  assign n28039 = n28033 & n28038 ;
  assign n28040 = ( n28002 & ~n28037 ) | ( n28002 & n28039 ) | ( ~n28037 & n28039 ) ;
  assign n28041 = n28002 | n28036 ;
  assign n28042 = ( n28002 & n28033 ) | ( n28002 & n28041 ) | ( n28033 & n28041 ) ;
  assign n28043 = n28037 & ~n28042 ;
  assign n28044 = n28040 | n28043 ;
  assign n28045 = n27618 | n27638 ;
  assign n28046 = ( n27618 & ~n27621 ) | ( n27618 & n28045 ) | ( ~n27621 & n28045 ) ;
  assign n28047 = ~n28044 & n28046 ;
  assign n28048 = n28044 & ~n28046 ;
  assign n28049 = n28047 | n28048 ;
  assign n28050 = x91 & n14045 ;
  assign n28051 = x90 & n14040 ;
  assign n28052 = x89 & ~n14039 ;
  assign n28053 = n14552 & n28052 ;
  assign n28054 = n28051 | n28053 ;
  assign n28055 = n28050 | n28054 ;
  assign n28056 = n14048 | n28050 ;
  assign n28057 = n28054 | n28056 ;
  assign n28058 = ( n3768 & n28055 ) | ( n3768 & n28057 ) | ( n28055 & n28057 ) ;
  assign n28059 = x56 & n28057 ;
  assign n28060 = x56 & n28050 ;
  assign n28061 = ( x56 & n28054 ) | ( x56 & n28060 ) | ( n28054 & n28060 ) ;
  assign n28062 = ( n3768 & n28059 ) | ( n3768 & n28061 ) | ( n28059 & n28061 ) ;
  assign n28063 = x56 & ~n28061 ;
  assign n28064 = x56 & ~n28057 ;
  assign n28065 = ( ~n3768 & n28063 ) | ( ~n3768 & n28064 ) | ( n28063 & n28064 ) ;
  assign n28066 = ( n28058 & ~n28062 ) | ( n28058 & n28065 ) | ( ~n28062 & n28065 ) ;
  assign n28067 = ~n28049 & n28066 ;
  assign n28068 = n28049 | n28067 ;
  assign n28070 = n27645 | n27664 ;
  assign n28071 = ( n27645 & ~n27647 ) | ( n27645 & n28070 ) | ( ~n27647 & n28070 ) ;
  assign n28069 = n28049 & n28066 ;
  assign n28072 = n28069 & n28071 ;
  assign n28073 = ( ~n28068 & n28071 ) | ( ~n28068 & n28072 ) | ( n28071 & n28072 ) ;
  assign n28074 = n28069 | n28071 ;
  assign n28075 = n28068 & ~n28074 ;
  assign n28076 = n28073 | n28075 ;
  assign n28077 = x94 & n12574 ;
  assign n28078 = x93 & n12569 ;
  assign n28079 = x92 & ~n12568 ;
  assign n28080 = n13076 & n28079 ;
  assign n28081 = n28078 | n28080 ;
  assign n28082 = n28077 | n28081 ;
  assign n28083 = n12577 | n28077 ;
  assign n28084 = n28081 | n28083 ;
  assign n28085 = ( n4583 & n28082 ) | ( n4583 & n28084 ) | ( n28082 & n28084 ) ;
  assign n28086 = x53 & n28084 ;
  assign n28087 = x53 & n28077 ;
  assign n28088 = ( x53 & n28081 ) | ( x53 & n28087 ) | ( n28081 & n28087 ) ;
  assign n28089 = ( n4583 & n28086 ) | ( n4583 & n28088 ) | ( n28086 & n28088 ) ;
  assign n28090 = x53 & ~n28088 ;
  assign n28091 = x53 & ~n28084 ;
  assign n28092 = ( ~n4583 & n28090 ) | ( ~n4583 & n28091 ) | ( n28090 & n28091 ) ;
  assign n28093 = ( n28085 & ~n28089 ) | ( n28085 & n28092 ) | ( ~n28089 & n28092 ) ;
  assign n28094 = ~n28076 & n28093 ;
  assign n28095 = n28076 | n28094 ;
  assign n28097 = n27667 & ~n27688 ;
  assign n28098 = ( n27668 & n27688 ) | ( n27668 & ~n28097 ) | ( n27688 & ~n28097 ) ;
  assign n28099 = ( n27669 & ~n27671 ) | ( n27669 & n28098 ) | ( ~n27671 & n28098 ) ;
  assign n28096 = n28076 & n28093 ;
  assign n28100 = n28096 & n28099 ;
  assign n28101 = ( ~n28095 & n28099 ) | ( ~n28095 & n28100 ) | ( n28099 & n28100 ) ;
  assign n28102 = n28096 | n28099 ;
  assign n28103 = n28095 & ~n28102 ;
  assign n28104 = n28101 | n28103 ;
  assign n28105 = ~n27691 & n27693 ;
  assign n28106 = n27691 | n28105 ;
  assign n28107 = x97 & n11205 ;
  assign n28108 = x96 & n11200 ;
  assign n28109 = x95 & ~n11199 ;
  assign n28110 = n11679 & n28109 ;
  assign n28111 = n28108 | n28110 ;
  assign n28112 = n28107 | n28111 ;
  assign n28113 = n11208 | n28107 ;
  assign n28114 = n28111 | n28113 ;
  assign n28115 = ( n5505 & n28112 ) | ( n5505 & n28114 ) | ( n28112 & n28114 ) ;
  assign n28116 = x50 & n28114 ;
  assign n28117 = x50 & n28107 ;
  assign n28118 = ( x50 & n28111 ) | ( x50 & n28117 ) | ( n28111 & n28117 ) ;
  assign n28119 = ( n5505 & n28116 ) | ( n5505 & n28118 ) | ( n28116 & n28118 ) ;
  assign n28120 = x50 & ~n28118 ;
  assign n28121 = x50 & ~n28114 ;
  assign n28122 = ( ~n5505 & n28120 ) | ( ~n5505 & n28121 ) | ( n28120 & n28121 ) ;
  assign n28123 = ( n28115 & ~n28119 ) | ( n28115 & n28122 ) | ( ~n28119 & n28122 ) ;
  assign n28124 = n27008 & n27586 ;
  assign n28125 = n27109 & n27586 ;
  assign n28126 = ( ~n27692 & n28124 ) | ( ~n27692 & n28125 ) | ( n28124 & n28125 ) ;
  assign n28127 = n27691 & n28126 ;
  assign n28128 = n27008 & n28123 ;
  assign n28129 = n27109 & n28123 ;
  assign n28130 = ( ~n27692 & n28128 ) | ( ~n27692 & n28129 ) | ( n28128 & n28129 ) ;
  assign n28131 = ~n27691 & n28130 ;
  assign n28132 = ( n28123 & n28127 ) | ( n28123 & n28131 ) | ( n28127 & n28131 ) ;
  assign n28133 = ( n27586 & n28123 ) | ( n27586 & n28130 ) | ( n28123 & n28130 ) ;
  assign n28134 = n27586 & n28123 ;
  assign n28135 = ( ~n27691 & n28133 ) | ( ~n27691 & n28134 ) | ( n28133 & n28134 ) ;
  assign n28136 = ( ~n28106 & n28132 ) | ( ~n28106 & n28135 ) | ( n28132 & n28135 ) ;
  assign n28137 = n27008 | n28123 ;
  assign n28138 = n27109 | n28123 ;
  assign n28139 = ( ~n27692 & n28137 ) | ( ~n27692 & n28138 ) | ( n28137 & n28138 ) ;
  assign n28140 = ( ~n27691 & n28123 ) | ( ~n27691 & n28139 ) | ( n28123 & n28139 ) ;
  assign n28141 = n28127 | n28140 ;
  assign n28142 = n27586 | n28139 ;
  assign n28143 = n27586 | n28123 ;
  assign n28144 = ( ~n27691 & n28142 ) | ( ~n27691 & n28143 ) | ( n28142 & n28143 ) ;
  assign n28145 = ( ~n28106 & n28141 ) | ( ~n28106 & n28144 ) | ( n28141 & n28144 ) ;
  assign n28146 = ~n28136 & n28145 ;
  assign n28147 = n28104 & n28146 ;
  assign n28148 = n28104 | n28146 ;
  assign n28149 = ~n28147 & n28148 ;
  assign n28150 = x100 & n9933 ;
  assign n28151 = x99 & n9928 ;
  assign n28152 = x98 & ~n9927 ;
  assign n28153 = n10379 & n28152 ;
  assign n28154 = n28151 | n28153 ;
  assign n28155 = n28150 | n28154 ;
  assign n28156 = n9936 | n28150 ;
  assign n28157 = n28154 | n28156 ;
  assign n28158 = ( n6483 & n28155 ) | ( n6483 & n28157 ) | ( n28155 & n28157 ) ;
  assign n28159 = x47 & n28157 ;
  assign n28160 = x47 & n28150 ;
  assign n28161 = ( x47 & n28154 ) | ( x47 & n28160 ) | ( n28154 & n28160 ) ;
  assign n28162 = ( n6483 & n28159 ) | ( n6483 & n28161 ) | ( n28159 & n28161 ) ;
  assign n28163 = x47 & ~n28161 ;
  assign n28164 = x47 & ~n28157 ;
  assign n28165 = ( ~n6483 & n28163 ) | ( ~n6483 & n28164 ) | ( n28163 & n28164 ) ;
  assign n28166 = ( n28158 & ~n28162 ) | ( n28158 & n28165 ) | ( ~n28162 & n28165 ) ;
  assign n28167 = ~n28149 & n28166 ;
  assign n28168 = n28149 & ~n28166 ;
  assign n28169 = n28167 | n28168 ;
  assign n28170 = ( n27701 & ~n27702 ) | ( n27701 & n27724 ) | ( ~n27702 & n27724 ) ;
  assign n28171 = n28169 & ~n28170 ;
  assign n28172 = ~n28169 & n28170 ;
  assign n28173 = n28171 | n28172 ;
  assign n28174 = x103 & n8724 ;
  assign n28175 = x102 & n8719 ;
  assign n28176 = x101 & ~n8718 ;
  assign n28177 = n9149 & n28176 ;
  assign n28178 = n28175 | n28177 ;
  assign n28179 = n28174 | n28178 ;
  assign n28180 = n8727 | n28174 ;
  assign n28181 = n28178 | n28180 ;
  assign n28182 = ( n7529 & n28179 ) | ( n7529 & n28181 ) | ( n28179 & n28181 ) ;
  assign n28183 = x44 & n28181 ;
  assign n28184 = x44 & n28174 ;
  assign n28185 = ( x44 & n28178 ) | ( x44 & n28184 ) | ( n28178 & n28184 ) ;
  assign n28186 = ( n7529 & n28183 ) | ( n7529 & n28185 ) | ( n28183 & n28185 ) ;
  assign n28187 = x44 & ~n28185 ;
  assign n28188 = x44 & ~n28181 ;
  assign n28189 = ( ~n7529 & n28187 ) | ( ~n7529 & n28188 ) | ( n28187 & n28188 ) ;
  assign n28190 = ( n28182 & ~n28186 ) | ( n28182 & n28189 ) | ( ~n28186 & n28189 ) ;
  assign n28191 = ~n28173 & n28190 ;
  assign n28192 = n28173 | n28191 ;
  assign n28193 = n28173 & n28190 ;
  assign n28194 = n28192 & ~n28193 ;
  assign n28195 = n27726 | n27728 ;
  assign n28196 = ~n27726 & n28195 ;
  assign n28197 = n27726 & ~n27728 ;
  assign n28198 = n27569 & ~n28197 ;
  assign n28199 = ~n28196 & n28198 ;
  assign n28200 = ( ~n27569 & n28195 ) | ( ~n27569 & n28199 ) | ( n28195 & n28199 ) ;
  assign n28201 = n28194 & ~n28200 ;
  assign n28202 = ~n28194 & n28200 ;
  assign n28203 = n28201 | n28202 ;
  assign n28204 = x106 & n7566 ;
  assign n28205 = x105 & n7561 ;
  assign n28206 = x104 & ~n7560 ;
  assign n28207 = n7953 & n28206 ;
  assign n28208 = n28205 | n28207 ;
  assign n28209 = n28204 | n28208 ;
  assign n28210 = n7569 | n28204 ;
  assign n28211 = n28208 | n28210 ;
  assign n28212 = ( n8656 & n28209 ) | ( n8656 & n28211 ) | ( n28209 & n28211 ) ;
  assign n28213 = x41 & n28211 ;
  assign n28214 = x41 & n28204 ;
  assign n28215 = ( x41 & n28208 ) | ( x41 & n28214 ) | ( n28208 & n28214 ) ;
  assign n28216 = ( n8656 & n28213 ) | ( n8656 & n28215 ) | ( n28213 & n28215 ) ;
  assign n28217 = x41 & ~n28215 ;
  assign n28218 = x41 & ~n28211 ;
  assign n28219 = ( ~n8656 & n28217 ) | ( ~n8656 & n28218 ) | ( n28217 & n28218 ) ;
  assign n28220 = ( n28212 & ~n28216 ) | ( n28212 & n28219 ) | ( ~n28216 & n28219 ) ;
  assign n28221 = n28203 & n28220 ;
  assign n28222 = n28203 | n28220 ;
  assign n28223 = ~n28221 & n28222 ;
  assign n28224 = n27733 | n27753 ;
  assign n28225 = ( n27733 & n27736 ) | ( n27733 & n28224 ) | ( n27736 & n28224 ) ;
  assign n28226 = n28223 | n28225 ;
  assign n28227 = n28223 & n28225 ;
  assign n28228 = n28226 & ~n28227 ;
  assign n28229 = x109 & n6536 ;
  assign n28230 = x108 & n6531 ;
  assign n28231 = x107 & ~n6530 ;
  assign n28232 = n6871 & n28231 ;
  assign n28233 = n28230 | n28232 ;
  assign n28234 = n28229 | n28233 ;
  assign n28235 = n6539 | n28229 ;
  assign n28236 = n28233 | n28235 ;
  assign n28237 = ( n9878 & n28234 ) | ( n9878 & n28236 ) | ( n28234 & n28236 ) ;
  assign n28238 = x38 & n28236 ;
  assign n28239 = x38 & n28229 ;
  assign n28240 = ( x38 & n28233 ) | ( x38 & n28239 ) | ( n28233 & n28239 ) ;
  assign n28241 = ( n9878 & n28238 ) | ( n9878 & n28240 ) | ( n28238 & n28240 ) ;
  assign n28242 = x38 & ~n28240 ;
  assign n28243 = x38 & ~n28236 ;
  assign n28244 = ( ~n9878 & n28242 ) | ( ~n9878 & n28243 ) | ( n28242 & n28243 ) ;
  assign n28245 = ( n28237 & ~n28241 ) | ( n28237 & n28244 ) | ( ~n28241 & n28244 ) ;
  assign n28246 = n28228 & n28245 ;
  assign n28247 = n28228 & ~n28246 ;
  assign n28249 = n27763 | n27783 ;
  assign n28250 = ( n27763 & n27766 ) | ( n27763 & n28249 ) | ( n27766 & n28249 ) ;
  assign n28248 = ~n28228 & n28245 ;
  assign n28251 = n28248 & n28250 ;
  assign n28252 = ( n28247 & n28250 ) | ( n28247 & n28251 ) | ( n28250 & n28251 ) ;
  assign n28253 = n28248 | n28250 ;
  assign n28254 = n28247 | n28253 ;
  assign n28255 = ~n28252 & n28254 ;
  assign n28256 = x112 & n5554 ;
  assign n28257 = x111 & n5549 ;
  assign n28258 = x110 & ~n5548 ;
  assign n28259 = n5893 & n28258 ;
  assign n28260 = n28257 | n28259 ;
  assign n28261 = n28256 | n28260 ;
  assign n28262 = n5557 | n28256 ;
  assign n28263 = n28260 | n28262 ;
  assign n28264 = ( n11172 & n28261 ) | ( n11172 & n28263 ) | ( n28261 & n28263 ) ;
  assign n28265 = x35 & n28263 ;
  assign n28266 = x35 & n28256 ;
  assign n28267 = ( x35 & n28260 ) | ( x35 & n28266 ) | ( n28260 & n28266 ) ;
  assign n28268 = ( n11172 & n28265 ) | ( n11172 & n28267 ) | ( n28265 & n28267 ) ;
  assign n28269 = x35 & ~n28267 ;
  assign n28270 = x35 & ~n28263 ;
  assign n28271 = ( ~n11172 & n28269 ) | ( ~n11172 & n28270 ) | ( n28269 & n28270 ) ;
  assign n28272 = ( n28264 & ~n28268 ) | ( n28264 & n28271 ) | ( ~n28268 & n28271 ) ;
  assign n28273 = n28255 & n28272 ;
  assign n28274 = n28255 & ~n28273 ;
  assign n28276 = n27788 | n27808 ;
  assign n28277 = ( n27786 & n27808 ) | ( n27786 & n28276 ) | ( n27808 & n28276 ) ;
  assign n28278 = ( n27789 & n27791 ) | ( n27789 & n28277 ) | ( n27791 & n28277 ) ;
  assign n28275 = ~n28255 & n28272 ;
  assign n28279 = n28275 & n28278 ;
  assign n28280 = ( n28274 & n28278 ) | ( n28274 & n28279 ) | ( n28278 & n28279 ) ;
  assign n28281 = n28275 | n28278 ;
  assign n28282 = n28274 | n28281 ;
  assign n28283 = ~n28280 & n28282 ;
  assign n28284 = ~n27979 & n28283 ;
  assign n28285 = n27979 & ~n28283 ;
  assign n28286 = n28284 | n28285 ;
  assign n28287 = n27960 & n28286 ;
  assign n28288 = n27960 & ~n28287 ;
  assign n28289 = ~n27960 & n28286 ;
  assign n28290 = n28288 | n28289 ;
  assign n28291 = ~n27927 & n28290 ;
  assign n28292 = n27927 & ~n28290 ;
  assign n28293 = n28291 | n28292 ;
  assign n28294 = n27905 & ~n28293 ;
  assign n28295 = n27905 | n28293 ;
  assign n28296 = ( ~n27905 & n28294 ) | ( ~n27905 & n28295 ) | ( n28294 & n28295 ) ;
  assign n28297 = n27438 | n27823 ;
  assign n28298 = ( n27438 & n27439 ) | ( n27438 & n28297 ) | ( n27439 & n28297 ) ;
  assign n28299 = ( n27876 & n28296 ) | ( n27876 & ~n28298 ) | ( n28296 & ~n28298 ) ;
  assign n28300 = ( ~n28296 & n28298 ) | ( ~n28296 & n28299 ) | ( n28298 & n28299 ) ;
  assign n28301 = ( ~n27876 & n28299 ) | ( ~n27876 & n28300 ) | ( n28299 & n28300 ) ;
  assign n28302 = ~n27859 & n28301 ;
  assign n28303 = n27859 & n28301 ;
  assign n28304 = n27859 & ~n28303 ;
  assign n28305 = n28302 | n28304 ;
  assign n28306 = n27839 | n27851 ;
  assign n28307 = n27839 | n27850 ;
  assign n28308 = ( n27389 & n28306 ) | ( n27389 & n28307 ) | ( n28306 & n28307 ) ;
  assign n28309 = ( n27839 & n27844 ) | ( n27839 & n28307 ) | ( n27844 & n28307 ) ;
  assign n28310 = ( n26022 & n28308 ) | ( n26022 & n28309 ) | ( n28308 & n28309 ) ;
  assign n28311 = ( n26490 & n28308 ) | ( n26490 & n28309 ) | ( n28308 & n28309 ) ;
  assign n28312 = ( n26949 & n28310 ) | ( n26949 & n28311 ) | ( n28310 & n28311 ) ;
  assign n28313 = n28305 & n28312 ;
  assign n28314 = n27839 & n28305 ;
  assign n28315 = ( n27852 & n28305 ) | ( n27852 & n28314 ) | ( n28305 & n28314 ) ;
  assign n28316 = ( n27851 & n28305 ) | ( n27851 & n28314 ) | ( n28305 & n28314 ) ;
  assign n28317 = ( n27383 & n28315 ) | ( n27383 & n28316 ) | ( n28315 & n28316 ) ;
  assign n28318 = ( n26030 & n28313 ) | ( n26030 & n28317 ) | ( n28313 & n28317 ) ;
  assign n28319 = n27839 | n27852 ;
  assign n28320 = ( n27383 & n28306 ) | ( n27383 & n28319 ) | ( n28306 & n28319 ) ;
  assign n28321 = ( n26030 & n28312 ) | ( n26030 & n28320 ) | ( n28312 & n28320 ) ;
  assign n28322 = ( n27859 & ~n28301 ) | ( n27859 & n28321 ) | ( ~n28301 & n28321 ) ;
  assign n28323 = ( n28302 & ~n28318 ) | ( n28302 & n28322 ) | ( ~n28318 & n28322 ) ;
  assign n28338 = n27900 | n28293 ;
  assign n28339 = ( n27900 & n27905 ) | ( n27900 & n28338 ) | ( n27905 & n28338 ) ;
  assign n28324 = x127 & n1854 ;
  assign n28325 = x126 & ~n1853 ;
  assign n28326 = n2037 & n28325 ;
  assign n28327 = n28324 | n28326 ;
  assign n28328 = n1862 | n28327 ;
  assign n28329 = ( n19328 & n28327 ) | ( n19328 & n28328 ) | ( n28327 & n28328 ) ;
  assign n28330 = x20 & n28327 ;
  assign n28331 = ( x20 & n3354 ) | ( x20 & n28327 ) | ( n3354 & n28327 ) ;
  assign n28332 = ( n19328 & n28330 ) | ( n19328 & n28331 ) | ( n28330 & n28331 ) ;
  assign n28333 = x20 & ~n3354 ;
  assign n28334 = ~n28327 & n28333 ;
  assign n28335 = x20 & ~n28327 ;
  assign n28336 = ( ~n19328 & n28334 ) | ( ~n19328 & n28335 ) | ( n28334 & n28335 ) ;
  assign n28337 = ( n28329 & ~n28332 ) | ( n28329 & n28336 ) | ( ~n28332 & n28336 ) ;
  assign n28340 = n28337 & n28339 ;
  assign n28341 = n28339 & ~n28340 ;
  assign n28342 = n28337 & ~n28339 ;
  assign n28343 = x122 & n3085 ;
  assign n28344 = x121 & n3080 ;
  assign n28345 = x120 & ~n3079 ;
  assign n28346 = n3309 & n28345 ;
  assign n28347 = n28344 | n28346 ;
  assign n28348 = n28343 | n28347 ;
  assign n28349 = n3088 | n28343 ;
  assign n28350 = n28347 | n28349 ;
  assign n28351 = ( n16043 & n28348 ) | ( n16043 & n28350 ) | ( n28348 & n28350 ) ;
  assign n28352 = x26 & n28350 ;
  assign n28353 = x26 & n28343 ;
  assign n28354 = ( x26 & n28347 ) | ( x26 & n28353 ) | ( n28347 & n28353 ) ;
  assign n28355 = ( n16043 & n28352 ) | ( n16043 & n28354 ) | ( n28352 & n28354 ) ;
  assign n28356 = x26 & ~n28354 ;
  assign n28357 = x26 & ~n28350 ;
  assign n28358 = ( ~n16043 & n28356 ) | ( ~n16043 & n28357 ) | ( n28356 & n28357 ) ;
  assign n28359 = ( n28351 & ~n28355 ) | ( n28351 & n28358 ) | ( ~n28355 & n28358 ) ;
  assign n28360 = ( n27954 & n28286 ) | ( n27954 & n28359 ) | ( n28286 & n28359 ) ;
  assign n28361 = n27950 & n28359 ;
  assign n28362 = n27953 & n28359 ;
  assign n28363 = ( n27932 & n28361 ) | ( n27932 & n28362 ) | ( n28361 & n28362 ) ;
  assign n28364 = ( n27960 & n28360 ) | ( n27960 & n28363 ) | ( n28360 & n28363 ) ;
  assign n28365 = n27950 | n28359 ;
  assign n28366 = n27953 | n28359 ;
  assign n28367 = ( n27932 & n28365 ) | ( n27932 & n28366 ) | ( n28365 & n28366 ) ;
  assign n28368 = n28286 | n28367 ;
  assign n28369 = ( n27960 & n28367 ) | ( n27960 & n28368 ) | ( n28367 & n28368 ) ;
  assign n28370 = ~n28364 & n28369 ;
  assign n28371 = x83 & n18290 ;
  assign n28372 = x63 & x82 ;
  assign n28373 = ~n18290 & n28372 ;
  assign n28374 = n28371 | n28373 ;
  assign n28375 = n27608 | n28025 ;
  assign n28376 = ( n28025 & ~n28027 ) | ( n28025 & n28375 ) | ( ~n28027 & n28375 ) ;
  assign n28377 = n28374 & ~n28376 ;
  assign n28378 = ~n28374 & n28376 ;
  assign n28379 = n28377 | n28378 ;
  assign n28380 = x85 & n17141 ;
  assign n28381 = x84 & ~n17140 ;
  assign n28382 = n17724 & n28381 ;
  assign n28383 = n28380 | n28382 ;
  assign n28384 = x86 & n17146 ;
  assign n28385 = n17149 | n28384 ;
  assign n28386 = n28383 | n28385 ;
  assign n28387 = x62 & ~n28386 ;
  assign n28388 = ~n28379 & n28387 ;
  assign n28389 = x62 & x86 ;
  assign n28390 = n17146 & n28389 ;
  assign n28391 = x62 & ~n28390 ;
  assign n28392 = ~n28383 & n28391 ;
  assign n28393 = ~n28379 & n28392 ;
  assign n28394 = ( ~n2606 & n28388 ) | ( ~n2606 & n28393 ) | ( n28388 & n28393 ) ;
  assign n28395 = ~x62 & n28386 ;
  assign n28396 = ~x62 & n28384 ;
  assign n28397 = ( ~x62 & n28383 ) | ( ~x62 & n28396 ) | ( n28383 & n28396 ) ;
  assign n28398 = ( n2606 & n28395 ) | ( n2606 & n28397 ) | ( n28395 & n28397 ) ;
  assign n28399 = ( ~n28379 & n28394 ) | ( ~n28379 & n28398 ) | ( n28394 & n28398 ) ;
  assign n28400 = n28379 & ~n28387 ;
  assign n28401 = n28379 & ~n28392 ;
  assign n28402 = ( n2606 & n28400 ) | ( n2606 & n28401 ) | ( n28400 & n28401 ) ;
  assign n28403 = ~n28398 & n28402 ;
  assign n28404 = n28399 | n28403 ;
  assign n28405 = n28031 | n28036 ;
  assign n28406 = ( n28031 & ~n28033 ) | ( n28031 & n28405 ) | ( ~n28033 & n28405 ) ;
  assign n28407 = ~n28404 & n28406 ;
  assign n28408 = n28404 & ~n28406 ;
  assign n28409 = n28407 | n28408 ;
  assign n28410 = x89 & n15552 ;
  assign n28411 = x88 & n15547 ;
  assign n28412 = x87 & ~n15546 ;
  assign n28413 = n16123 & n28412 ;
  assign n28414 = n28411 | n28413 ;
  assign n28415 = n28410 | n28414 ;
  assign n28416 = n15555 | n28410 ;
  assign n28417 = n28414 | n28416 ;
  assign n28418 = ( n3282 & n28415 ) | ( n3282 & n28417 ) | ( n28415 & n28417 ) ;
  assign n28419 = x59 & n28417 ;
  assign n28420 = x59 & n28410 ;
  assign n28421 = ( x59 & n28414 ) | ( x59 & n28420 ) | ( n28414 & n28420 ) ;
  assign n28422 = ( n3282 & n28419 ) | ( n3282 & n28421 ) | ( n28419 & n28421 ) ;
  assign n28423 = x59 & ~n28421 ;
  assign n28424 = x59 & ~n28417 ;
  assign n28425 = ( ~n3282 & n28423 ) | ( ~n3282 & n28424 ) | ( n28423 & n28424 ) ;
  assign n28426 = ( n28418 & ~n28422 ) | ( n28418 & n28425 ) | ( ~n28422 & n28425 ) ;
  assign n28427 = n28409 | n28426 ;
  assign n28428 = n28409 & ~n28426 ;
  assign n28429 = ( ~n28409 & n28427 ) | ( ~n28409 & n28428 ) | ( n28427 & n28428 ) ;
  assign n28430 = n28040 | n28047 ;
  assign n28431 = n28429 & n28430 ;
  assign n28432 = n28429 | n28430 ;
  assign n28433 = ~n28431 & n28432 ;
  assign n28434 = x92 & n14045 ;
  assign n28435 = x91 & n14040 ;
  assign n28436 = x90 & ~n14039 ;
  assign n28437 = n14552 & n28436 ;
  assign n28438 = n28435 | n28437 ;
  assign n28439 = n28434 | n28438 ;
  assign n28440 = n14048 | n28434 ;
  assign n28441 = n28438 | n28440 ;
  assign n28442 = ( n4040 & n28439 ) | ( n4040 & n28441 ) | ( n28439 & n28441 ) ;
  assign n28443 = x56 & n28441 ;
  assign n28444 = x56 & n28434 ;
  assign n28445 = ( x56 & n28438 ) | ( x56 & n28444 ) | ( n28438 & n28444 ) ;
  assign n28446 = ( n4040 & n28443 ) | ( n4040 & n28445 ) | ( n28443 & n28445 ) ;
  assign n28447 = x56 & ~n28445 ;
  assign n28448 = x56 & ~n28441 ;
  assign n28449 = ( ~n4040 & n28447 ) | ( ~n4040 & n28448 ) | ( n28447 & n28448 ) ;
  assign n28450 = ( n28442 & ~n28446 ) | ( n28442 & n28449 ) | ( ~n28446 & n28449 ) ;
  assign n28451 = n28433 & ~n28450 ;
  assign n28452 = ~n28433 & n28450 ;
  assign n28453 = n28451 | n28452 ;
  assign n28454 = n28067 | n28071 ;
  assign n28455 = ~n28067 & n28068 ;
  assign n28456 = ( n28072 & n28454 ) | ( n28072 & ~n28455 ) | ( n28454 & ~n28455 ) ;
  assign n28457 = ~n28453 & n28456 ;
  assign n28458 = n28453 & ~n28456 ;
  assign n28459 = n28457 | n28458 ;
  assign n28460 = x95 & n12574 ;
  assign n28461 = x94 & n12569 ;
  assign n28462 = x93 & ~n12568 ;
  assign n28463 = n13076 & n28462 ;
  assign n28464 = n28461 | n28463 ;
  assign n28465 = n28460 | n28464 ;
  assign n28466 = n12577 | n28460 ;
  assign n28467 = n28464 | n28466 ;
  assign n28468 = ( n4897 & n28465 ) | ( n4897 & n28467 ) | ( n28465 & n28467 ) ;
  assign n28469 = x53 & n28467 ;
  assign n28470 = x53 & n28460 ;
  assign n28471 = ( x53 & n28464 ) | ( x53 & n28470 ) | ( n28464 & n28470 ) ;
  assign n28472 = ( n4897 & n28469 ) | ( n4897 & n28471 ) | ( n28469 & n28471 ) ;
  assign n28473 = x53 & ~n28471 ;
  assign n28474 = x53 & ~n28467 ;
  assign n28475 = ( ~n4897 & n28473 ) | ( ~n4897 & n28474 ) | ( n28473 & n28474 ) ;
  assign n28476 = ( n28468 & ~n28472 ) | ( n28468 & n28475 ) | ( ~n28472 & n28475 ) ;
  assign n28477 = n28459 | n28476 ;
  assign n28478 = n28459 & ~n28476 ;
  assign n28479 = ( ~n28459 & n28477 ) | ( ~n28459 & n28478 ) | ( n28477 & n28478 ) ;
  assign n28480 = n28094 | n28099 ;
  assign n28481 = ~n28094 & n28095 ;
  assign n28482 = ( n28100 & n28480 ) | ( n28100 & ~n28481 ) | ( n28480 & ~n28481 ) ;
  assign n28483 = n28479 & ~n28482 ;
  assign n28484 = ~n28479 & n28482 ;
  assign n28485 = n28483 | n28484 ;
  assign n28486 = x98 & n11205 ;
  assign n28487 = x97 & n11200 ;
  assign n28488 = x96 & ~n11199 ;
  assign n28489 = n11679 & n28488 ;
  assign n28490 = n28487 | n28489 ;
  assign n28491 = n28486 | n28490 ;
  assign n28492 = n11208 | n28486 ;
  assign n28493 = n28490 | n28492 ;
  assign n28494 = ( ~n5850 & n28491 ) | ( ~n5850 & n28493 ) | ( n28491 & n28493 ) ;
  assign n28495 = n28491 & n28493 ;
  assign n28496 = ( n5834 & n28494 ) | ( n5834 & n28495 ) | ( n28494 & n28495 ) ;
  assign n28497 = x50 & n28493 ;
  assign n28498 = x50 & n28486 ;
  assign n28499 = ( x50 & n28490 ) | ( x50 & n28498 ) | ( n28490 & n28498 ) ;
  assign n28500 = ( ~n5850 & n28497 ) | ( ~n5850 & n28499 ) | ( n28497 & n28499 ) ;
  assign n28501 = n28497 & n28499 ;
  assign n28502 = ( n5834 & n28500 ) | ( n5834 & n28501 ) | ( n28500 & n28501 ) ;
  assign n28503 = x50 & ~n28499 ;
  assign n28504 = x50 & ~n28493 ;
  assign n28505 = ( n5850 & n28503 ) | ( n5850 & n28504 ) | ( n28503 & n28504 ) ;
  assign n28506 = n28503 | n28504 ;
  assign n28507 = ( ~n5834 & n28505 ) | ( ~n5834 & n28506 ) | ( n28505 & n28506 ) ;
  assign n28508 = ( n28496 & ~n28502 ) | ( n28496 & n28507 ) | ( ~n28502 & n28507 ) ;
  assign n28509 = n28485 & n28508 ;
  assign n28510 = n28479 & ~n28508 ;
  assign n28511 = ( n28482 & n28508 ) | ( n28482 & ~n28510 ) | ( n28508 & ~n28510 ) ;
  assign n28512 = n28483 | n28511 ;
  assign n28513 = ~n28509 & n28512 ;
  assign n28514 = n28104 & ~n28136 ;
  assign n28515 = ( n28136 & n28146 ) | ( n28136 & ~n28514 ) | ( n28146 & ~n28514 ) ;
  assign n28516 = n28513 & ~n28515 ;
  assign n28517 = ~n28513 & n28515 ;
  assign n28518 = n28516 | n28517 ;
  assign n28519 = x101 & n9933 ;
  assign n28520 = x100 & n9928 ;
  assign n28521 = x99 & ~n9927 ;
  assign n28522 = n10379 & n28521 ;
  assign n28523 = n28520 | n28522 ;
  assign n28524 = n28519 | n28523 ;
  assign n28525 = n9936 | n28519 ;
  assign n28526 = n28523 | n28525 ;
  assign n28527 = ( n6844 & n28524 ) | ( n6844 & n28526 ) | ( n28524 & n28526 ) ;
  assign n28528 = x47 & n28526 ;
  assign n28529 = x47 & n28519 ;
  assign n28530 = ( x47 & n28523 ) | ( x47 & n28529 ) | ( n28523 & n28529 ) ;
  assign n28531 = ( n6844 & n28528 ) | ( n6844 & n28530 ) | ( n28528 & n28530 ) ;
  assign n28532 = x47 & ~n28530 ;
  assign n28533 = x47 & ~n28526 ;
  assign n28534 = ( ~n6844 & n28532 ) | ( ~n6844 & n28533 ) | ( n28532 & n28533 ) ;
  assign n28535 = ( n28527 & ~n28531 ) | ( n28527 & n28534 ) | ( ~n28531 & n28534 ) ;
  assign n28536 = n28518 & ~n28535 ;
  assign n28537 = ~n28518 & n28535 ;
  assign n28538 = n28536 | n28537 ;
  assign n28539 = n28167 | n28170 ;
  assign n28540 = ( n28167 & ~n28169 ) | ( n28167 & n28539 ) | ( ~n28169 & n28539 ) ;
  assign n28541 = n28538 & n28540 ;
  assign n28542 = ~n28538 & n28540 ;
  assign n28543 = x104 & n8724 ;
  assign n28544 = x103 & n8719 ;
  assign n28545 = x102 & ~n8718 ;
  assign n28546 = n9149 & n28545 ;
  assign n28547 = n28544 | n28546 ;
  assign n28548 = n28543 | n28547 ;
  assign n28549 = n8727 | n28543 ;
  assign n28550 = n28547 | n28549 ;
  assign n28551 = ( n7911 & n28548 ) | ( n7911 & n28550 ) | ( n28548 & n28550 ) ;
  assign n28552 = x44 & n28550 ;
  assign n28553 = x44 & n28543 ;
  assign n28554 = ( x44 & n28547 ) | ( x44 & n28553 ) | ( n28547 & n28553 ) ;
  assign n28555 = ( n7911 & n28552 ) | ( n7911 & n28554 ) | ( n28552 & n28554 ) ;
  assign n28556 = x44 & ~n28554 ;
  assign n28557 = x44 & ~n28550 ;
  assign n28558 = ( ~n7911 & n28556 ) | ( ~n7911 & n28557 ) | ( n28556 & n28557 ) ;
  assign n28559 = ( n28551 & ~n28555 ) | ( n28551 & n28558 ) | ( ~n28555 & n28558 ) ;
  assign n28560 = n28538 & ~n28559 ;
  assign n28561 = ( n28542 & ~n28559 ) | ( n28542 & n28560 ) | ( ~n28559 & n28560 ) ;
  assign n28562 = ~n28541 & n28561 ;
  assign n28563 = n28538 | n28542 ;
  assign n28564 = n28541 & n28559 ;
  assign n28565 = ( n28559 & ~n28563 ) | ( n28559 & n28564 ) | ( ~n28563 & n28564 ) ;
  assign n28566 = n28562 | n28565 ;
  assign n28567 = ( n28173 & ~n28190 ) | ( n28173 & n28195 ) | ( ~n28190 & n28195 ) ;
  assign n28568 = ( n27569 & ~n28173 ) | ( n27569 & n28190 ) | ( ~n28173 & n28190 ) ;
  assign n28569 = ( n28199 & n28567 ) | ( n28199 & ~n28568 ) | ( n28567 & ~n28568 ) ;
  assign n28570 = n28566 | n28569 ;
  assign n28571 = n28566 & n28569 ;
  assign n28572 = n28570 & ~n28571 ;
  assign n28573 = x107 & n7566 ;
  assign n28574 = x106 & n7561 ;
  assign n28575 = x105 & ~n7560 ;
  assign n28576 = n7953 & n28575 ;
  assign n28577 = n28574 | n28576 ;
  assign n28578 = n28573 | n28577 ;
  assign n28579 = n7569 | n28573 ;
  assign n28580 = n28577 | n28579 ;
  assign n28581 = ( n9084 & n28578 ) | ( n9084 & n28580 ) | ( n28578 & n28580 ) ;
  assign n28582 = x41 & n28580 ;
  assign n28583 = x41 & n28573 ;
  assign n28584 = ( x41 & n28577 ) | ( x41 & n28583 ) | ( n28577 & n28583 ) ;
  assign n28585 = ( n9084 & n28582 ) | ( n9084 & n28584 ) | ( n28582 & n28584 ) ;
  assign n28586 = x41 & ~n28584 ;
  assign n28587 = x41 & ~n28580 ;
  assign n28588 = ( ~n9084 & n28586 ) | ( ~n9084 & n28587 ) | ( n28586 & n28587 ) ;
  assign n28589 = ( n28581 & ~n28585 ) | ( n28581 & n28588 ) | ( ~n28585 & n28588 ) ;
  assign n28590 = n28572 & ~n28589 ;
  assign n28591 = n28572 | n28589 ;
  assign n28592 = ( ~n28572 & n28590 ) | ( ~n28572 & n28591 ) | ( n28590 & n28591 ) ;
  assign n28593 = n28221 | n28225 ;
  assign n28594 = ( n28221 & n28223 ) | ( n28221 & n28593 ) | ( n28223 & n28593 ) ;
  assign n28595 = n28592 | n28594 ;
  assign n28596 = n28592 & n28594 ;
  assign n28597 = n28595 & ~n28596 ;
  assign n28598 = x110 & n6536 ;
  assign n28599 = x109 & n6531 ;
  assign n28600 = x108 & ~n6530 ;
  assign n28601 = n6871 & n28600 ;
  assign n28602 = n28599 | n28601 ;
  assign n28603 = n28598 | n28602 ;
  assign n28604 = n6539 | n28598 ;
  assign n28605 = n28602 | n28604 ;
  assign n28606 = ( n10330 & n28603 ) | ( n10330 & n28605 ) | ( n28603 & n28605 ) ;
  assign n28607 = x38 & n28605 ;
  assign n28608 = x38 & n28598 ;
  assign n28609 = ( x38 & n28602 ) | ( x38 & n28608 ) | ( n28602 & n28608 ) ;
  assign n28610 = ( n10330 & n28607 ) | ( n10330 & n28609 ) | ( n28607 & n28609 ) ;
  assign n28611 = x38 & ~n28609 ;
  assign n28612 = x38 & ~n28605 ;
  assign n28613 = ( ~n10330 & n28611 ) | ( ~n10330 & n28612 ) | ( n28611 & n28612 ) ;
  assign n28614 = ( n28606 & ~n28610 ) | ( n28606 & n28613 ) | ( ~n28610 & n28613 ) ;
  assign n28615 = ~n28597 & n28614 ;
  assign n28616 = n28592 | n28614 ;
  assign n28617 = ( n28594 & n28614 ) | ( n28594 & n28616 ) | ( n28614 & n28616 ) ;
  assign n28618 = n28595 & ~n28617 ;
  assign n28619 = n28615 | n28618 ;
  assign n28620 = n28246 | n28252 ;
  assign n28621 = n28619 | n28620 ;
  assign n28622 = n28619 & n28620 ;
  assign n28623 = n28621 & ~n28622 ;
  assign n28624 = x113 & n5554 ;
  assign n28625 = x112 & n5549 ;
  assign n28626 = x111 & ~n5548 ;
  assign n28627 = n5893 & n28626 ;
  assign n28628 = n28625 | n28627 ;
  assign n28629 = n28624 | n28628 ;
  assign n28630 = n5557 | n28624 ;
  assign n28631 = n28628 | n28630 ;
  assign n28632 = ( ~n11642 & n28629 ) | ( ~n11642 & n28631 ) | ( n28629 & n28631 ) ;
  assign n28633 = n28629 & n28631 ;
  assign n28634 = ( n11626 & n28632 ) | ( n11626 & n28633 ) | ( n28632 & n28633 ) ;
  assign n28635 = x35 & n28634 ;
  assign n28636 = x35 & ~n28634 ;
  assign n28637 = ( n28634 & ~n28635 ) | ( n28634 & n28636 ) | ( ~n28635 & n28636 ) ;
  assign n28638 = ~n28623 & n28637 ;
  assign n28639 = n28618 | n28637 ;
  assign n28640 = n28615 | n28639 ;
  assign n28641 = ( n28620 & n28637 ) | ( n28620 & n28640 ) | ( n28637 & n28640 ) ;
  assign n28642 = n28621 & ~n28641 ;
  assign n28643 = n28638 | n28642 ;
  assign n28644 = x119 & n3816 ;
  assign n28645 = x118 & n3811 ;
  assign n28646 = x117 & ~n3810 ;
  assign n28647 = n4067 & n28646 ;
  assign n28648 = n28645 | n28647 ;
  assign n28649 = n28644 | n28648 ;
  assign n28650 = n3819 | n28644 ;
  assign n28651 = n28648 | n28650 ;
  assign n28652 = ( n14496 & n28649 ) | ( n14496 & n28651 ) | ( n28649 & n28651 ) ;
  assign n28653 = x29 & n28651 ;
  assign n28654 = x29 & n28644 ;
  assign n28655 = ( x29 & n28648 ) | ( x29 & n28654 ) | ( n28648 & n28654 ) ;
  assign n28656 = ( n14496 & n28653 ) | ( n14496 & n28655 ) | ( n28653 & n28655 ) ;
  assign n28657 = x29 & ~n28655 ;
  assign n28658 = x29 & ~n28651 ;
  assign n28659 = ( ~n14496 & n28657 ) | ( ~n14496 & n28658 ) | ( n28657 & n28658 ) ;
  assign n28660 = ( n28652 & ~n28656 ) | ( n28652 & n28659 ) | ( ~n28656 & n28659 ) ;
  assign n28661 = n27974 | n28283 ;
  assign n28662 = ( n27976 & n28283 ) | ( n27976 & n28661 ) | ( n28283 & n28661 ) ;
  assign n28663 = n28660 | n28662 ;
  assign n28664 = n27977 | n28660 ;
  assign n28665 = ( n27979 & n28663 ) | ( n27979 & n28664 ) | ( n28663 & n28664 ) ;
  assign n28666 = n28660 & n28662 ;
  assign n28667 = n27977 & n28660 ;
  assign n28668 = ( n27979 & n28666 ) | ( n27979 & n28667 ) | ( n28666 & n28667 ) ;
  assign n28669 = n28665 & ~n28668 ;
  assign n28670 = x116 & n4631 ;
  assign n28671 = x115 & n4626 ;
  assign n28672 = x114 & ~n4625 ;
  assign n28673 = n4943 & n28672 ;
  assign n28674 = n28671 | n28673 ;
  assign n28675 = n28670 | n28674 ;
  assign n28676 = n4634 | n28670 ;
  assign n28677 = n28674 | n28676 ;
  assign n28678 = ( ~n13040 & n28675 ) | ( ~n13040 & n28677 ) | ( n28675 & n28677 ) ;
  assign n28679 = n28675 & n28677 ;
  assign n28680 = ( n13022 & n28678 ) | ( n13022 & n28679 ) | ( n28678 & n28679 ) ;
  assign n28681 = x32 & n28680 ;
  assign n28682 = x32 & ~n28680 ;
  assign n28683 = ( n28680 & ~n28681 ) | ( n28680 & n28682 ) | ( ~n28681 & n28682 ) ;
  assign n28684 = n28272 & n28683 ;
  assign n28685 = n28255 & n28684 ;
  assign n28686 = ( n28280 & n28683 ) | ( n28280 & n28685 ) | ( n28683 & n28685 ) ;
  assign n28687 = n28272 | n28683 ;
  assign n28688 = ( n28255 & n28683 ) | ( n28255 & n28687 ) | ( n28683 & n28687 ) ;
  assign n28689 = n28280 | n28688 ;
  assign n28690 = ~n28686 & n28689 ;
  assign n28691 = ( n28643 & n28669 ) | ( n28643 & ~n28690 ) | ( n28669 & ~n28690 ) ;
  assign n28692 = ( ~n28669 & n28690 ) | ( ~n28669 & n28691 ) | ( n28690 & n28691 ) ;
  assign n28693 = ( ~n28643 & n28691 ) | ( ~n28643 & n28692 ) | ( n28691 & n28692 ) ;
  assign n28694 = n28370 & n28693 ;
  assign n28695 = n28370 | n28693 ;
  assign n28696 = ~n28694 & n28695 ;
  assign n28697 = x125 & n2429 ;
  assign n28698 = x124 & n2424 ;
  assign n28699 = x123 & ~n2423 ;
  assign n28700 = n2631 & n28699 ;
  assign n28701 = n28698 | n28700 ;
  assign n28702 = n28697 | n28701 ;
  assign n28703 = n2432 | n28697 ;
  assign n28704 = n28701 | n28703 ;
  assign n28705 = ( n17670 & n28702 ) | ( n17670 & n28704 ) | ( n28702 & n28704 ) ;
  assign n28706 = x23 & n28704 ;
  assign n28707 = x23 & n28697 ;
  assign n28708 = ( x23 & n28701 ) | ( x23 & n28707 ) | ( n28701 & n28707 ) ;
  assign n28709 = ( n17670 & n28706 ) | ( n17670 & n28708 ) | ( n28706 & n28708 ) ;
  assign n28710 = x23 & ~n28708 ;
  assign n28711 = x23 & ~n28704 ;
  assign n28712 = ( ~n17670 & n28710 ) | ( ~n17670 & n28711 ) | ( n28710 & n28711 ) ;
  assign n28713 = ( n28705 & ~n28709 ) | ( n28705 & n28712 ) | ( ~n28709 & n28712 ) ;
  assign n28714 = n27925 | n28290 ;
  assign n28715 = ( n27925 & n27927 ) | ( n27925 & n28714 ) | ( n27927 & n28714 ) ;
  assign n28716 = n28713 | n28715 ;
  assign n28717 = n28713 & n28715 ;
  assign n28718 = n28716 & ~n28717 ;
  assign n28719 = n28696 & n28718 ;
  assign n28720 = n28718 & ~n28719 ;
  assign n28721 = ( n28696 & ~n28719 ) | ( n28696 & n28720 ) | ( ~n28719 & n28720 ) ;
  assign n28722 = n28342 | n28721 ;
  assign n28723 = n28341 | n28722 ;
  assign n28724 = n28342 & n28721 ;
  assign n28725 = ( n28341 & n28721 ) | ( n28341 & n28724 ) | ( n28721 & n28724 ) ;
  assign n28726 = n28723 & ~n28725 ;
  assign n28727 = n27431 & n27876 ;
  assign n28728 = n27436 & n28727 ;
  assign n28729 = ( n27823 & n27876 ) | ( n27823 & n28728 ) | ( n27876 & n28728 ) ;
  assign n28730 = n27876 & n28727 ;
  assign n28731 = n27436 & n28730 ;
  assign n28732 = ( n27439 & n28729 ) | ( n27439 & n28731 ) | ( n28729 & n28731 ) ;
  assign n28733 = n28298 & ~n28732 ;
  assign n28734 = n27876 & ~n28727 ;
  assign n28735 = ( ~n27436 & n27876 ) | ( ~n27436 & n28734 ) | ( n27876 & n28734 ) ;
  assign n28736 = ~n27823 & n28735 ;
  assign n28737 = ( ~n27439 & n28735 ) | ( ~n27439 & n28736 ) | ( n28735 & n28736 ) ;
  assign n28738 = n28296 & ~n28737 ;
  assign n28739 = ~n28733 & n28738 ;
  assign n28740 = ( n28296 & n28732 ) | ( n28296 & ~n28739 ) | ( n28732 & ~n28739 ) ;
  assign n28741 = n28726 & ~n28740 ;
  assign n28742 = ~n28726 & n28740 ;
  assign n28743 = n28741 | n28742 ;
  assign n28744 = n28303 | n28314 ;
  assign n28745 = n28302 | n28303 ;
  assign n28746 = n28304 | n28745 ;
  assign n28747 = ( n27851 & n28744 ) | ( n27851 & n28746 ) | ( n28744 & n28746 ) ;
  assign n28748 = n28743 & n28747 ;
  assign n28749 = n28743 & n28746 ;
  assign n28750 = n28743 & n28744 ;
  assign n28751 = ( n27852 & n28749 ) | ( n27852 & n28750 ) | ( n28749 & n28750 ) ;
  assign n28752 = ( n27383 & n28748 ) | ( n27383 & n28751 ) | ( n28748 & n28751 ) ;
  assign n28753 = n28303 & n28743 ;
  assign n28754 = ( n28312 & n28749 ) | ( n28312 & n28753 ) | ( n28749 & n28753 ) ;
  assign n28755 = ( n26030 & n28752 ) | ( n26030 & n28754 ) | ( n28752 & n28754 ) ;
  assign n28756 = ( n27852 & n28744 ) | ( n27852 & n28746 ) | ( n28744 & n28746 ) ;
  assign n28757 = ( n27383 & n28747 ) | ( n27383 & n28756 ) | ( n28747 & n28756 ) ;
  assign n28758 = ( n28303 & n28312 ) | ( n28303 & n28746 ) | ( n28312 & n28746 ) ;
  assign n28759 = ( n26030 & n28757 ) | ( n26030 & n28758 ) | ( n28757 & n28758 ) ;
  assign n28760 = ( ~n28726 & n28740 ) | ( ~n28726 & n28759 ) | ( n28740 & n28759 ) ;
  assign n28761 = ( n28741 & ~n28755 ) | ( n28741 & n28760 ) | ( ~n28755 & n28760 ) ;
  assign n28762 = n28696 | n28713 ;
  assign n28763 = ( n28696 & n28715 ) | ( n28696 & n28762 ) | ( n28715 & n28762 ) ;
  assign n28764 = ( n28717 & n28718 ) | ( n28717 & n28763 ) | ( n28718 & n28763 ) ;
  assign n28765 = x127 & ~n1853 ;
  assign n28766 = n2037 & n28765 ;
  assign n28767 = n1862 & n19877 ;
  assign n28768 = n28766 | n28767 ;
  assign n28769 = n1862 & n19880 ;
  assign n28770 = n28766 | n28769 ;
  assign n28771 = ( n18202 & n28768 ) | ( n18202 & n28770 ) | ( n28768 & n28770 ) ;
  assign n28772 = n28768 & n28770 ;
  assign n28773 = ( n18212 & n28771 ) | ( n18212 & n28772 ) | ( n28771 & n28772 ) ;
  assign n28774 = ( n18214 & n28771 ) | ( n18214 & n28772 ) | ( n28771 & n28772 ) ;
  assign n28775 = ( n14002 & n28773 ) | ( n14002 & n28774 ) | ( n28773 & n28774 ) ;
  assign n28776 = x20 & n28773 ;
  assign n28777 = x20 & n28774 ;
  assign n28778 = ( n14002 & n28776 ) | ( n14002 & n28777 ) | ( n28776 & n28777 ) ;
  assign n28779 = x20 & ~n28777 ;
  assign n28780 = x20 & ~n28776 ;
  assign n28781 = ( ~n14002 & n28779 ) | ( ~n14002 & n28780 ) | ( n28779 & n28780 ) ;
  assign n28782 = ( n28775 & ~n28778 ) | ( n28775 & n28781 ) | ( ~n28778 & n28781 ) ;
  assign n28783 = n28763 & n28782 ;
  assign n28784 = n28717 & n28782 ;
  assign n28785 = ( n28718 & n28783 ) | ( n28718 & n28784 ) | ( n28783 & n28784 ) ;
  assign n28786 = n28764 & ~n28785 ;
  assign n28787 = x126 & n2429 ;
  assign n28788 = x125 & n2424 ;
  assign n28789 = x124 & ~n2423 ;
  assign n28790 = n2631 & n28789 ;
  assign n28791 = n28788 | n28790 ;
  assign n28792 = n28787 | n28791 ;
  assign n28793 = n2432 | n28787 ;
  assign n28794 = n28791 | n28793 ;
  assign n28795 = ( n18220 & n28792 ) | ( n18220 & n28794 ) | ( n28792 & n28794 ) ;
  assign n28796 = x23 & n28794 ;
  assign n28797 = x23 & n28787 ;
  assign n28798 = ( x23 & n28791 ) | ( x23 & n28797 ) | ( n28791 & n28797 ) ;
  assign n28799 = ( n18220 & n28796 ) | ( n18220 & n28798 ) | ( n28796 & n28798 ) ;
  assign n28800 = x23 & ~n28798 ;
  assign n28801 = x23 & ~n28794 ;
  assign n28802 = ( ~n18220 & n28800 ) | ( ~n18220 & n28801 ) | ( n28800 & n28801 ) ;
  assign n28803 = ( n28795 & ~n28799 ) | ( n28795 & n28802 ) | ( ~n28799 & n28802 ) ;
  assign n28804 = n28364 | n28693 ;
  assign n28805 = ( n28364 & n28370 ) | ( n28364 & n28804 ) | ( n28370 & n28804 ) ;
  assign n28806 = ~n28803 & n28805 ;
  assign n28807 = x123 & n3085 ;
  assign n28808 = x122 & n3080 ;
  assign n28809 = x121 & ~n3079 ;
  assign n28810 = n3309 & n28809 ;
  assign n28811 = n28808 | n28810 ;
  assign n28812 = n28807 | n28811 ;
  assign n28813 = n3088 | n28807 ;
  assign n28814 = n28811 | n28813 ;
  assign n28815 = ( n16086 & n28812 ) | ( n16086 & n28814 ) | ( n28812 & n28814 ) ;
  assign n28816 = x26 & n28814 ;
  assign n28817 = x26 & n28807 ;
  assign n28818 = ( x26 & n28811 ) | ( x26 & n28817 ) | ( n28811 & n28817 ) ;
  assign n28819 = ( n16086 & n28816 ) | ( n16086 & n28818 ) | ( n28816 & n28818 ) ;
  assign n28820 = x26 & ~n28818 ;
  assign n28821 = x26 & ~n28814 ;
  assign n28822 = ( ~n16086 & n28820 ) | ( ~n16086 & n28821 ) | ( n28820 & n28821 ) ;
  assign n28823 = ( n28815 & ~n28819 ) | ( n28815 & n28822 ) | ( ~n28819 & n28822 ) ;
  assign n28824 = n28643 & n28690 ;
  assign n28825 = n28643 | n28690 ;
  assign n28826 = ~n28824 & n28825 ;
  assign n28827 = n28668 | n28826 ;
  assign n28828 = ( n28668 & n28669 ) | ( n28668 & n28827 ) | ( n28669 & n28827 ) ;
  assign n28829 = n28823 | n28828 ;
  assign n28830 = n28823 & n28828 ;
  assign n28831 = n28829 & ~n28830 ;
  assign n28849 = n28643 | n28686 ;
  assign n28850 = ( n28686 & n28690 ) | ( n28686 & n28849 ) | ( n28690 & n28849 ) ;
  assign n28832 = x120 & n3816 ;
  assign n28833 = x119 & n3811 ;
  assign n28834 = x118 & ~n3810 ;
  assign n28835 = n4067 & n28834 ;
  assign n28836 = n28833 | n28835 ;
  assign n28837 = n28832 | n28836 ;
  assign n28838 = n3819 | n28832 ;
  assign n28839 = n28836 | n28838 ;
  assign n28840 = ( n14991 & n28837 ) | ( n14991 & n28839 ) | ( n28837 & n28839 ) ;
  assign n28841 = x29 & n28839 ;
  assign n28842 = x29 & n28832 ;
  assign n28843 = ( x29 & n28836 ) | ( x29 & n28842 ) | ( n28836 & n28842 ) ;
  assign n28844 = ( n14991 & n28841 ) | ( n14991 & n28843 ) | ( n28841 & n28843 ) ;
  assign n28845 = x29 & ~n28843 ;
  assign n28846 = x29 & ~n28839 ;
  assign n28847 = ( ~n14991 & n28845 ) | ( ~n14991 & n28846 ) | ( n28845 & n28846 ) ;
  assign n28848 = ( n28840 & ~n28844 ) | ( n28840 & n28847 ) | ( ~n28844 & n28847 ) ;
  assign n28851 = n28848 & n28850 ;
  assign n28852 = n28850 & ~n28851 ;
  assign n28853 = x114 & n5554 ;
  assign n28854 = x113 & n5549 ;
  assign n28855 = x112 & ~n5548 ;
  assign n28856 = n5893 & n28855 ;
  assign n28857 = n28854 | n28856 ;
  assign n28858 = n28853 | n28857 ;
  assign n28859 = n5557 | n28853 ;
  assign n28860 = n28857 | n28859 ;
  assign n28861 = ( ~n12095 & n28858 ) | ( ~n12095 & n28860 ) | ( n28858 & n28860 ) ;
  assign n28862 = n28858 & n28860 ;
  assign n28863 = ( n12079 & n28861 ) | ( n12079 & n28862 ) | ( n28861 & n28862 ) ;
  assign n28864 = x35 & n28863 ;
  assign n28865 = x35 & ~n28863 ;
  assign n28866 = ( n28863 & ~n28864 ) | ( n28863 & n28865 ) | ( ~n28864 & n28865 ) ;
  assign n28867 = x117 & n4631 ;
  assign n28868 = x116 & n4626 ;
  assign n28869 = x115 & ~n4625 ;
  assign n28870 = n4943 & n28869 ;
  assign n28871 = n28868 | n28870 ;
  assign n28872 = n28867 | n28871 ;
  assign n28873 = n4634 | n28867 ;
  assign n28874 = n28871 | n28873 ;
  assign n28875 = ( ~n13522 & n28872 ) | ( ~n13522 & n28874 ) | ( n28872 & n28874 ) ;
  assign n28876 = n28872 & n28874 ;
  assign n28877 = ( n13503 & n28875 ) | ( n13503 & n28876 ) | ( n28875 & n28876 ) ;
  assign n28878 = x32 & n28877 ;
  assign n28879 = x32 & ~n28877 ;
  assign n28880 = ( n28877 & ~n28878 ) | ( n28877 & n28879 ) | ( ~n28878 & n28879 ) ;
  assign n28881 = n28641 & n28880 ;
  assign n28882 = n28622 & n28880 ;
  assign n28883 = ( n28623 & n28881 ) | ( n28623 & n28882 ) | ( n28881 & n28882 ) ;
  assign n28884 = n28641 | n28880 ;
  assign n28885 = n28622 | n28880 ;
  assign n28886 = ( n28623 & n28884 ) | ( n28623 & n28885 ) | ( n28884 & n28885 ) ;
  assign n28887 = ~n28883 & n28886 ;
  assign n28888 = n28542 | n28565 ;
  assign n28889 = x84 & n18290 ;
  assign n28890 = x63 & x83 ;
  assign n28891 = ~n18290 & n28890 ;
  assign n28892 = n28889 | n28891 ;
  assign n28893 = n28374 & ~n28892 ;
  assign n28894 = ~n28374 & n28892 ;
  assign n28895 = n28893 | n28894 ;
  assign n28897 = x86 & n17141 ;
  assign n28898 = x85 & ~n17140 ;
  assign n28899 = n17724 & n28898 ;
  assign n28900 = n28897 | n28899 ;
  assign n28896 = x87 & n17146 ;
  assign n28902 = n17149 | n28896 ;
  assign n28903 = n28900 | n28902 ;
  assign n28901 = n28896 | n28900 ;
  assign n28904 = n28901 & n28903 ;
  assign n28905 = ( n2816 & n28903 ) | ( n2816 & n28904 ) | ( n28903 & n28904 ) ;
  assign n28906 = x62 & n28904 ;
  assign n28907 = x62 & n28903 ;
  assign n28908 = ( n2816 & n28906 ) | ( n2816 & n28907 ) | ( n28906 & n28907 ) ;
  assign n28909 = x62 & ~n28904 ;
  assign n28910 = x62 & ~n28903 ;
  assign n28911 = ( ~n2816 & n28909 ) | ( ~n2816 & n28910 ) | ( n28909 & n28910 ) ;
  assign n28912 = ( n28905 & ~n28908 ) | ( n28905 & n28911 ) | ( ~n28908 & n28911 ) ;
  assign n28913 = ~n28895 & n28912 ;
  assign n28914 = n28895 & ~n28912 ;
  assign n28915 = n28913 | n28914 ;
  assign n28916 = n28378 | n28398 ;
  assign n28917 = ~n28378 & n28379 ;
  assign n28918 = ( n28394 & n28916 ) | ( n28394 & ~n28917 ) | ( n28916 & ~n28917 ) ;
  assign n28919 = ~n28915 & n28918 ;
  assign n28920 = n28915 & ~n28918 ;
  assign n28921 = n28919 | n28920 ;
  assign n28922 = x90 & n15552 ;
  assign n28923 = x89 & n15547 ;
  assign n28924 = x88 & ~n15546 ;
  assign n28925 = n16123 & n28924 ;
  assign n28926 = n28923 | n28925 ;
  assign n28927 = n28922 | n28926 ;
  assign n28928 = n15555 | n28922 ;
  assign n28929 = n28926 | n28928 ;
  assign n28930 = ( n3519 & n28927 ) | ( n3519 & n28929 ) | ( n28927 & n28929 ) ;
  assign n28931 = x59 & n28929 ;
  assign n28932 = x59 & n28922 ;
  assign n28933 = ( x59 & n28926 ) | ( x59 & n28932 ) | ( n28926 & n28932 ) ;
  assign n28934 = ( n3519 & n28931 ) | ( n3519 & n28933 ) | ( n28931 & n28933 ) ;
  assign n28935 = x59 & ~n28933 ;
  assign n28936 = x59 & ~n28929 ;
  assign n28937 = ( ~n3519 & n28935 ) | ( ~n3519 & n28936 ) | ( n28935 & n28936 ) ;
  assign n28938 = ( n28930 & ~n28934 ) | ( n28930 & n28937 ) | ( ~n28934 & n28937 ) ;
  assign n28939 = ~n28921 & n28938 ;
  assign n28940 = n28921 & ~n28938 ;
  assign n28941 = n28939 | n28940 ;
  assign n28942 = n28404 & ~n28426 ;
  assign n28943 = ( n28406 & n28426 ) | ( n28406 & ~n28942 ) | ( n28426 & ~n28942 ) ;
  assign n28944 = ( n28407 & ~n28409 ) | ( n28407 & n28943 ) | ( ~n28409 & n28943 ) ;
  assign n28945 = ~n28941 & n28944 ;
  assign n28946 = n28941 & ~n28944 ;
  assign n28947 = n28945 | n28946 ;
  assign n28948 = x93 & n14045 ;
  assign n28949 = x92 & n14040 ;
  assign n28950 = x91 & ~n14039 ;
  assign n28951 = n14552 & n28950 ;
  assign n28952 = n28949 | n28951 ;
  assign n28953 = n28948 | n28952 ;
  assign n28954 = n14048 | n28948 ;
  assign n28955 = n28952 | n28954 ;
  assign n28956 = ( n4305 & n28953 ) | ( n4305 & n28955 ) | ( n28953 & n28955 ) ;
  assign n28957 = x56 & n28955 ;
  assign n28958 = x56 & n28948 ;
  assign n28959 = ( x56 & n28952 ) | ( x56 & n28958 ) | ( n28952 & n28958 ) ;
  assign n28960 = ( n4305 & n28957 ) | ( n4305 & n28959 ) | ( n28957 & n28959 ) ;
  assign n28961 = x56 & ~n28959 ;
  assign n28962 = x56 & ~n28955 ;
  assign n28963 = ( ~n4305 & n28961 ) | ( ~n4305 & n28962 ) | ( n28961 & n28962 ) ;
  assign n28964 = ( n28956 & ~n28960 ) | ( n28956 & n28963 ) | ( ~n28960 & n28963 ) ;
  assign n28965 = n28947 | n28964 ;
  assign n28966 = n28947 & ~n28964 ;
  assign n28967 = ( ~n28947 & n28965 ) | ( ~n28947 & n28966 ) | ( n28965 & n28966 ) ;
  assign n28968 = ( ~n28429 & n28430 ) | ( ~n28429 & n28450 ) | ( n28430 & n28450 ) ;
  assign n28969 = ~n28967 & n28968 ;
  assign n28970 = n28967 | n28969 ;
  assign n28971 = x96 & n12574 ;
  assign n28972 = x95 & n12569 ;
  assign n28973 = x94 & ~n12568 ;
  assign n28974 = n13076 & n28973 ;
  assign n28975 = n28972 | n28974 ;
  assign n28976 = n28971 | n28975 ;
  assign n28977 = n12577 | n28971 ;
  assign n28978 = n28975 | n28977 ;
  assign n28979 = ( n5202 & n28976 ) | ( n5202 & n28978 ) | ( n28976 & n28978 ) ;
  assign n28980 = x53 & n28978 ;
  assign n28981 = x53 & n28971 ;
  assign n28982 = ( x53 & n28975 ) | ( x53 & n28981 ) | ( n28975 & n28981 ) ;
  assign n28983 = ( n5202 & n28980 ) | ( n5202 & n28982 ) | ( n28980 & n28982 ) ;
  assign n28984 = x53 & ~n28982 ;
  assign n28985 = x53 & ~n28978 ;
  assign n28986 = ( ~n5202 & n28984 ) | ( ~n5202 & n28985 ) | ( n28984 & n28985 ) ;
  assign n28987 = ( n28979 & ~n28983 ) | ( n28979 & n28986 ) | ( ~n28983 & n28986 ) ;
  assign n28988 = n28968 & ~n28987 ;
  assign n28989 = n28967 & n28988 ;
  assign n28990 = ( n28970 & n28987 ) | ( n28970 & ~n28989 ) | ( n28987 & ~n28989 ) ;
  assign n28991 = ~n28968 & n28987 ;
  assign n28992 = ( ~n28967 & n28987 ) | ( ~n28967 & n28991 ) | ( n28987 & n28991 ) ;
  assign n28993 = n28970 & n28992 ;
  assign n28994 = n28990 & ~n28993 ;
  assign n28995 = n28457 | n28476 ;
  assign n28996 = ( n28457 & ~n28459 ) | ( n28457 & n28995 ) | ( ~n28459 & n28995 ) ;
  assign n28997 = ~n28994 & n28996 ;
  assign n28998 = n28994 & ~n28996 ;
  assign n28999 = n28997 | n28998 ;
  assign n29000 = x99 & n11205 ;
  assign n29001 = x98 & n11200 ;
  assign n29002 = x97 & ~n11199 ;
  assign n29003 = n11679 & n29002 ;
  assign n29004 = n29001 | n29003 ;
  assign n29005 = n29000 | n29004 ;
  assign n29006 = n11208 | n29000 ;
  assign n29007 = n29004 | n29006 ;
  assign n29008 = ( n6164 & n29005 ) | ( n6164 & n29007 ) | ( n29005 & n29007 ) ;
  assign n29009 = x50 & n29007 ;
  assign n29010 = x50 & n29000 ;
  assign n29011 = ( x50 & n29004 ) | ( x50 & n29010 ) | ( n29004 & n29010 ) ;
  assign n29012 = ( n6164 & n29009 ) | ( n6164 & n29011 ) | ( n29009 & n29011 ) ;
  assign n29013 = x50 & ~n29011 ;
  assign n29014 = x50 & ~n29007 ;
  assign n29015 = ( ~n6164 & n29013 ) | ( ~n6164 & n29014 ) | ( n29013 & n29014 ) ;
  assign n29016 = ( n29008 & ~n29012 ) | ( n29008 & n29015 ) | ( ~n29012 & n29015 ) ;
  assign n29017 = ~n28999 & n29016 ;
  assign n29018 = n28999 & ~n29016 ;
  assign n29019 = n29017 | n29018 ;
  assign n29020 = ( n28484 & ~n28485 ) | ( n28484 & n28511 ) | ( ~n28485 & n28511 ) ;
  assign n29021 = ~n29019 & n29020 ;
  assign n29022 = n29019 & ~n29020 ;
  assign n29023 = n29021 | n29022 ;
  assign n29024 = x102 & n9933 ;
  assign n29025 = x101 & n9928 ;
  assign n29026 = x100 & ~n9927 ;
  assign n29027 = n10379 & n29026 ;
  assign n29028 = n29025 | n29027 ;
  assign n29029 = n29024 | n29028 ;
  assign n29030 = n9936 | n29024 ;
  assign n29031 = n29028 | n29030 ;
  assign n29032 = ( n7178 & n29029 ) | ( n7178 & n29031 ) | ( n29029 & n29031 ) ;
  assign n29033 = x47 & n29031 ;
  assign n29034 = x47 & n29024 ;
  assign n29035 = ( x47 & n29028 ) | ( x47 & n29034 ) | ( n29028 & n29034 ) ;
  assign n29036 = ( n7178 & n29033 ) | ( n7178 & n29035 ) | ( n29033 & n29035 ) ;
  assign n29037 = x47 & ~n29035 ;
  assign n29038 = x47 & ~n29031 ;
  assign n29039 = ( ~n7178 & n29037 ) | ( ~n7178 & n29038 ) | ( n29037 & n29038 ) ;
  assign n29040 = ( n29032 & ~n29036 ) | ( n29032 & n29039 ) | ( ~n29036 & n29039 ) ;
  assign n29041 = ~n29023 & n29040 ;
  assign n29042 = n29023 & ~n29040 ;
  assign n29043 = n29041 | n29042 ;
  assign n29044 = n28517 | n28535 ;
  assign n29045 = ( n28517 & ~n28518 ) | ( n28517 & n29044 ) | ( ~n28518 & n29044 ) ;
  assign n29046 = ~n29043 & n29045 ;
  assign n29047 = n29043 & ~n29045 ;
  assign n29048 = n29046 | n29047 ;
  assign n29049 = x105 & n8724 ;
  assign n29050 = x104 & n8719 ;
  assign n29051 = x103 & ~n8718 ;
  assign n29052 = n9149 & n29051 ;
  assign n29053 = n29050 | n29052 ;
  assign n29054 = n29049 | n29053 ;
  assign n29055 = n8727 | n29049 ;
  assign n29056 = n29053 | n29055 ;
  assign n29057 = ( n8273 & n29054 ) | ( n8273 & n29056 ) | ( n29054 & n29056 ) ;
  assign n29058 = x44 & n29056 ;
  assign n29059 = x44 & n29049 ;
  assign n29060 = ( x44 & n29053 ) | ( x44 & n29059 ) | ( n29053 & n29059 ) ;
  assign n29061 = ( n8273 & n29058 ) | ( n8273 & n29060 ) | ( n29058 & n29060 ) ;
  assign n29062 = x44 & ~n29060 ;
  assign n29063 = x44 & ~n29056 ;
  assign n29064 = ( ~n8273 & n29062 ) | ( ~n8273 & n29063 ) | ( n29062 & n29063 ) ;
  assign n29065 = ( n29057 & ~n29061 ) | ( n29057 & n29064 ) | ( ~n29061 & n29064 ) ;
  assign n29066 = ~n29048 & n29065 ;
  assign n29067 = n29048 & ~n29065 ;
  assign n29068 = n29066 | n29067 ;
  assign n29069 = n28888 & ~n29068 ;
  assign n29070 = ~n28888 & n29068 ;
  assign n29071 = n29069 | n29070 ;
  assign n29072 = x108 & n7566 ;
  assign n29073 = x107 & n7561 ;
  assign n29074 = x106 & ~n7560 ;
  assign n29075 = n7953 & n29074 ;
  assign n29076 = n29073 | n29075 ;
  assign n29077 = n29072 | n29076 ;
  assign n29078 = n7569 | n29072 ;
  assign n29079 = n29076 | n29078 ;
  assign n29080 = ( n9479 & n29077 ) | ( n9479 & n29079 ) | ( n29077 & n29079 ) ;
  assign n29081 = x41 & n29079 ;
  assign n29082 = x41 & n29072 ;
  assign n29083 = ( x41 & n29076 ) | ( x41 & n29082 ) | ( n29076 & n29082 ) ;
  assign n29084 = ( n9479 & n29081 ) | ( n9479 & n29083 ) | ( n29081 & n29083 ) ;
  assign n29085 = x41 & ~n29083 ;
  assign n29086 = x41 & ~n29079 ;
  assign n29087 = ( ~n9479 & n29085 ) | ( ~n9479 & n29086 ) | ( n29085 & n29086 ) ;
  assign n29088 = ( n29080 & ~n29084 ) | ( n29080 & n29087 ) | ( ~n29084 & n29087 ) ;
  assign n29089 = ~n29071 & n29088 ;
  assign n29090 = n29071 & ~n29088 ;
  assign n29091 = n29089 | n29090 ;
  assign n29092 = n28569 & ~n28589 ;
  assign n29093 = ( n28566 & ~n28589 ) | ( n28566 & n29092 ) | ( ~n28589 & n29092 ) ;
  assign n29094 = ( n28570 & ~n28572 ) | ( n28570 & n29093 ) | ( ~n28572 & n29093 ) ;
  assign n29095 = n29091 | n29094 ;
  assign n29096 = n29091 & n29094 ;
  assign n29097 = n29095 & ~n29096 ;
  assign n29098 = x111 & n6536 ;
  assign n29099 = x110 & n6531 ;
  assign n29100 = x109 & ~n6530 ;
  assign n29101 = n6871 & n29100 ;
  assign n29102 = n29099 | n29101 ;
  assign n29103 = n29098 | n29102 ;
  assign n29104 = n6539 | n29098 ;
  assign n29105 = n29102 | n29104 ;
  assign n29106 = ( n10749 & n29103 ) | ( n10749 & n29105 ) | ( n29103 & n29105 ) ;
  assign n29107 = x38 & n29105 ;
  assign n29108 = x38 & n29098 ;
  assign n29109 = ( x38 & n29102 ) | ( x38 & n29108 ) | ( n29102 & n29108 ) ;
  assign n29110 = ( n10749 & n29107 ) | ( n10749 & n29109 ) | ( n29107 & n29109 ) ;
  assign n29111 = x38 & ~n29109 ;
  assign n29112 = x38 & ~n29105 ;
  assign n29113 = ( ~n10749 & n29111 ) | ( ~n10749 & n29112 ) | ( n29111 & n29112 ) ;
  assign n29114 = ( n29106 & ~n29110 ) | ( n29106 & n29113 ) | ( ~n29110 & n29113 ) ;
  assign n29115 = n29097 & ~n29114 ;
  assign n29116 = n29097 | n29114 ;
  assign n29117 = ( ~n29097 & n29115 ) | ( ~n29097 & n29116 ) | ( n29115 & n29116 ) ;
  assign n29118 = ( n28596 & n28597 ) | ( n28596 & n28617 ) | ( n28597 & n28617 ) ;
  assign n29119 = n29117 | n29118 ;
  assign n29120 = n29117 & n29118 ;
  assign n29121 = n29119 & ~n29120 ;
  assign n29122 = ( n28866 & n28887 ) | ( n28866 & ~n29121 ) | ( n28887 & ~n29121 ) ;
  assign n29123 = ( ~n28887 & n29121 ) | ( ~n28887 & n29122 ) | ( n29121 & n29122 ) ;
  assign n29124 = ( ~n28866 & n29122 ) | ( ~n28866 & n29123 ) | ( n29122 & n29123 ) ;
  assign n29125 = n28848 & ~n28850 ;
  assign n29126 = ~n29124 & n29125 ;
  assign n29127 = ( n28852 & ~n29124 ) | ( n28852 & n29126 ) | ( ~n29124 & n29126 ) ;
  assign n29128 = n29124 & ~n29125 ;
  assign n29129 = ~n28852 & n29128 ;
  assign n29130 = n29127 | n29129 ;
  assign n29131 = ~n28831 & n29130 ;
  assign n29132 = n28831 & ~n29130 ;
  assign n29133 = n29131 | n29132 ;
  assign n29134 = n28364 & n28803 ;
  assign n29135 = ( n28693 & n28803 ) | ( n28693 & n29134 ) | ( n28803 & n29134 ) ;
  assign n29136 = ( n28370 & n29134 ) | ( n28370 & n29135 ) | ( n29134 & n29135 ) ;
  assign n29137 = n29133 | n29136 ;
  assign n29138 = n28803 & ~n29133 ;
  assign n29139 = ( n28806 & ~n29137 ) | ( n28806 & n29138 ) | ( ~n29137 & n29138 ) ;
  assign n29140 = n29133 & n29136 ;
  assign n29141 = ~n28803 & n29133 ;
  assign n29142 = ( ~n28806 & n29140 ) | ( ~n28806 & n29141 ) | ( n29140 & n29141 ) ;
  assign n29143 = n29139 | n29142 ;
  assign n29144 = n28782 & n29143 ;
  assign n29145 = ~n28764 & n29144 ;
  assign n29146 = ( n28786 & n29143 ) | ( n28786 & n29145 ) | ( n29143 & n29145 ) ;
  assign n29147 = n28782 | n29143 ;
  assign n29148 = ( ~n28764 & n29143 ) | ( ~n28764 & n29147 ) | ( n29143 & n29147 ) ;
  assign n29149 = n28786 | n29148 ;
  assign n29150 = ~n29146 & n29149 ;
  assign n29151 = n28340 | n28721 ;
  assign n29152 = n28340 | n28341 ;
  assign n29153 = ( n28724 & n29151 ) | ( n28724 & n29152 ) | ( n29151 & n29152 ) ;
  assign n29154 = n29150 & n29153 ;
  assign n29155 = n29150 | n29153 ;
  assign n29156 = ~n29154 & n29155 ;
  assign n29157 = n28726 & n28740 ;
  assign n29158 = n28751 | n29157 ;
  assign n29159 = n28743 | n29157 ;
  assign n29160 = ( n28747 & n29157 ) | ( n28747 & n29159 ) | ( n29157 & n29159 ) ;
  assign n29161 = ( n27383 & n29158 ) | ( n27383 & n29160 ) | ( n29158 & n29160 ) ;
  assign n29162 = n28753 | n29157 ;
  assign n29163 = ( n28746 & n29157 ) | ( n28746 & n29159 ) | ( n29157 & n29159 ) ;
  assign n29164 = ( n28312 & n29162 ) | ( n28312 & n29163 ) | ( n29162 & n29163 ) ;
  assign n29165 = ( n26030 & n29161 ) | ( n26030 & n29164 ) | ( n29161 & n29164 ) ;
  assign n29166 = n29156 | n29165 ;
  assign n29167 = n29156 & n29157 ;
  assign n29168 = ( n28751 & n29156 ) | ( n28751 & n29167 ) | ( n29156 & n29167 ) ;
  assign n29169 = n29156 & n29159 ;
  assign n29170 = ( n28747 & n29167 ) | ( n28747 & n29169 ) | ( n29167 & n29169 ) ;
  assign n29171 = ( n27383 & n29168 ) | ( n27383 & n29170 ) | ( n29168 & n29170 ) ;
  assign n29172 = ( n28746 & n29167 ) | ( n28746 & n29169 ) | ( n29167 & n29169 ) ;
  assign n29173 = ( n28753 & n29156 ) | ( n28753 & n29167 ) | ( n29156 & n29167 ) ;
  assign n29174 = ( n28312 & n29172 ) | ( n28312 & n29173 ) | ( n29172 & n29173 ) ;
  assign n29175 = ( n26030 & n29171 ) | ( n26030 & n29174 ) | ( n29171 & n29174 ) ;
  assign n29176 = n29166 & ~n29175 ;
  assign n29177 = x124 & n3085 ;
  assign n29178 = x123 & n3080 ;
  assign n29179 = x122 & ~n3079 ;
  assign n29180 = n3309 & n29179 ;
  assign n29181 = n29178 | n29180 ;
  assign n29182 = n29177 | n29181 ;
  assign n29183 = n3088 | n29177 ;
  assign n29184 = n29181 | n29183 ;
  assign n29185 = ( n17084 & n29182 ) | ( n17084 & n29184 ) | ( n29182 & n29184 ) ;
  assign n29186 = x26 & n29184 ;
  assign n29187 = x26 & n29177 ;
  assign n29188 = ( x26 & n29181 ) | ( x26 & n29187 ) | ( n29181 & n29187 ) ;
  assign n29189 = ( n17084 & n29186 ) | ( n17084 & n29188 ) | ( n29186 & n29188 ) ;
  assign n29190 = x26 & ~n29188 ;
  assign n29191 = x26 & ~n29184 ;
  assign n29192 = ( ~n17084 & n29190 ) | ( ~n17084 & n29191 ) | ( n29190 & n29191 ) ;
  assign n29193 = ( n29185 & ~n29189 ) | ( n29185 & n29192 ) | ( ~n29189 & n29192 ) ;
  assign n29194 = n28830 | n29130 ;
  assign n29195 = ( n28830 & n28831 ) | ( n28830 & n29194 ) | ( n28831 & n29194 ) ;
  assign n29196 = n29193 | n29195 ;
  assign n29197 = n29193 & n29195 ;
  assign n29198 = n29196 & ~n29197 ;
  assign n29199 = ( n28803 & n28806 ) | ( n28803 & ~n29136 ) | ( n28806 & ~n29136 ) ;
  assign n29200 = ( n29136 & n29137 ) | ( n29136 & n29199 ) | ( n29137 & n29199 ) ;
  assign n29201 = x127 & n2429 ;
  assign n29202 = x126 & n2424 ;
  assign n29203 = x125 & ~n2423 ;
  assign n29204 = n2631 & n29203 ;
  assign n29205 = n29202 | n29204 ;
  assign n29206 = n29201 | n29205 ;
  assign n29207 = n2432 | n29201 ;
  assign n29208 = n29205 | n29207 ;
  assign n29209 = ( n18763 & n29206 ) | ( n18763 & n29208 ) | ( n29206 & n29208 ) ;
  assign n29210 = x23 & n29208 ;
  assign n29211 = x23 & n29201 ;
  assign n29212 = ( x23 & n29205 ) | ( x23 & n29211 ) | ( n29205 & n29211 ) ;
  assign n29213 = ( n18763 & n29210 ) | ( n18763 & n29212 ) | ( n29210 & n29212 ) ;
  assign n29214 = x23 & ~n29212 ;
  assign n29215 = x23 & ~n29208 ;
  assign n29216 = ( ~n18763 & n29214 ) | ( ~n18763 & n29215 ) | ( n29214 & n29215 ) ;
  assign n29217 = ( n29209 & ~n29213 ) | ( n29209 & n29216 ) | ( ~n29213 & n29216 ) ;
  assign n29218 = n29133 & n29217 ;
  assign n29219 = ( n29136 & n29217 ) | ( n29136 & n29218 ) | ( n29217 & n29218 ) ;
  assign n29220 = n29134 & n29217 ;
  assign n29221 = n28370 & n29217 ;
  assign n29222 = ( n29135 & n29220 ) | ( n29135 & n29221 ) | ( n29220 & n29221 ) ;
  assign n29223 = ( n29199 & n29219 ) | ( n29199 & n29222 ) | ( n29219 & n29222 ) ;
  assign n29224 = n29200 & ~n29223 ;
  assign n29232 = x85 & n18290 ;
  assign n29233 = x63 & x84 ;
  assign n29234 = ~n18290 & n29233 ;
  assign n29235 = n29232 | n29234 ;
  assign n29236 = ~x20 & n29235 ;
  assign n29237 = x20 & ~n29235 ;
  assign n29238 = n29236 | n29237 ;
  assign n29239 = n28892 & ~n29238 ;
  assign n29240 = ~n28892 & n29238 ;
  assign n29241 = n29239 | n29240 ;
  assign n29242 = x87 & n17141 ;
  assign n29243 = x86 & ~n17140 ;
  assign n29244 = n17724 & n29243 ;
  assign n29245 = n29242 | n29244 ;
  assign n29246 = x88 & n17146 ;
  assign n29247 = n17149 | n29246 ;
  assign n29248 = n29245 | n29247 ;
  assign n29249 = ~x62 & n29248 ;
  assign n29250 = ~x62 & n29246 ;
  assign n29251 = ( ~x62 & n29245 ) | ( ~x62 & n29250 ) | ( n29245 & n29250 ) ;
  assign n29252 = ( ~n3039 & n29249 ) | ( ~n3039 & n29251 ) | ( n29249 & n29251 ) ;
  assign n29253 = n29249 & n29251 ;
  assign n29254 = ( n3023 & n29252 ) | ( n3023 & n29253 ) | ( n29252 & n29253 ) ;
  assign n29255 = x62 & ~n29248 ;
  assign n29256 = x62 & x88 ;
  assign n29257 = n17146 & n29256 ;
  assign n29258 = x62 & ~n29257 ;
  assign n29259 = ~n29245 & n29258 ;
  assign n29260 = ( n3039 & n29255 ) | ( n3039 & n29259 ) | ( n29255 & n29259 ) ;
  assign n29261 = n29255 | n29259 ;
  assign n29262 = ( ~n3023 & n29260 ) | ( ~n3023 & n29261 ) | ( n29260 & n29261 ) ;
  assign n29263 = n29254 | n29262 ;
  assign n29264 = ~n29241 & n29263 ;
  assign n29265 = n29241 & ~n29263 ;
  assign n29266 = n29264 | n29265 ;
  assign n29267 = ~n28893 & n28895 ;
  assign n29268 = ( n28893 & n28912 ) | ( n28893 & ~n29267 ) | ( n28912 & ~n29267 ) ;
  assign n29269 = ~n29266 & n29268 ;
  assign n29270 = n29266 | n29269 ;
  assign n29271 = x91 & n15552 ;
  assign n29272 = x90 & n15547 ;
  assign n29273 = x89 & ~n15546 ;
  assign n29274 = n16123 & n29273 ;
  assign n29275 = n29272 | n29274 ;
  assign n29276 = n29271 | n29275 ;
  assign n29277 = n15555 | n29271 ;
  assign n29278 = n29275 | n29277 ;
  assign n29279 = ( n3768 & n29276 ) | ( n3768 & n29278 ) | ( n29276 & n29278 ) ;
  assign n29280 = x59 & n29278 ;
  assign n29281 = x59 & n29271 ;
  assign n29282 = ( x59 & n29275 ) | ( x59 & n29281 ) | ( n29275 & n29281 ) ;
  assign n29283 = ( n3768 & n29280 ) | ( n3768 & n29282 ) | ( n29280 & n29282 ) ;
  assign n29284 = x59 & ~n29282 ;
  assign n29285 = x59 & ~n29278 ;
  assign n29286 = ( ~n3768 & n29284 ) | ( ~n3768 & n29285 ) | ( n29284 & n29285 ) ;
  assign n29287 = ( n29279 & ~n29283 ) | ( n29279 & n29286 ) | ( ~n29283 & n29286 ) ;
  assign n29288 = n29268 & n29287 ;
  assign n29289 = n29266 & n29288 ;
  assign n29290 = ( ~n29270 & n29287 ) | ( ~n29270 & n29289 ) | ( n29287 & n29289 ) ;
  assign n29291 = n29268 | n29287 ;
  assign n29292 = ( n29266 & n29287 ) | ( n29266 & n29291 ) | ( n29287 & n29291 ) ;
  assign n29293 = n29270 & ~n29292 ;
  assign n29294 = n29290 | n29293 ;
  assign n29295 = n28918 | n28938 ;
  assign n29296 = ( ~n28915 & n28938 ) | ( ~n28915 & n29295 ) | ( n28938 & n29295 ) ;
  assign n29297 = ( n28919 & ~n28921 ) | ( n28919 & n29296 ) | ( ~n28921 & n29296 ) ;
  assign n29298 = n29294 & ~n29297 ;
  assign n29299 = ~n29294 & n29297 ;
  assign n29300 = n29298 | n29299 ;
  assign n29301 = x94 & n14045 ;
  assign n29302 = x93 & n14040 ;
  assign n29303 = x92 & ~n14039 ;
  assign n29304 = n14552 & n29303 ;
  assign n29305 = n29302 | n29304 ;
  assign n29306 = n29301 | n29305 ;
  assign n29307 = n14048 | n29301 ;
  assign n29308 = n29305 | n29307 ;
  assign n29309 = ( n4583 & n29306 ) | ( n4583 & n29308 ) | ( n29306 & n29308 ) ;
  assign n29310 = x56 & n29308 ;
  assign n29311 = x56 & n29301 ;
  assign n29312 = ( x56 & n29305 ) | ( x56 & n29311 ) | ( n29305 & n29311 ) ;
  assign n29313 = ( n4583 & n29310 ) | ( n4583 & n29312 ) | ( n29310 & n29312 ) ;
  assign n29314 = x56 & ~n29312 ;
  assign n29315 = x56 & ~n29308 ;
  assign n29316 = ( ~n4583 & n29314 ) | ( ~n4583 & n29315 ) | ( n29314 & n29315 ) ;
  assign n29317 = ( n29309 & ~n29313 ) | ( n29309 & n29316 ) | ( ~n29313 & n29316 ) ;
  assign n29318 = ~n29300 & n29317 ;
  assign n29319 = n29300 | n29318 ;
  assign n29321 = n28945 | n28964 ;
  assign n29322 = ( n28945 & ~n28947 ) | ( n28945 & n29321 ) | ( ~n28947 & n29321 ) ;
  assign n29320 = n29300 & n29317 ;
  assign n29323 = n29320 & n29322 ;
  assign n29324 = ( ~n29319 & n29322 ) | ( ~n29319 & n29323 ) | ( n29322 & n29323 ) ;
  assign n29325 = n29320 | n29322 ;
  assign n29326 = n29319 & ~n29325 ;
  assign n29327 = n29324 | n29326 ;
  assign n29328 = x97 & n12574 ;
  assign n29329 = x96 & n12569 ;
  assign n29330 = x95 & ~n12568 ;
  assign n29331 = n13076 & n29330 ;
  assign n29332 = n29329 | n29331 ;
  assign n29333 = n29328 | n29332 ;
  assign n29334 = n12577 | n29328 ;
  assign n29335 = n29332 | n29334 ;
  assign n29336 = ( n5505 & n29333 ) | ( n5505 & n29335 ) | ( n29333 & n29335 ) ;
  assign n29337 = x53 & n29335 ;
  assign n29338 = x53 & n29328 ;
  assign n29339 = ( x53 & n29332 ) | ( x53 & n29338 ) | ( n29332 & n29338 ) ;
  assign n29340 = ( n5505 & n29337 ) | ( n5505 & n29339 ) | ( n29337 & n29339 ) ;
  assign n29341 = x53 & ~n29339 ;
  assign n29342 = x53 & ~n29335 ;
  assign n29343 = ( ~n5505 & n29341 ) | ( ~n5505 & n29342 ) | ( n29341 & n29342 ) ;
  assign n29344 = ( n29336 & ~n29340 ) | ( n29336 & n29343 ) | ( ~n29340 & n29343 ) ;
  assign n29345 = n28967 & n28968 ;
  assign n29346 = n28968 | n28987 ;
  assign n29347 = ( ~n28967 & n28987 ) | ( ~n28967 & n29346 ) | ( n28987 & n29346 ) ;
  assign n29348 = ( n28969 & n29345 ) | ( n28969 & n29347 ) | ( n29345 & n29347 ) ;
  assign n29349 = n28969 | n29347 ;
  assign n29350 = ( ~n28970 & n29348 ) | ( ~n28970 & n29349 ) | ( n29348 & n29349 ) ;
  assign n29351 = n29344 & n29350 ;
  assign n29352 = n29344 | n29350 ;
  assign n29353 = ~n29351 & n29352 ;
  assign n29354 = n29327 & n29353 ;
  assign n29355 = n29327 | n29353 ;
  assign n29356 = ~n29354 & n29355 ;
  assign n29357 = x100 & n11205 ;
  assign n29358 = x99 & n11200 ;
  assign n29359 = x98 & ~n11199 ;
  assign n29360 = n11679 & n29359 ;
  assign n29361 = n29358 | n29360 ;
  assign n29362 = n29357 | n29361 ;
  assign n29363 = n11208 | n29357 ;
  assign n29364 = n29361 | n29363 ;
  assign n29365 = ( n6483 & n29362 ) | ( n6483 & n29364 ) | ( n29362 & n29364 ) ;
  assign n29366 = x50 & n29364 ;
  assign n29367 = x50 & n29357 ;
  assign n29368 = ( x50 & n29361 ) | ( x50 & n29367 ) | ( n29361 & n29367 ) ;
  assign n29369 = ( n6483 & n29366 ) | ( n6483 & n29368 ) | ( n29366 & n29368 ) ;
  assign n29370 = x50 & ~n29368 ;
  assign n29371 = x50 & ~n29364 ;
  assign n29372 = ( ~n6483 & n29370 ) | ( ~n6483 & n29371 ) | ( n29370 & n29371 ) ;
  assign n29373 = ( n29365 & ~n29369 ) | ( n29365 & n29372 ) | ( ~n29369 & n29372 ) ;
  assign n29374 = ~n29356 & n29373 ;
  assign n29375 = n29356 & ~n29373 ;
  assign n29376 = n29374 | n29375 ;
  assign n29377 = n28997 | n29016 ;
  assign n29378 = ( n28997 & ~n28999 ) | ( n28997 & n29377 ) | ( ~n28999 & n29377 ) ;
  assign n29379 = n29376 & ~n29378 ;
  assign n29380 = ~n29376 & n29378 ;
  assign n29381 = n29379 | n29380 ;
  assign n29382 = x103 & n9933 ;
  assign n29383 = x102 & n9928 ;
  assign n29384 = x101 & ~n9927 ;
  assign n29385 = n10379 & n29384 ;
  assign n29386 = n29383 | n29385 ;
  assign n29387 = n29382 | n29386 ;
  assign n29388 = n9936 | n29382 ;
  assign n29389 = n29386 | n29388 ;
  assign n29390 = ( n7529 & n29387 ) | ( n7529 & n29389 ) | ( n29387 & n29389 ) ;
  assign n29391 = x47 & n29389 ;
  assign n29392 = x47 & n29382 ;
  assign n29393 = ( x47 & n29386 ) | ( x47 & n29392 ) | ( n29386 & n29392 ) ;
  assign n29394 = ( n7529 & n29391 ) | ( n7529 & n29393 ) | ( n29391 & n29393 ) ;
  assign n29395 = x47 & ~n29393 ;
  assign n29396 = x47 & ~n29389 ;
  assign n29397 = ( ~n7529 & n29395 ) | ( ~n7529 & n29396 ) | ( n29395 & n29396 ) ;
  assign n29398 = ( n29390 & ~n29394 ) | ( n29390 & n29397 ) | ( ~n29394 & n29397 ) ;
  assign n29399 = ~n29381 & n29398 ;
  assign n29400 = n29381 | n29399 ;
  assign n29401 = n29381 & n29398 ;
  assign n29402 = n29019 & ~n29040 ;
  assign n29403 = ( n29020 & n29040 ) | ( n29020 & ~n29402 ) | ( n29040 & ~n29402 ) ;
  assign n29404 = ( n29021 & ~n29023 ) | ( n29021 & n29403 ) | ( ~n29023 & n29403 ) ;
  assign n29405 = n29401 | n29404 ;
  assign n29406 = n29400 & ~n29405 ;
  assign n29407 = n29401 & n29404 ;
  assign n29408 = ( ~n29400 & n29404 ) | ( ~n29400 & n29407 ) | ( n29404 & n29407 ) ;
  assign n29409 = n29406 | n29408 ;
  assign n29410 = x106 & n8724 ;
  assign n29411 = x105 & n8719 ;
  assign n29412 = x104 & ~n8718 ;
  assign n29413 = n9149 & n29412 ;
  assign n29414 = n29411 | n29413 ;
  assign n29415 = n29410 | n29414 ;
  assign n29416 = n8727 | n29410 ;
  assign n29417 = n29414 | n29416 ;
  assign n29418 = ( n8656 & n29415 ) | ( n8656 & n29417 ) | ( n29415 & n29417 ) ;
  assign n29419 = x44 & n29417 ;
  assign n29420 = x44 & n29410 ;
  assign n29421 = ( x44 & n29414 ) | ( x44 & n29420 ) | ( n29414 & n29420 ) ;
  assign n29422 = ( n8656 & n29419 ) | ( n8656 & n29421 ) | ( n29419 & n29421 ) ;
  assign n29423 = x44 & ~n29421 ;
  assign n29424 = x44 & ~n29417 ;
  assign n29425 = ( ~n8656 & n29423 ) | ( ~n8656 & n29424 ) | ( n29423 & n29424 ) ;
  assign n29426 = ( n29418 & ~n29422 ) | ( n29418 & n29425 ) | ( ~n29422 & n29425 ) ;
  assign n29427 = ~n29409 & n29426 ;
  assign n29428 = n29409 | n29427 ;
  assign n29429 = n29409 & n29426 ;
  assign n29430 = n29046 | n29065 ;
  assign n29431 = ( n29046 & ~n29048 ) | ( n29046 & n29430 ) | ( ~n29048 & n29430 ) ;
  assign n29432 = n29429 | n29431 ;
  assign n29433 = n29428 & ~n29432 ;
  assign n29434 = n29429 & n29431 ;
  assign n29435 = ( ~n29428 & n29431 ) | ( ~n29428 & n29434 ) | ( n29431 & n29434 ) ;
  assign n29436 = n29433 | n29435 ;
  assign n29437 = x109 & n7566 ;
  assign n29438 = x108 & n7561 ;
  assign n29439 = x107 & ~n7560 ;
  assign n29440 = n7953 & n29439 ;
  assign n29441 = n29438 | n29440 ;
  assign n29442 = n29437 | n29441 ;
  assign n29443 = n7569 | n29437 ;
  assign n29444 = n29441 | n29443 ;
  assign n29445 = ( n9878 & n29442 ) | ( n9878 & n29444 ) | ( n29442 & n29444 ) ;
  assign n29446 = x41 & n29444 ;
  assign n29447 = x41 & n29437 ;
  assign n29448 = ( x41 & n29441 ) | ( x41 & n29447 ) | ( n29441 & n29447 ) ;
  assign n29449 = ( n9878 & n29446 ) | ( n9878 & n29448 ) | ( n29446 & n29448 ) ;
  assign n29450 = x41 & ~n29448 ;
  assign n29451 = x41 & ~n29444 ;
  assign n29452 = ( ~n9878 & n29450 ) | ( ~n9878 & n29451 ) | ( n29450 & n29451 ) ;
  assign n29453 = ( n29445 & ~n29449 ) | ( n29445 & n29452 ) | ( ~n29449 & n29452 ) ;
  assign n29454 = ~n29436 & n29453 ;
  assign n29455 = n29436 | n29454 ;
  assign n29456 = n29436 & n29453 ;
  assign n29457 = n29455 & ~n29456 ;
  assign n29458 = n29068 & ~n29088 ;
  assign n29459 = ( n28888 & n29088 ) | ( n28888 & ~n29458 ) | ( n29088 & ~n29458 ) ;
  assign n29460 = ( n29069 & ~n29071 ) | ( n29069 & n29459 ) | ( ~n29071 & n29459 ) ;
  assign n29461 = n29457 & ~n29460 ;
  assign n29462 = ~n29457 & n29460 ;
  assign n29463 = n29461 | n29462 ;
  assign n29464 = x112 & n6536 ;
  assign n29465 = x111 & n6531 ;
  assign n29466 = x110 & ~n6530 ;
  assign n29467 = n6871 & n29466 ;
  assign n29468 = n29465 | n29467 ;
  assign n29469 = n29464 | n29468 ;
  assign n29470 = n6539 | n29464 ;
  assign n29471 = n29468 | n29470 ;
  assign n29472 = ( n11172 & n29469 ) | ( n11172 & n29471 ) | ( n29469 & n29471 ) ;
  assign n29473 = x38 & n29471 ;
  assign n29474 = x38 & n29464 ;
  assign n29475 = ( x38 & n29468 ) | ( x38 & n29474 ) | ( n29468 & n29474 ) ;
  assign n29476 = ( n11172 & n29473 ) | ( n11172 & n29475 ) | ( n29473 & n29475 ) ;
  assign n29477 = x38 & ~n29475 ;
  assign n29478 = x38 & ~n29471 ;
  assign n29479 = ( ~n11172 & n29477 ) | ( ~n11172 & n29478 ) | ( n29477 & n29478 ) ;
  assign n29480 = ( n29472 & ~n29476 ) | ( n29472 & n29479 ) | ( ~n29476 & n29479 ) ;
  assign n29481 = ~n29463 & n29480 ;
  assign n29482 = n29463 | n29481 ;
  assign n29484 = n29094 & ~n29114 ;
  assign n29485 = ( n29091 & ~n29114 ) | ( n29091 & n29484 ) | ( ~n29114 & n29484 ) ;
  assign n29486 = ( n29095 & ~n29097 ) | ( n29095 & n29485 ) | ( ~n29097 & n29485 ) ;
  assign n29483 = n29463 & n29480 ;
  assign n29487 = n29483 & ~n29486 ;
  assign n29488 = ( n29482 & n29486 ) | ( n29482 & ~n29487 ) | ( n29486 & ~n29487 ) ;
  assign n29489 = ~n29483 & n29486 ;
  assign n29490 = n29482 & n29489 ;
  assign n29491 = n29488 & ~n29490 ;
  assign n29492 = x115 & n5554 ;
  assign n29493 = x114 & n5549 ;
  assign n29494 = x113 & ~n5548 ;
  assign n29495 = n5893 & n29494 ;
  assign n29496 = n29493 | n29495 ;
  assign n29497 = n29492 | n29496 ;
  assign n29498 = n5557 | n29492 ;
  assign n29499 = n29496 | n29498 ;
  assign n29500 = ( ~n12550 & n29497 ) | ( ~n12550 & n29499 ) | ( n29497 & n29499 ) ;
  assign n29501 = n29497 & n29499 ;
  assign n29502 = ( n12532 & n29500 ) | ( n12532 & n29501 ) | ( n29500 & n29501 ) ;
  assign n29503 = x35 & n29502 ;
  assign n29504 = x35 & ~n29502 ;
  assign n29505 = ( n29502 & ~n29503 ) | ( n29502 & n29504 ) | ( ~n29503 & n29504 ) ;
  assign n29506 = n29491 & n29505 ;
  assign n29507 = n29491 | n29505 ;
  assign n29508 = ~n29506 & n29507 ;
  assign n29509 = n28866 | n29120 ;
  assign n29510 = ( n29120 & n29121 ) | ( n29120 & n29509 ) | ( n29121 & n29509 ) ;
  assign n29511 = n29508 & n29510 ;
  assign n29512 = n29508 & ~n29511 ;
  assign n29513 = ~n29508 & n29510 ;
  assign n29514 = n29512 | n29513 ;
  assign n29515 = x121 & n3816 ;
  assign n29516 = x120 & n3811 ;
  assign n29517 = x119 & ~n3810 ;
  assign n29518 = n4067 & n29517 ;
  assign n29519 = n29516 | n29518 ;
  assign n29520 = n29515 | n29519 ;
  assign n29521 = n3819 | n29515 ;
  assign n29522 = n29519 | n29521 ;
  assign n29523 = ( n15501 & n29520 ) | ( n15501 & n29522 ) | ( n29520 & n29522 ) ;
  assign n29524 = x29 & n29522 ;
  assign n29525 = x29 & n29515 ;
  assign n29526 = ( x29 & n29519 ) | ( x29 & n29525 ) | ( n29519 & n29525 ) ;
  assign n29527 = ( n15501 & n29524 ) | ( n15501 & n29526 ) | ( n29524 & n29526 ) ;
  assign n29528 = x29 & ~n29526 ;
  assign n29529 = x29 & ~n29522 ;
  assign n29530 = ( ~n15501 & n29528 ) | ( ~n15501 & n29529 ) | ( n29528 & n29529 ) ;
  assign n29531 = ( n29523 & ~n29527 ) | ( n29523 & n29530 ) | ( ~n29527 & n29530 ) ;
  assign n29532 = ( n28848 & n28850 ) | ( n28848 & n29122 ) | ( n28850 & n29122 ) ;
  assign n29533 = ( n28848 & n28850 ) | ( n28848 & ~n28866 ) | ( n28850 & ~n28866 ) ;
  assign n29534 = ( n29123 & n29532 ) | ( n29123 & n29533 ) | ( n29532 & n29533 ) ;
  assign n29535 = ~n29531 & n29534 ;
  assign n29536 = n29531 & ~n29534 ;
  assign n29537 = n29535 | n29536 ;
  assign n29538 = x118 & n4631 ;
  assign n29539 = x117 & n4626 ;
  assign n29540 = x116 & ~n4625 ;
  assign n29541 = n4943 & n29540 ;
  assign n29542 = n29539 | n29541 ;
  assign n29543 = n29538 | n29542 ;
  assign n29544 = n4634 | n29538 ;
  assign n29545 = n29542 | n29544 ;
  assign n29546 = ( ~n14002 & n29543 ) | ( ~n14002 & n29545 ) | ( n29543 & n29545 ) ;
  assign n29547 = n29543 & n29545 ;
  assign n29548 = ( n13981 & n29546 ) | ( n13981 & n29547 ) | ( n29546 & n29547 ) ;
  assign n29549 = x32 & n29548 ;
  assign n29550 = x32 & ~n29548 ;
  assign n29551 = ( n29548 & ~n29549 ) | ( n29548 & n29550 ) | ( ~n29549 & n29550 ) ;
  assign n29552 = n28866 & n29121 ;
  assign n29553 = n28866 | n29121 ;
  assign n29554 = ~n29552 & n29553 ;
  assign n29555 = n28883 | n29554 ;
  assign n29556 = ( n28883 & n28887 ) | ( n28883 & n29555 ) | ( n28887 & n29555 ) ;
  assign n29557 = n29551 | n29556 ;
  assign n29558 = n29551 & n29556 ;
  assign n29559 = n29557 & ~n29558 ;
  assign n29560 = ( n29514 & n29537 ) | ( n29514 & ~n29559 ) | ( n29537 & ~n29559 ) ;
  assign n29561 = ( ~n29537 & n29559 ) | ( ~n29537 & n29560 ) | ( n29559 & n29560 ) ;
  assign n29562 = ( ~n29514 & n29560 ) | ( ~n29514 & n29561 ) | ( n29560 & n29561 ) ;
  assign n29563 = n29198 & n29562 ;
  assign n29225 = ~n29133 & n29217 ;
  assign n29226 = ~n29136 & n29225 ;
  assign n29227 = ~n29134 & n29217 ;
  assign n29228 = ~n28370 & n29217 ;
  assign n29229 = ( ~n29135 & n29227 ) | ( ~n29135 & n29228 ) | ( n29227 & n29228 ) ;
  assign n29230 = ( ~n29199 & n29226 ) | ( ~n29199 & n29229 ) | ( n29226 & n29229 ) ;
  assign n29564 = ( n29198 & ~n29230 ) | ( n29198 & n29562 ) | ( ~n29230 & n29562 ) ;
  assign n29565 = ( ~n29224 & n29563 ) | ( ~n29224 & n29564 ) | ( n29563 & n29564 ) ;
  assign n29231 = n29224 | n29230 ;
  assign n29566 = ( n29231 & ~n29562 ) | ( n29231 & n29565 ) | ( ~n29562 & n29565 ) ;
  assign n29567 = ( ~n29198 & n29565 ) | ( ~n29198 & n29566 ) | ( n29565 & n29566 ) ;
  assign n29568 = n28785 | n29145 ;
  assign n29569 = n28785 | n29143 ;
  assign n29570 = ( n28786 & n29568 ) | ( n28786 & n29569 ) | ( n29568 & n29569 ) ;
  assign n29571 = n29567 | n29570 ;
  assign n29572 = n29567 & n29570 ;
  assign n29573 = n29571 & ~n29572 ;
  assign n29574 = n29154 | n29167 ;
  assign n29575 = n29154 | n29156 ;
  assign n29576 = ( n28751 & n29574 ) | ( n28751 & n29575 ) | ( n29574 & n29575 ) ;
  assign n29577 = n29154 | n29169 ;
  assign n29578 = ( n28747 & n29574 ) | ( n28747 & n29577 ) | ( n29574 & n29577 ) ;
  assign n29579 = ( n27383 & n29576 ) | ( n27383 & n29578 ) | ( n29576 & n29578 ) ;
  assign n29580 = n29154 | n29172 ;
  assign n29581 = ( n28753 & n29574 ) | ( n28753 & n29575 ) | ( n29574 & n29575 ) ;
  assign n29582 = ( n28312 & n29580 ) | ( n28312 & n29581 ) | ( n29580 & n29581 ) ;
  assign n29583 = ( n26030 & n29579 ) | ( n26030 & n29582 ) | ( n29579 & n29582 ) ;
  assign n29584 = n29573 | n29583 ;
  assign n29585 = n29573 & n29579 ;
  assign n29586 = n29573 & n29581 ;
  assign n29587 = n29154 & n29573 ;
  assign n29588 = ( n29172 & n29573 ) | ( n29172 & n29587 ) | ( n29573 & n29587 ) ;
  assign n29589 = ( n28312 & n29586 ) | ( n28312 & n29588 ) | ( n29586 & n29588 ) ;
  assign n29590 = ( n26030 & n29585 ) | ( n26030 & n29589 ) | ( n29585 & n29589 ) ;
  assign n29591 = n29584 & ~n29590 ;
  assign n29592 = n29327 & ~n29344 ;
  assign n29593 = ( n29327 & ~n29350 ) | ( n29327 & n29592 ) | ( ~n29350 & n29592 ) ;
  assign n29594 = ( n29351 & n29353 ) | ( n29351 & ~n29593 ) | ( n29353 & ~n29593 ) ;
  assign n29595 = n29318 | n29324 ;
  assign n29596 = x86 & n18290 ;
  assign n29597 = x63 & x85 ;
  assign n29598 = ~n18290 & n29597 ;
  assign n29599 = n29596 | n29598 ;
  assign n29600 = n28892 | n29236 ;
  assign n29601 = ( n29236 & ~n29238 ) | ( n29236 & n29600 ) | ( ~n29238 & n29600 ) ;
  assign n29602 = n29599 & ~n29601 ;
  assign n29603 = ~n29599 & n29601 ;
  assign n29604 = n29602 | n29603 ;
  assign n29606 = x88 & n17141 ;
  assign n29607 = x87 & ~n17140 ;
  assign n29608 = n17724 & n29607 ;
  assign n29609 = n29606 | n29608 ;
  assign n29605 = x89 & n17146 ;
  assign n29611 = n17149 | n29605 ;
  assign n29612 = n29609 | n29611 ;
  assign n29610 = n29605 | n29609 ;
  assign n29613 = n29610 & n29612 ;
  assign n29614 = ( n3282 & n29612 ) | ( n3282 & n29613 ) | ( n29612 & n29613 ) ;
  assign n29615 = x62 & n29613 ;
  assign n29616 = x62 & n29612 ;
  assign n29617 = ( n3282 & n29615 ) | ( n3282 & n29616 ) | ( n29615 & n29616 ) ;
  assign n29618 = x62 & ~n29613 ;
  assign n29619 = x62 & ~n29612 ;
  assign n29620 = ( ~n3282 & n29618 ) | ( ~n3282 & n29619 ) | ( n29618 & n29619 ) ;
  assign n29621 = ( n29614 & ~n29617 ) | ( n29614 & n29620 ) | ( ~n29617 & n29620 ) ;
  assign n29622 = ~n29604 & n29621 ;
  assign n29623 = n29604 & ~n29621 ;
  assign n29624 = n29622 | n29623 ;
  assign n29625 = n29264 | n29268 ;
  assign n29626 = ( n29264 & ~n29266 ) | ( n29264 & n29625 ) | ( ~n29266 & n29625 ) ;
  assign n29627 = ~n29624 & n29626 ;
  assign n29628 = n29624 & ~n29626 ;
  assign n29629 = n29627 | n29628 ;
  assign n29630 = x92 & n15552 ;
  assign n29631 = x91 & n15547 ;
  assign n29632 = x90 & ~n15546 ;
  assign n29633 = n16123 & n29632 ;
  assign n29634 = n29631 | n29633 ;
  assign n29635 = n29630 | n29634 ;
  assign n29636 = n15555 | n29630 ;
  assign n29637 = n29634 | n29636 ;
  assign n29638 = ( n4040 & n29635 ) | ( n4040 & n29637 ) | ( n29635 & n29637 ) ;
  assign n29639 = x59 & n29637 ;
  assign n29640 = x59 & n29630 ;
  assign n29641 = ( x59 & n29634 ) | ( x59 & n29640 ) | ( n29634 & n29640 ) ;
  assign n29642 = ( n4040 & n29639 ) | ( n4040 & n29641 ) | ( n29639 & n29641 ) ;
  assign n29643 = x59 & ~n29641 ;
  assign n29644 = x59 & ~n29637 ;
  assign n29645 = ( ~n4040 & n29643 ) | ( ~n4040 & n29644 ) | ( n29643 & n29644 ) ;
  assign n29646 = ( n29638 & ~n29642 ) | ( n29638 & n29645 ) | ( ~n29642 & n29645 ) ;
  assign n29647 = ~n29629 & n29646 ;
  assign n29648 = n29629 & ~n29646 ;
  assign n29649 = n29647 | n29648 ;
  assign n29650 = n29290 | n29297 ;
  assign n29651 = ( n29290 & ~n29294 ) | ( n29290 & n29650 ) | ( ~n29294 & n29650 ) ;
  assign n29652 = ~n29649 & n29651 ;
  assign n29653 = n29649 & ~n29651 ;
  assign n29654 = n29652 | n29653 ;
  assign n29655 = x95 & n14045 ;
  assign n29656 = x94 & n14040 ;
  assign n29657 = x93 & ~n14039 ;
  assign n29658 = n14552 & n29657 ;
  assign n29659 = n29656 | n29658 ;
  assign n29660 = n29655 | n29659 ;
  assign n29661 = n14048 | n29655 ;
  assign n29662 = n29659 | n29661 ;
  assign n29663 = ( n4897 & n29660 ) | ( n4897 & n29662 ) | ( n29660 & n29662 ) ;
  assign n29664 = x56 & n29662 ;
  assign n29665 = x56 & n29655 ;
  assign n29666 = ( x56 & n29659 ) | ( x56 & n29665 ) | ( n29659 & n29665 ) ;
  assign n29667 = ( n4897 & n29664 ) | ( n4897 & n29666 ) | ( n29664 & n29666 ) ;
  assign n29668 = x56 & ~n29666 ;
  assign n29669 = x56 & ~n29662 ;
  assign n29670 = ( ~n4897 & n29668 ) | ( ~n4897 & n29669 ) | ( n29668 & n29669 ) ;
  assign n29671 = ( n29663 & ~n29667 ) | ( n29663 & n29670 ) | ( ~n29667 & n29670 ) ;
  assign n29672 = n29654 | n29671 ;
  assign n29673 = n29654 & ~n29671 ;
  assign n29674 = ( ~n29654 & n29672 ) | ( ~n29654 & n29673 ) | ( n29672 & n29673 ) ;
  assign n29675 = ~n29595 & n29674 ;
  assign n29676 = n29595 & ~n29674 ;
  assign n29677 = n29675 | n29676 ;
  assign n29678 = x98 & n12574 ;
  assign n29679 = x97 & n12569 ;
  assign n29680 = x96 & ~n12568 ;
  assign n29681 = n13076 & n29680 ;
  assign n29682 = n29679 | n29681 ;
  assign n29683 = n29678 | n29682 ;
  assign n29684 = n12577 | n29678 ;
  assign n29685 = n29682 | n29684 ;
  assign n29686 = ( ~n5850 & n29683 ) | ( ~n5850 & n29685 ) | ( n29683 & n29685 ) ;
  assign n29687 = n29683 & n29685 ;
  assign n29688 = ( n5834 & n29686 ) | ( n5834 & n29687 ) | ( n29686 & n29687 ) ;
  assign n29689 = x53 & n29685 ;
  assign n29690 = x53 & n29678 ;
  assign n29691 = ( x53 & n29682 ) | ( x53 & n29690 ) | ( n29682 & n29690 ) ;
  assign n29692 = ( ~n5850 & n29689 ) | ( ~n5850 & n29691 ) | ( n29689 & n29691 ) ;
  assign n29693 = n29689 & n29691 ;
  assign n29694 = ( n5834 & n29692 ) | ( n5834 & n29693 ) | ( n29692 & n29693 ) ;
  assign n29695 = x53 & ~n29691 ;
  assign n29696 = x53 & ~n29685 ;
  assign n29697 = ( n5850 & n29695 ) | ( n5850 & n29696 ) | ( n29695 & n29696 ) ;
  assign n29698 = n29695 | n29696 ;
  assign n29699 = ( ~n5834 & n29697 ) | ( ~n5834 & n29698 ) | ( n29697 & n29698 ) ;
  assign n29700 = ( n29688 & ~n29694 ) | ( n29688 & n29699 ) | ( ~n29694 & n29699 ) ;
  assign n29701 = n29677 & n29700 ;
  assign n29702 = n29594 & n29701 ;
  assign n29703 = n29674 & ~n29700 ;
  assign n29704 = ( n29595 & n29700 ) | ( n29595 & ~n29703 ) | ( n29700 & ~n29703 ) ;
  assign n29705 = n29675 | n29704 ;
  assign n29706 = ( n29594 & n29702 ) | ( n29594 & ~n29705 ) | ( n29702 & ~n29705 ) ;
  assign n29707 = x101 & n11205 ;
  assign n29708 = x100 & n11200 ;
  assign n29709 = x99 & ~n11199 ;
  assign n29710 = n11679 & n29709 ;
  assign n29711 = n29708 | n29710 ;
  assign n29712 = n29707 | n29711 ;
  assign n29713 = n11208 | n29707 ;
  assign n29714 = n29711 | n29713 ;
  assign n29715 = ( n6844 & n29712 ) | ( n6844 & n29714 ) | ( n29712 & n29714 ) ;
  assign n29716 = x50 & n29714 ;
  assign n29717 = x50 & n29707 ;
  assign n29718 = ( x50 & n29711 ) | ( x50 & n29717 ) | ( n29711 & n29717 ) ;
  assign n29719 = ( n6844 & n29716 ) | ( n6844 & n29718 ) | ( n29716 & n29718 ) ;
  assign n29720 = x50 & ~n29718 ;
  assign n29721 = x50 & ~n29714 ;
  assign n29722 = ( ~n6844 & n29720 ) | ( ~n6844 & n29721 ) | ( n29720 & n29721 ) ;
  assign n29723 = ( n29715 & ~n29719 ) | ( n29715 & n29722 ) | ( ~n29719 & n29722 ) ;
  assign n29724 = ~n29701 & n29705 ;
  assign n29725 = ~n29594 & n29724 ;
  assign n29726 = ~n29723 & n29725 ;
  assign n29727 = ( n29706 & ~n29723 ) | ( n29706 & n29726 ) | ( ~n29723 & n29726 ) ;
  assign n29728 = n29723 & ~n29725 ;
  assign n29729 = ~n29706 & n29728 ;
  assign n29730 = n29727 | n29729 ;
  assign n29731 = n29374 | n29378 ;
  assign n29732 = ( n29374 & ~n29376 ) | ( n29374 & n29731 ) | ( ~n29376 & n29731 ) ;
  assign n29733 = n29730 & n29732 ;
  assign n29734 = ~n29730 & n29732 ;
  assign n29735 = x104 & n9933 ;
  assign n29736 = x103 & n9928 ;
  assign n29737 = x102 & ~n9927 ;
  assign n29738 = n10379 & n29737 ;
  assign n29739 = n29736 | n29738 ;
  assign n29740 = n29735 | n29739 ;
  assign n29741 = n9936 | n29735 ;
  assign n29742 = n29739 | n29741 ;
  assign n29743 = ( n7911 & n29740 ) | ( n7911 & n29742 ) | ( n29740 & n29742 ) ;
  assign n29744 = x47 & n29742 ;
  assign n29745 = x47 & n29735 ;
  assign n29746 = ( x47 & n29739 ) | ( x47 & n29745 ) | ( n29739 & n29745 ) ;
  assign n29747 = ( n7911 & n29744 ) | ( n7911 & n29746 ) | ( n29744 & n29746 ) ;
  assign n29748 = x47 & ~n29746 ;
  assign n29749 = x47 & ~n29742 ;
  assign n29750 = ( ~n7911 & n29748 ) | ( ~n7911 & n29749 ) | ( n29748 & n29749 ) ;
  assign n29751 = ( n29743 & ~n29747 ) | ( n29743 & n29750 ) | ( ~n29747 & n29750 ) ;
  assign n29752 = n29730 & ~n29751 ;
  assign n29753 = ( n29734 & ~n29751 ) | ( n29734 & n29752 ) | ( ~n29751 & n29752 ) ;
  assign n29754 = ~n29733 & n29753 ;
  assign n29755 = n29730 | n29734 ;
  assign n29756 = n29733 & n29751 ;
  assign n29757 = ( n29751 & ~n29755 ) | ( n29751 & n29756 ) | ( ~n29755 & n29756 ) ;
  assign n29758 = n29754 | n29757 ;
  assign n29759 = n29399 | n29408 ;
  assign n29760 = ~n29758 & n29759 ;
  assign n29761 = n29758 & ~n29759 ;
  assign n29762 = n29760 | n29761 ;
  assign n29763 = x107 & n8724 ;
  assign n29764 = x106 & n8719 ;
  assign n29765 = x105 & ~n8718 ;
  assign n29766 = n9149 & n29765 ;
  assign n29767 = n29764 | n29766 ;
  assign n29768 = n29763 | n29767 ;
  assign n29769 = n8727 | n29763 ;
  assign n29770 = n29767 | n29769 ;
  assign n29771 = ( n9084 & n29768 ) | ( n9084 & n29770 ) | ( n29768 & n29770 ) ;
  assign n29772 = x44 & n29770 ;
  assign n29773 = x44 & n29763 ;
  assign n29774 = ( x44 & n29767 ) | ( x44 & n29773 ) | ( n29767 & n29773 ) ;
  assign n29775 = ( n9084 & n29772 ) | ( n9084 & n29774 ) | ( n29772 & n29774 ) ;
  assign n29776 = x44 & ~n29774 ;
  assign n29777 = x44 & ~n29770 ;
  assign n29778 = ( ~n9084 & n29776 ) | ( ~n9084 & n29777 ) | ( n29776 & n29777 ) ;
  assign n29779 = ( n29771 & ~n29775 ) | ( n29771 & n29778 ) | ( ~n29775 & n29778 ) ;
  assign n29780 = n29762 | n29779 ;
  assign n29781 = n29762 & ~n29779 ;
  assign n29782 = ( ~n29762 & n29780 ) | ( ~n29762 & n29781 ) | ( n29780 & n29781 ) ;
  assign n29783 = n29427 | n29435 ;
  assign n29784 = n29782 & ~n29783 ;
  assign n29785 = ~n29782 & n29783 ;
  assign n29786 = n29784 | n29785 ;
  assign n29787 = x110 & n7566 ;
  assign n29788 = x109 & n7561 ;
  assign n29789 = x108 & ~n7560 ;
  assign n29790 = n7953 & n29789 ;
  assign n29791 = n29788 | n29790 ;
  assign n29792 = n29787 | n29791 ;
  assign n29793 = n7569 | n29787 ;
  assign n29794 = n29791 | n29793 ;
  assign n29795 = ( n10330 & n29792 ) | ( n10330 & n29794 ) | ( n29792 & n29794 ) ;
  assign n29796 = x41 & n29794 ;
  assign n29797 = x41 & n29787 ;
  assign n29798 = ( x41 & n29791 ) | ( x41 & n29797 ) | ( n29791 & n29797 ) ;
  assign n29799 = ( n10330 & n29796 ) | ( n10330 & n29798 ) | ( n29796 & n29798 ) ;
  assign n29800 = x41 & ~n29798 ;
  assign n29801 = x41 & ~n29794 ;
  assign n29802 = ( ~n10330 & n29800 ) | ( ~n10330 & n29801 ) | ( n29800 & n29801 ) ;
  assign n29803 = ( n29795 & ~n29799 ) | ( n29795 & n29802 ) | ( ~n29799 & n29802 ) ;
  assign n29804 = n29786 & n29803 ;
  assign n29805 = n29785 | n29803 ;
  assign n29806 = n29784 | n29805 ;
  assign n29807 = ~n29804 & n29806 ;
  assign n29808 = n29454 | n29460 ;
  assign n29809 = ( n29454 & ~n29457 ) | ( n29454 & n29808 ) | ( ~n29457 & n29808 ) ;
  assign n29810 = n29807 & ~n29809 ;
  assign n29811 = ~n29807 & n29809 ;
  assign n29812 = n29810 | n29811 ;
  assign n29813 = x113 & n6536 ;
  assign n29814 = x112 & n6531 ;
  assign n29815 = x111 & ~n6530 ;
  assign n29816 = n6871 & n29815 ;
  assign n29817 = n29814 | n29816 ;
  assign n29818 = n29813 | n29817 ;
  assign n29819 = n6539 | n29813 ;
  assign n29820 = n29817 | n29819 ;
  assign n29821 = ( ~n11642 & n29818 ) | ( ~n11642 & n29820 ) | ( n29818 & n29820 ) ;
  assign n29822 = n29818 & n29820 ;
  assign n29823 = ( n11626 & n29821 ) | ( n11626 & n29822 ) | ( n29821 & n29822 ) ;
  assign n29824 = x38 & n29823 ;
  assign n29825 = x38 & ~n29823 ;
  assign n29826 = ( n29823 & ~n29824 ) | ( n29823 & n29825 ) | ( ~n29824 & n29825 ) ;
  assign n29827 = n29812 & n29826 ;
  assign n29828 = n29811 | n29826 ;
  assign n29829 = n29810 | n29828 ;
  assign n29830 = ~n29827 & n29829 ;
  assign n29831 = ~n29481 & n29488 ;
  assign n29832 = n29830 & n29831 ;
  assign n29833 = n29830 | n29831 ;
  assign n29834 = ~n29832 & n29833 ;
  assign n29835 = x116 & n5554 ;
  assign n29836 = x115 & n5549 ;
  assign n29837 = x114 & ~n5548 ;
  assign n29838 = n5893 & n29837 ;
  assign n29839 = n29836 | n29838 ;
  assign n29840 = n29835 | n29839 ;
  assign n29841 = n5557 | n29835 ;
  assign n29842 = n29839 | n29841 ;
  assign n29843 = ( ~n13040 & n29840 ) | ( ~n13040 & n29842 ) | ( n29840 & n29842 ) ;
  assign n29844 = n29840 & n29842 ;
  assign n29845 = ( n13022 & n29843 ) | ( n13022 & n29844 ) | ( n29843 & n29844 ) ;
  assign n29846 = x35 & n29845 ;
  assign n29847 = x35 & ~n29845 ;
  assign n29848 = ( n29845 & ~n29846 ) | ( n29845 & n29847 ) | ( ~n29846 & n29847 ) ;
  assign n29849 = ~n29834 & n29848 ;
  assign n29850 = n29830 & ~n29848 ;
  assign n29851 = ( n29831 & ~n29848 ) | ( n29831 & n29850 ) | ( ~n29848 & n29850 ) ;
  assign n29852 = ~n29832 & n29851 ;
  assign n29853 = n29849 | n29852 ;
  assign n29855 = x121 & n3811 ;
  assign n29856 = x120 & ~n3810 ;
  assign n29857 = n4067 & n29856 ;
  assign n29858 = n29855 | n29857 ;
  assign n29854 = x122 & n3816 ;
  assign n29860 = n3819 | n29854 ;
  assign n29861 = n29858 | n29860 ;
  assign n29859 = n29854 | n29858 ;
  assign n29862 = n29859 & n29861 ;
  assign n29863 = ( n16043 & n29861 ) | ( n16043 & n29862 ) | ( n29861 & n29862 ) ;
  assign n29864 = x29 & n29862 ;
  assign n29865 = x29 & n29861 ;
  assign n29866 = ( n16043 & n29864 ) | ( n16043 & n29865 ) | ( n29864 & n29865 ) ;
  assign n29867 = x29 & ~n29862 ;
  assign n29868 = x29 & ~n29861 ;
  assign n29869 = ( ~n16043 & n29867 ) | ( ~n16043 & n29868 ) | ( n29867 & n29868 ) ;
  assign n29870 = ( n29863 & ~n29866 ) | ( n29863 & n29869 ) | ( ~n29866 & n29869 ) ;
  assign n29871 = n29514 | n29558 ;
  assign n29872 = ( n29558 & n29559 ) | ( n29558 & n29871 ) | ( n29559 & n29871 ) ;
  assign n29873 = n29870 & n29872 ;
  assign n29874 = n29870 | n29872 ;
  assign n29875 = ~n29873 & n29874 ;
  assign n29893 = n29506 | n29510 ;
  assign n29894 = ( n29506 & n29508 ) | ( n29506 & n29893 ) | ( n29508 & n29893 ) ;
  assign n29876 = x119 & n4631 ;
  assign n29877 = x118 & n4626 ;
  assign n29878 = x117 & ~n4625 ;
  assign n29879 = n4943 & n29878 ;
  assign n29880 = n29877 | n29879 ;
  assign n29881 = n29876 | n29880 ;
  assign n29882 = n4634 | n29876 ;
  assign n29883 = n29880 | n29882 ;
  assign n29884 = ( n14496 & n29881 ) | ( n14496 & n29883 ) | ( n29881 & n29883 ) ;
  assign n29885 = x32 & n29883 ;
  assign n29886 = x32 & n29876 ;
  assign n29887 = ( x32 & n29880 ) | ( x32 & n29886 ) | ( n29880 & n29886 ) ;
  assign n29888 = ( n14496 & n29885 ) | ( n14496 & n29887 ) | ( n29885 & n29887 ) ;
  assign n29889 = x32 & ~n29887 ;
  assign n29890 = x32 & ~n29883 ;
  assign n29891 = ( ~n14496 & n29889 ) | ( ~n14496 & n29890 ) | ( n29889 & n29890 ) ;
  assign n29892 = ( n29884 & ~n29888 ) | ( n29884 & n29891 ) | ( ~n29888 & n29891 ) ;
  assign n29895 = n29892 | n29894 ;
  assign n29896 = ~n29892 & n29894 ;
  assign n29897 = ( ~n29894 & n29895 ) | ( ~n29894 & n29896 ) | ( n29895 & n29896 ) ;
  assign n29898 = ( n29853 & n29875 ) | ( n29853 & ~n29897 ) | ( n29875 & ~n29897 ) ;
  assign n29899 = ( ~n29875 & n29897 ) | ( ~n29875 & n29898 ) | ( n29897 & n29898 ) ;
  assign n29900 = ( ~n29853 & n29898 ) | ( ~n29853 & n29899 ) | ( n29898 & n29899 ) ;
  assign n29901 = x127 & n2424 ;
  assign n29902 = x126 & ~n2423 ;
  assign n29903 = n2631 & n29902 ;
  assign n29904 = n29901 | n29903 ;
  assign n29905 = n2432 | n29904 ;
  assign n29906 = ( n19328 & n29904 ) | ( n19328 & n29905 ) | ( n29904 & n29905 ) ;
  assign n29907 = x23 & n29904 ;
  assign n29908 = ( x23 & n4112 ) | ( x23 & n29904 ) | ( n4112 & n29904 ) ;
  assign n29909 = ( n19328 & n29907 ) | ( n19328 & n29908 ) | ( n29907 & n29908 ) ;
  assign n29910 = x23 & ~n4112 ;
  assign n29911 = ~n29904 & n29910 ;
  assign n29912 = x23 & ~n29904 ;
  assign n29913 = ( ~n19328 & n29911 ) | ( ~n19328 & n29912 ) | ( n29911 & n29912 ) ;
  assign n29914 = ( n29906 & ~n29909 ) | ( n29906 & n29913 ) | ( ~n29909 & n29913 ) ;
  assign n29915 = n29197 | n29562 ;
  assign n29916 = ( n29197 & n29198 ) | ( n29197 & n29915 ) | ( n29198 & n29915 ) ;
  assign n29917 = n29914 & n29916 ;
  assign n29918 = n29914 | n29916 ;
  assign n29919 = ~n29917 & n29918 ;
  assign n29920 = n29514 & n29559 ;
  assign n29921 = n29514 | n29559 ;
  assign n29922 = ~n29920 & n29921 ;
  assign n29923 = x125 & n3085 ;
  assign n29924 = x124 & n3080 ;
  assign n29925 = x123 & ~n3079 ;
  assign n29926 = n3309 & n29925 ;
  assign n29927 = n29924 | n29926 ;
  assign n29928 = n29923 | n29927 ;
  assign n29929 = n3088 | n29923 ;
  assign n29930 = n29927 | n29929 ;
  assign n29931 = ( n17670 & n29928 ) | ( n17670 & n29930 ) | ( n29928 & n29930 ) ;
  assign n29932 = x26 & n29930 ;
  assign n29933 = x26 & n29923 ;
  assign n29934 = ( x26 & n29927 ) | ( x26 & n29933 ) | ( n29927 & n29933 ) ;
  assign n29935 = ( n17670 & n29932 ) | ( n17670 & n29934 ) | ( n29932 & n29934 ) ;
  assign n29936 = x26 & ~n29934 ;
  assign n29937 = x26 & ~n29930 ;
  assign n29938 = ( ~n17670 & n29936 ) | ( ~n17670 & n29937 ) | ( n29936 & n29937 ) ;
  assign n29939 = ( n29931 & ~n29935 ) | ( n29931 & n29938 ) | ( ~n29935 & n29938 ) ;
  assign n29940 = n29534 & n29939 ;
  assign n29941 = n29531 & n29939 ;
  assign n29942 = ( n29922 & n29940 ) | ( n29922 & n29941 ) | ( n29940 & n29941 ) ;
  assign n29943 = n29534 | n29939 ;
  assign n29944 = n29531 | n29939 ;
  assign n29945 = ( n29922 & n29943 ) | ( n29922 & n29944 ) | ( n29943 & n29944 ) ;
  assign n29946 = ~n29942 & n29945 ;
  assign n29947 = ( n29900 & n29919 ) | ( n29900 & ~n29946 ) | ( n29919 & ~n29946 ) ;
  assign n29948 = ( ~n29919 & n29946 ) | ( ~n29919 & n29947 ) | ( n29946 & n29947 ) ;
  assign n29949 = ( ~n29900 & n29947 ) | ( ~n29900 & n29948 ) | ( n29947 & n29948 ) ;
  assign n29950 = n29198 | n29562 ;
  assign n29951 = n29230 & n29950 ;
  assign n29952 = ( n29224 & n29950 ) | ( n29224 & n29951 ) | ( n29950 & n29951 ) ;
  assign n29953 = ~n29223 & n29563 ;
  assign n29954 = ( n29223 & n29952 ) | ( n29223 & ~n29953 ) | ( n29952 & ~n29953 ) ;
  assign n29955 = n29949 | n29954 ;
  assign n29956 = n29949 & n29954 ;
  assign n29957 = n29955 & ~n29956 ;
  assign n29958 = n29572 | n29573 ;
  assign n29959 = ( n29572 & n29579 ) | ( n29572 & n29958 ) | ( n29579 & n29958 ) ;
  assign n29960 = n29572 | n29587 ;
  assign n29961 = ( n29172 & n29958 ) | ( n29172 & n29960 ) | ( n29958 & n29960 ) ;
  assign n29962 = ( n29572 & n29581 ) | ( n29572 & n29958 ) | ( n29581 & n29958 ) ;
  assign n29963 = ( n28312 & n29961 ) | ( n28312 & n29962 ) | ( n29961 & n29962 ) ;
  assign n29964 = ( n26030 & n29959 ) | ( n26030 & n29963 ) | ( n29959 & n29963 ) ;
  assign n29965 = n29957 | n29964 ;
  assign n29966 = n29572 & n29957 ;
  assign n29967 = ( n29573 & n29957 ) | ( n29573 & n29966 ) | ( n29957 & n29966 ) ;
  assign n29968 = ( n29579 & n29966 ) | ( n29579 & n29967 ) | ( n29966 & n29967 ) ;
  assign n29969 = n29957 & n29960 ;
  assign n29970 = n29957 & n29958 ;
  assign n29971 = ( n29172 & n29969 ) | ( n29172 & n29970 ) | ( n29969 & n29970 ) ;
  assign n29972 = ( n29581 & n29966 ) | ( n29581 & n29970 ) | ( n29966 & n29970 ) ;
  assign n29973 = ( n28312 & n29971 ) | ( n28312 & n29972 ) | ( n29971 & n29972 ) ;
  assign n29974 = ( n26030 & n29968 ) | ( n26030 & n29973 ) | ( n29968 & n29973 ) ;
  assign n29975 = n29965 & ~n29974 ;
  assign n29976 = n29898 & n29946 ;
  assign n29977 = ~n29853 & n29946 ;
  assign n29978 = ( n29899 & n29976 ) | ( n29899 & n29977 ) | ( n29976 & n29977 ) ;
  assign n29979 = n29898 | n29946 ;
  assign n29980 = n29853 & ~n29946 ;
  assign n29981 = ( n29899 & n29979 ) | ( n29899 & ~n29980 ) | ( n29979 & ~n29980 ) ;
  assign n29982 = ~n29978 & n29981 ;
  assign n29983 = n29914 | n29982 ;
  assign n29984 = ( n29916 & n29982 ) | ( n29916 & n29983 ) | ( n29982 & n29983 ) ;
  assign n29985 = ( n29917 & n29919 ) | ( n29917 & n29984 ) | ( n29919 & n29984 ) ;
  assign n29986 = x126 & n3085 ;
  assign n29987 = x125 & n3080 ;
  assign n29988 = x124 & ~n3079 ;
  assign n29989 = n3309 & n29988 ;
  assign n29990 = n29987 | n29989 ;
  assign n29991 = n29986 | n29990 ;
  assign n29992 = n3088 | n29986 ;
  assign n29993 = n29990 | n29992 ;
  assign n29994 = ( n18220 & n29991 ) | ( n18220 & n29993 ) | ( n29991 & n29993 ) ;
  assign n29995 = x26 & n29993 ;
  assign n29996 = x26 & n29986 ;
  assign n29997 = ( x26 & n29990 ) | ( x26 & n29996 ) | ( n29990 & n29996 ) ;
  assign n29998 = ( n18220 & n29995 ) | ( n18220 & n29997 ) | ( n29995 & n29997 ) ;
  assign n29999 = x26 & ~n29997 ;
  assign n30000 = x26 & ~n29993 ;
  assign n30001 = ( ~n18220 & n29999 ) | ( ~n18220 & n30000 ) | ( n29999 & n30000 ) ;
  assign n30002 = ( n29994 & ~n29998 ) | ( n29994 & n30001 ) | ( ~n29998 & n30001 ) ;
  assign n30003 = n29853 & n29897 ;
  assign n30004 = n29853 | n29897 ;
  assign n30005 = ~n30003 & n30004 ;
  assign n30006 = n29870 | n30005 ;
  assign n30007 = ( n29872 & n30005 ) | ( n29872 & n30006 ) | ( n30005 & n30006 ) ;
  assign n30008 = n30002 & n30007 ;
  assign n30009 = n29873 & n30002 ;
  assign n30010 = ( n29875 & n30008 ) | ( n29875 & n30009 ) | ( n30008 & n30009 ) ;
  assign n30011 = n30002 | n30007 ;
  assign n30012 = n29873 | n30002 ;
  assign n30013 = ( n29875 & n30011 ) | ( n29875 & n30012 ) | ( n30011 & n30012 ) ;
  assign n30014 = ~n30010 & n30013 ;
  assign n30015 = x123 & n3816 ;
  assign n30016 = x122 & n3811 ;
  assign n30017 = x121 & ~n3810 ;
  assign n30018 = n4067 & n30017 ;
  assign n30019 = n30016 | n30018 ;
  assign n30020 = n30015 | n30019 ;
  assign n30021 = n3819 | n30015 ;
  assign n30022 = n30019 | n30021 ;
  assign n30023 = ( n16086 & n30020 ) | ( n16086 & n30022 ) | ( n30020 & n30022 ) ;
  assign n30024 = x29 & n30022 ;
  assign n30025 = x29 & n30015 ;
  assign n30026 = ( x29 & n30019 ) | ( x29 & n30025 ) | ( n30019 & n30025 ) ;
  assign n30027 = ( n16086 & n30024 ) | ( n16086 & n30026 ) | ( n30024 & n30026 ) ;
  assign n30028 = x29 & ~n30026 ;
  assign n30029 = x29 & ~n30022 ;
  assign n30030 = ( ~n16086 & n30028 ) | ( ~n16086 & n30029 ) | ( n30028 & n30029 ) ;
  assign n30031 = ( n30023 & ~n30027 ) | ( n30023 & n30030 ) | ( ~n30027 & n30030 ) ;
  assign n30032 = ( n29506 & n29510 ) | ( n29506 & n29892 ) | ( n29510 & n29892 ) ;
  assign n30033 = n29505 & n29892 ;
  assign n30034 = n29491 & n30033 ;
  assign n30035 = ( n29508 & n30032 ) | ( n29508 & n30034 ) | ( n30032 & n30034 ) ;
  assign n30036 = n29853 | n30035 ;
  assign n30037 = ( n29897 & n30035 ) | ( n29897 & n30036 ) | ( n30035 & n30036 ) ;
  assign n30038 = ~n30031 & n30037 ;
  assign n30039 = x120 & n4631 ;
  assign n30040 = x119 & n4626 ;
  assign n30041 = x118 & ~n4625 ;
  assign n30042 = n4943 & n30041 ;
  assign n30043 = n30040 | n30042 ;
  assign n30044 = n30039 | n30043 ;
  assign n30045 = n4634 | n30039 ;
  assign n30046 = n30043 | n30045 ;
  assign n30047 = ( n14991 & n30044 ) | ( n14991 & n30046 ) | ( n30044 & n30046 ) ;
  assign n30048 = x32 & n30046 ;
  assign n30049 = x32 & n30039 ;
  assign n30050 = ( x32 & n30043 ) | ( x32 & n30049 ) | ( n30043 & n30049 ) ;
  assign n30051 = ( n14991 & n30048 ) | ( n14991 & n30050 ) | ( n30048 & n30050 ) ;
  assign n30052 = x32 & ~n30050 ;
  assign n30053 = x32 & ~n30046 ;
  assign n30054 = ( ~n14991 & n30052 ) | ( ~n14991 & n30053 ) | ( n30052 & n30053 ) ;
  assign n30055 = ( n30047 & ~n30051 ) | ( n30047 & n30054 ) | ( ~n30051 & n30054 ) ;
  assign n30056 = ~n29851 & n30055 ;
  assign n30057 = ~n29833 & n30055 ;
  assign n30058 = ( n29834 & n30056 ) | ( n29834 & n30057 ) | ( n30056 & n30057 ) ;
  assign n30059 = n29851 & ~n30055 ;
  assign n30060 = n29833 & ~n30055 ;
  assign n30061 = ( ~n29834 & n30059 ) | ( ~n29834 & n30060 ) | ( n30059 & n30060 ) ;
  assign n30062 = n30058 | n30061 ;
  assign n30281 = ( n29811 & ~n29812 ) | ( n29811 & n29828 ) | ( ~n29812 & n29828 ) ;
  assign n30063 = n29734 | n29757 ;
  assign n30064 = x105 & n9933 ;
  assign n30065 = x104 & n9928 ;
  assign n30066 = x103 & ~n9927 ;
  assign n30067 = n10379 & n30066 ;
  assign n30068 = n30065 | n30067 ;
  assign n30069 = n30064 | n30068 ;
  assign n30070 = n9936 | n30064 ;
  assign n30071 = n30068 | n30070 ;
  assign n30072 = ( n8273 & n30069 ) | ( n8273 & n30071 ) | ( n30069 & n30071 ) ;
  assign n30073 = x47 & n30071 ;
  assign n30074 = x47 & n30064 ;
  assign n30075 = ( x47 & n30068 ) | ( x47 & n30074 ) | ( n30068 & n30074 ) ;
  assign n30076 = ( n8273 & n30073 ) | ( n8273 & n30075 ) | ( n30073 & n30075 ) ;
  assign n30077 = x47 & ~n30075 ;
  assign n30078 = x47 & ~n30071 ;
  assign n30079 = ( ~n8273 & n30077 ) | ( ~n8273 & n30078 ) | ( n30077 & n30078 ) ;
  assign n30080 = ( n30072 & ~n30076 ) | ( n30072 & n30079 ) | ( ~n30076 & n30079 ) ;
  assign n30081 = x87 & n18290 ;
  assign n30082 = x63 & x86 ;
  assign n30083 = ~n18290 & n30082 ;
  assign n30084 = n30081 | n30083 ;
  assign n30085 = n29599 & ~n30084 ;
  assign n30086 = ~n29599 & n30084 ;
  assign n30087 = n30085 | n30086 ;
  assign n30089 = x89 & n17141 ;
  assign n30090 = x88 & ~n17140 ;
  assign n30091 = n17724 & n30090 ;
  assign n30092 = n30089 | n30091 ;
  assign n30088 = x90 & n17146 ;
  assign n30094 = n17149 | n30088 ;
  assign n30095 = n30092 | n30094 ;
  assign n30093 = n30088 | n30092 ;
  assign n30096 = n30093 & n30095 ;
  assign n30097 = ( n3519 & n30095 ) | ( n3519 & n30096 ) | ( n30095 & n30096 ) ;
  assign n30098 = x62 & n30096 ;
  assign n30099 = x62 & n30095 ;
  assign n30100 = ( n3519 & n30098 ) | ( n3519 & n30099 ) | ( n30098 & n30099 ) ;
  assign n30101 = x62 & ~n30096 ;
  assign n30102 = x62 & ~n30095 ;
  assign n30103 = ( ~n3519 & n30101 ) | ( ~n3519 & n30102 ) | ( n30101 & n30102 ) ;
  assign n30104 = ( n30097 & ~n30100 ) | ( n30097 & n30103 ) | ( ~n30100 & n30103 ) ;
  assign n30105 = ~n30087 & n30104 ;
  assign n30106 = n30087 & ~n30104 ;
  assign n30107 = n30105 | n30106 ;
  assign n30108 = ~n29603 & n29604 ;
  assign n30109 = ( n29603 & n29621 ) | ( n29603 & ~n30108 ) | ( n29621 & ~n30108 ) ;
  assign n30110 = ~n30107 & n30109 ;
  assign n30111 = n30107 & ~n30109 ;
  assign n30112 = n30110 | n30111 ;
  assign n30113 = x93 & n15552 ;
  assign n30114 = x92 & n15547 ;
  assign n30115 = x91 & ~n15546 ;
  assign n30116 = n16123 & n30115 ;
  assign n30117 = n30114 | n30116 ;
  assign n30118 = n30113 | n30117 ;
  assign n30119 = n15555 | n30113 ;
  assign n30120 = n30117 | n30119 ;
  assign n30121 = ( n4305 & n30118 ) | ( n4305 & n30120 ) | ( n30118 & n30120 ) ;
  assign n30122 = x59 & n30120 ;
  assign n30123 = x59 & n30113 ;
  assign n30124 = ( x59 & n30117 ) | ( x59 & n30123 ) | ( n30117 & n30123 ) ;
  assign n30125 = ( n4305 & n30122 ) | ( n4305 & n30124 ) | ( n30122 & n30124 ) ;
  assign n30126 = x59 & ~n30124 ;
  assign n30127 = x59 & ~n30120 ;
  assign n30128 = ( ~n4305 & n30126 ) | ( ~n4305 & n30127 ) | ( n30126 & n30127 ) ;
  assign n30129 = ( n30121 & ~n30125 ) | ( n30121 & n30128 ) | ( ~n30125 & n30128 ) ;
  assign n30130 = n30112 | n30129 ;
  assign n30131 = n30112 & ~n30129 ;
  assign n30132 = ( ~n30112 & n30130 ) | ( ~n30112 & n30131 ) | ( n30130 & n30131 ) ;
  assign n30133 = n29627 | n29646 ;
  assign n30134 = ( n29627 & ~n29629 ) | ( n29627 & n30133 ) | ( ~n29629 & n30133 ) ;
  assign n30135 = n30132 & ~n30134 ;
  assign n30136 = ~n30132 & n30134 ;
  assign n30137 = n30135 | n30136 ;
  assign n30138 = x96 & n14045 ;
  assign n30139 = x95 & n14040 ;
  assign n30140 = x94 & ~n14039 ;
  assign n30141 = n14552 & n30140 ;
  assign n30142 = n30139 | n30141 ;
  assign n30143 = n30138 | n30142 ;
  assign n30144 = n14048 | n30138 ;
  assign n30145 = n30142 | n30144 ;
  assign n30146 = ( n5202 & n30143 ) | ( n5202 & n30145 ) | ( n30143 & n30145 ) ;
  assign n30147 = x56 & n30145 ;
  assign n30148 = x56 & n30138 ;
  assign n30149 = ( x56 & n30142 ) | ( x56 & n30148 ) | ( n30142 & n30148 ) ;
  assign n30150 = ( n5202 & n30147 ) | ( n5202 & n30149 ) | ( n30147 & n30149 ) ;
  assign n30151 = x56 & ~n30149 ;
  assign n30152 = x56 & ~n30145 ;
  assign n30153 = ( ~n5202 & n30151 ) | ( ~n5202 & n30152 ) | ( n30151 & n30152 ) ;
  assign n30154 = ( n30146 & ~n30150 ) | ( n30146 & n30153 ) | ( ~n30150 & n30153 ) ;
  assign n30155 = n30137 & ~n30154 ;
  assign n30156 = ~n30137 & n30154 ;
  assign n30157 = n30155 | n30156 ;
  assign n30158 = n29652 | n29671 ;
  assign n30159 = ( n29652 & ~n29654 ) | ( n29652 & n30158 ) | ( ~n29654 & n30158 ) ;
  assign n30160 = ~n30157 & n30159 ;
  assign n30161 = n30157 & ~n30159 ;
  assign n30162 = n30160 | n30161 ;
  assign n30163 = x99 & n12574 ;
  assign n30164 = x98 & n12569 ;
  assign n30165 = x97 & ~n12568 ;
  assign n30166 = n13076 & n30165 ;
  assign n30167 = n30164 | n30166 ;
  assign n30168 = n30163 | n30167 ;
  assign n30169 = n12577 | n30163 ;
  assign n30170 = n30167 | n30169 ;
  assign n30171 = ( n6164 & n30168 ) | ( n6164 & n30170 ) | ( n30168 & n30170 ) ;
  assign n30172 = x53 & n30170 ;
  assign n30173 = x53 & n30163 ;
  assign n30174 = ( x53 & n30167 ) | ( x53 & n30173 ) | ( n30167 & n30173 ) ;
  assign n30175 = ( n6164 & n30172 ) | ( n6164 & n30174 ) | ( n30172 & n30174 ) ;
  assign n30176 = x53 & ~n30174 ;
  assign n30177 = x53 & ~n30170 ;
  assign n30178 = ( ~n6164 & n30176 ) | ( ~n6164 & n30177 ) | ( n30176 & n30177 ) ;
  assign n30179 = ( n30171 & ~n30175 ) | ( n30171 & n30178 ) | ( ~n30175 & n30178 ) ;
  assign n30180 = ~n30162 & n30179 ;
  assign n30181 = n30162 & ~n30179 ;
  assign n30182 = n30180 | n30181 ;
  assign n30183 = ( n29676 & ~n29677 ) | ( n29676 & n29704 ) | ( ~n29677 & n29704 ) ;
  assign n30184 = ~n30182 & n30183 ;
  assign n30185 = n30182 & ~n30183 ;
  assign n30186 = n30184 | n30185 ;
  assign n30187 = x102 & n11205 ;
  assign n30188 = x101 & n11200 ;
  assign n30189 = x100 & ~n11199 ;
  assign n30190 = n11679 & n30189 ;
  assign n30191 = n30188 | n30190 ;
  assign n30192 = n30187 | n30191 ;
  assign n30193 = n11208 | n30187 ;
  assign n30194 = n30191 | n30193 ;
  assign n30195 = ( n7178 & n30192 ) | ( n7178 & n30194 ) | ( n30192 & n30194 ) ;
  assign n30196 = x50 & n30194 ;
  assign n30197 = x50 & n30187 ;
  assign n30198 = ( x50 & n30191 ) | ( x50 & n30197 ) | ( n30191 & n30197 ) ;
  assign n30199 = ( n7178 & n30196 ) | ( n7178 & n30198 ) | ( n30196 & n30198 ) ;
  assign n30200 = x50 & ~n30198 ;
  assign n30201 = x50 & ~n30194 ;
  assign n30202 = ( ~n7178 & n30200 ) | ( ~n7178 & n30201 ) | ( n30200 & n30201 ) ;
  assign n30203 = ( n30195 & ~n30199 ) | ( n30195 & n30202 ) | ( ~n30199 & n30202 ) ;
  assign n30204 = n30186 | n30203 ;
  assign n30205 = n30186 & ~n30203 ;
  assign n30206 = ( ~n30186 & n30204 ) | ( ~n30186 & n30205 ) | ( n30204 & n30205 ) ;
  assign n30207 = n29706 | n29729 ;
  assign n30208 = ( n30080 & n30206 ) | ( n30080 & ~n30207 ) | ( n30206 & ~n30207 ) ;
  assign n30209 = ( ~n30206 & n30207 ) | ( ~n30206 & n30208 ) | ( n30207 & n30208 ) ;
  assign n30210 = ( ~n30080 & n30208 ) | ( ~n30080 & n30209 ) | ( n30208 & n30209 ) ;
  assign n30211 = n30063 & ~n30210 ;
  assign n30212 = ~n30063 & n30210 ;
  assign n30213 = n30211 | n30212 ;
  assign n30214 = x108 & n8724 ;
  assign n30215 = x107 & n8719 ;
  assign n30216 = x106 & ~n8718 ;
  assign n30217 = n9149 & n30216 ;
  assign n30218 = n30215 | n30217 ;
  assign n30219 = n30214 | n30218 ;
  assign n30220 = n8727 | n30214 ;
  assign n30221 = n30218 | n30220 ;
  assign n30222 = ( n9479 & n30219 ) | ( n9479 & n30221 ) | ( n30219 & n30221 ) ;
  assign n30223 = x44 & n30221 ;
  assign n30224 = x44 & n30214 ;
  assign n30225 = ( x44 & n30218 ) | ( x44 & n30224 ) | ( n30218 & n30224 ) ;
  assign n30226 = ( n9479 & n30223 ) | ( n9479 & n30225 ) | ( n30223 & n30225 ) ;
  assign n30227 = x44 & ~n30225 ;
  assign n30228 = x44 & ~n30221 ;
  assign n30229 = ( ~n9479 & n30227 ) | ( ~n9479 & n30228 ) | ( n30227 & n30228 ) ;
  assign n30230 = ( n30222 & ~n30226 ) | ( n30222 & n30229 ) | ( ~n30226 & n30229 ) ;
  assign n30231 = ~n30213 & n30230 ;
  assign n30232 = n30213 & ~n30230 ;
  assign n30233 = n30231 | n30232 ;
  assign n30234 = n29758 & ~n29779 ;
  assign n30235 = ( n29759 & n29779 ) | ( n29759 & ~n30234 ) | ( n29779 & ~n30234 ) ;
  assign n30236 = ( n29760 & ~n29762 ) | ( n29760 & n30235 ) | ( ~n29762 & n30235 ) ;
  assign n30237 = ~n30233 & n30236 ;
  assign n30238 = n30233 & ~n30236 ;
  assign n30239 = n30237 | n30238 ;
  assign n30240 = x111 & n7566 ;
  assign n30241 = x110 & n7561 ;
  assign n30242 = x109 & ~n7560 ;
  assign n30243 = n7953 & n30242 ;
  assign n30244 = n30241 | n30243 ;
  assign n30245 = n30240 | n30244 ;
  assign n30246 = n7569 | n30240 ;
  assign n30247 = n30244 | n30246 ;
  assign n30248 = ( n10749 & n30245 ) | ( n10749 & n30247 ) | ( n30245 & n30247 ) ;
  assign n30249 = x41 & n30247 ;
  assign n30250 = x41 & n30240 ;
  assign n30251 = ( x41 & n30244 ) | ( x41 & n30250 ) | ( n30244 & n30250 ) ;
  assign n30252 = ( n10749 & n30249 ) | ( n10749 & n30251 ) | ( n30249 & n30251 ) ;
  assign n30253 = x41 & ~n30251 ;
  assign n30254 = x41 & ~n30247 ;
  assign n30255 = ( ~n10749 & n30253 ) | ( ~n10749 & n30254 ) | ( n30253 & n30254 ) ;
  assign n30256 = ( n30248 & ~n30252 ) | ( n30248 & n30255 ) | ( ~n30252 & n30255 ) ;
  assign n30257 = n30239 | n30256 ;
  assign n30258 = n30239 & ~n30256 ;
  assign n30259 = ( ~n30239 & n30257 ) | ( ~n30239 & n30258 ) | ( n30257 & n30258 ) ;
  assign n30260 = ( n29785 & ~n29786 ) | ( n29785 & n29805 ) | ( ~n29786 & n29805 ) ;
  assign n30261 = n30259 & ~n30260 ;
  assign n30262 = ~n30259 & n30260 ;
  assign n30263 = n30261 | n30262 ;
  assign n30264 = x114 & n6536 ;
  assign n30265 = x113 & n6531 ;
  assign n30266 = x112 & ~n6530 ;
  assign n30267 = n6871 & n30266 ;
  assign n30268 = n30265 | n30267 ;
  assign n30269 = n30264 | n30268 ;
  assign n30270 = n6539 | n30264 ;
  assign n30271 = n30268 | n30270 ;
  assign n30272 = ( ~n12095 & n30269 ) | ( ~n12095 & n30271 ) | ( n30269 & n30271 ) ;
  assign n30273 = n30269 & n30271 ;
  assign n30274 = ( n12079 & n30272 ) | ( n12079 & n30273 ) | ( n30272 & n30273 ) ;
  assign n30275 = x38 & n30274 ;
  assign n30276 = x38 & ~n30274 ;
  assign n30277 = ( n30274 & ~n30275 ) | ( n30274 & n30276 ) | ( ~n30275 & n30276 ) ;
  assign n30278 = n30263 & ~n30277 ;
  assign n30279 = ~n30263 & n30277 ;
  assign n30280 = n30278 | n30279 ;
  assign n30282 = ~n30280 & n30281 ;
  assign n30283 = n30281 & ~n30282 ;
  assign n30284 = n30280 | n30282 ;
  assign n30285 = ~n30283 & n30284 ;
  assign n30286 = x117 & n5554 ;
  assign n30287 = x116 & n5549 ;
  assign n30288 = x115 & ~n5548 ;
  assign n30289 = n5893 & n30288 ;
  assign n30290 = n30287 | n30289 ;
  assign n30291 = n30286 | n30290 ;
  assign n30292 = n5557 | n30286 ;
  assign n30293 = n30290 | n30292 ;
  assign n30294 = ( ~n13522 & n30291 ) | ( ~n13522 & n30293 ) | ( n30291 & n30293 ) ;
  assign n30295 = n30291 & n30293 ;
  assign n30296 = ( n13503 & n30294 ) | ( n13503 & n30295 ) | ( n30294 & n30295 ) ;
  assign n30297 = x35 & n30296 ;
  assign n30298 = x35 & ~n30296 ;
  assign n30299 = ( n30296 & ~n30297 ) | ( n30296 & n30298 ) | ( ~n30297 & n30298 ) ;
  assign n30300 = n30285 & n30299 ;
  assign n30301 = n30285 | n30299 ;
  assign n30302 = ~n30300 & n30301 ;
  assign n30303 = n30062 & ~n30302 ;
  assign n30304 = ~n30058 & n30302 ;
  assign n30305 = ~n30061 & n30304 ;
  assign n30306 = n30303 | n30305 ;
  assign n30307 = n30031 & n30035 ;
  assign n30308 = ( n29853 & n30031 ) | ( n29853 & n30307 ) | ( n30031 & n30307 ) ;
  assign n30309 = ( n29897 & n30307 ) | ( n29897 & n30308 ) | ( n30307 & n30308 ) ;
  assign n30310 = n30306 | n30309 ;
  assign n30311 = n30031 & ~n30306 ;
  assign n30312 = ( n30038 & ~n30310 ) | ( n30038 & n30311 ) | ( ~n30310 & n30311 ) ;
  assign n30313 = n30306 & n30309 ;
  assign n30314 = ~n30031 & n30306 ;
  assign n30315 = ( ~n30038 & n30313 ) | ( ~n30038 & n30314 ) | ( n30313 & n30314 ) ;
  assign n30316 = n30312 | n30315 ;
  assign n30317 = ~n30014 & n30316 ;
  assign n30318 = n30014 & ~n30316 ;
  assign n30319 = n30317 | n30318 ;
  assign n30320 = x127 & ~n2423 ;
  assign n30321 = n2631 & n30320 ;
  assign n30322 = n2432 & n19877 ;
  assign n30323 = n30321 | n30322 ;
  assign n30324 = n2432 & n19880 ;
  assign n30325 = n30321 | n30324 ;
  assign n30326 = ( n18202 & n30323 ) | ( n18202 & n30325 ) | ( n30323 & n30325 ) ;
  assign n30327 = n30323 & n30325 ;
  assign n30328 = ( n18212 & n30326 ) | ( n18212 & n30327 ) | ( n30326 & n30327 ) ;
  assign n30329 = ( n18214 & n30326 ) | ( n18214 & n30327 ) | ( n30326 & n30327 ) ;
  assign n30330 = ( n14002 & n30328 ) | ( n14002 & n30329 ) | ( n30328 & n30329 ) ;
  assign n30331 = x23 & n30328 ;
  assign n30332 = x23 & n30329 ;
  assign n30333 = ( n14002 & n30331 ) | ( n14002 & n30332 ) | ( n30331 & n30332 ) ;
  assign n30334 = x23 & ~n30332 ;
  assign n30335 = x23 & ~n30331 ;
  assign n30336 = ( ~n14002 & n30334 ) | ( ~n14002 & n30335 ) | ( n30334 & n30335 ) ;
  assign n30337 = ( n30330 & ~n30333 ) | ( n30330 & n30336 ) | ( ~n30333 & n30336 ) ;
  assign n30338 = n29942 | n29978 ;
  assign n30339 = ( n30319 & n30337 ) | ( n30319 & ~n30338 ) | ( n30337 & ~n30338 ) ;
  assign n30340 = ( n30319 & ~n30337 ) | ( n30319 & n30338 ) | ( ~n30337 & n30338 ) ;
  assign n30341 = ( ~n30319 & n30339 ) | ( ~n30319 & n30340 ) | ( n30339 & n30340 ) ;
  assign n30342 = n29984 & n30341 ;
  assign n30343 = n29917 & n30341 ;
  assign n30344 = ( n29919 & n30342 ) | ( n29919 & n30343 ) | ( n30342 & n30343 ) ;
  assign n30345 = n29985 & ~n30344 ;
  assign n30346 = ~n29984 & n30341 ;
  assign n30347 = ~n29917 & n30341 ;
  assign n30348 = ( ~n29919 & n30346 ) | ( ~n29919 & n30347 ) | ( n30346 & n30347 ) ;
  assign n30349 = n30345 | n30348 ;
  assign n30350 = n29956 & n30349 ;
  assign n30351 = ( n29967 & n30349 ) | ( n29967 & n30350 ) | ( n30349 & n30350 ) ;
  assign n30352 = ( n29966 & n30349 ) | ( n29966 & n30350 ) | ( n30349 & n30350 ) ;
  assign n30353 = ( n29579 & n30351 ) | ( n29579 & n30352 ) | ( n30351 & n30352 ) ;
  assign n30354 = n29956 | n29969 ;
  assign n30355 = n30349 & n30354 ;
  assign n30356 = n29956 | n29970 ;
  assign n30357 = n30349 & n30356 ;
  assign n30358 = ( n29172 & n30355 ) | ( n29172 & n30357 ) | ( n30355 & n30357 ) ;
  assign n30359 = n29956 | n29966 ;
  assign n30360 = n30349 & n30359 ;
  assign n30361 = ( n29581 & n30357 ) | ( n29581 & n30360 ) | ( n30357 & n30360 ) ;
  assign n30362 = ( n28312 & n30358 ) | ( n28312 & n30361 ) | ( n30358 & n30361 ) ;
  assign n30363 = ( n26030 & n30353 ) | ( n26030 & n30362 ) | ( n30353 & n30362 ) ;
  assign n30364 = n29956 | n29967 ;
  assign n30365 = ( n29579 & n30359 ) | ( n29579 & n30364 ) | ( n30359 & n30364 ) ;
  assign n30366 = ( n29172 & n30354 ) | ( n29172 & n30356 ) | ( n30354 & n30356 ) ;
  assign n30367 = ( n29581 & n30356 ) | ( n29581 & n30359 ) | ( n30356 & n30359 ) ;
  assign n30368 = ( n28312 & n30366 ) | ( n28312 & n30367 ) | ( n30366 & n30367 ) ;
  assign n30369 = ( n26030 & n30365 ) | ( n26030 & n30368 ) | ( n30365 & n30368 ) ;
  assign n30370 = ~n30363 & n30369 ;
  assign n30371 = ( n30349 & ~n30363 ) | ( n30349 & n30370 ) | ( ~n30363 & n30370 ) ;
  assign n30372 = x88 & n18290 ;
  assign n30373 = x63 & x87 ;
  assign n30374 = ~n18290 & n30373 ;
  assign n30375 = n30372 | n30374 ;
  assign n30376 = ~x23 & n30375 ;
  assign n30377 = x23 & ~n30375 ;
  assign n30378 = n30376 | n30377 ;
  assign n30379 = n30084 & ~n30378 ;
  assign n30380 = ~n30084 & n30378 ;
  assign n30381 = n30379 | n30380 ;
  assign n30382 = x90 & n17141 ;
  assign n30383 = x89 & ~n17140 ;
  assign n30384 = n17724 & n30383 ;
  assign n30385 = n30382 | n30384 ;
  assign n30386 = x91 & n17146 ;
  assign n30387 = n17149 | n30386 ;
  assign n30388 = n30385 | n30387 ;
  assign n30389 = ~x62 & n30388 ;
  assign n30390 = ~x62 & n30386 ;
  assign n30391 = ( ~x62 & n30385 ) | ( ~x62 & n30390 ) | ( n30385 & n30390 ) ;
  assign n30392 = ( n3768 & n30389 ) | ( n3768 & n30391 ) | ( n30389 & n30391 ) ;
  assign n30393 = x62 & ~n30388 ;
  assign n30394 = x62 & x91 ;
  assign n30395 = n17146 & n30394 ;
  assign n30396 = x62 & ~n30395 ;
  assign n30397 = ~n30385 & n30396 ;
  assign n30398 = ( ~n3768 & n30393 ) | ( ~n3768 & n30397 ) | ( n30393 & n30397 ) ;
  assign n30399 = n30392 | n30398 ;
  assign n30400 = ~n30381 & n30399 ;
  assign n30401 = n30381 & ~n30399 ;
  assign n30402 = n30400 | n30401 ;
  assign n30403 = ~n30085 & n30087 ;
  assign n30404 = ( n30085 & n30104 ) | ( n30085 & ~n30403 ) | ( n30104 & ~n30403 ) ;
  assign n30405 = n30402 & n30404 ;
  assign n30406 = n30402 | n30404 ;
  assign n30407 = ~n30405 & n30406 ;
  assign n30408 = x94 & n15552 ;
  assign n30409 = x93 & n15547 ;
  assign n30410 = x92 & ~n15546 ;
  assign n30411 = n16123 & n30410 ;
  assign n30412 = n30409 | n30411 ;
  assign n30413 = n30408 | n30412 ;
  assign n30414 = n15555 | n30408 ;
  assign n30415 = n30412 | n30414 ;
  assign n30416 = ( n4583 & n30413 ) | ( n4583 & n30415 ) | ( n30413 & n30415 ) ;
  assign n30417 = x59 & n30415 ;
  assign n30418 = x59 & n30408 ;
  assign n30419 = ( x59 & n30412 ) | ( x59 & n30418 ) | ( n30412 & n30418 ) ;
  assign n30420 = ( n4583 & n30417 ) | ( n4583 & n30419 ) | ( n30417 & n30419 ) ;
  assign n30421 = x59 & ~n30419 ;
  assign n30422 = x59 & ~n30415 ;
  assign n30423 = ( ~n4583 & n30421 ) | ( ~n4583 & n30422 ) | ( n30421 & n30422 ) ;
  assign n30424 = ( n30416 & ~n30420 ) | ( n30416 & n30423 ) | ( ~n30420 & n30423 ) ;
  assign n30425 = ~n30407 & n30424 ;
  assign n30426 = n30407 & ~n30424 ;
  assign n30427 = n30425 | n30426 ;
  assign n30428 = n30109 | n30129 ;
  assign n30429 = ( ~n30107 & n30129 ) | ( ~n30107 & n30428 ) | ( n30129 & n30428 ) ;
  assign n30430 = ( n30110 & ~n30112 ) | ( n30110 & n30429 ) | ( ~n30112 & n30429 ) ;
  assign n30431 = n30427 & ~n30430 ;
  assign n30432 = ~n30427 & n30430 ;
  assign n30433 = n30431 | n30432 ;
  assign n30434 = x97 & n14045 ;
  assign n30435 = x96 & n14040 ;
  assign n30436 = x95 & ~n14039 ;
  assign n30437 = n14552 & n30436 ;
  assign n30438 = n30435 | n30437 ;
  assign n30439 = n30434 | n30438 ;
  assign n30440 = n14048 | n30434 ;
  assign n30441 = n30438 | n30440 ;
  assign n30442 = ( n5505 & n30439 ) | ( n5505 & n30441 ) | ( n30439 & n30441 ) ;
  assign n30443 = x56 & n30441 ;
  assign n30444 = x56 & n30434 ;
  assign n30445 = ( x56 & n30438 ) | ( x56 & n30444 ) | ( n30438 & n30444 ) ;
  assign n30446 = ( n5505 & n30443 ) | ( n5505 & n30445 ) | ( n30443 & n30445 ) ;
  assign n30447 = x56 & ~n30445 ;
  assign n30448 = x56 & ~n30441 ;
  assign n30449 = ( ~n5505 & n30447 ) | ( ~n5505 & n30448 ) | ( n30447 & n30448 ) ;
  assign n30450 = ( n30442 & ~n30446 ) | ( n30442 & n30449 ) | ( ~n30446 & n30449 ) ;
  assign n30451 = n30134 | n30154 ;
  assign n30452 = ( ~n30132 & n30154 ) | ( ~n30132 & n30451 ) | ( n30154 & n30451 ) ;
  assign n30453 = n30450 & n30452 ;
  assign n30454 = n30136 & n30450 ;
  assign n30455 = ( ~n30137 & n30453 ) | ( ~n30137 & n30454 ) | ( n30453 & n30454 ) ;
  assign n30456 = n30450 | n30452 ;
  assign n30457 = n30136 | n30450 ;
  assign n30458 = ( ~n30137 & n30456 ) | ( ~n30137 & n30457 ) | ( n30456 & n30457 ) ;
  assign n30459 = ~n30455 & n30458 ;
  assign n30460 = ~n30433 & n30459 ;
  assign n30461 = n30433 & ~n30459 ;
  assign n30462 = n30460 | n30461 ;
  assign n30463 = x100 & n12574 ;
  assign n30464 = x99 & n12569 ;
  assign n30465 = x98 & ~n12568 ;
  assign n30466 = n13076 & n30465 ;
  assign n30467 = n30464 | n30466 ;
  assign n30468 = n30463 | n30467 ;
  assign n30469 = n12577 | n30463 ;
  assign n30470 = n30467 | n30469 ;
  assign n30471 = ( n6483 & n30468 ) | ( n6483 & n30470 ) | ( n30468 & n30470 ) ;
  assign n30472 = x53 & n30470 ;
  assign n30473 = x53 & n30463 ;
  assign n30474 = ( x53 & n30467 ) | ( x53 & n30473 ) | ( n30467 & n30473 ) ;
  assign n30475 = ( n6483 & n30472 ) | ( n6483 & n30474 ) | ( n30472 & n30474 ) ;
  assign n30476 = x53 & ~n30474 ;
  assign n30477 = x53 & ~n30470 ;
  assign n30478 = ( ~n6483 & n30476 ) | ( ~n6483 & n30477 ) | ( n30476 & n30477 ) ;
  assign n30479 = ( n30471 & ~n30475 ) | ( n30471 & n30478 ) | ( ~n30475 & n30478 ) ;
  assign n30480 = ~n30462 & n30479 ;
  assign n30481 = n30462 | n30480 ;
  assign n30483 = n30159 | n30179 ;
  assign n30484 = ( ~n30157 & n30179 ) | ( ~n30157 & n30483 ) | ( n30179 & n30483 ) ;
  assign n30485 = ( n30160 & ~n30162 ) | ( n30160 & n30484 ) | ( ~n30162 & n30484 ) ;
  assign n30482 = n30462 & n30479 ;
  assign n30486 = n30482 & n30485 ;
  assign n30487 = ( ~n30481 & n30485 ) | ( ~n30481 & n30486 ) | ( n30485 & n30486 ) ;
  assign n30488 = n30482 | n30485 ;
  assign n30489 = n30481 & ~n30488 ;
  assign n30490 = n30487 | n30489 ;
  assign n30491 = x103 & n11205 ;
  assign n30492 = x102 & n11200 ;
  assign n30493 = x101 & ~n11199 ;
  assign n30494 = n11679 & n30493 ;
  assign n30495 = n30492 | n30494 ;
  assign n30496 = n30491 | n30495 ;
  assign n30497 = n11208 | n30491 ;
  assign n30498 = n30495 | n30497 ;
  assign n30499 = ( n7529 & n30496 ) | ( n7529 & n30498 ) | ( n30496 & n30498 ) ;
  assign n30500 = x50 & n30498 ;
  assign n30501 = x50 & n30491 ;
  assign n30502 = ( x50 & n30495 ) | ( x50 & n30501 ) | ( n30495 & n30501 ) ;
  assign n30503 = ( n7529 & n30500 ) | ( n7529 & n30502 ) | ( n30500 & n30502 ) ;
  assign n30504 = x50 & ~n30502 ;
  assign n30505 = x50 & ~n30498 ;
  assign n30506 = ( ~n7529 & n30504 ) | ( ~n7529 & n30505 ) | ( n30504 & n30505 ) ;
  assign n30507 = ( n30499 & ~n30503 ) | ( n30499 & n30506 ) | ( ~n30503 & n30506 ) ;
  assign n30508 = ~n30490 & n30507 ;
  assign n30509 = n30490 | n30508 ;
  assign n30511 = n30184 | n30203 ;
  assign n30512 = ( n30184 & ~n30186 ) | ( n30184 & n30511 ) | ( ~n30186 & n30511 ) ;
  assign n30510 = n30490 & n30507 ;
  assign n30513 = n30510 & n30512 ;
  assign n30514 = ( ~n30509 & n30512 ) | ( ~n30509 & n30513 ) | ( n30512 & n30513 ) ;
  assign n30515 = n30510 | n30512 ;
  assign n30516 = n30509 & ~n30515 ;
  assign n30517 = n30514 | n30516 ;
  assign n30518 = x106 & n9933 ;
  assign n30519 = x105 & n9928 ;
  assign n30520 = x104 & ~n9927 ;
  assign n30521 = n10379 & n30520 ;
  assign n30522 = n30519 | n30521 ;
  assign n30523 = n30518 | n30522 ;
  assign n30524 = n9936 | n30518 ;
  assign n30525 = n30522 | n30524 ;
  assign n30526 = ( n8656 & n30523 ) | ( n8656 & n30525 ) | ( n30523 & n30525 ) ;
  assign n30527 = x47 & n30525 ;
  assign n30528 = x47 & n30518 ;
  assign n30529 = ( x47 & n30522 ) | ( x47 & n30528 ) | ( n30522 & n30528 ) ;
  assign n30530 = ( n8656 & n30527 ) | ( n8656 & n30529 ) | ( n30527 & n30529 ) ;
  assign n30531 = x47 & ~n30529 ;
  assign n30532 = x47 & ~n30525 ;
  assign n30533 = ( ~n8656 & n30531 ) | ( ~n8656 & n30532 ) | ( n30531 & n30532 ) ;
  assign n30534 = ( n30526 & ~n30530 ) | ( n30526 & n30533 ) | ( ~n30530 & n30533 ) ;
  assign n30535 = ~n30517 & n30534 ;
  assign n30536 = n30517 | n30535 ;
  assign n30537 = n30517 & n30534 ;
  assign n30538 = ~n30206 & n30207 ;
  assign n30539 = n30206 | n30207 ;
  assign n30540 = n30080 & ~n30206 ;
  assign n30541 = ( n30080 & ~n30207 ) | ( n30080 & n30540 ) | ( ~n30207 & n30540 ) ;
  assign n30542 = n30539 & n30541 ;
  assign n30543 = ( n30080 & n30538 ) | ( n30080 & ~n30542 ) | ( n30538 & ~n30542 ) ;
  assign n30544 = ~n30537 & n30543 ;
  assign n30545 = n30536 & n30544 ;
  assign n30546 = n30537 & ~n30543 ;
  assign n30547 = ( n30536 & n30543 ) | ( n30536 & ~n30546 ) | ( n30543 & ~n30546 ) ;
  assign n30548 = ~n30545 & n30547 ;
  assign n30549 = x109 & n8724 ;
  assign n30550 = x108 & n8719 ;
  assign n30551 = x107 & ~n8718 ;
  assign n30552 = n9149 & n30551 ;
  assign n30553 = n30550 | n30552 ;
  assign n30554 = n30549 | n30553 ;
  assign n30555 = n8727 | n30549 ;
  assign n30556 = n30553 | n30555 ;
  assign n30557 = ( n9878 & n30554 ) | ( n9878 & n30556 ) | ( n30554 & n30556 ) ;
  assign n30558 = x44 & n30556 ;
  assign n30559 = x44 & n30549 ;
  assign n30560 = ( x44 & n30553 ) | ( x44 & n30559 ) | ( n30553 & n30559 ) ;
  assign n30561 = ( n9878 & n30558 ) | ( n9878 & n30560 ) | ( n30558 & n30560 ) ;
  assign n30562 = x44 & ~n30560 ;
  assign n30563 = x44 & ~n30556 ;
  assign n30564 = ( ~n9878 & n30562 ) | ( ~n9878 & n30563 ) | ( n30562 & n30563 ) ;
  assign n30565 = ( n30557 & ~n30561 ) | ( n30557 & n30564 ) | ( ~n30561 & n30564 ) ;
  assign n30566 = ~n30548 & n30565 ;
  assign n30567 = n30548 & ~n30565 ;
  assign n30568 = n30566 | n30567 ;
  assign n30569 = n30210 & ~n30230 ;
  assign n30570 = ( n30063 & n30230 ) | ( n30063 & ~n30569 ) | ( n30230 & ~n30569 ) ;
  assign n30571 = ( n30211 & ~n30213 ) | ( n30211 & n30570 ) | ( ~n30213 & n30570 ) ;
  assign n30572 = n30568 & ~n30571 ;
  assign n30573 = ~n30568 & n30571 ;
  assign n30574 = n30572 | n30573 ;
  assign n30575 = x112 & n7566 ;
  assign n30576 = x111 & n7561 ;
  assign n30577 = x110 & ~n7560 ;
  assign n30578 = n7953 & n30577 ;
  assign n30579 = n30576 | n30578 ;
  assign n30580 = n30575 | n30579 ;
  assign n30581 = n7569 | n30575 ;
  assign n30582 = n30579 | n30581 ;
  assign n30583 = ( n11172 & n30580 ) | ( n11172 & n30582 ) | ( n30580 & n30582 ) ;
  assign n30584 = x41 & n30582 ;
  assign n30585 = x41 & n30575 ;
  assign n30586 = ( x41 & n30579 ) | ( x41 & n30585 ) | ( n30579 & n30585 ) ;
  assign n30587 = ( n11172 & n30584 ) | ( n11172 & n30586 ) | ( n30584 & n30586 ) ;
  assign n30588 = x41 & ~n30586 ;
  assign n30589 = x41 & ~n30582 ;
  assign n30590 = ( ~n11172 & n30588 ) | ( ~n11172 & n30589 ) | ( n30588 & n30589 ) ;
  assign n30591 = ( n30583 & ~n30587 ) | ( n30583 & n30590 ) | ( ~n30587 & n30590 ) ;
  assign n30592 = ~n30574 & n30591 ;
  assign n30593 = n30574 | n30592 ;
  assign n30595 = n30237 | n30256 ;
  assign n30596 = ( n30237 & ~n30239 ) | ( n30237 & n30595 ) | ( ~n30239 & n30595 ) ;
  assign n30594 = n30574 & n30591 ;
  assign n30597 = n30594 & n30596 ;
  assign n30598 = ( ~n30593 & n30596 ) | ( ~n30593 & n30597 ) | ( n30596 & n30597 ) ;
  assign n30599 = n30594 | n30596 ;
  assign n30600 = n30593 & ~n30599 ;
  assign n30601 = n30598 | n30600 ;
  assign n30602 = x115 & n6536 ;
  assign n30603 = x114 & n6531 ;
  assign n30604 = x113 & ~n6530 ;
  assign n30605 = n6871 & n30604 ;
  assign n30606 = n30603 | n30605 ;
  assign n30607 = n30602 | n30606 ;
  assign n30608 = n6539 | n30602 ;
  assign n30609 = n30606 | n30608 ;
  assign n30610 = ( ~n12550 & n30607 ) | ( ~n12550 & n30609 ) | ( n30607 & n30609 ) ;
  assign n30611 = n30607 & n30609 ;
  assign n30612 = ( n12532 & n30610 ) | ( n12532 & n30611 ) | ( n30610 & n30611 ) ;
  assign n30613 = x38 & n30612 ;
  assign n30614 = x38 & ~n30612 ;
  assign n30615 = ( n30612 & ~n30613 ) | ( n30612 & n30614 ) | ( ~n30613 & n30614 ) ;
  assign n30616 = ~n30601 & n30615 ;
  assign n30617 = n30601 & ~n30615 ;
  assign n30618 = n30616 | n30617 ;
  assign n30619 = n30262 | n30277 ;
  assign n30620 = ( n30262 & ~n30263 ) | ( n30262 & n30619 ) | ( ~n30263 & n30619 ) ;
  assign n30621 = ~n30618 & n30620 ;
  assign n30622 = n30618 | n30621 ;
  assign n30623 = x118 & n5554 ;
  assign n30624 = x117 & n5549 ;
  assign n30625 = x116 & ~n5548 ;
  assign n30626 = n5893 & n30625 ;
  assign n30627 = n30624 | n30626 ;
  assign n30628 = n30623 | n30627 ;
  assign n30629 = n5557 | n30623 ;
  assign n30630 = n30627 | n30629 ;
  assign n30631 = ( ~n14002 & n30628 ) | ( ~n14002 & n30630 ) | ( n30628 & n30630 ) ;
  assign n30632 = n30628 & n30630 ;
  assign n30633 = ( n13981 & n30631 ) | ( n13981 & n30632 ) | ( n30631 & n30632 ) ;
  assign n30634 = x35 & n30633 ;
  assign n30635 = x35 & ~n30633 ;
  assign n30636 = ( n30633 & ~n30634 ) | ( n30633 & n30635 ) | ( ~n30634 & n30635 ) ;
  assign n30637 = n30620 | n30636 ;
  assign n30638 = ( n30618 & n30636 ) | ( n30618 & n30637 ) | ( n30636 & n30637 ) ;
  assign n30639 = n30622 & ~n30638 ;
  assign n30640 = n30620 & n30636 ;
  assign n30641 = n30618 & n30640 ;
  assign n30642 = ( ~n30622 & n30636 ) | ( ~n30622 & n30641 ) | ( n30636 & n30641 ) ;
  assign n30643 = n30639 | n30642 ;
  assign n30644 = n30282 | n30299 ;
  assign n30645 = ( n30282 & ~n30285 ) | ( n30282 & n30644 ) | ( ~n30285 & n30644 ) ;
  assign n30646 = ~n30643 & n30645 ;
  assign n30647 = n30643 & ~n30645 ;
  assign n30648 = n30646 | n30647 ;
  assign n30649 = x121 & n4631 ;
  assign n30650 = x120 & n4626 ;
  assign n30651 = x119 & ~n4625 ;
  assign n30652 = n4943 & n30651 ;
  assign n30653 = n30650 | n30652 ;
  assign n30654 = n30649 | n30653 ;
  assign n30655 = n4634 | n30649 ;
  assign n30656 = n30653 | n30655 ;
  assign n30657 = ( n15501 & n30654 ) | ( n15501 & n30656 ) | ( n30654 & n30656 ) ;
  assign n30658 = x32 & n30656 ;
  assign n30659 = x32 & n30649 ;
  assign n30660 = ( x32 & n30653 ) | ( x32 & n30659 ) | ( n30653 & n30659 ) ;
  assign n30661 = ( n15501 & n30658 ) | ( n15501 & n30660 ) | ( n30658 & n30660 ) ;
  assign n30662 = x32 & ~n30660 ;
  assign n30663 = x32 & ~n30656 ;
  assign n30664 = ( ~n15501 & n30662 ) | ( ~n15501 & n30663 ) | ( n30662 & n30663 ) ;
  assign n30665 = ( n30657 & ~n30661 ) | ( n30657 & n30664 ) | ( ~n30661 & n30664 ) ;
  assign n30666 = ( ~n30058 & n30062 ) | ( ~n30058 & n30304 ) | ( n30062 & n30304 ) ;
  assign n30667 = ~n30665 & n30666 ;
  assign n30668 = n30665 & ~n30666 ;
  assign n30669 = n30667 | n30668 ;
  assign n30670 = ( n30031 & n30038 ) | ( n30031 & ~n30309 ) | ( n30038 & ~n30309 ) ;
  assign n30671 = ( n30309 & n30310 ) | ( n30309 & n30670 ) | ( n30310 & n30670 ) ;
  assign n30672 = x124 & n3816 ;
  assign n30673 = x123 & n3811 ;
  assign n30674 = x122 & ~n3810 ;
  assign n30675 = n4067 & n30674 ;
  assign n30676 = n30673 | n30675 ;
  assign n30677 = n30672 | n30676 ;
  assign n30678 = n3819 | n30672 ;
  assign n30679 = n30676 | n30678 ;
  assign n30680 = ( n17084 & n30677 ) | ( n17084 & n30679 ) | ( n30677 & n30679 ) ;
  assign n30681 = x29 & n30679 ;
  assign n30682 = x29 & n30672 ;
  assign n30683 = ( x29 & n30676 ) | ( x29 & n30682 ) | ( n30676 & n30682 ) ;
  assign n30684 = ( n17084 & n30681 ) | ( n17084 & n30683 ) | ( n30681 & n30683 ) ;
  assign n30685 = x29 & ~n30683 ;
  assign n30686 = x29 & ~n30679 ;
  assign n30687 = ( ~n17084 & n30685 ) | ( ~n17084 & n30686 ) | ( n30685 & n30686 ) ;
  assign n30688 = ( n30680 & ~n30684 ) | ( n30680 & n30687 ) | ( ~n30684 & n30687 ) ;
  assign n30689 = n30310 & n30688 ;
  assign n30690 = n30309 & n30688 ;
  assign n30691 = ( n30670 & n30689 ) | ( n30670 & n30690 ) | ( n30689 & n30690 ) ;
  assign n30692 = ~n30310 & n30688 ;
  assign n30693 = ~n30309 & n30688 ;
  assign n30694 = ( ~n30670 & n30692 ) | ( ~n30670 & n30693 ) | ( n30692 & n30693 ) ;
  assign n30695 = ( n30671 & ~n30691 ) | ( n30671 & n30694 ) | ( ~n30691 & n30694 ) ;
  assign n30696 = ( n30648 & ~n30669 ) | ( n30648 & n30695 ) | ( ~n30669 & n30695 ) ;
  assign n30697 = ( n30669 & ~n30695 ) | ( n30669 & n30696 ) | ( ~n30695 & n30696 ) ;
  assign n30698 = ( ~n30648 & n30696 ) | ( ~n30648 & n30697 ) | ( n30696 & n30697 ) ;
  assign n30699 = x127 & n3085 ;
  assign n30700 = x126 & n3080 ;
  assign n30701 = x125 & ~n3079 ;
  assign n30702 = n3309 & n30701 ;
  assign n30703 = n30700 | n30702 ;
  assign n30704 = n30699 | n30703 ;
  assign n30705 = n3088 | n30699 ;
  assign n30706 = n30703 | n30705 ;
  assign n30707 = ( n18763 & n30704 ) | ( n18763 & n30706 ) | ( n30704 & n30706 ) ;
  assign n30708 = x26 & n30706 ;
  assign n30709 = x26 & n30699 ;
  assign n30710 = ( x26 & n30703 ) | ( x26 & n30709 ) | ( n30703 & n30709 ) ;
  assign n30711 = ( n18763 & n30708 ) | ( n18763 & n30710 ) | ( n30708 & n30710 ) ;
  assign n30712 = x26 & ~n30710 ;
  assign n30713 = x26 & ~n30706 ;
  assign n30714 = ( ~n18763 & n30712 ) | ( ~n18763 & n30713 ) | ( n30712 & n30713 ) ;
  assign n30715 = ( n30707 & ~n30711 ) | ( n30707 & n30714 ) | ( ~n30711 & n30714 ) ;
  assign n30716 = n30010 | n30316 ;
  assign n30717 = ( n30010 & n30014 ) | ( n30010 & n30716 ) | ( n30014 & n30716 ) ;
  assign n30718 = ( n30698 & n30715 ) | ( n30698 & ~n30717 ) | ( n30715 & ~n30717 ) ;
  assign n30719 = ( ~n30715 & n30717 ) | ( ~n30715 & n30718 ) | ( n30717 & n30718 ) ;
  assign n30720 = ( ~n30698 & n30718 ) | ( ~n30698 & n30719 ) | ( n30718 & n30719 ) ;
  assign n30721 = ~n29942 & n30337 ;
  assign n30722 = ~n29978 & n30721 ;
  assign n30723 = n30319 & ~n30722 ;
  assign n30724 = n29942 & n30337 ;
  assign n30725 = ( n29978 & n30337 ) | ( n29978 & n30724 ) | ( n30337 & n30724 ) ;
  assign n30726 = n30338 & ~n30725 ;
  assign n30727 = ( n30319 & n30725 ) | ( n30319 & n30726 ) | ( n30725 & n30726 ) ;
  assign n30728 = n30319 | n30725 ;
  assign n30729 = ( ~n30723 & n30727 ) | ( ~n30723 & n30728 ) | ( n30727 & n30728 ) ;
  assign n30730 = n30720 & ~n30729 ;
  assign n30731 = n30344 | n30358 ;
  assign n30732 = n30344 | n30361 ;
  assign n30733 = ( n28312 & n30731 ) | ( n28312 & n30732 ) | ( n30731 & n30732 ) ;
  assign n30734 = n30344 | n30350 ;
  assign n30735 = n30344 | n30349 ;
  assign n30736 = ( n29967 & n30734 ) | ( n29967 & n30735 ) | ( n30734 & n30735 ) ;
  assign n30737 = ( n29966 & n30734 ) | ( n29966 & n30735 ) | ( n30734 & n30735 ) ;
  assign n30738 = ( n29576 & n30736 ) | ( n29576 & n30737 ) | ( n30736 & n30737 ) ;
  assign n30739 = ( n29578 & n30736 ) | ( n29578 & n30737 ) | ( n30736 & n30737 ) ;
  assign n30740 = ( n27383 & n30738 ) | ( n27383 & n30739 ) | ( n30738 & n30739 ) ;
  assign n30741 = ( n25496 & n30733 ) | ( n25496 & n30740 ) | ( n30733 & n30740 ) ;
  assign n30742 = n30733 | n30740 ;
  assign n30743 = ( n25522 & n30741 ) | ( n25522 & n30742 ) | ( n30741 & n30742 ) ;
  assign n30744 = ( n25519 & n30741 ) | ( n25519 & n30742 ) | ( n30741 & n30742 ) ;
  assign n30745 = ( n22794 & n30743 ) | ( n22794 & n30744 ) | ( n30743 & n30744 ) ;
  assign n30746 = ( ~n30720 & n30729 ) | ( ~n30720 & n30745 ) | ( n30729 & n30745 ) ;
  assign n30747 = n30720 & n30729 ;
  assign n30748 = n30729 & ~n30747 ;
  assign n30749 = n30730 | n30748 ;
  assign n30750 = n30742 & n30749 ;
  assign n30751 = n30741 & n30749 ;
  assign n30752 = ( n25522 & n30750 ) | ( n25522 & n30751 ) | ( n30750 & n30751 ) ;
  assign n30753 = ( n25519 & n30750 ) | ( n25519 & n30751 ) | ( n30750 & n30751 ) ;
  assign n30754 = ( n22794 & n30752 ) | ( n22794 & n30753 ) | ( n30752 & n30753 ) ;
  assign n30755 = ( n30730 & n30746 ) | ( n30730 & ~n30754 ) | ( n30746 & ~n30754 ) ;
  assign n31101 = n30715 & n30717 ;
  assign n31102 = n30717 & ~n31101 ;
  assign n31103 = n30696 & n30715 ;
  assign n31104 = ~n30648 & n30715 ;
  assign n31105 = ( n30697 & n31103 ) | ( n30697 & n31104 ) | ( n31103 & n31104 ) ;
  assign n31106 = ~n30717 & n31105 ;
  assign n31107 = n31101 | n31106 ;
  assign n31108 = n30698 | n31101 ;
  assign n31109 = ( n31102 & n31107 ) | ( n31102 & n31108 ) | ( n31107 & n31108 ) ;
  assign n30770 = n30648 | n30669 ;
  assign n30771 = n30648 & n30669 ;
  assign n30772 = n30770 & ~n30771 ;
  assign n30773 = n30691 | n30772 ;
  assign n30774 = ( n30691 & n30695 ) | ( n30691 & n30773 ) | ( n30695 & n30773 ) ;
  assign n30756 = x127 & n3080 ;
  assign n30757 = x126 & ~n3079 ;
  assign n30758 = n3309 & n30757 ;
  assign n30759 = n30756 | n30758 ;
  assign n30760 = n3088 | n30759 ;
  assign n30761 = ( n19328 & n30759 ) | ( n19328 & n30760 ) | ( n30759 & n30760 ) ;
  assign n30762 = x26 & n30759 ;
  assign n30763 = ( x26 & n4990 ) | ( x26 & n30759 ) | ( n4990 & n30759 ) ;
  assign n30764 = ( n19328 & n30762 ) | ( n19328 & n30763 ) | ( n30762 & n30763 ) ;
  assign n30765 = x26 & ~n4990 ;
  assign n30766 = ~n30759 & n30765 ;
  assign n30767 = x26 & ~n30759 ;
  assign n30768 = ( ~n19328 & n30766 ) | ( ~n19328 & n30767 ) | ( n30766 & n30767 ) ;
  assign n30769 = ( n30761 & ~n30764 ) | ( n30761 & n30768 ) | ( ~n30764 & n30768 ) ;
  assign n30775 = n30769 & n30774 ;
  assign n30776 = n30774 & ~n30775 ;
  assign n30777 = n30769 & ~n30774 ;
  assign n30778 = n30648 & ~n30665 ;
  assign n30779 = ( n30648 & n30666 ) | ( n30648 & n30778 ) | ( n30666 & n30778 ) ;
  assign n30780 = ( ~n30668 & n30669 ) | ( ~n30668 & n30779 ) | ( n30669 & n30779 ) ;
  assign n30781 = x125 & n3816 ;
  assign n30782 = x124 & n3811 ;
  assign n30783 = x123 & ~n3810 ;
  assign n30784 = n4067 & n30783 ;
  assign n30785 = n30782 | n30784 ;
  assign n30786 = n30781 | n30785 ;
  assign n30787 = n3819 | n30781 ;
  assign n30788 = n30785 | n30787 ;
  assign n30789 = ( n17670 & n30786 ) | ( n17670 & n30788 ) | ( n30786 & n30788 ) ;
  assign n30790 = x29 & n30788 ;
  assign n30791 = x29 & n30781 ;
  assign n30792 = ( x29 & n30785 ) | ( x29 & n30791 ) | ( n30785 & n30791 ) ;
  assign n30793 = ( n17670 & n30790 ) | ( n17670 & n30792 ) | ( n30790 & n30792 ) ;
  assign n30794 = x29 & ~n30792 ;
  assign n30795 = x29 & ~n30788 ;
  assign n30796 = ( ~n17670 & n30794 ) | ( ~n17670 & n30795 ) | ( n30794 & n30795 ) ;
  assign n30797 = ( n30789 & ~n30793 ) | ( n30789 & n30796 ) | ( ~n30793 & n30796 ) ;
  assign n30798 = ~n30779 & n30797 ;
  assign n30799 = n30668 & n30797 ;
  assign n30800 = ( ~n30669 & n30798 ) | ( ~n30669 & n30799 ) | ( n30798 & n30799 ) ;
  assign n30801 = n30780 | n30800 ;
  assign n30803 = x121 & n4626 ;
  assign n30804 = x120 & ~n4625 ;
  assign n30805 = n4943 & n30804 ;
  assign n30806 = n30803 | n30805 ;
  assign n30802 = x122 & n4631 ;
  assign n30808 = n4634 | n30802 ;
  assign n30809 = n30806 | n30808 ;
  assign n30807 = n30802 | n30806 ;
  assign n30810 = n30807 & n30809 ;
  assign n30811 = ( n16043 & n30809 ) | ( n16043 & n30810 ) | ( n30809 & n30810 ) ;
  assign n30812 = x32 & n30810 ;
  assign n30813 = x32 & n30809 ;
  assign n30814 = ( n16043 & n30812 ) | ( n16043 & n30813 ) | ( n30812 & n30813 ) ;
  assign n30815 = x32 & ~n30810 ;
  assign n30816 = x32 & ~n30809 ;
  assign n30817 = ( ~n16043 & n30815 ) | ( ~n16043 & n30816 ) | ( n30815 & n30816 ) ;
  assign n30818 = ( n30811 & ~n30814 ) | ( n30811 & n30817 ) | ( ~n30814 & n30817 ) ;
  assign n30819 = n30641 & n30818 ;
  assign n30820 = n30636 & n30818 ;
  assign n30821 = ( ~n30622 & n30819 ) | ( ~n30622 & n30820 ) | ( n30819 & n30820 ) ;
  assign n30822 = ( n30646 & n30818 ) | ( n30646 & n30821 ) | ( n30818 & n30821 ) ;
  assign n30823 = n30641 | n30818 ;
  assign n30824 = n30636 | n30818 ;
  assign n30825 = ( ~n30622 & n30823 ) | ( ~n30622 & n30824 ) | ( n30823 & n30824 ) ;
  assign n30826 = n30646 | n30825 ;
  assign n30827 = ~n30822 & n30826 ;
  assign n31060 = n30616 | n30620 ;
  assign n31061 = ( n30616 & ~n30618 ) | ( n30616 & n31060 ) | ( ~n30618 & n31060 ) ;
  assign n30828 = n30592 | n30598 ;
  assign n31014 = n30566 | n30571 ;
  assign n31015 = ( n30566 & ~n30568 ) | ( n30566 & n31014 ) | ( ~n30568 & n31014 ) ;
  assign n30829 = n30508 | n30514 ;
  assign n30830 = n30480 | n30487 ;
  assign n30831 = x89 & n18290 ;
  assign n30832 = x63 & x88 ;
  assign n30833 = ~n18290 & n30832 ;
  assign n30834 = n30831 | n30833 ;
  assign n30835 = n30084 | n30376 ;
  assign n30836 = ( n30376 & ~n30378 ) | ( n30376 & n30835 ) | ( ~n30378 & n30835 ) ;
  assign n30837 = n30834 & ~n30836 ;
  assign n30838 = ~n30834 & n30836 ;
  assign n30839 = n30837 | n30838 ;
  assign n30841 = x91 & n17141 ;
  assign n30842 = x90 & ~n17140 ;
  assign n30843 = n17724 & n30842 ;
  assign n30844 = n30841 | n30843 ;
  assign n30840 = x92 & n17146 ;
  assign n30846 = n17149 | n30840 ;
  assign n30847 = n30844 | n30846 ;
  assign n30845 = n30840 | n30844 ;
  assign n30848 = n30845 & n30847 ;
  assign n30849 = ( n4040 & n30847 ) | ( n4040 & n30848 ) | ( n30847 & n30848 ) ;
  assign n30850 = x62 & n30848 ;
  assign n30851 = x62 & n30847 ;
  assign n30852 = ( n4040 & n30850 ) | ( n4040 & n30851 ) | ( n30850 & n30851 ) ;
  assign n30853 = x62 & ~n30848 ;
  assign n30854 = x62 & ~n30847 ;
  assign n30855 = ( ~n4040 & n30853 ) | ( ~n4040 & n30854 ) | ( n30853 & n30854 ) ;
  assign n30856 = ( n30849 & ~n30852 ) | ( n30849 & n30855 ) | ( ~n30852 & n30855 ) ;
  assign n30857 = ~n30839 & n30856 ;
  assign n30858 = n30839 & ~n30856 ;
  assign n30859 = n30857 | n30858 ;
  assign n30860 = n30400 | n30404 ;
  assign n30861 = ( n30400 & ~n30402 ) | ( n30400 & n30860 ) | ( ~n30402 & n30860 ) ;
  assign n30862 = ~n30859 & n30861 ;
  assign n30863 = n30859 & ~n30861 ;
  assign n30864 = n30862 | n30863 ;
  assign n30865 = x95 & n15552 ;
  assign n30866 = x94 & n15547 ;
  assign n30867 = x93 & ~n15546 ;
  assign n30868 = n16123 & n30867 ;
  assign n30869 = n30866 | n30868 ;
  assign n30870 = n30865 | n30869 ;
  assign n30871 = n15555 | n30865 ;
  assign n30872 = n30869 | n30871 ;
  assign n30873 = ( n4897 & n30870 ) | ( n4897 & n30872 ) | ( n30870 & n30872 ) ;
  assign n30874 = x59 & n30872 ;
  assign n30875 = x59 & n30865 ;
  assign n30876 = ( x59 & n30869 ) | ( x59 & n30875 ) | ( n30869 & n30875 ) ;
  assign n30877 = ( n4897 & n30874 ) | ( n4897 & n30876 ) | ( n30874 & n30876 ) ;
  assign n30878 = x59 & ~n30876 ;
  assign n30879 = x59 & ~n30872 ;
  assign n30880 = ( ~n4897 & n30878 ) | ( ~n4897 & n30879 ) | ( n30878 & n30879 ) ;
  assign n30881 = ( n30873 & ~n30877 ) | ( n30873 & n30880 ) | ( ~n30877 & n30880 ) ;
  assign n30882 = n30864 | n30881 ;
  assign n30883 = n30864 & ~n30881 ;
  assign n30884 = ( ~n30864 & n30882 ) | ( ~n30864 & n30883 ) | ( n30882 & n30883 ) ;
  assign n30885 = n30425 | n30430 ;
  assign n30886 = ( n30425 & ~n30427 ) | ( n30425 & n30885 ) | ( ~n30427 & n30885 ) ;
  assign n30887 = n30884 & ~n30886 ;
  assign n30888 = ~n30884 & n30886 ;
  assign n30889 = n30887 | n30888 ;
  assign n30890 = x98 & n14045 ;
  assign n30891 = x97 & n14040 ;
  assign n30892 = x96 & ~n14039 ;
  assign n30893 = n14552 & n30892 ;
  assign n30894 = n30891 | n30893 ;
  assign n30895 = n30890 | n30894 ;
  assign n30896 = n14048 | n30890 ;
  assign n30897 = n30894 | n30896 ;
  assign n30898 = ( ~n5850 & n30895 ) | ( ~n5850 & n30897 ) | ( n30895 & n30897 ) ;
  assign n30899 = n30895 & n30897 ;
  assign n30900 = ( n5834 & n30898 ) | ( n5834 & n30899 ) | ( n30898 & n30899 ) ;
  assign n30901 = x56 & n30897 ;
  assign n30902 = x56 & n30890 ;
  assign n30903 = ( x56 & n30894 ) | ( x56 & n30902 ) | ( n30894 & n30902 ) ;
  assign n30904 = ( ~n5850 & n30901 ) | ( ~n5850 & n30903 ) | ( n30901 & n30903 ) ;
  assign n30905 = n30901 & n30903 ;
  assign n30906 = ( n5834 & n30904 ) | ( n5834 & n30905 ) | ( n30904 & n30905 ) ;
  assign n30907 = x56 & ~n30903 ;
  assign n30908 = x56 & ~n30897 ;
  assign n30909 = ( n5850 & n30907 ) | ( n5850 & n30908 ) | ( n30907 & n30908 ) ;
  assign n30910 = n30907 | n30908 ;
  assign n30911 = ( ~n5834 & n30909 ) | ( ~n5834 & n30910 ) | ( n30909 & n30910 ) ;
  assign n30912 = ( n30900 & ~n30906 ) | ( n30900 & n30911 ) | ( ~n30906 & n30911 ) ;
  assign n30913 = n30889 & n30912 ;
  assign n30914 = n30888 | n30912 ;
  assign n30915 = n30887 | n30914 ;
  assign n30916 = ~n30913 & n30915 ;
  assign n30917 = n30433 & ~n30455 ;
  assign n30918 = ( n30455 & n30459 ) | ( n30455 & ~n30917 ) | ( n30459 & ~n30917 ) ;
  assign n30919 = n30916 & ~n30918 ;
  assign n30920 = ~n30916 & n30918 ;
  assign n30921 = n30919 | n30920 ;
  assign n30922 = x101 & n12574 ;
  assign n30923 = x100 & n12569 ;
  assign n30924 = x99 & ~n12568 ;
  assign n30925 = n13076 & n30924 ;
  assign n30926 = n30923 | n30925 ;
  assign n30927 = n30922 | n30926 ;
  assign n30928 = n12577 | n30922 ;
  assign n30929 = n30926 | n30928 ;
  assign n30930 = ( n6844 & n30927 ) | ( n6844 & n30929 ) | ( n30927 & n30929 ) ;
  assign n30931 = x53 & n30929 ;
  assign n30932 = x53 & n30922 ;
  assign n30933 = ( x53 & n30926 ) | ( x53 & n30932 ) | ( n30926 & n30932 ) ;
  assign n30934 = ( n6844 & n30931 ) | ( n6844 & n30933 ) | ( n30931 & n30933 ) ;
  assign n30935 = x53 & ~n30933 ;
  assign n30936 = x53 & ~n30929 ;
  assign n30937 = ( ~n6844 & n30935 ) | ( ~n6844 & n30936 ) | ( n30935 & n30936 ) ;
  assign n30938 = ( n30930 & ~n30934 ) | ( n30930 & n30937 ) | ( ~n30934 & n30937 ) ;
  assign n30939 = n30921 & ~n30938 ;
  assign n30940 = ~n30921 & n30938 ;
  assign n30941 = n30939 | n30940 ;
  assign n30942 = n30830 & ~n30941 ;
  assign n30943 = n30830 & ~n30942 ;
  assign n30944 = x104 & n11205 ;
  assign n30945 = x103 & n11200 ;
  assign n30946 = x102 & ~n11199 ;
  assign n30947 = n11679 & n30946 ;
  assign n30948 = n30945 | n30947 ;
  assign n30949 = n30944 | n30948 ;
  assign n30950 = n11208 | n30944 ;
  assign n30951 = n30948 | n30950 ;
  assign n30952 = ( n7911 & n30949 ) | ( n7911 & n30951 ) | ( n30949 & n30951 ) ;
  assign n30953 = x50 & n30951 ;
  assign n30954 = x50 & n30944 ;
  assign n30955 = ( x50 & n30948 ) | ( x50 & n30954 ) | ( n30948 & n30954 ) ;
  assign n30956 = ( n7911 & n30953 ) | ( n7911 & n30955 ) | ( n30953 & n30955 ) ;
  assign n30957 = x50 & ~n30955 ;
  assign n30958 = x50 & ~n30951 ;
  assign n30959 = ( ~n7911 & n30957 ) | ( ~n7911 & n30958 ) | ( n30957 & n30958 ) ;
  assign n30960 = ( n30952 & ~n30956 ) | ( n30952 & n30959 ) | ( ~n30956 & n30959 ) ;
  assign n30961 = n30941 & ~n30960 ;
  assign n30962 = ( n30830 & ~n30960 ) | ( n30830 & n30961 ) | ( ~n30960 & n30961 ) ;
  assign n30963 = ~n30943 & n30962 ;
  assign n30964 = ( n30830 & ~n30941 ) | ( n30830 & n30960 ) | ( ~n30941 & n30960 ) ;
  assign n30965 = ~n30942 & n30964 ;
  assign n30966 = n30963 | n30965 ;
  assign n30967 = n30829 & ~n30966 ;
  assign n30968 = ~n30829 & n30966 ;
  assign n30969 = n30967 | n30968 ;
  assign n30970 = x107 & n9933 ;
  assign n30971 = x106 & n9928 ;
  assign n30972 = x105 & ~n9927 ;
  assign n30973 = n10379 & n30972 ;
  assign n30974 = n30971 | n30973 ;
  assign n30975 = n30970 | n30974 ;
  assign n30976 = n9936 | n30970 ;
  assign n30977 = n30974 | n30976 ;
  assign n30978 = ( n9084 & n30975 ) | ( n9084 & n30977 ) | ( n30975 & n30977 ) ;
  assign n30979 = x47 & n30977 ;
  assign n30980 = x47 & n30970 ;
  assign n30981 = ( x47 & n30974 ) | ( x47 & n30980 ) | ( n30974 & n30980 ) ;
  assign n30982 = ( n9084 & n30979 ) | ( n9084 & n30981 ) | ( n30979 & n30981 ) ;
  assign n30983 = x47 & ~n30981 ;
  assign n30984 = x47 & ~n30977 ;
  assign n30985 = ( ~n9084 & n30983 ) | ( ~n9084 & n30984 ) | ( n30983 & n30984 ) ;
  assign n30986 = ( n30978 & ~n30982 ) | ( n30978 & n30985 ) | ( ~n30982 & n30985 ) ;
  assign n30987 = n30969 | n30986 ;
  assign n30988 = n30969 & ~n30986 ;
  assign n30989 = ( ~n30969 & n30987 ) | ( ~n30969 & n30988 ) | ( n30987 & n30988 ) ;
  assign n30990 = ( ~n30517 & n30534 ) | ( ~n30517 & n30538 ) | ( n30534 & n30538 ) ;
  assign n30991 = ( n30080 & ~n30517 ) | ( n30080 & n30534 ) | ( ~n30517 & n30534 ) ;
  assign n30992 = ( ~n30542 & n30990 ) | ( ~n30542 & n30991 ) | ( n30990 & n30991 ) ;
  assign n30993 = n30989 & ~n30992 ;
  assign n30994 = ~n30989 & n30992 ;
  assign n30995 = n30993 | n30994 ;
  assign n30996 = x110 & n8724 ;
  assign n30997 = x109 & n8719 ;
  assign n30998 = x108 & ~n8718 ;
  assign n30999 = n9149 & n30998 ;
  assign n31000 = n30997 | n30999 ;
  assign n31001 = n30996 | n31000 ;
  assign n31002 = n8727 | n30996 ;
  assign n31003 = n31000 | n31002 ;
  assign n31004 = ( n10330 & n31001 ) | ( n10330 & n31003 ) | ( n31001 & n31003 ) ;
  assign n31005 = x44 & n31003 ;
  assign n31006 = x44 & n30996 ;
  assign n31007 = ( x44 & n31000 ) | ( x44 & n31006 ) | ( n31000 & n31006 ) ;
  assign n31008 = ( n10330 & n31005 ) | ( n10330 & n31007 ) | ( n31005 & n31007 ) ;
  assign n31009 = x44 & ~n31007 ;
  assign n31010 = x44 & ~n31003 ;
  assign n31011 = ( ~n10330 & n31009 ) | ( ~n10330 & n31010 ) | ( n31009 & n31010 ) ;
  assign n31012 = ( n31004 & ~n31008 ) | ( n31004 & n31011 ) | ( ~n31008 & n31011 ) ;
  assign n31013 = n30995 & n31012 ;
  assign n31016 = n31013 & n31015 ;
  assign n31017 = n30992 | n31012 ;
  assign n31018 = ( ~n30989 & n31012 ) | ( ~n30989 & n31017 ) | ( n31012 & n31017 ) ;
  assign n31019 = n30993 | n31018 ;
  assign n31020 = ( n31015 & n31016 ) | ( n31015 & ~n31019 ) | ( n31016 & ~n31019 ) ;
  assign n31021 = ~n31013 & n31019 ;
  assign n31022 = ~n31015 & n31021 ;
  assign n31023 = n31020 | n31022 ;
  assign n31024 = x113 & n7566 ;
  assign n31025 = x112 & n7561 ;
  assign n31026 = x111 & ~n7560 ;
  assign n31027 = n7953 & n31026 ;
  assign n31028 = n31025 | n31027 ;
  assign n31029 = n31024 | n31028 ;
  assign n31030 = n7569 | n31024 ;
  assign n31031 = n31028 | n31030 ;
  assign n31032 = ( ~n11642 & n31029 ) | ( ~n11642 & n31031 ) | ( n31029 & n31031 ) ;
  assign n31033 = n31029 & n31031 ;
  assign n31034 = ( n11626 & n31032 ) | ( n11626 & n31033 ) | ( n31032 & n31033 ) ;
  assign n31035 = x41 & n31034 ;
  assign n31036 = x41 & ~n31034 ;
  assign n31037 = ( n31034 & ~n31035 ) | ( n31034 & n31036 ) | ( ~n31035 & n31036 ) ;
  assign n31038 = n31022 | n31037 ;
  assign n31039 = n31020 | n31038 ;
  assign n31040 = n31022 & ~n31037 ;
  assign n31041 = ( n31020 & ~n31037 ) | ( n31020 & n31040 ) | ( ~n31037 & n31040 ) ;
  assign n31042 = ( ~n31023 & n31039 ) | ( ~n31023 & n31041 ) | ( n31039 & n31041 ) ;
  assign n31043 = ~n30828 & n31042 ;
  assign n31044 = n30828 & ~n31042 ;
  assign n31045 = n31043 | n31044 ;
  assign n31046 = x116 & n6536 ;
  assign n31047 = x115 & n6531 ;
  assign n31048 = x114 & ~n6530 ;
  assign n31049 = n6871 & n31048 ;
  assign n31050 = n31047 | n31049 ;
  assign n31051 = n31046 | n31050 ;
  assign n31052 = n6539 | n31046 ;
  assign n31053 = n31050 | n31052 ;
  assign n31054 = ( ~n13040 & n31051 ) | ( ~n13040 & n31053 ) | ( n31051 & n31053 ) ;
  assign n31055 = n31051 & n31053 ;
  assign n31056 = ( n13022 & n31054 ) | ( n13022 & n31055 ) | ( n31054 & n31055 ) ;
  assign n31057 = x38 & n31056 ;
  assign n31058 = x38 & ~n31056 ;
  assign n31059 = ( n31056 & ~n31057 ) | ( n31056 & n31058 ) | ( ~n31057 & n31058 ) ;
  assign n31062 = ( n31045 & ~n31059 ) | ( n31045 & n31061 ) | ( ~n31059 & n31061 ) ;
  assign n31063 = ( ~n31045 & n31059 ) | ( ~n31045 & n31061 ) | ( n31059 & n31061 ) ;
  assign n31064 = ( ~n31061 & n31062 ) | ( ~n31061 & n31063 ) | ( n31062 & n31063 ) ;
  assign n31065 = x119 & n5554 ;
  assign n31066 = x118 & n5549 ;
  assign n31067 = x117 & ~n5548 ;
  assign n31068 = n5893 & n31067 ;
  assign n31069 = n31066 | n31068 ;
  assign n31070 = n31065 | n31069 ;
  assign n31071 = n5557 | n31065 ;
  assign n31072 = n31069 | n31071 ;
  assign n31073 = ( n14496 & n31070 ) | ( n14496 & n31072 ) | ( n31070 & n31072 ) ;
  assign n31074 = x35 & n31072 ;
  assign n31075 = x35 & n31065 ;
  assign n31076 = ( x35 & n31069 ) | ( x35 & n31075 ) | ( n31069 & n31075 ) ;
  assign n31077 = ( n14496 & n31074 ) | ( n14496 & n31076 ) | ( n31074 & n31076 ) ;
  assign n31078 = x35 & ~n31076 ;
  assign n31079 = x35 & ~n31072 ;
  assign n31080 = ( ~n14496 & n31078 ) | ( ~n14496 & n31079 ) | ( n31078 & n31079 ) ;
  assign n31081 = ( n31073 & ~n31077 ) | ( n31073 & n31080 ) | ( ~n31077 & n31080 ) ;
  assign n31082 = ~n31064 & n31081 ;
  assign n31083 = n31064 & ~n31081 ;
  assign n31084 = n31082 | n31083 ;
  assign n31085 = n30827 & ~n31084 ;
  assign n31086 = ~n30827 & n31084 ;
  assign n31087 = n31085 | n31086 ;
  assign n31088 = n30779 & n30797 ;
  assign n31089 = ~n30668 & n30797 ;
  assign n31090 = ( n30669 & n31088 ) | ( n30669 & n31089 ) | ( n31088 & n31089 ) ;
  assign n31091 = ~n31087 & n31090 ;
  assign n31092 = ( n30801 & n31087 ) | ( n30801 & ~n31091 ) | ( n31087 & ~n31091 ) ;
  assign n31093 = n31087 & ~n31090 ;
  assign n31094 = n30801 & n31093 ;
  assign n31095 = n31092 & ~n31094 ;
  assign n31096 = n30777 | n31095 ;
  assign n31097 = n30776 | n31096 ;
  assign n31098 = n30777 & n31095 ;
  assign n31099 = ( n30776 & n31095 ) | ( n30776 & n31098 ) | ( n31095 & n31098 ) ;
  assign n31100 = n31097 & ~n31099 ;
  assign n31110 = n31100 & n31109 ;
  assign n31111 = n31109 & ~n31110 ;
  assign n31112 = n30747 | n30754 ;
  assign n31113 = n31100 & ~n31109 ;
  assign n31114 = n31112 | n31113 ;
  assign n31115 = n31111 | n31114 ;
  assign n31116 = n31111 | n31113 ;
  assign n31117 = n30747 & n31113 ;
  assign n31118 = ( n30747 & n31111 ) | ( n30747 & n31117 ) | ( n31111 & n31117 ) ;
  assign n31119 = ( n30754 & n31116 ) | ( n30754 & n31118 ) | ( n31116 & n31118 ) ;
  assign n31120 = n31115 & ~n31119 ;
  assign n31121 = n30775 | n31099 ;
  assign n31122 = ~n30800 & n31092 ;
  assign n31123 = x127 & ~n3079 ;
  assign n31124 = n3309 & n31123 ;
  assign n31125 = n3088 & n19877 ;
  assign n31126 = n31124 | n31125 ;
  assign n31127 = n3088 & n19880 ;
  assign n31128 = n31124 | n31127 ;
  assign n31129 = ( n18202 & n31126 ) | ( n18202 & n31128 ) | ( n31126 & n31128 ) ;
  assign n31130 = n31126 & n31128 ;
  assign n31131 = ( n18212 & n31129 ) | ( n18212 & n31130 ) | ( n31129 & n31130 ) ;
  assign n31132 = ( n18214 & n31129 ) | ( n18214 & n31130 ) | ( n31129 & n31130 ) ;
  assign n31133 = ( n14002 & n31131 ) | ( n14002 & n31132 ) | ( n31131 & n31132 ) ;
  assign n31134 = x26 & n31131 ;
  assign n31135 = x26 & n31132 ;
  assign n31136 = ( n14002 & n31134 ) | ( n14002 & n31135 ) | ( n31134 & n31135 ) ;
  assign n31137 = x26 & ~n31135 ;
  assign n31138 = x26 & ~n31134 ;
  assign n31139 = ( ~n14002 & n31137 ) | ( ~n14002 & n31138 ) | ( n31137 & n31138 ) ;
  assign n31140 = ( n31133 & ~n31136 ) | ( n31133 & n31139 ) | ( ~n31136 & n31139 ) ;
  assign n31141 = n30797 & n31140 ;
  assign n31142 = ~n30779 & n31141 ;
  assign n31143 = n30668 & n31141 ;
  assign n31144 = ( ~n30669 & n31142 ) | ( ~n30669 & n31143 ) | ( n31142 & n31143 ) ;
  assign n31145 = ( ~n31092 & n31140 ) | ( ~n31092 & n31144 ) | ( n31140 & n31144 ) ;
  assign n31146 = n31122 | n31145 ;
  assign n31147 = x126 & n3816 ;
  assign n31148 = x125 & n3811 ;
  assign n31149 = x124 & ~n3810 ;
  assign n31150 = n4067 & n31149 ;
  assign n31151 = n31148 | n31150 ;
  assign n31152 = n31147 | n31151 ;
  assign n31153 = n3819 | n31147 ;
  assign n31154 = n31151 | n31153 ;
  assign n31155 = ( n18220 & n31152 ) | ( n18220 & n31154 ) | ( n31152 & n31154 ) ;
  assign n31156 = x29 & n31154 ;
  assign n31157 = x29 & n31147 ;
  assign n31158 = ( x29 & n31151 ) | ( x29 & n31157 ) | ( n31151 & n31157 ) ;
  assign n31159 = ( n18220 & n31156 ) | ( n18220 & n31158 ) | ( n31156 & n31158 ) ;
  assign n31160 = x29 & ~n31158 ;
  assign n31161 = x29 & ~n31154 ;
  assign n31162 = ( ~n18220 & n31160 ) | ( ~n18220 & n31161 ) | ( n31160 & n31161 ) ;
  assign n31163 = ( n31155 & ~n31159 ) | ( n31155 & n31162 ) | ( ~n31159 & n31162 ) ;
  assign n31164 = ~n30822 & n31084 ;
  assign n31165 = ( n30822 & n30827 ) | ( n30822 & ~n31164 ) | ( n30827 & ~n31164 ) ;
  assign n31166 = n31163 | n31165 ;
  assign n31167 = n31163 & n31165 ;
  assign n31168 = n31166 & ~n31167 ;
  assign n31169 = x123 & n4631 ;
  assign n31170 = x122 & n4626 ;
  assign n31171 = x121 & ~n4625 ;
  assign n31172 = n4943 & n31171 ;
  assign n31173 = n31170 | n31172 ;
  assign n31174 = n31169 | n31173 ;
  assign n31175 = n4634 | n31169 ;
  assign n31176 = n31173 | n31175 ;
  assign n31177 = ( n16086 & n31174 ) | ( n16086 & n31176 ) | ( n31174 & n31176 ) ;
  assign n31178 = x32 & n31176 ;
  assign n31179 = x32 & n31169 ;
  assign n31180 = ( x32 & n31173 ) | ( x32 & n31179 ) | ( n31173 & n31179 ) ;
  assign n31181 = ( n16086 & n31178 ) | ( n16086 & n31180 ) | ( n31178 & n31180 ) ;
  assign n31182 = x32 & ~n31180 ;
  assign n31183 = x32 & ~n31176 ;
  assign n31184 = ( ~n16086 & n31182 ) | ( ~n16086 & n31183 ) | ( n31182 & n31183 ) ;
  assign n31185 = ( n31177 & ~n31181 ) | ( n31177 & n31184 ) | ( ~n31181 & n31184 ) ;
  assign n31186 = ~n31045 & n31059 ;
  assign n31187 = n31045 | n31186 ;
  assign n31188 = n31045 & n31059 ;
  assign n31189 = n31061 & n31188 ;
  assign n31190 = ( n31061 & ~n31187 ) | ( n31061 & n31189 ) | ( ~n31187 & n31189 ) ;
  assign n31191 = n31185 & n31190 ;
  assign n31192 = ( n31082 & n31185 ) | ( n31082 & n31191 ) | ( n31185 & n31191 ) ;
  assign n31193 = n31185 | n31190 ;
  assign n31194 = n31082 | n31193 ;
  assign n31195 = ~n31192 & n31194 ;
  assign n31196 = n30942 | n30965 ;
  assign n31299 = n30920 | n30938 ;
  assign n31300 = ( n30920 & ~n30921 ) | ( n30920 & n31299 ) | ( ~n30921 & n31299 ) ;
  assign n31197 = x90 & n18290 ;
  assign n31198 = x63 & x89 ;
  assign n31199 = ~n18290 & n31198 ;
  assign n31200 = n31197 | n31199 ;
  assign n31201 = n30834 & ~n31200 ;
  assign n31202 = ~n30834 & n31200 ;
  assign n31203 = n31201 | n31202 ;
  assign n31205 = x92 & n17141 ;
  assign n31206 = x91 & ~n17140 ;
  assign n31207 = n17724 & n31206 ;
  assign n31208 = n31205 | n31207 ;
  assign n31204 = x93 & n17146 ;
  assign n31210 = n17149 | n31204 ;
  assign n31211 = n31208 | n31210 ;
  assign n31209 = n31204 | n31208 ;
  assign n31212 = n31209 & n31211 ;
  assign n31213 = ( n4305 & n31211 ) | ( n4305 & n31212 ) | ( n31211 & n31212 ) ;
  assign n31214 = x62 & n31212 ;
  assign n31215 = x62 & n31211 ;
  assign n31216 = ( n4305 & n31214 ) | ( n4305 & n31215 ) | ( n31214 & n31215 ) ;
  assign n31217 = x62 & ~n31212 ;
  assign n31218 = x62 & ~n31211 ;
  assign n31219 = ( ~n4305 & n31217 ) | ( ~n4305 & n31218 ) | ( n31217 & n31218 ) ;
  assign n31220 = ( n31213 & ~n31216 ) | ( n31213 & n31219 ) | ( ~n31216 & n31219 ) ;
  assign n31221 = ~n31203 & n31220 ;
  assign n31222 = n31203 & ~n31220 ;
  assign n31223 = n31221 | n31222 ;
  assign n31224 = ~n30838 & n30839 ;
  assign n31225 = ( n30838 & n30856 ) | ( n30838 & ~n31224 ) | ( n30856 & ~n31224 ) ;
  assign n31226 = ~n31223 & n31225 ;
  assign n31227 = n31223 & ~n31225 ;
  assign n31228 = n31226 | n31227 ;
  assign n31229 = x96 & n15552 ;
  assign n31230 = x95 & n15547 ;
  assign n31231 = x94 & ~n15546 ;
  assign n31232 = n16123 & n31231 ;
  assign n31233 = n31230 | n31232 ;
  assign n31234 = n31229 | n31233 ;
  assign n31235 = n15555 | n31229 ;
  assign n31236 = n31233 | n31235 ;
  assign n31237 = ( n5202 & n31234 ) | ( n5202 & n31236 ) | ( n31234 & n31236 ) ;
  assign n31238 = x59 & n31236 ;
  assign n31239 = x59 & n31229 ;
  assign n31240 = ( x59 & n31233 ) | ( x59 & n31239 ) | ( n31233 & n31239 ) ;
  assign n31241 = ( n5202 & n31238 ) | ( n5202 & n31240 ) | ( n31238 & n31240 ) ;
  assign n31242 = x59 & ~n31240 ;
  assign n31243 = x59 & ~n31236 ;
  assign n31244 = ( ~n5202 & n31242 ) | ( ~n5202 & n31243 ) | ( n31242 & n31243 ) ;
  assign n31245 = ( n31237 & ~n31241 ) | ( n31237 & n31244 ) | ( ~n31241 & n31244 ) ;
  assign n31246 = ~n31228 & n31245 ;
  assign n31247 = n31228 & ~n31245 ;
  assign n31248 = n31246 | n31247 ;
  assign n31249 = n30859 & ~n30881 ;
  assign n31250 = ( n30861 & n30881 ) | ( n30861 & ~n31249 ) | ( n30881 & ~n31249 ) ;
  assign n31251 = ( n30862 & ~n30864 ) | ( n30862 & n31250 ) | ( ~n30864 & n31250 ) ;
  assign n31252 = ~n31248 & n31251 ;
  assign n31253 = n31248 & ~n31251 ;
  assign n31254 = n31252 | n31253 ;
  assign n31255 = x99 & n14045 ;
  assign n31256 = x98 & n14040 ;
  assign n31257 = x97 & ~n14039 ;
  assign n31258 = n14552 & n31257 ;
  assign n31259 = n31256 | n31258 ;
  assign n31260 = n31255 | n31259 ;
  assign n31261 = n14048 | n31255 ;
  assign n31262 = n31259 | n31261 ;
  assign n31263 = ( n6164 & n31260 ) | ( n6164 & n31262 ) | ( n31260 & n31262 ) ;
  assign n31264 = x56 & n31262 ;
  assign n31265 = x56 & n31255 ;
  assign n31266 = ( x56 & n31259 ) | ( x56 & n31265 ) | ( n31259 & n31265 ) ;
  assign n31267 = ( n6164 & n31264 ) | ( n6164 & n31266 ) | ( n31264 & n31266 ) ;
  assign n31268 = x56 & ~n31266 ;
  assign n31269 = x56 & ~n31262 ;
  assign n31270 = ( ~n6164 & n31268 ) | ( ~n6164 & n31269 ) | ( n31268 & n31269 ) ;
  assign n31271 = ( n31263 & ~n31267 ) | ( n31263 & n31270 ) | ( ~n31267 & n31270 ) ;
  assign n31272 = ~n31254 & n31271 ;
  assign n31273 = n31254 & ~n31271 ;
  assign n31274 = n31272 | n31273 ;
  assign n31275 = ( n30888 & ~n30889 ) | ( n30888 & n30914 ) | ( ~n30889 & n30914 ) ;
  assign n31276 = ~n31274 & n31275 ;
  assign n31277 = n31274 & ~n31275 ;
  assign n31278 = n31276 | n31277 ;
  assign n31279 = x102 & n12574 ;
  assign n31280 = x101 & n12569 ;
  assign n31281 = x100 & ~n12568 ;
  assign n31282 = n13076 & n31281 ;
  assign n31283 = n31280 | n31282 ;
  assign n31284 = n31279 | n31283 ;
  assign n31285 = n12577 | n31279 ;
  assign n31286 = n31283 | n31285 ;
  assign n31287 = ( n7178 & n31284 ) | ( n7178 & n31286 ) | ( n31284 & n31286 ) ;
  assign n31288 = x53 & n31286 ;
  assign n31289 = x53 & n31279 ;
  assign n31290 = ( x53 & n31283 ) | ( x53 & n31289 ) | ( n31283 & n31289 ) ;
  assign n31291 = ( n7178 & n31288 ) | ( n7178 & n31290 ) | ( n31288 & n31290 ) ;
  assign n31292 = x53 & ~n31290 ;
  assign n31293 = x53 & ~n31286 ;
  assign n31294 = ( ~n7178 & n31292 ) | ( ~n7178 & n31293 ) | ( n31292 & n31293 ) ;
  assign n31295 = ( n31287 & ~n31291 ) | ( n31287 & n31294 ) | ( ~n31291 & n31294 ) ;
  assign n31296 = n31278 | n31295 ;
  assign n31297 = n31278 & ~n31295 ;
  assign n31298 = ( ~n31278 & n31296 ) | ( ~n31278 & n31297 ) | ( n31296 & n31297 ) ;
  assign n31301 = ~n31298 & n31300 ;
  assign n31302 = n31300 & ~n31301 ;
  assign n31303 = x105 & n11205 ;
  assign n31304 = x104 & n11200 ;
  assign n31305 = x103 & ~n11199 ;
  assign n31306 = n11679 & n31305 ;
  assign n31307 = n31304 | n31306 ;
  assign n31308 = n31303 | n31307 ;
  assign n31309 = n11208 | n31303 ;
  assign n31310 = n31307 | n31309 ;
  assign n31311 = ( n8273 & n31308 ) | ( n8273 & n31310 ) | ( n31308 & n31310 ) ;
  assign n31312 = x50 & n31310 ;
  assign n31313 = x50 & n31303 ;
  assign n31314 = ( x50 & n31307 ) | ( x50 & n31313 ) | ( n31307 & n31313 ) ;
  assign n31315 = ( n8273 & n31312 ) | ( n8273 & n31314 ) | ( n31312 & n31314 ) ;
  assign n31316 = x50 & ~n31314 ;
  assign n31317 = x50 & ~n31310 ;
  assign n31318 = ( ~n8273 & n31316 ) | ( ~n8273 & n31317 ) | ( n31316 & n31317 ) ;
  assign n31319 = ( n31311 & ~n31315 ) | ( n31311 & n31318 ) | ( ~n31315 & n31318 ) ;
  assign n31320 = n31298 | n31300 ;
  assign n31321 = n31319 | n31320 ;
  assign n31322 = ( ~n31302 & n31319 ) | ( ~n31302 & n31321 ) | ( n31319 & n31321 ) ;
  assign n31323 = n31319 & n31320 ;
  assign n31324 = ~n31302 & n31323 ;
  assign n31325 = n31322 & ~n31324 ;
  assign n31326 = n31196 & ~n31325 ;
  assign n31327 = ~n31196 & n31325 ;
  assign n31328 = n31326 | n31327 ;
  assign n31329 = x108 & n9933 ;
  assign n31330 = x107 & n9928 ;
  assign n31331 = x106 & ~n9927 ;
  assign n31332 = n10379 & n31331 ;
  assign n31333 = n31330 | n31332 ;
  assign n31334 = n31329 | n31333 ;
  assign n31335 = n9936 | n31329 ;
  assign n31336 = n31333 | n31335 ;
  assign n31337 = ( n9479 & n31334 ) | ( n9479 & n31336 ) | ( n31334 & n31336 ) ;
  assign n31338 = x47 & n31336 ;
  assign n31339 = x47 & n31329 ;
  assign n31340 = ( x47 & n31333 ) | ( x47 & n31339 ) | ( n31333 & n31339 ) ;
  assign n31341 = ( n9479 & n31338 ) | ( n9479 & n31340 ) | ( n31338 & n31340 ) ;
  assign n31342 = x47 & ~n31340 ;
  assign n31343 = x47 & ~n31336 ;
  assign n31344 = ( ~n9479 & n31342 ) | ( ~n9479 & n31343 ) | ( n31342 & n31343 ) ;
  assign n31345 = ( n31337 & ~n31341 ) | ( n31337 & n31344 ) | ( ~n31341 & n31344 ) ;
  assign n31346 = ~n31328 & n31345 ;
  assign n31347 = n31328 & ~n31345 ;
  assign n31348 = n31346 | n31347 ;
  assign n31349 = n30967 | n30986 ;
  assign n31350 = ( n30967 & ~n30969 ) | ( n30967 & n31349 ) | ( ~n30969 & n31349 ) ;
  assign n31351 = ~n31348 & n31350 ;
  assign n31352 = n31348 & ~n31350 ;
  assign n31353 = n31351 | n31352 ;
  assign n31354 = x111 & n8724 ;
  assign n31355 = x110 & n8719 ;
  assign n31356 = x109 & ~n8718 ;
  assign n31357 = n9149 & n31356 ;
  assign n31358 = n31355 | n31357 ;
  assign n31359 = n31354 | n31358 ;
  assign n31360 = n8727 | n31354 ;
  assign n31361 = n31358 | n31360 ;
  assign n31362 = ( n10749 & n31359 ) | ( n10749 & n31361 ) | ( n31359 & n31361 ) ;
  assign n31363 = x44 & n31361 ;
  assign n31364 = x44 & n31354 ;
  assign n31365 = ( x44 & n31358 ) | ( x44 & n31364 ) | ( n31358 & n31364 ) ;
  assign n31366 = ( n10749 & n31363 ) | ( n10749 & n31365 ) | ( n31363 & n31365 ) ;
  assign n31367 = x44 & ~n31365 ;
  assign n31368 = x44 & ~n31361 ;
  assign n31369 = ( ~n10749 & n31367 ) | ( ~n10749 & n31368 ) | ( n31367 & n31368 ) ;
  assign n31370 = ( n31362 & ~n31366 ) | ( n31362 & n31369 ) | ( ~n31366 & n31369 ) ;
  assign n31371 = n31353 | n31370 ;
  assign n31372 = n31353 & ~n31370 ;
  assign n31373 = ( ~n31353 & n31371 ) | ( ~n31353 & n31372 ) | ( n31371 & n31372 ) ;
  assign n31374 = ( n30994 & ~n30995 ) | ( n30994 & n31018 ) | ( ~n30995 & n31018 ) ;
  assign n31375 = n31373 & ~n31374 ;
  assign n31376 = ~n31373 & n31374 ;
  assign n31377 = n31375 | n31376 ;
  assign n31378 = x114 & n7566 ;
  assign n31379 = x113 & n7561 ;
  assign n31380 = x112 & ~n7560 ;
  assign n31381 = n7953 & n31380 ;
  assign n31382 = n31379 | n31381 ;
  assign n31383 = n31378 | n31382 ;
  assign n31384 = n7569 | n31378 ;
  assign n31385 = n31382 | n31384 ;
  assign n31386 = ( ~n12095 & n31383 ) | ( ~n12095 & n31385 ) | ( n31383 & n31385 ) ;
  assign n31387 = n31383 & n31385 ;
  assign n31388 = ( n12079 & n31386 ) | ( n12079 & n31387 ) | ( n31386 & n31387 ) ;
  assign n31389 = x41 & n31388 ;
  assign n31390 = x41 & ~n31388 ;
  assign n31391 = ( n31388 & ~n31389 ) | ( n31388 & n31390 ) | ( ~n31389 & n31390 ) ;
  assign n31392 = n31377 & ~n31391 ;
  assign n31393 = ~n31377 & n31391 ;
  assign n31394 = n31392 | n31393 ;
  assign n31395 = n31015 | n31037 ;
  assign n31396 = n31019 & ~n31037 ;
  assign n31397 = ( n31016 & n31395 ) | ( n31016 & ~n31396 ) | ( n31395 & ~n31396 ) ;
  assign n31398 = ( n31020 & ~n31023 ) | ( n31020 & n31397 ) | ( ~n31023 & n31397 ) ;
  assign n31399 = n31394 & n31398 ;
  assign n31400 = ~n31394 & n31398 ;
  assign n31401 = x117 & n6536 ;
  assign n31402 = x116 & n6531 ;
  assign n31403 = x115 & ~n6530 ;
  assign n31404 = n6871 & n31403 ;
  assign n31405 = n31402 | n31404 ;
  assign n31406 = n31401 | n31405 ;
  assign n31407 = n6539 | n31401 ;
  assign n31408 = n31405 | n31407 ;
  assign n31409 = ( ~n13522 & n31406 ) | ( ~n13522 & n31408 ) | ( n31406 & n31408 ) ;
  assign n31410 = n31406 & n31408 ;
  assign n31411 = ( n13503 & n31409 ) | ( n13503 & n31410 ) | ( n31409 & n31410 ) ;
  assign n31412 = x38 & n31411 ;
  assign n31413 = x38 & ~n31411 ;
  assign n31414 = ( n31411 & ~n31412 ) | ( n31411 & n31413 ) | ( ~n31412 & n31413 ) ;
  assign n31415 = n31394 & ~n31414 ;
  assign n31416 = ( n31400 & ~n31414 ) | ( n31400 & n31415 ) | ( ~n31414 & n31415 ) ;
  assign n31417 = ~n31399 & n31416 ;
  assign n31418 = n31394 | n31398 ;
  assign n31419 = n31394 & n31414 ;
  assign n31420 = n31398 & n31419 ;
  assign n31421 = ( n31414 & ~n31418 ) | ( n31414 & n31420 ) | ( ~n31418 & n31420 ) ;
  assign n31422 = n31417 | n31421 ;
  assign n31423 = n31042 & ~n31059 ;
  assign n31424 = ( n30828 & n31059 ) | ( n30828 & ~n31423 ) | ( n31059 & ~n31423 ) ;
  assign n31425 = ( n31044 & ~n31045 ) | ( n31044 & n31424 ) | ( ~n31045 & n31424 ) ;
  assign n31426 = ~n31422 & n31425 ;
  assign n31427 = n31422 & ~n31425 ;
  assign n31428 = n31426 | n31427 ;
  assign n31429 = x120 & n5554 ;
  assign n31430 = x119 & n5549 ;
  assign n31431 = x118 & ~n5548 ;
  assign n31432 = n5893 & n31431 ;
  assign n31433 = n31430 | n31432 ;
  assign n31434 = n31429 | n31433 ;
  assign n31435 = n5557 | n31429 ;
  assign n31436 = n31433 | n31435 ;
  assign n31437 = ( n14991 & n31434 ) | ( n14991 & n31436 ) | ( n31434 & n31436 ) ;
  assign n31438 = x35 & n31436 ;
  assign n31439 = x35 & n31429 ;
  assign n31440 = ( x35 & n31433 ) | ( x35 & n31439 ) | ( n31433 & n31439 ) ;
  assign n31441 = ( n14991 & n31438 ) | ( n14991 & n31440 ) | ( n31438 & n31440 ) ;
  assign n31442 = x35 & ~n31440 ;
  assign n31443 = x35 & ~n31436 ;
  assign n31444 = ( ~n14991 & n31442 ) | ( ~n14991 & n31443 ) | ( n31442 & n31443 ) ;
  assign n31445 = ( n31437 & ~n31441 ) | ( n31437 & n31444 ) | ( ~n31441 & n31444 ) ;
  assign n31446 = n31428 | n31445 ;
  assign n31447 = n31428 & ~n31445 ;
  assign n31448 = ( ~n31428 & n31446 ) | ( ~n31428 & n31447 ) | ( n31446 & n31447 ) ;
  assign n31449 = n31195 | n31448 ;
  assign n31450 = ~n31192 & n31448 ;
  assign n31451 = n31194 & n31450 ;
  assign n31452 = n31449 & ~n31451 ;
  assign n31453 = ~n31168 & n31452 ;
  assign n31454 = n31168 & ~n31452 ;
  assign n31455 = n31453 | n31454 ;
  assign n31456 = ~n30797 & n31140 ;
  assign n31457 = ( n30779 & n31140 ) | ( n30779 & n31456 ) | ( n31140 & n31456 ) ;
  assign n31458 = ( ~n30668 & n31140 ) | ( ~n30668 & n31456 ) | ( n31140 & n31456 ) ;
  assign n31459 = ( n30669 & n31457 ) | ( n30669 & n31458 ) | ( n31457 & n31458 ) ;
  assign n31460 = ~n31455 & n31459 ;
  assign n31461 = n31092 & n31460 ;
  assign n31462 = ( n31146 & n31455 ) | ( n31146 & ~n31461 ) | ( n31455 & ~n31461 ) ;
  assign n31463 = n31455 & ~n31459 ;
  assign n31464 = ( ~n31092 & n31455 ) | ( ~n31092 & n31463 ) | ( n31455 & n31463 ) ;
  assign n31465 = n31146 & n31464 ;
  assign n31466 = n31462 & ~n31465 ;
  assign n31467 = n31121 & n31466 ;
  assign n31468 = n31121 | n31466 ;
  assign n31469 = ~n31467 & n31468 ;
  assign n31470 = n31110 | n31118 ;
  assign n31471 = n31110 | n31113 ;
  assign n31472 = n31111 | n31471 ;
  assign n31473 = ( n30754 & n31470 ) | ( n30754 & n31472 ) | ( n31470 & n31472 ) ;
  assign n31474 = n31469 | n31473 ;
  assign n31475 = n31469 & n31472 ;
  assign n31476 = n31110 & n31469 ;
  assign n31477 = ( n31118 & n31469 ) | ( n31118 & n31476 ) | ( n31469 & n31476 ) ;
  assign n31478 = ( n30754 & n31475 ) | ( n30754 & n31477 ) | ( n31475 & n31477 ) ;
  assign n31479 = n31474 & ~n31478 ;
  assign n31480 = x127 & n3816 ;
  assign n31481 = x126 & n3811 ;
  assign n31482 = x125 & ~n3810 ;
  assign n31483 = n4067 & n31482 ;
  assign n31484 = n31481 | n31483 ;
  assign n31485 = n31480 | n31484 ;
  assign n31486 = n3819 | n31480 ;
  assign n31487 = n31484 | n31486 ;
  assign n31488 = ( n18763 & n31485 ) | ( n18763 & n31487 ) | ( n31485 & n31487 ) ;
  assign n31489 = x29 & n31487 ;
  assign n31490 = x29 & n31480 ;
  assign n31491 = ( x29 & n31484 ) | ( x29 & n31490 ) | ( n31484 & n31490 ) ;
  assign n31492 = ( n18763 & n31489 ) | ( n18763 & n31491 ) | ( n31489 & n31491 ) ;
  assign n31493 = x29 & ~n31491 ;
  assign n31494 = x29 & ~n31487 ;
  assign n31495 = ( ~n18763 & n31493 ) | ( ~n18763 & n31494 ) | ( n31493 & n31494 ) ;
  assign n31496 = ( n31488 & ~n31492 ) | ( n31488 & n31495 ) | ( ~n31492 & n31495 ) ;
  assign n31497 = n31163 & n31496 ;
  assign n31498 = n31165 & n31497 ;
  assign n31499 = ( ~n31452 & n31496 ) | ( ~n31452 & n31498 ) | ( n31496 & n31498 ) ;
  assign n31500 = n31496 & n31497 ;
  assign n31501 = n31165 & n31500 ;
  assign n31502 = ( n31168 & n31499 ) | ( n31168 & n31501 ) | ( n31499 & n31501 ) ;
  assign n31503 = ~n31167 & n31452 ;
  assign n31504 = ( n31167 & n31168 ) | ( n31167 & ~n31503 ) | ( n31168 & ~n31503 ) ;
  assign n31505 = ~n31502 & n31504 ;
  assign n31506 = n31400 | n31421 ;
  assign n31507 = x97 & n15552 ;
  assign n31508 = x96 & n15547 ;
  assign n31509 = x95 & ~n15546 ;
  assign n31510 = n16123 & n31509 ;
  assign n31511 = n31508 | n31510 ;
  assign n31512 = n31507 | n31511 ;
  assign n31513 = n15555 | n31507 ;
  assign n31514 = n31511 | n31513 ;
  assign n31515 = ( n5505 & n31512 ) | ( n5505 & n31514 ) | ( n31512 & n31514 ) ;
  assign n31516 = x59 & n31514 ;
  assign n31517 = x59 & n31507 ;
  assign n31518 = ( x59 & n31511 ) | ( x59 & n31517 ) | ( n31511 & n31517 ) ;
  assign n31519 = ( n5505 & n31516 ) | ( n5505 & n31518 ) | ( n31516 & n31518 ) ;
  assign n31520 = x59 & ~n31518 ;
  assign n31521 = x59 & ~n31514 ;
  assign n31522 = ( ~n5505 & n31520 ) | ( ~n5505 & n31521 ) | ( n31520 & n31521 ) ;
  assign n31523 = ( n31515 & ~n31519 ) | ( n31515 & n31522 ) | ( ~n31519 & n31522 ) ;
  assign n31524 = n31225 | n31245 ;
  assign n31525 = ( ~n31223 & n31245 ) | ( ~n31223 & n31524 ) | ( n31245 & n31524 ) ;
  assign n31526 = n31523 | n31525 ;
  assign n31527 = n31226 | n31523 ;
  assign n31528 = ( ~n31228 & n31526 ) | ( ~n31228 & n31527 ) | ( n31526 & n31527 ) ;
  assign n31529 = n31523 & n31525 ;
  assign n31530 = n31226 & n31523 ;
  assign n31531 = ( ~n31228 & n31529 ) | ( ~n31228 & n31530 ) | ( n31529 & n31530 ) ;
  assign n31532 = n31528 & ~n31531 ;
  assign n31533 = x91 & n18290 ;
  assign n31534 = x63 & x90 ;
  assign n31535 = ~n18290 & n31534 ;
  assign n31536 = n31533 | n31535 ;
  assign n31537 = ~x26 & n31536 ;
  assign n31538 = x26 & ~n31536 ;
  assign n31539 = n31537 | n31538 ;
  assign n31540 = n31200 & ~n31539 ;
  assign n31541 = ~n31200 & n31539 ;
  assign n31542 = n31540 | n31541 ;
  assign n31543 = ( ~n31201 & n31203 ) | ( ~n31201 & n31542 ) | ( n31203 & n31542 ) ;
  assign n31544 = n31201 & ~n31542 ;
  assign n31545 = ( n31220 & ~n31543 ) | ( n31220 & n31544 ) | ( ~n31543 & n31544 ) ;
  assign n31546 = ~n31201 & n31203 ;
  assign n31547 = n31542 & n31546 ;
  assign n31548 = ~n31201 & n31542 ;
  assign n31549 = ( ~n31220 & n31547 ) | ( ~n31220 & n31548 ) | ( n31547 & n31548 ) ;
  assign n31550 = n31545 | n31549 ;
  assign n31551 = x94 & n17146 ;
  assign n31552 = x93 & n17141 ;
  assign n31553 = x92 & ~n17140 ;
  assign n31554 = n17724 & n31553 ;
  assign n31555 = n31552 | n31554 ;
  assign n31556 = n31551 | n31555 ;
  assign n31557 = n17149 | n31551 ;
  assign n31558 = n31555 | n31557 ;
  assign n31559 = ( n4583 & n31556 ) | ( n4583 & n31558 ) | ( n31556 & n31558 ) ;
  assign n31560 = x62 & n31558 ;
  assign n31561 = x62 & n31551 ;
  assign n31562 = ( x62 & n31555 ) | ( x62 & n31561 ) | ( n31555 & n31561 ) ;
  assign n31563 = ( n4583 & n31560 ) | ( n4583 & n31562 ) | ( n31560 & n31562 ) ;
  assign n31564 = x62 & ~n31562 ;
  assign n31565 = x62 & ~n31558 ;
  assign n31566 = ( ~n4583 & n31564 ) | ( ~n4583 & n31565 ) | ( n31564 & n31565 ) ;
  assign n31567 = ( n31559 & ~n31563 ) | ( n31559 & n31566 ) | ( ~n31563 & n31566 ) ;
  assign n31568 = ~n31550 & n31567 ;
  assign n31569 = n31550 | n31568 ;
  assign n31570 = n31550 & n31567 ;
  assign n31571 = n31569 & ~n31570 ;
  assign n31572 = ~n31532 & n31571 ;
  assign n31573 = n31532 & ~n31571 ;
  assign n31574 = n31572 | n31573 ;
  assign n31575 = x100 & n14045 ;
  assign n31576 = x99 & n14040 ;
  assign n31577 = x98 & ~n14039 ;
  assign n31578 = n14552 & n31577 ;
  assign n31579 = n31576 | n31578 ;
  assign n31580 = n31575 | n31579 ;
  assign n31581 = n14048 | n31575 ;
  assign n31582 = n31579 | n31581 ;
  assign n31583 = ( n6483 & n31580 ) | ( n6483 & n31582 ) | ( n31580 & n31582 ) ;
  assign n31584 = x56 & n31582 ;
  assign n31585 = x56 & n31575 ;
  assign n31586 = ( x56 & n31579 ) | ( x56 & n31585 ) | ( n31579 & n31585 ) ;
  assign n31587 = ( n6483 & n31584 ) | ( n6483 & n31586 ) | ( n31584 & n31586 ) ;
  assign n31588 = x56 & ~n31586 ;
  assign n31589 = x56 & ~n31582 ;
  assign n31590 = ( ~n6483 & n31588 ) | ( ~n6483 & n31589 ) | ( n31588 & n31589 ) ;
  assign n31591 = ( n31583 & ~n31587 ) | ( n31583 & n31590 ) | ( ~n31587 & n31590 ) ;
  assign n31592 = ~n31574 & n31591 ;
  assign n31593 = n31574 | n31592 ;
  assign n31595 = n31252 | n31271 ;
  assign n31596 = ( n31252 & ~n31254 ) | ( n31252 & n31595 ) | ( ~n31254 & n31595 ) ;
  assign n31594 = n31574 & n31591 ;
  assign n31597 = n31594 & n31596 ;
  assign n31598 = ( ~n31593 & n31596 ) | ( ~n31593 & n31597 ) | ( n31596 & n31597 ) ;
  assign n31599 = n31594 | n31596 ;
  assign n31600 = n31593 & ~n31599 ;
  assign n31601 = n31598 | n31600 ;
  assign n31602 = x103 & n12574 ;
  assign n31603 = x102 & n12569 ;
  assign n31604 = x101 & ~n12568 ;
  assign n31605 = n13076 & n31604 ;
  assign n31606 = n31603 | n31605 ;
  assign n31607 = n31602 | n31606 ;
  assign n31608 = n12577 | n31602 ;
  assign n31609 = n31606 | n31608 ;
  assign n31610 = ( n7529 & n31607 ) | ( n7529 & n31609 ) | ( n31607 & n31609 ) ;
  assign n31611 = x53 & n31609 ;
  assign n31612 = x53 & n31602 ;
  assign n31613 = ( x53 & n31606 ) | ( x53 & n31612 ) | ( n31606 & n31612 ) ;
  assign n31614 = ( n7529 & n31611 ) | ( n7529 & n31613 ) | ( n31611 & n31613 ) ;
  assign n31615 = x53 & ~n31613 ;
  assign n31616 = x53 & ~n31609 ;
  assign n31617 = ( ~n7529 & n31615 ) | ( ~n7529 & n31616 ) | ( n31615 & n31616 ) ;
  assign n31618 = ( n31610 & ~n31614 ) | ( n31610 & n31617 ) | ( ~n31614 & n31617 ) ;
  assign n31619 = ~n31601 & n31618 ;
  assign n31620 = n31601 | n31619 ;
  assign n31622 = n31276 | n31295 ;
  assign n31623 = ( n31276 & ~n31278 ) | ( n31276 & n31622 ) | ( ~n31278 & n31622 ) ;
  assign n31621 = n31601 & n31618 ;
  assign n31624 = n31621 & n31623 ;
  assign n31625 = ( ~n31620 & n31623 ) | ( ~n31620 & n31624 ) | ( n31623 & n31624 ) ;
  assign n31626 = n31621 | n31623 ;
  assign n31627 = n31620 & ~n31626 ;
  assign n31628 = n31625 | n31627 ;
  assign n31629 = x106 & n11205 ;
  assign n31630 = x105 & n11200 ;
  assign n31631 = x104 & ~n11199 ;
  assign n31632 = n11679 & n31631 ;
  assign n31633 = n31630 | n31632 ;
  assign n31634 = n31629 | n31633 ;
  assign n31635 = n11208 | n31629 ;
  assign n31636 = n31633 | n31635 ;
  assign n31637 = ( n8656 & n31634 ) | ( n8656 & n31636 ) | ( n31634 & n31636 ) ;
  assign n31638 = x50 & n31636 ;
  assign n31639 = x50 & n31629 ;
  assign n31640 = ( x50 & n31633 ) | ( x50 & n31639 ) | ( n31633 & n31639 ) ;
  assign n31641 = ( n8656 & n31638 ) | ( n8656 & n31640 ) | ( n31638 & n31640 ) ;
  assign n31642 = x50 & ~n31640 ;
  assign n31643 = x50 & ~n31636 ;
  assign n31644 = ( ~n8656 & n31642 ) | ( ~n8656 & n31643 ) | ( n31642 & n31643 ) ;
  assign n31645 = ( n31637 & ~n31641 ) | ( n31637 & n31644 ) | ( ~n31641 & n31644 ) ;
  assign n31646 = ~n31628 & n31645 ;
  assign n31647 = n31628 | n31646 ;
  assign n31648 = ( ~n31298 & n31300 ) | ( ~n31298 & n31319 ) | ( n31300 & n31319 ) ;
  assign n31649 = n31645 & ~n31648 ;
  assign n31650 = n31628 & n31649 ;
  assign n31651 = ( n31647 & n31648 ) | ( n31647 & ~n31650 ) | ( n31648 & ~n31650 ) ;
  assign n31652 = ~n31645 & n31648 ;
  assign n31653 = ( ~n31628 & n31648 ) | ( ~n31628 & n31652 ) | ( n31648 & n31652 ) ;
  assign n31654 = n31647 & n31653 ;
  assign n31655 = n31651 & ~n31654 ;
  assign n31656 = x109 & n9933 ;
  assign n31657 = x108 & n9928 ;
  assign n31658 = x107 & ~n9927 ;
  assign n31659 = n10379 & n31658 ;
  assign n31660 = n31657 | n31659 ;
  assign n31661 = n31656 | n31660 ;
  assign n31662 = n9936 | n31656 ;
  assign n31663 = n31660 | n31662 ;
  assign n31664 = ( n9878 & n31661 ) | ( n9878 & n31663 ) | ( n31661 & n31663 ) ;
  assign n31665 = x47 & n31663 ;
  assign n31666 = x47 & n31656 ;
  assign n31667 = ( x47 & n31660 ) | ( x47 & n31666 ) | ( n31660 & n31666 ) ;
  assign n31668 = ( n9878 & n31665 ) | ( n9878 & n31667 ) | ( n31665 & n31667 ) ;
  assign n31669 = x47 & ~n31667 ;
  assign n31670 = x47 & ~n31663 ;
  assign n31671 = ( ~n9878 & n31669 ) | ( ~n9878 & n31670 ) | ( n31669 & n31670 ) ;
  assign n31672 = ( n31664 & ~n31668 ) | ( n31664 & n31671 ) | ( ~n31668 & n31671 ) ;
  assign n31673 = ~n31655 & n31672 ;
  assign n31674 = n31655 & ~n31672 ;
  assign n31675 = n31673 | n31674 ;
  assign n31676 = n31325 & ~n31345 ;
  assign n31677 = ( n31196 & n31345 ) | ( n31196 & ~n31676 ) | ( n31345 & ~n31676 ) ;
  assign n31678 = ( n31326 & ~n31328 ) | ( n31326 & n31677 ) | ( ~n31328 & n31677 ) ;
  assign n31679 = n31675 & ~n31678 ;
  assign n31680 = ~n31675 & n31678 ;
  assign n31681 = n31679 | n31680 ;
  assign n31682 = x112 & n8724 ;
  assign n31683 = x111 & n8719 ;
  assign n31684 = x110 & ~n8718 ;
  assign n31685 = n9149 & n31684 ;
  assign n31686 = n31683 | n31685 ;
  assign n31687 = n31682 | n31686 ;
  assign n31688 = n8727 | n31682 ;
  assign n31689 = n31686 | n31688 ;
  assign n31690 = ( n11172 & n31687 ) | ( n11172 & n31689 ) | ( n31687 & n31689 ) ;
  assign n31691 = x44 & n31689 ;
  assign n31692 = x44 & n31682 ;
  assign n31693 = ( x44 & n31686 ) | ( x44 & n31692 ) | ( n31686 & n31692 ) ;
  assign n31694 = ( n11172 & n31691 ) | ( n11172 & n31693 ) | ( n31691 & n31693 ) ;
  assign n31695 = x44 & ~n31693 ;
  assign n31696 = x44 & ~n31689 ;
  assign n31697 = ( ~n11172 & n31695 ) | ( ~n11172 & n31696 ) | ( n31695 & n31696 ) ;
  assign n31698 = ( n31690 & ~n31694 ) | ( n31690 & n31697 ) | ( ~n31694 & n31697 ) ;
  assign n31699 = ~n31681 & n31698 ;
  assign n31700 = n31681 | n31699 ;
  assign n31701 = n31681 & n31698 ;
  assign n31702 = n31700 & ~n31701 ;
  assign n31703 = n31351 | n31370 ;
  assign n31704 = ( n31351 & ~n31353 ) | ( n31351 & n31703 ) | ( ~n31353 & n31703 ) ;
  assign n31705 = n31702 & ~n31704 ;
  assign n31706 = ~n31702 & n31704 ;
  assign n31707 = n31705 | n31706 ;
  assign n31708 = x115 & n7566 ;
  assign n31709 = x114 & n7561 ;
  assign n31710 = x113 & ~n7560 ;
  assign n31711 = n7953 & n31710 ;
  assign n31712 = n31709 | n31711 ;
  assign n31713 = n31708 | n31712 ;
  assign n31714 = n7569 | n31708 ;
  assign n31715 = n31712 | n31714 ;
  assign n31716 = ( ~n12550 & n31713 ) | ( ~n12550 & n31715 ) | ( n31713 & n31715 ) ;
  assign n31717 = n31713 & n31715 ;
  assign n31718 = ( n12532 & n31716 ) | ( n12532 & n31717 ) | ( n31716 & n31717 ) ;
  assign n31719 = x41 & n31718 ;
  assign n31720 = x41 & ~n31718 ;
  assign n31721 = ( n31718 & ~n31719 ) | ( n31718 & n31720 ) | ( ~n31719 & n31720 ) ;
  assign n31722 = ~n31707 & n31721 ;
  assign n31723 = n31707 & ~n31721 ;
  assign n31724 = n31722 | n31723 ;
  assign n31725 = n31376 | n31391 ;
  assign n31726 = ( n31376 & ~n31377 ) | ( n31376 & n31725 ) | ( ~n31377 & n31725 ) ;
  assign n31727 = ~n31724 & n31726 ;
  assign n31728 = n31724 | n31727 ;
  assign n31729 = x118 & n6536 ;
  assign n31730 = x117 & n6531 ;
  assign n31731 = x116 & ~n6530 ;
  assign n31732 = n6871 & n31731 ;
  assign n31733 = n31730 | n31732 ;
  assign n31734 = n31729 | n31733 ;
  assign n31735 = n6539 | n31729 ;
  assign n31736 = n31733 | n31735 ;
  assign n31737 = ( ~n14002 & n31734 ) | ( ~n14002 & n31736 ) | ( n31734 & n31736 ) ;
  assign n31738 = n31734 & n31736 ;
  assign n31739 = ( n13981 & n31737 ) | ( n13981 & n31738 ) | ( n31737 & n31738 ) ;
  assign n31740 = x38 & n31739 ;
  assign n31741 = x38 & ~n31739 ;
  assign n31742 = ( n31739 & ~n31740 ) | ( n31739 & n31741 ) | ( ~n31740 & n31741 ) ;
  assign n31743 = n31726 & n31742 ;
  assign n31744 = n31724 & n31743 ;
  assign n31745 = ( ~n31728 & n31742 ) | ( ~n31728 & n31744 ) | ( n31742 & n31744 ) ;
  assign n31746 = n31726 | n31742 ;
  assign n31747 = ( n31724 & n31742 ) | ( n31724 & n31746 ) | ( n31742 & n31746 ) ;
  assign n31748 = n31728 & ~n31747 ;
  assign n31749 = n31745 | n31748 ;
  assign n31750 = n31506 & ~n31749 ;
  assign n31751 = ~n31506 & n31749 ;
  assign n31752 = n31750 | n31751 ;
  assign n31753 = x121 & n5554 ;
  assign n31754 = x120 & n5549 ;
  assign n31755 = x119 & ~n5548 ;
  assign n31756 = n5893 & n31755 ;
  assign n31757 = n31754 | n31756 ;
  assign n31758 = n31753 | n31757 ;
  assign n31759 = n5557 | n31753 ;
  assign n31760 = n31757 | n31759 ;
  assign n31761 = ( n15501 & n31758 ) | ( n15501 & n31760 ) | ( n31758 & n31760 ) ;
  assign n31762 = x35 & n31760 ;
  assign n31763 = x35 & n31753 ;
  assign n31764 = ( x35 & n31757 ) | ( x35 & n31763 ) | ( n31757 & n31763 ) ;
  assign n31765 = ( n15501 & n31762 ) | ( n15501 & n31764 ) | ( n31762 & n31764 ) ;
  assign n31766 = x35 & ~n31764 ;
  assign n31767 = x35 & ~n31760 ;
  assign n31768 = ( ~n15501 & n31766 ) | ( ~n15501 & n31767 ) | ( n31766 & n31767 ) ;
  assign n31769 = ( n31761 & ~n31765 ) | ( n31761 & n31768 ) | ( ~n31765 & n31768 ) ;
  assign n31770 = ~n31752 & n31769 ;
  assign n31771 = n31752 | n31770 ;
  assign n31773 = n31426 | n31445 ;
  assign n31774 = ( n31426 & ~n31428 ) | ( n31426 & n31773 ) | ( ~n31428 & n31773 ) ;
  assign n31772 = n31752 & n31769 ;
  assign n31775 = n31772 & n31774 ;
  assign n31776 = ( ~n31771 & n31774 ) | ( ~n31771 & n31775 ) | ( n31774 & n31775 ) ;
  assign n31777 = n31772 | n31774 ;
  assign n31778 = n31771 & ~n31777 ;
  assign n31779 = n31776 | n31778 ;
  assign n31780 = x124 & n4631 ;
  assign n31781 = x123 & n4626 ;
  assign n31782 = x122 & ~n4625 ;
  assign n31783 = n4943 & n31782 ;
  assign n31784 = n31781 | n31783 ;
  assign n31785 = n31780 | n31784 ;
  assign n31786 = n4634 | n31780 ;
  assign n31787 = n31784 | n31786 ;
  assign n31788 = ( n17084 & n31785 ) | ( n17084 & n31787 ) | ( n31785 & n31787 ) ;
  assign n31789 = x32 & n31787 ;
  assign n31790 = x32 & n31780 ;
  assign n31791 = ( x32 & n31784 ) | ( x32 & n31790 ) | ( n31784 & n31790 ) ;
  assign n31792 = ( n17084 & n31789 ) | ( n17084 & n31791 ) | ( n31789 & n31791 ) ;
  assign n31793 = x32 & ~n31791 ;
  assign n31794 = x32 & ~n31787 ;
  assign n31795 = ( ~n17084 & n31793 ) | ( ~n17084 & n31794 ) | ( n31793 & n31794 ) ;
  assign n31796 = ( n31788 & ~n31792 ) | ( n31788 & n31795 ) | ( ~n31792 & n31795 ) ;
  assign n31797 = ( n31192 & n31195 ) | ( n31192 & ~n31450 ) | ( n31195 & ~n31450 ) ;
  assign n31798 = n31796 | n31797 ;
  assign n31799 = n31796 & n31797 ;
  assign n31800 = n31798 & ~n31799 ;
  assign n31801 = n31779 | n31800 ;
  assign n31802 = n31779 & n31800 ;
  assign n31803 = n31801 & ~n31802 ;
  assign n31804 = n31496 & ~n31497 ;
  assign n31805 = ( ~n31165 & n31496 ) | ( ~n31165 & n31804 ) | ( n31496 & n31804 ) ;
  assign n31806 = n31452 & n31805 ;
  assign n31807 = ( ~n31168 & n31805 ) | ( ~n31168 & n31806 ) | ( n31805 & n31806 ) ;
  assign n31808 = ~n31803 & n31807 ;
  assign n31809 = ( n31505 & ~n31803 ) | ( n31505 & n31808 ) | ( ~n31803 & n31808 ) ;
  assign n31810 = n31803 & ~n31807 ;
  assign n31811 = ~n31505 & n31810 ;
  assign n31812 = n31809 | n31811 ;
  assign n31813 = n31145 & ~n31812 ;
  assign n31814 = ( n31462 & n31812 ) | ( n31462 & ~n31813 ) | ( n31812 & ~n31813 ) ;
  assign n31815 = ~n31145 & n31812 ;
  assign n31816 = n31462 & n31815 ;
  assign n31817 = n31814 & ~n31816 ;
  assign n31818 = n31467 | n31476 ;
  assign n31819 = n31467 | n31469 ;
  assign n31820 = ( n31118 & n31818 ) | ( n31118 & n31819 ) | ( n31818 & n31819 ) ;
  assign n31821 = ( n31467 & n31472 ) | ( n31467 & n31819 ) | ( n31472 & n31819 ) ;
  assign n31822 = ( n30754 & n31820 ) | ( n30754 & n31821 ) | ( n31820 & n31821 ) ;
  assign n31823 = n31817 | n31822 ;
  assign n31824 = n31817 & n31820 ;
  assign n31825 = n31467 & n31817 ;
  assign n31826 = ( n31469 & n31817 ) | ( n31469 & n31825 ) | ( n31817 & n31825 ) ;
  assign n31827 = ( n31472 & n31825 ) | ( n31472 & n31826 ) | ( n31825 & n31826 ) ;
  assign n31828 = ( n30754 & n31824 ) | ( n30754 & n31827 ) | ( n31824 & n31827 ) ;
  assign n31829 = n31823 & ~n31828 ;
  assign n31830 = n31502 | n31809 ;
  assign n31831 = x125 & n4631 ;
  assign n31832 = x124 & n4626 ;
  assign n31833 = x123 & ~n4625 ;
  assign n31834 = n4943 & n31833 ;
  assign n31835 = n31832 | n31834 ;
  assign n31836 = n31831 | n31835 ;
  assign n31837 = n4634 | n31831 ;
  assign n31838 = n31835 | n31837 ;
  assign n31839 = ( n17670 & n31836 ) | ( n17670 & n31838 ) | ( n31836 & n31838 ) ;
  assign n31840 = x32 & n31838 ;
  assign n31841 = x32 & n31831 ;
  assign n31842 = ( x32 & n31835 ) | ( x32 & n31841 ) | ( n31835 & n31841 ) ;
  assign n31843 = ( n17670 & n31840 ) | ( n17670 & n31842 ) | ( n31840 & n31842 ) ;
  assign n31844 = x32 & ~n31842 ;
  assign n31845 = x32 & ~n31838 ;
  assign n31846 = ( ~n17670 & n31844 ) | ( ~n17670 & n31845 ) | ( n31844 & n31845 ) ;
  assign n31847 = ( n31839 & ~n31843 ) | ( n31839 & n31846 ) | ( ~n31843 & n31846 ) ;
  assign n31848 = n31769 & n31847 ;
  assign n31849 = ~n31752 & n31848 ;
  assign n31850 = ( n31774 & n31847 ) | ( n31774 & n31849 ) | ( n31847 & n31849 ) ;
  assign n31851 = ( ~n31771 & n31847 ) | ( ~n31771 & n31849 ) | ( n31847 & n31849 ) ;
  assign n31852 = ( n31775 & n31850 ) | ( n31775 & n31851 ) | ( n31850 & n31851 ) ;
  assign n31853 = n31769 | n31847 ;
  assign n31854 = ( ~n31752 & n31847 ) | ( ~n31752 & n31853 ) | ( n31847 & n31853 ) ;
  assign n31855 = n31774 | n31854 ;
  assign n31856 = n31771 & ~n31854 ;
  assign n31857 = ( n31775 & n31855 ) | ( n31775 & ~n31856 ) | ( n31855 & ~n31856 ) ;
  assign n31858 = ~n31852 & n31857 ;
  assign n31859 = n31745 | n31750 ;
  assign n31860 = n31673 | n31680 ;
  assign n31861 = ( ~n31628 & n31645 ) | ( ~n31628 & n31648 ) | ( n31645 & n31648 ) ;
  assign n31862 = x101 & n14045 ;
  assign n31863 = x100 & n14040 ;
  assign n31864 = x99 & ~n14039 ;
  assign n31865 = n14552 & n31864 ;
  assign n31866 = n31863 | n31865 ;
  assign n31867 = n31862 | n31866 ;
  assign n31868 = n14048 | n31862 ;
  assign n31869 = n31866 | n31868 ;
  assign n31870 = ( n6844 & n31867 ) | ( n6844 & n31869 ) | ( n31867 & n31869 ) ;
  assign n31871 = x56 & n31869 ;
  assign n31872 = x56 & n31862 ;
  assign n31873 = ( x56 & n31866 ) | ( x56 & n31872 ) | ( n31866 & n31872 ) ;
  assign n31874 = ( n6844 & n31871 ) | ( n6844 & n31873 ) | ( n31871 & n31873 ) ;
  assign n31875 = x56 & ~n31873 ;
  assign n31876 = x56 & ~n31869 ;
  assign n31877 = ( ~n6844 & n31875 ) | ( ~n6844 & n31876 ) | ( n31875 & n31876 ) ;
  assign n31878 = ( n31870 & ~n31874 ) | ( n31870 & n31877 ) | ( ~n31874 & n31877 ) ;
  assign n31879 = x92 & n18290 ;
  assign n31880 = x63 & x91 ;
  assign n31881 = ~n18290 & n31880 ;
  assign n31882 = n31879 | n31881 ;
  assign n31883 = n31200 | n31537 ;
  assign n31884 = ( n31537 & ~n31539 ) | ( n31537 & n31883 ) | ( ~n31539 & n31883 ) ;
  assign n31885 = n31882 & ~n31884 ;
  assign n31886 = ~n31882 & n31884 ;
  assign n31887 = n31885 | n31886 ;
  assign n31888 = x94 & n17141 ;
  assign n31889 = x93 & ~n17140 ;
  assign n31890 = n17724 & n31889 ;
  assign n31891 = n31888 | n31890 ;
  assign n31892 = x95 & n17146 ;
  assign n31893 = n17149 | n31892 ;
  assign n31894 = n31891 | n31893 ;
  assign n31895 = x62 & ~n31894 ;
  assign n31896 = ~n31887 & n31895 ;
  assign n31897 = x62 & x95 ;
  assign n31898 = n17146 & n31897 ;
  assign n31899 = x62 & ~n31898 ;
  assign n31900 = ~n31891 & n31899 ;
  assign n31901 = ~n31887 & n31900 ;
  assign n31902 = ( ~n4897 & n31896 ) | ( ~n4897 & n31901 ) | ( n31896 & n31901 ) ;
  assign n31903 = ~x62 & n31894 ;
  assign n31904 = ~x62 & n31892 ;
  assign n31905 = ( ~x62 & n31891 ) | ( ~x62 & n31904 ) | ( n31891 & n31904 ) ;
  assign n31906 = ( n4897 & n31903 ) | ( n4897 & n31905 ) | ( n31903 & n31905 ) ;
  assign n31907 = ( ~n31887 & n31902 ) | ( ~n31887 & n31906 ) | ( n31902 & n31906 ) ;
  assign n31908 = n31887 & ~n31895 ;
  assign n31909 = n31887 & ~n31900 ;
  assign n31910 = ( n4897 & n31908 ) | ( n4897 & n31909 ) | ( n31908 & n31909 ) ;
  assign n31911 = ~n31906 & n31910 ;
  assign n31912 = n31907 | n31911 ;
  assign n31913 = n31545 | n31567 ;
  assign n31914 = ( n31545 & ~n31550 ) | ( n31545 & n31913 ) | ( ~n31550 & n31913 ) ;
  assign n31915 = ~n31912 & n31914 ;
  assign n31916 = n31912 & ~n31914 ;
  assign n31917 = n31915 | n31916 ;
  assign n31918 = x98 & n15552 ;
  assign n31919 = x97 & n15547 ;
  assign n31920 = x96 & ~n15546 ;
  assign n31921 = n16123 & n31920 ;
  assign n31922 = n31919 | n31921 ;
  assign n31923 = n31918 | n31922 ;
  assign n31924 = n15555 | n31918 ;
  assign n31925 = n31922 | n31924 ;
  assign n31926 = ( ~n5850 & n31923 ) | ( ~n5850 & n31925 ) | ( n31923 & n31925 ) ;
  assign n31927 = n31923 & n31925 ;
  assign n31928 = ( n5834 & n31926 ) | ( n5834 & n31927 ) | ( n31926 & n31927 ) ;
  assign n31929 = x59 & n31925 ;
  assign n31930 = x59 & n31918 ;
  assign n31931 = ( x59 & n31922 ) | ( x59 & n31930 ) | ( n31922 & n31930 ) ;
  assign n31932 = ( ~n5850 & n31929 ) | ( ~n5850 & n31931 ) | ( n31929 & n31931 ) ;
  assign n31933 = n31929 & n31931 ;
  assign n31934 = ( n5834 & n31932 ) | ( n5834 & n31933 ) | ( n31932 & n31933 ) ;
  assign n31935 = x59 & ~n31931 ;
  assign n31936 = x59 & ~n31925 ;
  assign n31937 = ( n5850 & n31935 ) | ( n5850 & n31936 ) | ( n31935 & n31936 ) ;
  assign n31938 = n31935 | n31936 ;
  assign n31939 = ( ~n5834 & n31937 ) | ( ~n5834 & n31938 ) | ( n31937 & n31938 ) ;
  assign n31940 = ( n31928 & ~n31934 ) | ( n31928 & n31939 ) | ( ~n31934 & n31939 ) ;
  assign n31941 = n31917 | n31940 ;
  assign n31942 = n31917 & ~n31940 ;
  assign n31943 = ( ~n31917 & n31941 ) | ( ~n31917 & n31942 ) | ( n31941 & n31942 ) ;
  assign n31944 = ~n31531 & n31571 ;
  assign n31945 = ( n31531 & n31532 ) | ( n31531 & ~n31944 ) | ( n31532 & ~n31944 ) ;
  assign n31946 = ( n31878 & n31943 ) | ( n31878 & ~n31945 ) | ( n31943 & ~n31945 ) ;
  assign n31947 = ( ~n31943 & n31945 ) | ( ~n31943 & n31946 ) | ( n31945 & n31946 ) ;
  assign n31948 = ( ~n31878 & n31946 ) | ( ~n31878 & n31947 ) | ( n31946 & n31947 ) ;
  assign n31950 = x104 & n12574 ;
  assign n31951 = x103 & n12569 ;
  assign n31952 = x102 & ~n12568 ;
  assign n31953 = n13076 & n31952 ;
  assign n31954 = n31951 | n31953 ;
  assign n31955 = n31950 | n31954 ;
  assign n31956 = n12577 | n31950 ;
  assign n31957 = n31954 | n31956 ;
  assign n31958 = ( n7911 & n31955 ) | ( n7911 & n31957 ) | ( n31955 & n31957 ) ;
  assign n31959 = x53 & n31957 ;
  assign n31960 = x53 & n31950 ;
  assign n31961 = ( x53 & n31954 ) | ( x53 & n31960 ) | ( n31954 & n31960 ) ;
  assign n31962 = ( n7911 & n31959 ) | ( n7911 & n31961 ) | ( n31959 & n31961 ) ;
  assign n31963 = x53 & ~n31961 ;
  assign n31964 = x53 & ~n31957 ;
  assign n31965 = ( ~n7911 & n31963 ) | ( ~n7911 & n31964 ) | ( n31963 & n31964 ) ;
  assign n31966 = ( n31958 & ~n31962 ) | ( n31958 & n31965 ) | ( ~n31962 & n31965 ) ;
  assign n31967 = ( ~n31592 & n31948 ) | ( ~n31592 & n31966 ) | ( n31948 & n31966 ) ;
  assign n31968 = n31946 & n31966 ;
  assign n31969 = ~n31878 & n31966 ;
  assign n31970 = ( n31947 & n31968 ) | ( n31947 & n31969 ) | ( n31968 & n31969 ) ;
  assign n31971 = ( ~n31598 & n31967 ) | ( ~n31598 & n31970 ) | ( n31967 & n31970 ) ;
  assign n31949 = n31592 | n31598 ;
  assign n31972 = ( n31949 & ~n31966 ) | ( n31949 & n31971 ) | ( ~n31966 & n31971 ) ;
  assign n31973 = ( ~n31948 & n31971 ) | ( ~n31948 & n31972 ) | ( n31971 & n31972 ) ;
  assign n31974 = n31619 & ~n31973 ;
  assign n31975 = ( n31625 & ~n31973 ) | ( n31625 & n31974 ) | ( ~n31973 & n31974 ) ;
  assign n31976 = ~n31619 & n31973 ;
  assign n31977 = ~n31625 & n31976 ;
  assign n31978 = n31975 | n31977 ;
  assign n31979 = x107 & n11205 ;
  assign n31980 = x106 & n11200 ;
  assign n31981 = x105 & ~n11199 ;
  assign n31982 = n11679 & n31981 ;
  assign n31983 = n31980 | n31982 ;
  assign n31984 = n31979 | n31983 ;
  assign n31985 = n11208 | n31979 ;
  assign n31986 = n31983 | n31985 ;
  assign n31987 = ( n9084 & n31984 ) | ( n9084 & n31986 ) | ( n31984 & n31986 ) ;
  assign n31988 = x50 & n31986 ;
  assign n31989 = x50 & n31979 ;
  assign n31990 = ( x50 & n31983 ) | ( x50 & n31989 ) | ( n31983 & n31989 ) ;
  assign n31991 = ( n9084 & n31988 ) | ( n9084 & n31990 ) | ( n31988 & n31990 ) ;
  assign n31992 = x50 & ~n31990 ;
  assign n31993 = x50 & ~n31986 ;
  assign n31994 = ( ~n9084 & n31992 ) | ( ~n9084 & n31993 ) | ( n31992 & n31993 ) ;
  assign n31995 = ( n31987 & ~n31991 ) | ( n31987 & n31994 ) | ( ~n31991 & n31994 ) ;
  assign n31996 = n31978 | n31995 ;
  assign n31997 = n31978 & ~n31995 ;
  assign n31998 = ( ~n31978 & n31996 ) | ( ~n31978 & n31997 ) | ( n31996 & n31997 ) ;
  assign n31999 = ~n31861 & n31998 ;
  assign n32000 = x110 & n9933 ;
  assign n32001 = x109 & n9928 ;
  assign n32002 = x108 & ~n9927 ;
  assign n32003 = n10379 & n32002 ;
  assign n32004 = n32001 | n32003 ;
  assign n32005 = n32000 | n32004 ;
  assign n32006 = n9936 | n32000 ;
  assign n32007 = n32004 | n32006 ;
  assign n32008 = ( n10330 & n32005 ) | ( n10330 & n32007 ) | ( n32005 & n32007 ) ;
  assign n32009 = x47 & n32007 ;
  assign n32010 = x47 & n32000 ;
  assign n32011 = ( x47 & n32004 ) | ( x47 & n32010 ) | ( n32004 & n32010 ) ;
  assign n32012 = ( n10330 & n32009 ) | ( n10330 & n32011 ) | ( n32009 & n32011 ) ;
  assign n32013 = x47 & ~n32011 ;
  assign n32014 = x47 & ~n32007 ;
  assign n32015 = ( ~n10330 & n32013 ) | ( ~n10330 & n32014 ) | ( n32013 & n32014 ) ;
  assign n32016 = ( n32008 & ~n32012 ) | ( n32008 & n32015 ) | ( ~n32012 & n32015 ) ;
  assign n32017 = n31648 | n32016 ;
  assign n32018 = n31645 | n32016 ;
  assign n32019 = ( ~n31628 & n32017 ) | ( ~n31628 & n32018 ) | ( n32017 & n32018 ) ;
  assign n32020 = ( ~n31998 & n32016 ) | ( ~n31998 & n32019 ) | ( n32016 & n32019 ) ;
  assign n32021 = n31999 | n32020 ;
  assign n32022 = n31861 & ~n31998 ;
  assign n32023 = n31999 | n32022 ;
  assign n32024 = n32016 & n32023 ;
  assign n32025 = n31673 & n32024 ;
  assign n32026 = ( n31680 & n32024 ) | ( n31680 & n32025 ) | ( n32024 & n32025 ) ;
  assign n32027 = ( n31860 & ~n32021 ) | ( n31860 & n32026 ) | ( ~n32021 & n32026 ) ;
  assign n32028 = n31673 | n32024 ;
  assign n32029 = n31680 | n32028 ;
  assign n32030 = n32021 & ~n32029 ;
  assign n32031 = n32027 | n32030 ;
  assign n32032 = x113 & n8724 ;
  assign n32033 = x112 & n8719 ;
  assign n32034 = x111 & ~n8718 ;
  assign n32035 = n9149 & n32034 ;
  assign n32036 = n32033 | n32035 ;
  assign n32037 = n32032 | n32036 ;
  assign n32038 = n8727 | n32032 ;
  assign n32039 = n32036 | n32038 ;
  assign n32040 = ( ~n11642 & n32037 ) | ( ~n11642 & n32039 ) | ( n32037 & n32039 ) ;
  assign n32041 = n32037 & n32039 ;
  assign n32042 = ( n11626 & n32040 ) | ( n11626 & n32041 ) | ( n32040 & n32041 ) ;
  assign n32043 = x44 & n32042 ;
  assign n32044 = x44 & ~n32042 ;
  assign n32045 = ( n32042 & ~n32043 ) | ( n32042 & n32044 ) | ( ~n32043 & n32044 ) ;
  assign n32046 = n32031 | n32045 ;
  assign n32047 = n32031 & ~n32045 ;
  assign n32048 = ( ~n32031 & n32046 ) | ( ~n32031 & n32047 ) | ( n32046 & n32047 ) ;
  assign n32049 = n31699 | n31704 ;
  assign n32050 = ( n31699 & ~n31702 ) | ( n31699 & n32049 ) | ( ~n31702 & n32049 ) ;
  assign n32051 = n32048 & ~n32050 ;
  assign n32052 = ~n32048 & n32050 ;
  assign n32053 = n32051 | n32052 ;
  assign n32054 = x116 & n7566 ;
  assign n32055 = x115 & n7561 ;
  assign n32056 = x114 & ~n7560 ;
  assign n32057 = n7953 & n32056 ;
  assign n32058 = n32055 | n32057 ;
  assign n32059 = n32054 | n32058 ;
  assign n32060 = n7569 | n32054 ;
  assign n32061 = n32058 | n32060 ;
  assign n32062 = ( ~n13040 & n32059 ) | ( ~n13040 & n32061 ) | ( n32059 & n32061 ) ;
  assign n32063 = n32059 & n32061 ;
  assign n32064 = ( n13022 & n32062 ) | ( n13022 & n32063 ) | ( n32062 & n32063 ) ;
  assign n32065 = x41 & n32064 ;
  assign n32066 = x41 & ~n32064 ;
  assign n32067 = ( n32064 & ~n32065 ) | ( n32064 & n32066 ) | ( ~n32065 & n32066 ) ;
  assign n32068 = n32053 & n32067 ;
  assign n32069 = n32052 | n32067 ;
  assign n32070 = n32051 | n32069 ;
  assign n32071 = ~n32068 & n32070 ;
  assign n32072 = n31722 | n31726 ;
  assign n32073 = ( n31722 & ~n31724 ) | ( n31722 & n32072 ) | ( ~n31724 & n32072 ) ;
  assign n32074 = n32071 & n32073 ;
  assign n32075 = n32071 | n32073 ;
  assign n32076 = ~n32074 & n32075 ;
  assign n32077 = x119 & n6536 ;
  assign n32078 = x118 & n6531 ;
  assign n32079 = x117 & ~n6530 ;
  assign n32080 = n6871 & n32079 ;
  assign n32081 = n32078 | n32080 ;
  assign n32082 = n32077 | n32081 ;
  assign n32083 = n6539 | n32077 ;
  assign n32084 = n32081 | n32083 ;
  assign n32085 = ( n14496 & n32082 ) | ( n14496 & n32084 ) | ( n32082 & n32084 ) ;
  assign n32086 = x38 & n32084 ;
  assign n32087 = x38 & n32077 ;
  assign n32088 = ( x38 & n32081 ) | ( x38 & n32087 ) | ( n32081 & n32087 ) ;
  assign n32089 = ( n14496 & n32086 ) | ( n14496 & n32088 ) | ( n32086 & n32088 ) ;
  assign n32090 = x38 & ~n32088 ;
  assign n32091 = x38 & ~n32084 ;
  assign n32092 = ( ~n14496 & n32090 ) | ( ~n14496 & n32091 ) | ( n32090 & n32091 ) ;
  assign n32093 = ( n32085 & ~n32089 ) | ( n32085 & n32092 ) | ( ~n32089 & n32092 ) ;
  assign n32094 = ~n32076 & n32093 ;
  assign n32095 = n32076 & ~n32093 ;
  assign n32096 = n32094 | n32095 ;
  assign n32097 = n31859 & ~n32096 ;
  assign n32098 = ~n31859 & n32096 ;
  assign n32099 = n32097 | n32098 ;
  assign n32100 = x122 & n5554 ;
  assign n32101 = x121 & n5549 ;
  assign n32102 = x120 & ~n5548 ;
  assign n32103 = n5893 & n32102 ;
  assign n32104 = n32101 | n32103 ;
  assign n32105 = n32100 | n32104 ;
  assign n32106 = n5557 | n32100 ;
  assign n32107 = n32104 | n32106 ;
  assign n32108 = ( n16043 & n32105 ) | ( n16043 & n32107 ) | ( n32105 & n32107 ) ;
  assign n32109 = x35 & n32107 ;
  assign n32110 = x35 & n32100 ;
  assign n32111 = ( x35 & n32104 ) | ( x35 & n32110 ) | ( n32104 & n32110 ) ;
  assign n32112 = ( n16043 & n32109 ) | ( n16043 & n32111 ) | ( n32109 & n32111 ) ;
  assign n32113 = x35 & ~n32111 ;
  assign n32114 = x35 & ~n32107 ;
  assign n32115 = ( ~n16043 & n32113 ) | ( ~n16043 & n32114 ) | ( n32113 & n32114 ) ;
  assign n32116 = ( n32108 & ~n32112 ) | ( n32108 & n32115 ) | ( ~n32112 & n32115 ) ;
  assign n32117 = n32099 | n32116 ;
  assign n32118 = n32099 & ~n32116 ;
  assign n32119 = ( ~n32099 & n32117 ) | ( ~n32099 & n32118 ) | ( n32117 & n32118 ) ;
  assign n32120 = n31858 & ~n32119 ;
  assign n32121 = ~n31858 & n32119 ;
  assign n32122 = n32120 | n32121 ;
  assign n32123 = ( ~n31779 & n31796 ) | ( ~n31779 & n31797 ) | ( n31796 & n31797 ) ;
  assign n32124 = x127 & n3811 ;
  assign n32125 = x126 & ~n3810 ;
  assign n32126 = n4067 & n32125 ;
  assign n32127 = n32124 | n32126 ;
  assign n32128 = n3819 | n32127 ;
  assign n32129 = ( n19328 & n32127 ) | ( n19328 & n32128 ) | ( n32127 & n32128 ) ;
  assign n32130 = x29 & n32127 ;
  assign n32131 = ( x29 & n5940 ) | ( x29 & n32127 ) | ( n5940 & n32127 ) ;
  assign n32132 = ( n19328 & n32130 ) | ( n19328 & n32131 ) | ( n32130 & n32131 ) ;
  assign n32133 = x29 & ~n5940 ;
  assign n32134 = ~n32127 & n32133 ;
  assign n32135 = x29 & ~n32127 ;
  assign n32136 = ( ~n19328 & n32134 ) | ( ~n19328 & n32135 ) | ( n32134 & n32135 ) ;
  assign n32137 = ( n32129 & ~n32132 ) | ( n32129 & n32136 ) | ( ~n32132 & n32136 ) ;
  assign n32138 = n32123 | n32137 ;
  assign n32139 = n32123 & n32137 ;
  assign n32140 = n32138 & ~n32139 ;
  assign n32141 = n32122 | n32140 ;
  assign n32142 = ~n32140 & n32141 ;
  assign n32143 = ( ~n32122 & n32141 ) | ( ~n32122 & n32142 ) | ( n32141 & n32142 ) ;
  assign n32144 = ~n31830 & n32143 ;
  assign n32145 = n31830 & ~n32143 ;
  assign n32146 = n32144 | n32145 ;
  assign n32147 = n31814 & ~n31817 ;
  assign n32148 = ( n31814 & ~n31820 ) | ( n31814 & n32147 ) | ( ~n31820 & n32147 ) ;
  assign n32149 = n31814 & ~n31826 ;
  assign n32150 = ( ~n31467 & n31814 ) | ( ~n31467 & n32147 ) | ( n31814 & n32147 ) ;
  assign n32151 = ( ~n31472 & n32149 ) | ( ~n31472 & n32150 ) | ( n32149 & n32150 ) ;
  assign n32152 = ( ~n30754 & n32148 ) | ( ~n30754 & n32151 ) | ( n32148 & n32151 ) ;
  assign n32153 = n32146 & n32152 ;
  assign n32154 = n32146 | n32151 ;
  assign n32155 = n31814 | n32146 ;
  assign n32156 = ( ~n31817 & n32146 ) | ( ~n31817 & n32155 ) | ( n32146 & n32155 ) ;
  assign n32157 = ( ~n31820 & n32155 ) | ( ~n31820 & n32156 ) | ( n32155 & n32156 ) ;
  assign n32158 = ( ~n30754 & n32154 ) | ( ~n30754 & n32157 ) | ( n32154 & n32157 ) ;
  assign n32159 = ~n32153 & n32158 ;
  assign n32160 = ~n32145 & n32156 ;
  assign n32161 = ~n32145 & n32155 ;
  assign n32162 = ( ~n31820 & n32160 ) | ( ~n31820 & n32161 ) | ( n32160 & n32161 ) ;
  assign n32163 = ~n32145 & n32146 ;
  assign n32164 = ( ~n32145 & n32151 ) | ( ~n32145 & n32163 ) | ( n32151 & n32163 ) ;
  assign n32165 = ( ~n30754 & n32162 ) | ( ~n30754 & n32164 ) | ( n32162 & n32164 ) ;
  assign n32166 = x126 & n4631 ;
  assign n32167 = x125 & n4626 ;
  assign n32168 = x124 & ~n4625 ;
  assign n32169 = n4943 & n32168 ;
  assign n32170 = n32167 | n32169 ;
  assign n32171 = n32166 | n32170 ;
  assign n32172 = n4634 | n32166 ;
  assign n32173 = n32170 | n32172 ;
  assign n32174 = ( n18220 & n32171 ) | ( n18220 & n32173 ) | ( n32171 & n32173 ) ;
  assign n32175 = x32 & n32173 ;
  assign n32176 = x32 & n32166 ;
  assign n32177 = ( x32 & n32170 ) | ( x32 & n32176 ) | ( n32170 & n32176 ) ;
  assign n32178 = ( n18220 & n32175 ) | ( n18220 & n32177 ) | ( n32175 & n32177 ) ;
  assign n32179 = x32 & ~n32177 ;
  assign n32180 = x32 & ~n32173 ;
  assign n32181 = ( ~n18220 & n32179 ) | ( ~n18220 & n32180 ) | ( n32179 & n32180 ) ;
  assign n32182 = ( n32174 & ~n32178 ) | ( n32174 & n32181 ) | ( ~n32178 & n32181 ) ;
  assign n32183 = n32096 & ~n32116 ;
  assign n32184 = ( n31859 & n32116 ) | ( n31859 & ~n32183 ) | ( n32116 & ~n32183 ) ;
  assign n32185 = n32182 | n32184 ;
  assign n32186 = n32097 | n32182 ;
  assign n32187 = ( ~n32099 & n32185 ) | ( ~n32099 & n32186 ) | ( n32185 & n32186 ) ;
  assign n32188 = n32182 & n32184 ;
  assign n32189 = n32097 & n32182 ;
  assign n32190 = ( ~n32099 & n32188 ) | ( ~n32099 & n32189 ) | ( n32188 & n32189 ) ;
  assign n32191 = n32187 & ~n32190 ;
  assign n32274 = n31878 & ~n31943 ;
  assign n32275 = ( n31878 & ~n31945 ) | ( n31878 & n32274 ) | ( ~n31945 & n32274 ) ;
  assign n32276 = ~n31943 & n31945 ;
  assign n32277 = n31943 | n31945 ;
  assign n32278 = ( n31878 & n32276 ) | ( n31878 & ~n32277 ) | ( n32276 & ~n32277 ) ;
  assign n32279 = n31878 | n32276 ;
  assign n32280 = ( ~n32275 & n32278 ) | ( ~n32275 & n32279 ) | ( n32278 & n32279 ) ;
  assign n32192 = n31886 | n31907 ;
  assign n32193 = x93 & n18290 ;
  assign n32194 = x63 & x92 ;
  assign n32195 = ~n18290 & n32194 ;
  assign n32196 = n32193 | n32195 ;
  assign n32197 = ~n31882 & n32196 ;
  assign n32198 = n31882 & ~n32196 ;
  assign n32199 = n32197 | n32198 ;
  assign n32200 = n31882 | n32199 ;
  assign n32201 = n31884 & ~n32200 ;
  assign n32202 = ( n31907 & ~n32199 ) | ( n31907 & n32201 ) | ( ~n32199 & n32201 ) ;
  assign n32203 = n32192 & ~n32202 ;
  assign n32204 = x96 & n17146 ;
  assign n32205 = x95 & n17141 ;
  assign n32206 = x94 & ~n17140 ;
  assign n32207 = n17724 & n32206 ;
  assign n32208 = n32205 | n32207 ;
  assign n32209 = n32204 | n32208 ;
  assign n32210 = n17149 | n32204 ;
  assign n32211 = n32208 | n32210 ;
  assign n32212 = ( n5202 & n32209 ) | ( n5202 & n32211 ) | ( n32209 & n32211 ) ;
  assign n32213 = x62 & n32211 ;
  assign n32214 = x62 & n32204 ;
  assign n32215 = ( x62 & n32208 ) | ( x62 & n32214 ) | ( n32208 & n32214 ) ;
  assign n32216 = ( n5202 & n32213 ) | ( n5202 & n32215 ) | ( n32213 & n32215 ) ;
  assign n32217 = x62 & ~n32215 ;
  assign n32218 = x62 & ~n32211 ;
  assign n32219 = ( ~n5202 & n32217 ) | ( ~n5202 & n32218 ) | ( n32217 & n32218 ) ;
  assign n32220 = ( n32212 & ~n32216 ) | ( n32212 & n32219 ) | ( ~n32216 & n32219 ) ;
  assign n32221 = n32199 | n32201 ;
  assign n32222 = n31907 | n32221 ;
  assign n32223 = n32220 | n32222 ;
  assign n32224 = ( ~n32203 & n32220 ) | ( ~n32203 & n32223 ) | ( n32220 & n32223 ) ;
  assign n32225 = n32220 & n32222 ;
  assign n32226 = ~n32203 & n32225 ;
  assign n32227 = n32224 & ~n32226 ;
  assign n32228 = x99 & n15552 ;
  assign n32229 = x98 & n15547 ;
  assign n32230 = x97 & ~n15546 ;
  assign n32231 = n16123 & n32230 ;
  assign n32232 = n32229 | n32231 ;
  assign n32233 = n32228 | n32232 ;
  assign n32234 = n15555 | n32228 ;
  assign n32235 = n32232 | n32234 ;
  assign n32236 = ( n6164 & n32233 ) | ( n6164 & n32235 ) | ( n32233 & n32235 ) ;
  assign n32237 = x59 & n32235 ;
  assign n32238 = x59 & n32228 ;
  assign n32239 = ( x59 & n32232 ) | ( x59 & n32238 ) | ( n32232 & n32238 ) ;
  assign n32240 = ( n6164 & n32237 ) | ( n6164 & n32239 ) | ( n32237 & n32239 ) ;
  assign n32241 = x59 & ~n32239 ;
  assign n32242 = x59 & ~n32235 ;
  assign n32243 = ( ~n6164 & n32241 ) | ( ~n6164 & n32242 ) | ( n32241 & n32242 ) ;
  assign n32244 = ( n32236 & ~n32240 ) | ( n32236 & n32243 ) | ( ~n32240 & n32243 ) ;
  assign n32245 = ~n32227 & n32244 ;
  assign n32246 = n32227 & ~n32244 ;
  assign n32247 = n32245 | n32246 ;
  assign n32248 = n31912 & ~n31940 ;
  assign n32249 = ( n31914 & n31940 ) | ( n31914 & ~n32248 ) | ( n31940 & ~n32248 ) ;
  assign n32250 = ( n31915 & ~n31917 ) | ( n31915 & n32249 ) | ( ~n31917 & n32249 ) ;
  assign n32251 = ~n32247 & n32250 ;
  assign n32252 = n32247 & ~n32250 ;
  assign n32253 = n32251 | n32252 ;
  assign n32254 = x102 & n14045 ;
  assign n32255 = x101 & n14040 ;
  assign n32256 = x100 & ~n14039 ;
  assign n32257 = n14552 & n32256 ;
  assign n32258 = n32255 | n32257 ;
  assign n32259 = n32254 | n32258 ;
  assign n32260 = n14048 | n32254 ;
  assign n32261 = n32258 | n32260 ;
  assign n32262 = ( n7178 & n32259 ) | ( n7178 & n32261 ) | ( n32259 & n32261 ) ;
  assign n32263 = x56 & n32261 ;
  assign n32264 = x56 & n32254 ;
  assign n32265 = ( x56 & n32258 ) | ( x56 & n32264 ) | ( n32258 & n32264 ) ;
  assign n32266 = ( n7178 & n32263 ) | ( n7178 & n32265 ) | ( n32263 & n32265 ) ;
  assign n32267 = x56 & ~n32265 ;
  assign n32268 = x56 & ~n32261 ;
  assign n32269 = ( ~n7178 & n32267 ) | ( ~n7178 & n32268 ) | ( n32267 & n32268 ) ;
  assign n32270 = ( n32262 & ~n32266 ) | ( n32262 & n32269 ) | ( ~n32266 & n32269 ) ;
  assign n32271 = n32253 | n32270 ;
  assign n32272 = n32253 & ~n32270 ;
  assign n32273 = ( ~n32253 & n32271 ) | ( ~n32253 & n32272 ) | ( n32271 & n32272 ) ;
  assign n32281 = ~n32273 & n32280 ;
  assign n32282 = n32280 & ~n32281 ;
  assign n32283 = x105 & n12574 ;
  assign n32284 = x104 & n12569 ;
  assign n32285 = x103 & ~n12568 ;
  assign n32286 = n13076 & n32285 ;
  assign n32287 = n32284 | n32286 ;
  assign n32288 = n32283 | n32287 ;
  assign n32289 = n12577 | n32283 ;
  assign n32290 = n32287 | n32289 ;
  assign n32291 = ( n8273 & n32288 ) | ( n8273 & n32290 ) | ( n32288 & n32290 ) ;
  assign n32292 = x53 & n32290 ;
  assign n32293 = x53 & n32283 ;
  assign n32294 = ( x53 & n32287 ) | ( x53 & n32293 ) | ( n32287 & n32293 ) ;
  assign n32295 = ( n8273 & n32292 ) | ( n8273 & n32294 ) | ( n32292 & n32294 ) ;
  assign n32296 = x53 & ~n32294 ;
  assign n32297 = x53 & ~n32290 ;
  assign n32298 = ( ~n8273 & n32296 ) | ( ~n8273 & n32297 ) | ( n32296 & n32297 ) ;
  assign n32299 = ( n32291 & ~n32295 ) | ( n32291 & n32298 ) | ( ~n32295 & n32298 ) ;
  assign n32300 = n32273 | n32280 ;
  assign n32301 = n32299 | n32300 ;
  assign n32302 = ( ~n32282 & n32299 ) | ( ~n32282 & n32301 ) | ( n32299 & n32301 ) ;
  assign n32303 = n32299 & n32300 ;
  assign n32304 = ~n32282 & n32303 ;
  assign n32305 = n32302 & ~n32304 ;
  assign n32306 = n31592 & ~n31948 ;
  assign n32307 = ( n31598 & ~n31948 ) | ( n31598 & n32306 ) | ( ~n31948 & n32306 ) ;
  assign n32308 = n31949 & ~n32307 ;
  assign n32309 = n31948 | n32307 ;
  assign n32310 = ~n32308 & n32309 ;
  assign n32311 = n31966 | n32307 ;
  assign n32312 = ( n32307 & ~n32310 ) | ( n32307 & n32311 ) | ( ~n32310 & n32311 ) ;
  assign n32313 = ~n32305 & n32312 ;
  assign n32314 = n32305 & ~n32312 ;
  assign n32315 = n32313 | n32314 ;
  assign n32316 = x108 & n11205 ;
  assign n32317 = x107 & n11200 ;
  assign n32318 = x106 & ~n11199 ;
  assign n32319 = n11679 & n32318 ;
  assign n32320 = n32317 | n32319 ;
  assign n32321 = n32316 | n32320 ;
  assign n32322 = n11208 | n32316 ;
  assign n32323 = n32320 | n32322 ;
  assign n32324 = ( n9479 & n32321 ) | ( n9479 & n32323 ) | ( n32321 & n32323 ) ;
  assign n32325 = x50 & n32323 ;
  assign n32326 = x50 & n32316 ;
  assign n32327 = ( x50 & n32320 ) | ( x50 & n32326 ) | ( n32320 & n32326 ) ;
  assign n32328 = ( n9479 & n32325 ) | ( n9479 & n32327 ) | ( n32325 & n32327 ) ;
  assign n32329 = x50 & ~n32327 ;
  assign n32330 = x50 & ~n32323 ;
  assign n32331 = ( ~n9479 & n32329 ) | ( ~n9479 & n32330 ) | ( n32329 & n32330 ) ;
  assign n32332 = ( n32324 & ~n32328 ) | ( n32324 & n32331 ) | ( ~n32328 & n32331 ) ;
  assign n32333 = ~n32315 & n32332 ;
  assign n32334 = n32315 & ~n32332 ;
  assign n32335 = n32333 | n32334 ;
  assign n32336 = n31975 | n31995 ;
  assign n32337 = ( n31975 & ~n31978 ) | ( n31975 & n32336 ) | ( ~n31978 & n32336 ) ;
  assign n32338 = ~n32335 & n32337 ;
  assign n32339 = n32335 & ~n32337 ;
  assign n32340 = n32338 | n32339 ;
  assign n32341 = x111 & n9933 ;
  assign n32342 = x110 & n9928 ;
  assign n32343 = x109 & ~n9927 ;
  assign n32344 = n10379 & n32343 ;
  assign n32345 = n32342 | n32344 ;
  assign n32346 = n32341 | n32345 ;
  assign n32347 = n9936 | n32341 ;
  assign n32348 = n32345 | n32347 ;
  assign n32349 = ( n10749 & n32346 ) | ( n10749 & n32348 ) | ( n32346 & n32348 ) ;
  assign n32350 = x47 & n32348 ;
  assign n32351 = x47 & n32341 ;
  assign n32352 = ( x47 & n32345 ) | ( x47 & n32351 ) | ( n32345 & n32351 ) ;
  assign n32353 = ( n10749 & n32350 ) | ( n10749 & n32352 ) | ( n32350 & n32352 ) ;
  assign n32354 = x47 & ~n32352 ;
  assign n32355 = x47 & ~n32348 ;
  assign n32356 = ( ~n10749 & n32354 ) | ( ~n10749 & n32355 ) | ( n32354 & n32355 ) ;
  assign n32357 = ( n32349 & ~n32353 ) | ( n32349 & n32356 ) | ( ~n32353 & n32356 ) ;
  assign n32358 = n32340 | n32357 ;
  assign n32359 = n32340 & ~n32357 ;
  assign n32360 = ( ~n32340 & n32358 ) | ( ~n32340 & n32359 ) | ( n32358 & n32359 ) ;
  assign n32361 = ( n32020 & n32022 ) | ( n32020 & ~n32023 ) | ( n32022 & ~n32023 ) ;
  assign n32362 = n32360 & ~n32361 ;
  assign n32363 = ~n32360 & n32361 ;
  assign n32364 = n32362 | n32363 ;
  assign n32365 = x114 & n8724 ;
  assign n32366 = x113 & n8719 ;
  assign n32367 = x112 & ~n8718 ;
  assign n32368 = n9149 & n32367 ;
  assign n32369 = n32366 | n32368 ;
  assign n32370 = n32365 | n32369 ;
  assign n32371 = n8727 | n32365 ;
  assign n32372 = n32369 | n32371 ;
  assign n32373 = ( ~n12095 & n32370 ) | ( ~n12095 & n32372 ) | ( n32370 & n32372 ) ;
  assign n32374 = n32370 & n32372 ;
  assign n32375 = ( n12079 & n32373 ) | ( n12079 & n32374 ) | ( n32373 & n32374 ) ;
  assign n32376 = x44 & n32375 ;
  assign n32377 = x44 & ~n32375 ;
  assign n32378 = ( n32375 & ~n32376 ) | ( n32375 & n32377 ) | ( ~n32376 & n32377 ) ;
  assign n32379 = n32364 & ~n32378 ;
  assign n32380 = ~n32364 & n32378 ;
  assign n32381 = n32379 | n32380 ;
  assign n32382 = n32027 | n32045 ;
  assign n32383 = ( n32027 & ~n32031 ) | ( n32027 & n32382 ) | ( ~n32031 & n32382 ) ;
  assign n32384 = n32381 & n32383 ;
  assign n32385 = ~n32381 & n32383 ;
  assign n32386 = x117 & n7566 ;
  assign n32387 = x116 & n7561 ;
  assign n32388 = x115 & ~n7560 ;
  assign n32389 = n7953 & n32388 ;
  assign n32390 = n32387 | n32389 ;
  assign n32391 = n32386 | n32390 ;
  assign n32392 = n7569 | n32386 ;
  assign n32393 = n32390 | n32392 ;
  assign n32394 = ( ~n13522 & n32391 ) | ( ~n13522 & n32393 ) | ( n32391 & n32393 ) ;
  assign n32395 = n32391 & n32393 ;
  assign n32396 = ( n13503 & n32394 ) | ( n13503 & n32395 ) | ( n32394 & n32395 ) ;
  assign n32397 = x41 & n32396 ;
  assign n32398 = x41 & ~n32396 ;
  assign n32399 = ( n32396 & ~n32397 ) | ( n32396 & n32398 ) | ( ~n32397 & n32398 ) ;
  assign n32400 = n32381 & ~n32399 ;
  assign n32401 = ( n32385 & ~n32399 ) | ( n32385 & n32400 ) | ( ~n32399 & n32400 ) ;
  assign n32402 = ~n32384 & n32401 ;
  assign n32403 = n32381 | n32385 ;
  assign n32404 = n32384 & n32399 ;
  assign n32405 = ( n32399 & ~n32403 ) | ( n32399 & n32404 ) | ( ~n32403 & n32404 ) ;
  assign n32406 = n32402 | n32405 ;
  assign n32407 = ( n32052 & ~n32053 ) | ( n32052 & n32069 ) | ( ~n32053 & n32069 ) ;
  assign n32408 = ~n32406 & n32407 ;
  assign n32409 = n32406 & ~n32407 ;
  assign n32410 = n32408 | n32409 ;
  assign n32411 = x120 & n6536 ;
  assign n32412 = x119 & n6531 ;
  assign n32413 = x118 & ~n6530 ;
  assign n32414 = n6871 & n32413 ;
  assign n32415 = n32412 | n32414 ;
  assign n32416 = n32411 | n32415 ;
  assign n32417 = n6539 | n32411 ;
  assign n32418 = n32415 | n32417 ;
  assign n32419 = ( n14991 & n32416 ) | ( n14991 & n32418 ) | ( n32416 & n32418 ) ;
  assign n32420 = x38 & n32418 ;
  assign n32421 = x38 & n32411 ;
  assign n32422 = ( x38 & n32415 ) | ( x38 & n32421 ) | ( n32415 & n32421 ) ;
  assign n32423 = ( n14991 & n32420 ) | ( n14991 & n32422 ) | ( n32420 & n32422 ) ;
  assign n32424 = x38 & ~n32422 ;
  assign n32425 = x38 & ~n32418 ;
  assign n32426 = ( ~n14991 & n32424 ) | ( ~n14991 & n32425 ) | ( n32424 & n32425 ) ;
  assign n32427 = ( n32419 & ~n32423 ) | ( n32419 & n32426 ) | ( ~n32423 & n32426 ) ;
  assign n32428 = ~n32410 & n32427 ;
  assign n32429 = n32410 & ~n32427 ;
  assign n32430 = n32428 | n32429 ;
  assign n32431 = ( ~n32071 & n32073 ) | ( ~n32071 & n32093 ) | ( n32073 & n32093 ) ;
  assign n32432 = ~n32430 & n32431 ;
  assign n32433 = n32430 & ~n32431 ;
  assign n32434 = n32432 | n32433 ;
  assign n32435 = x123 & n5554 ;
  assign n32436 = x122 & n5549 ;
  assign n32437 = x121 & ~n5548 ;
  assign n32438 = n5893 & n32437 ;
  assign n32439 = n32436 | n32438 ;
  assign n32440 = n32435 | n32439 ;
  assign n32441 = n5557 | n32435 ;
  assign n32442 = n32439 | n32441 ;
  assign n32443 = ( n16086 & n32440 ) | ( n16086 & n32442 ) | ( n32440 & n32442 ) ;
  assign n32444 = x35 & n32442 ;
  assign n32445 = x35 & n32435 ;
  assign n32446 = ( x35 & n32439 ) | ( x35 & n32445 ) | ( n32439 & n32445 ) ;
  assign n32447 = ( n16086 & n32444 ) | ( n16086 & n32446 ) | ( n32444 & n32446 ) ;
  assign n32448 = x35 & ~n32446 ;
  assign n32449 = x35 & ~n32442 ;
  assign n32450 = ( ~n16086 & n32448 ) | ( ~n16086 & n32449 ) | ( n32448 & n32449 ) ;
  assign n32451 = ( n32443 & ~n32447 ) | ( n32443 & n32450 ) | ( ~n32447 & n32450 ) ;
  assign n32452 = n32434 | n32451 ;
  assign n32453 = n32434 & ~n32451 ;
  assign n32454 = ( ~n32434 & n32452 ) | ( ~n32434 & n32453 ) | ( n32452 & n32453 ) ;
  assign n32455 = ~n32191 & n32454 ;
  assign n32456 = n32191 & ~n32454 ;
  assign n32457 = n32455 | n32456 ;
  assign n32458 = x127 & ~n3810 ;
  assign n32459 = n4067 & n32458 ;
  assign n32460 = n3819 & n19877 ;
  assign n32461 = n32459 | n32460 ;
  assign n32462 = n3819 & n19880 ;
  assign n32463 = n32459 | n32462 ;
  assign n32464 = ( n18202 & n32461 ) | ( n18202 & n32463 ) | ( n32461 & n32463 ) ;
  assign n32465 = n32461 & n32463 ;
  assign n32466 = ( n18212 & n32464 ) | ( n18212 & n32465 ) | ( n32464 & n32465 ) ;
  assign n32467 = ( n18214 & n32464 ) | ( n18214 & n32465 ) | ( n32464 & n32465 ) ;
  assign n32468 = ( n14002 & n32466 ) | ( n14002 & n32467 ) | ( n32466 & n32467 ) ;
  assign n32469 = x29 & n32466 ;
  assign n32470 = x29 & n32467 ;
  assign n32471 = ( n14002 & n32469 ) | ( n14002 & n32470 ) | ( n32469 & n32470 ) ;
  assign n32472 = x29 & ~n32470 ;
  assign n32473 = x29 & ~n32469 ;
  assign n32474 = ( ~n14002 & n32472 ) | ( ~n14002 & n32473 ) | ( n32472 & n32473 ) ;
  assign n32475 = ( n32468 & ~n32471 ) | ( n32468 & n32474 ) | ( ~n32471 & n32474 ) ;
  assign n32476 = n31848 & n32475 ;
  assign n32477 = n32475 & ~n32476 ;
  assign n32478 = ( n31752 & n32475 ) | ( n31752 & n32477 ) | ( n32475 & n32477 ) ;
  assign n32479 = ~n31847 & n32475 ;
  assign n32480 = ( ~n31774 & n32478 ) | ( ~n31774 & n32479 ) | ( n32478 & n32479 ) ;
  assign n32481 = ( n31771 & n32478 ) | ( n31771 & n32479 ) | ( n32478 & n32479 ) ;
  assign n32482 = ( ~n31775 & n32480 ) | ( ~n31775 & n32481 ) | ( n32480 & n32481 ) ;
  assign n32483 = n32119 & n32482 ;
  assign n32484 = ( ~n31858 & n32482 ) | ( ~n31858 & n32483 ) | ( n32482 & n32483 ) ;
  assign n32485 = ~n32457 & n32484 ;
  assign n32486 = n31847 & n32475 ;
  assign n32487 = ~n31752 & n32476 ;
  assign n32488 = ( n31774 & n32486 ) | ( n31774 & n32487 ) | ( n32486 & n32487 ) ;
  assign n32489 = ( ~n31771 & n32486 ) | ( ~n31771 & n32487 ) | ( n32486 & n32487 ) ;
  assign n32490 = ( n31775 & n32488 ) | ( n31775 & n32489 ) | ( n32488 & n32489 ) ;
  assign n32491 = ( ~n32119 & n32475 ) | ( ~n32119 & n32490 ) | ( n32475 & n32490 ) ;
  assign n32492 = n32475 & n32490 ;
  assign n32493 = ( n31858 & n32491 ) | ( n31858 & n32492 ) | ( n32491 & n32492 ) ;
  assign n32494 = ( n31852 & n32120 ) | ( n31852 & ~n32493 ) | ( n32120 & ~n32493 ) ;
  assign n32495 = ( ~n32457 & n32485 ) | ( ~n32457 & n32494 ) | ( n32485 & n32494 ) ;
  assign n32496 = n32457 & ~n32484 ;
  assign n32497 = ~n32494 & n32496 ;
  assign n32498 = n32495 | n32497 ;
  assign n32499 = n32122 & ~n32139 ;
  assign n32500 = ( n32139 & n32140 ) | ( n32139 & ~n32499 ) | ( n32140 & ~n32499 ) ;
  assign n32501 = n32498 | n32500 ;
  assign n32502 = n32165 & n32501 ;
  assign n32503 = n32498 & n32500 ;
  assign n32504 = n32502 & ~n32503 ;
  assign n32505 = n32501 & ~n32503 ;
  assign n32506 = n32143 | n32505 ;
  assign n32507 = n31830 & ~n32506 ;
  assign n32508 = ( n32156 & n32505 ) | ( n32156 & ~n32507 ) | ( n32505 & ~n32507 ) ;
  assign n32509 = ( n32155 & n32505 ) | ( n32155 & ~n32507 ) | ( n32505 & ~n32507 ) ;
  assign n32510 = ( ~n31820 & n32508 ) | ( ~n31820 & n32509 ) | ( n32508 & n32509 ) ;
  assign n32511 = ( n32146 & n32505 ) | ( n32146 & ~n32507 ) | ( n32505 & ~n32507 ) ;
  assign n32512 = ( n32151 & ~n32507 ) | ( n32151 & n32511 ) | ( ~n32507 & n32511 ) ;
  assign n32513 = ( ~n30754 & n32510 ) | ( ~n30754 & n32512 ) | ( n32510 & n32512 ) ;
  assign n32514 = ~n32504 & n32513 ;
  assign n32515 = n32385 | n32405 ;
  assign n32516 = x97 & n17146 ;
  assign n32517 = x96 & n17141 ;
  assign n32518 = x95 & ~n17140 ;
  assign n32519 = n17724 & n32518 ;
  assign n32520 = n32517 | n32519 ;
  assign n32521 = n32516 | n32520 ;
  assign n32522 = n17149 | n32516 ;
  assign n32523 = n32520 | n32522 ;
  assign n32524 = ( n5505 & n32521 ) | ( n5505 & n32523 ) | ( n32521 & n32523 ) ;
  assign n32525 = x62 & n32523 ;
  assign n32526 = x62 & n32516 ;
  assign n32527 = ( x62 & n32520 ) | ( x62 & n32526 ) | ( n32520 & n32526 ) ;
  assign n32528 = ( n5505 & n32525 ) | ( n5505 & n32527 ) | ( n32525 & n32527 ) ;
  assign n32529 = x62 & ~n32527 ;
  assign n32530 = x62 & ~n32523 ;
  assign n32531 = ( ~n5505 & n32529 ) | ( ~n5505 & n32530 ) | ( n32529 & n32530 ) ;
  assign n32532 = ( n32524 & ~n32528 ) | ( n32524 & n32531 ) | ( ~n32528 & n32531 ) ;
  assign n32533 = n32198 | n32201 ;
  assign n32534 = ~n32198 & n32199 ;
  assign n32535 = ( n31907 & n32533 ) | ( n31907 & ~n32534 ) | ( n32533 & ~n32534 ) ;
  assign n32536 = x94 & n18290 ;
  assign n32537 = x63 & x93 ;
  assign n32538 = ~n18290 & n32537 ;
  assign n32539 = n32536 | n32538 ;
  assign n32540 = ~x29 & n32539 ;
  assign n32541 = x29 & ~n32539 ;
  assign n32542 = n32540 | n32541 ;
  assign n32543 = n32196 | n32542 ;
  assign n32544 = ~n32542 & n32543 ;
  assign n32545 = ( ~n32196 & n32543 ) | ( ~n32196 & n32544 ) | ( n32543 & n32544 ) ;
  assign n32546 = n32533 & ~n32545 ;
  assign n32547 = n32534 | n32543 ;
  assign n32548 = n32196 & n32198 ;
  assign n32549 = ( n32196 & ~n32199 ) | ( n32196 & n32548 ) | ( ~n32199 & n32548 ) ;
  assign n32550 = ( n32544 & n32547 ) | ( n32544 & ~n32549 ) | ( n32547 & ~n32549 ) ;
  assign n32551 = ( n31907 & n32546 ) | ( n31907 & ~n32550 ) | ( n32546 & ~n32550 ) ;
  assign n32552 = n32535 & ~n32551 ;
  assign n32553 = n32533 | n32545 ;
  assign n32554 = n32534 & ~n32543 ;
  assign n32555 = n32196 & n32534 ;
  assign n32556 = ( ~n32544 & n32554 ) | ( ~n32544 & n32555 ) | ( n32554 & n32555 ) ;
  assign n32557 = ( n31907 & n32553 ) | ( n31907 & ~n32556 ) | ( n32553 & ~n32556 ) ;
  assign n32558 = n32532 & n32557 ;
  assign n32559 = ~n32552 & n32558 ;
  assign n32560 = n32532 & ~n32559 ;
  assign n32561 = x100 & n15552 ;
  assign n32562 = x99 & n15547 ;
  assign n32563 = x98 & ~n15546 ;
  assign n32564 = n16123 & n32563 ;
  assign n32565 = n32562 | n32564 ;
  assign n32566 = n32561 | n32565 ;
  assign n32567 = n15555 | n32561 ;
  assign n32568 = n32565 | n32567 ;
  assign n32569 = ( n6483 & n32566 ) | ( n6483 & n32568 ) | ( n32566 & n32568 ) ;
  assign n32570 = x59 & n32568 ;
  assign n32571 = x59 & n32561 ;
  assign n32572 = ( x59 & n32565 ) | ( x59 & n32571 ) | ( n32565 & n32571 ) ;
  assign n32573 = ( n6483 & n32570 ) | ( n6483 & n32572 ) | ( n32570 & n32572 ) ;
  assign n32574 = x59 & ~n32572 ;
  assign n32575 = x59 & ~n32568 ;
  assign n32576 = ( ~n6483 & n32574 ) | ( ~n6483 & n32575 ) | ( n32574 & n32575 ) ;
  assign n32577 = ( n32569 & ~n32573 ) | ( n32569 & n32576 ) | ( ~n32573 & n32576 ) ;
  assign n32578 = n32559 & n32577 ;
  assign n32579 = ~n32557 & n32577 ;
  assign n32580 = ( n32552 & n32577 ) | ( n32552 & n32579 ) | ( n32577 & n32579 ) ;
  assign n32581 = ( ~n32560 & n32578 ) | ( ~n32560 & n32580 ) | ( n32578 & n32580 ) ;
  assign n32582 = n32559 | n32577 ;
  assign n32583 = n32557 & ~n32577 ;
  assign n32584 = ~n32552 & n32583 ;
  assign n32585 = ( n32560 & ~n32582 ) | ( n32560 & n32584 ) | ( ~n32582 & n32584 ) ;
  assign n32586 = n32581 | n32585 ;
  assign n32587 = ( n32220 & ~n32222 ) | ( n32220 & n32244 ) | ( ~n32222 & n32244 ) ;
  assign n32588 = n32220 | n32244 ;
  assign n32589 = ( n32203 & n32587 ) | ( n32203 & n32588 ) | ( n32587 & n32588 ) ;
  assign n32590 = ~n32586 & n32589 ;
  assign n32591 = n32586 & ~n32589 ;
  assign n32592 = n32590 | n32591 ;
  assign n32593 = x103 & n14045 ;
  assign n32594 = x102 & n14040 ;
  assign n32595 = x101 & ~n14039 ;
  assign n32596 = n14552 & n32595 ;
  assign n32597 = n32594 | n32596 ;
  assign n32598 = n32593 | n32597 ;
  assign n32599 = n14048 | n32593 ;
  assign n32600 = n32597 | n32599 ;
  assign n32601 = ( n7529 & n32598 ) | ( n7529 & n32600 ) | ( n32598 & n32600 ) ;
  assign n32602 = x56 & n32600 ;
  assign n32603 = x56 & n32593 ;
  assign n32604 = ( x56 & n32597 ) | ( x56 & n32603 ) | ( n32597 & n32603 ) ;
  assign n32605 = ( n7529 & n32602 ) | ( n7529 & n32604 ) | ( n32602 & n32604 ) ;
  assign n32606 = x56 & ~n32604 ;
  assign n32607 = x56 & ~n32600 ;
  assign n32608 = ( ~n7529 & n32606 ) | ( ~n7529 & n32607 ) | ( n32606 & n32607 ) ;
  assign n32609 = ( n32601 & ~n32605 ) | ( n32601 & n32608 ) | ( ~n32605 & n32608 ) ;
  assign n32610 = ~n32592 & n32609 ;
  assign n32611 = n32592 | n32610 ;
  assign n32613 = n32251 | n32270 ;
  assign n32614 = ( n32251 & ~n32253 ) | ( n32251 & n32613 ) | ( ~n32253 & n32613 ) ;
  assign n32612 = n32592 & n32609 ;
  assign n32615 = n32612 & n32614 ;
  assign n32616 = ( ~n32611 & n32614 ) | ( ~n32611 & n32615 ) | ( n32614 & n32615 ) ;
  assign n32617 = n32612 | n32614 ;
  assign n32618 = n32611 & ~n32617 ;
  assign n32619 = n32616 | n32618 ;
  assign n32620 = x106 & n12574 ;
  assign n32621 = x105 & n12569 ;
  assign n32622 = x104 & ~n12568 ;
  assign n32623 = n13076 & n32622 ;
  assign n32624 = n32621 | n32623 ;
  assign n32625 = n32620 | n32624 ;
  assign n32626 = n12577 | n32620 ;
  assign n32627 = n32624 | n32626 ;
  assign n32628 = ( n8656 & n32625 ) | ( n8656 & n32627 ) | ( n32625 & n32627 ) ;
  assign n32629 = x53 & n32627 ;
  assign n32630 = x53 & n32620 ;
  assign n32631 = ( x53 & n32624 ) | ( x53 & n32630 ) | ( n32624 & n32630 ) ;
  assign n32632 = ( n8656 & n32629 ) | ( n8656 & n32631 ) | ( n32629 & n32631 ) ;
  assign n32633 = x53 & ~n32631 ;
  assign n32634 = x53 & ~n32627 ;
  assign n32635 = ( ~n8656 & n32633 ) | ( ~n8656 & n32634 ) | ( n32633 & n32634 ) ;
  assign n32636 = ( n32628 & ~n32632 ) | ( n32628 & n32635 ) | ( ~n32632 & n32635 ) ;
  assign n32637 = ~n32619 & n32636 ;
  assign n32638 = n32619 | n32637 ;
  assign n32639 = ( ~n32273 & n32280 ) | ( ~n32273 & n32299 ) | ( n32280 & n32299 ) ;
  assign n32640 = n32636 & ~n32639 ;
  assign n32641 = n32619 & n32640 ;
  assign n32642 = ( n32638 & n32639 ) | ( n32638 & ~n32641 ) | ( n32639 & ~n32641 ) ;
  assign n32643 = ~n32636 & n32639 ;
  assign n32644 = ( ~n32619 & n32639 ) | ( ~n32619 & n32643 ) | ( n32639 & n32643 ) ;
  assign n32645 = n32638 & n32644 ;
  assign n32646 = n32642 & ~n32645 ;
  assign n32647 = x109 & n11205 ;
  assign n32648 = x108 & n11200 ;
  assign n32649 = x107 & ~n11199 ;
  assign n32650 = n11679 & n32649 ;
  assign n32651 = n32648 | n32650 ;
  assign n32652 = n32647 | n32651 ;
  assign n32653 = n11208 | n32647 ;
  assign n32654 = n32651 | n32653 ;
  assign n32655 = ( n9878 & n32652 ) | ( n9878 & n32654 ) | ( n32652 & n32654 ) ;
  assign n32656 = x50 & n32654 ;
  assign n32657 = x50 & n32647 ;
  assign n32658 = ( x50 & n32651 ) | ( x50 & n32657 ) | ( n32651 & n32657 ) ;
  assign n32659 = ( n9878 & n32656 ) | ( n9878 & n32658 ) | ( n32656 & n32658 ) ;
  assign n32660 = x50 & ~n32658 ;
  assign n32661 = x50 & ~n32654 ;
  assign n32662 = ( ~n9878 & n32660 ) | ( ~n9878 & n32661 ) | ( n32660 & n32661 ) ;
  assign n32663 = ( n32655 & ~n32659 ) | ( n32655 & n32662 ) | ( ~n32659 & n32662 ) ;
  assign n32664 = ~n32646 & n32663 ;
  assign n32665 = n32646 & ~n32663 ;
  assign n32666 = n32664 | n32665 ;
  assign n32667 = n32305 & ~n32332 ;
  assign n32668 = ( n32312 & n32332 ) | ( n32312 & ~n32667 ) | ( n32332 & ~n32667 ) ;
  assign n32669 = ( n32313 & ~n32315 ) | ( n32313 & n32668 ) | ( ~n32315 & n32668 ) ;
  assign n32670 = n32666 & ~n32669 ;
  assign n32671 = ~n32666 & n32669 ;
  assign n32672 = n32670 | n32671 ;
  assign n32673 = x112 & n9933 ;
  assign n32674 = x111 & n9928 ;
  assign n32675 = x110 & ~n9927 ;
  assign n32676 = n10379 & n32675 ;
  assign n32677 = n32674 | n32676 ;
  assign n32678 = n32673 | n32677 ;
  assign n32679 = n9936 | n32673 ;
  assign n32680 = n32677 | n32679 ;
  assign n32681 = ( n11172 & n32678 ) | ( n11172 & n32680 ) | ( n32678 & n32680 ) ;
  assign n32682 = x47 & n32680 ;
  assign n32683 = x47 & n32673 ;
  assign n32684 = ( x47 & n32677 ) | ( x47 & n32683 ) | ( n32677 & n32683 ) ;
  assign n32685 = ( n11172 & n32682 ) | ( n11172 & n32684 ) | ( n32682 & n32684 ) ;
  assign n32686 = x47 & ~n32684 ;
  assign n32687 = x47 & ~n32680 ;
  assign n32688 = ( ~n11172 & n32686 ) | ( ~n11172 & n32687 ) | ( n32686 & n32687 ) ;
  assign n32689 = ( n32681 & ~n32685 ) | ( n32681 & n32688 ) | ( ~n32685 & n32688 ) ;
  assign n32690 = ~n32672 & n32689 ;
  assign n32691 = n32672 | n32690 ;
  assign n32692 = n32672 & n32689 ;
  assign n32693 = n32691 & ~n32692 ;
  assign n32694 = n32337 | n32357 ;
  assign n32695 = ( ~n32335 & n32357 ) | ( ~n32335 & n32694 ) | ( n32357 & n32694 ) ;
  assign n32696 = ( n32338 & ~n32340 ) | ( n32338 & n32695 ) | ( ~n32340 & n32695 ) ;
  assign n32697 = n32693 & ~n32696 ;
  assign n32698 = ~n32693 & n32696 ;
  assign n32699 = n32697 | n32698 ;
  assign n32700 = x115 & n8724 ;
  assign n32701 = x114 & n8719 ;
  assign n32702 = x113 & ~n8718 ;
  assign n32703 = n9149 & n32702 ;
  assign n32704 = n32701 | n32703 ;
  assign n32705 = n32700 | n32704 ;
  assign n32706 = n8727 | n32700 ;
  assign n32707 = n32704 | n32706 ;
  assign n32708 = ( ~n12550 & n32705 ) | ( ~n12550 & n32707 ) | ( n32705 & n32707 ) ;
  assign n32709 = n32705 & n32707 ;
  assign n32710 = ( n12532 & n32708 ) | ( n12532 & n32709 ) | ( n32708 & n32709 ) ;
  assign n32711 = x44 & n32710 ;
  assign n32712 = x44 & ~n32710 ;
  assign n32713 = ( n32710 & ~n32711 ) | ( n32710 & n32712 ) | ( ~n32711 & n32712 ) ;
  assign n32714 = ~n32699 & n32713 ;
  assign n32715 = n32699 & ~n32713 ;
  assign n32716 = n32714 | n32715 ;
  assign n32717 = n32361 | n32378 ;
  assign n32718 = ( ~n32360 & n32378 ) | ( ~n32360 & n32717 ) | ( n32378 & n32717 ) ;
  assign n32719 = ( n32363 & ~n32364 ) | ( n32363 & n32718 ) | ( ~n32364 & n32718 ) ;
  assign n32720 = ~n32716 & n32719 ;
  assign n32721 = n32716 | n32720 ;
  assign n32722 = x118 & n7566 ;
  assign n32723 = x117 & n7561 ;
  assign n32724 = x116 & ~n7560 ;
  assign n32725 = n7953 & n32724 ;
  assign n32726 = n32723 | n32725 ;
  assign n32727 = n32722 | n32726 ;
  assign n32728 = n7569 | n32722 ;
  assign n32729 = n32726 | n32728 ;
  assign n32730 = ( ~n14002 & n32727 ) | ( ~n14002 & n32729 ) | ( n32727 & n32729 ) ;
  assign n32731 = n32727 & n32729 ;
  assign n32732 = ( n13981 & n32730 ) | ( n13981 & n32731 ) | ( n32730 & n32731 ) ;
  assign n32733 = x41 & n32732 ;
  assign n32734 = x41 & ~n32732 ;
  assign n32735 = ( n32732 & ~n32733 ) | ( n32732 & n32734 ) | ( ~n32733 & n32734 ) ;
  assign n32736 = n32719 & n32735 ;
  assign n32737 = n32716 & n32736 ;
  assign n32738 = ( ~n32721 & n32735 ) | ( ~n32721 & n32737 ) | ( n32735 & n32737 ) ;
  assign n32739 = n32719 | n32735 ;
  assign n32740 = ( n32716 & n32735 ) | ( n32716 & n32739 ) | ( n32735 & n32739 ) ;
  assign n32741 = n32721 & ~n32740 ;
  assign n32742 = n32738 | n32741 ;
  assign n32743 = n32515 & ~n32742 ;
  assign n32744 = ~n32515 & n32742 ;
  assign n32745 = n32743 | n32744 ;
  assign n32746 = x121 & n6536 ;
  assign n32747 = x120 & n6531 ;
  assign n32748 = x119 & ~n6530 ;
  assign n32749 = n6871 & n32748 ;
  assign n32750 = n32747 | n32749 ;
  assign n32751 = n32746 | n32750 ;
  assign n32752 = n6539 | n32746 ;
  assign n32753 = n32750 | n32752 ;
  assign n32754 = ( n15501 & n32751 ) | ( n15501 & n32753 ) | ( n32751 & n32753 ) ;
  assign n32755 = x38 & n32753 ;
  assign n32756 = x38 & n32746 ;
  assign n32757 = ( x38 & n32750 ) | ( x38 & n32756 ) | ( n32750 & n32756 ) ;
  assign n32758 = ( n15501 & n32755 ) | ( n15501 & n32757 ) | ( n32755 & n32757 ) ;
  assign n32759 = x38 & ~n32757 ;
  assign n32760 = x38 & ~n32753 ;
  assign n32761 = ( ~n15501 & n32759 ) | ( ~n15501 & n32760 ) | ( n32759 & n32760 ) ;
  assign n32762 = ( n32754 & ~n32758 ) | ( n32754 & n32761 ) | ( ~n32758 & n32761 ) ;
  assign n32763 = ~n32745 & n32762 ;
  assign n32764 = n32745 | n32763 ;
  assign n32766 = n32408 | n32427 ;
  assign n32767 = ( n32408 & ~n32410 ) | ( n32408 & n32766 ) | ( ~n32410 & n32766 ) ;
  assign n32765 = n32745 & n32762 ;
  assign n32768 = n32765 & n32767 ;
  assign n32769 = ( ~n32764 & n32767 ) | ( ~n32764 & n32768 ) | ( n32767 & n32768 ) ;
  assign n32770 = n32765 | n32767 ;
  assign n32771 = n32764 & ~n32770 ;
  assign n32772 = n32769 | n32771 ;
  assign n32773 = x124 & n5554 ;
  assign n32774 = x123 & n5549 ;
  assign n32775 = x122 & ~n5548 ;
  assign n32776 = n5893 & n32775 ;
  assign n32777 = n32774 | n32776 ;
  assign n32778 = n32773 | n32777 ;
  assign n32779 = n5557 | n32773 ;
  assign n32780 = n32777 | n32779 ;
  assign n32781 = ( n17084 & n32778 ) | ( n17084 & n32780 ) | ( n32778 & n32780 ) ;
  assign n32782 = x35 & n32780 ;
  assign n32783 = x35 & n32773 ;
  assign n32784 = ( x35 & n32777 ) | ( x35 & n32783 ) | ( n32777 & n32783 ) ;
  assign n32785 = ( n17084 & n32782 ) | ( n17084 & n32784 ) | ( n32782 & n32784 ) ;
  assign n32786 = x35 & ~n32784 ;
  assign n32787 = x35 & ~n32780 ;
  assign n32788 = ( ~n17084 & n32786 ) | ( ~n17084 & n32787 ) | ( n32786 & n32787 ) ;
  assign n32789 = ( n32781 & ~n32785 ) | ( n32781 & n32788 ) | ( ~n32785 & n32788 ) ;
  assign n32790 = ~n32772 & n32789 ;
  assign n32791 = n32772 | n32790 ;
  assign n32792 = n32431 | n32451 ;
  assign n32793 = ( ~n32430 & n32451 ) | ( ~n32430 & n32792 ) | ( n32451 & n32792 ) ;
  assign n32794 = ( n32432 & ~n32434 ) | ( n32432 & n32793 ) | ( ~n32434 & n32793 ) ;
  assign n32795 = n32772 & n32789 ;
  assign n32796 = n32794 & n32795 ;
  assign n32797 = ( ~n32791 & n32794 ) | ( ~n32791 & n32796 ) | ( n32794 & n32796 ) ;
  assign n32798 = n32794 | n32795 ;
  assign n32799 = n32791 & ~n32798 ;
  assign n32800 = n32797 | n32799 ;
  assign n32818 = ~n32190 & n32454 ;
  assign n32819 = ( n32190 & n32191 ) | ( n32190 & ~n32818 ) | ( n32191 & ~n32818 ) ;
  assign n32801 = x127 & n4631 ;
  assign n32802 = x126 & n4626 ;
  assign n32803 = x125 & ~n4625 ;
  assign n32804 = n4943 & n32803 ;
  assign n32805 = n32802 | n32804 ;
  assign n32806 = n32801 | n32805 ;
  assign n32807 = n4634 | n32801 ;
  assign n32808 = n32805 | n32807 ;
  assign n32809 = ( n18763 & n32806 ) | ( n18763 & n32808 ) | ( n32806 & n32808 ) ;
  assign n32810 = x32 & n32808 ;
  assign n32811 = x32 & n32801 ;
  assign n32812 = ( x32 & n32805 ) | ( x32 & n32811 ) | ( n32805 & n32811 ) ;
  assign n32813 = ( n18763 & n32810 ) | ( n18763 & n32812 ) | ( n32810 & n32812 ) ;
  assign n32814 = x32 & ~n32812 ;
  assign n32815 = x32 & ~n32808 ;
  assign n32816 = ( ~n18763 & n32814 ) | ( ~n18763 & n32815 ) | ( n32814 & n32815 ) ;
  assign n32817 = ( n32809 & ~n32813 ) | ( n32809 & n32816 ) | ( ~n32813 & n32816 ) ;
  assign n32820 = n32817 & n32819 ;
  assign n32821 = n32819 & ~n32820 ;
  assign n32822 = ~n32800 & n32817 ;
  assign n32823 = ~n32819 & n32822 ;
  assign n32824 = ( ~n32800 & n32821 ) | ( ~n32800 & n32823 ) | ( n32821 & n32823 ) ;
  assign n32825 = n32800 & ~n32817 ;
  assign n32826 = ( n32800 & n32819 ) | ( n32800 & n32825 ) | ( n32819 & n32825 ) ;
  assign n32827 = ~n32821 & n32826 ;
  assign n32828 = n32824 | n32827 ;
  assign n32829 = n32493 | n32494 ;
  assign n32830 = n32457 & ~n32493 ;
  assign n32831 = ( n32485 & n32829 ) | ( n32485 & ~n32830 ) | ( n32829 & ~n32830 ) ;
  assign n32832 = ~n32828 & n32831 ;
  assign n32833 = n32828 & ~n32831 ;
  assign n32834 = n32832 | n32833 ;
  assign n32835 = ~n32498 & n32500 ;
  assign n32836 = n32511 & ~n32835 ;
  assign n32837 = n32507 | n32835 ;
  assign n32838 = ( n32151 & n32836 ) | ( n32151 & ~n32837 ) | ( n32836 & ~n32837 ) ;
  assign n32839 = n32505 & ~n32835 ;
  assign n32840 = ( n32156 & ~n32837 ) | ( n32156 & n32839 ) | ( ~n32837 & n32839 ) ;
  assign n32841 = ( n32155 & ~n32837 ) | ( n32155 & n32839 ) | ( ~n32837 & n32839 ) ;
  assign n32842 = ( ~n31818 & n32840 ) | ( ~n31818 & n32841 ) | ( n32840 & n32841 ) ;
  assign n32843 = ( ~n31819 & n32840 ) | ( ~n31819 & n32841 ) | ( n32840 & n32841 ) ;
  assign n32844 = ( ~n31118 & n32842 ) | ( ~n31118 & n32843 ) | ( n32842 & n32843 ) ;
  assign n32845 = ( ~n30754 & n32838 ) | ( ~n30754 & n32844 ) | ( n32838 & n32844 ) ;
  assign n32846 = n32834 & n32845 ;
  assign n32847 = n32834 | n32844 ;
  assign n32848 = ~n32834 & n32835 ;
  assign n32849 = ( n32511 & n32834 ) | ( n32511 & ~n32848 ) | ( n32834 & ~n32848 ) ;
  assign n32850 = ( n32507 & ~n32834 ) | ( n32507 & n32848 ) | ( ~n32834 & n32848 ) ;
  assign n32851 = ( n32151 & n32849 ) | ( n32151 & ~n32850 ) | ( n32849 & ~n32850 ) ;
  assign n32852 = ( ~n30754 & n32847 ) | ( ~n30754 & n32851 ) | ( n32847 & n32851 ) ;
  assign n32853 = ~n32846 & n32852 ;
  assign n33140 = n32820 | n32823 ;
  assign n33141 = ( n32800 & ~n32819 ) | ( n32800 & n32825 ) | ( ~n32819 & n32825 ) ;
  assign n33142 = ( n32821 & n33140 ) | ( n32821 & ~n33141 ) | ( n33140 & ~n33141 ) ;
  assign n32854 = x125 & n5554 ;
  assign n32855 = x124 & n5549 ;
  assign n32856 = x123 & ~n5548 ;
  assign n32857 = n5893 & n32856 ;
  assign n32858 = n32855 | n32857 ;
  assign n32859 = n32854 | n32858 ;
  assign n32860 = n5557 | n32854 ;
  assign n32861 = n32858 | n32860 ;
  assign n32862 = ( n17670 & n32859 ) | ( n17670 & n32861 ) | ( n32859 & n32861 ) ;
  assign n32863 = x35 & n32861 ;
  assign n32864 = x35 & n32854 ;
  assign n32865 = ( x35 & n32858 ) | ( x35 & n32864 ) | ( n32858 & n32864 ) ;
  assign n32866 = ( n17670 & n32863 ) | ( n17670 & n32865 ) | ( n32863 & n32865 ) ;
  assign n32867 = x35 & ~n32865 ;
  assign n32868 = x35 & ~n32861 ;
  assign n32869 = ( ~n17670 & n32867 ) | ( ~n17670 & n32868 ) | ( n32867 & n32868 ) ;
  assign n32870 = ( n32862 & ~n32866 ) | ( n32862 & n32869 ) | ( ~n32866 & n32869 ) ;
  assign n32871 = x127 & n4626 ;
  assign n32872 = x126 & ~n4625 ;
  assign n32873 = n4943 & n32872 ;
  assign n32874 = n32871 | n32873 ;
  assign n32875 = n4634 | n32874 ;
  assign n32876 = ( n19328 & n32874 ) | ( n19328 & n32875 ) | ( n32874 & n32875 ) ;
  assign n32877 = x32 & n32874 ;
  assign n32878 = ( x32 & n6918 ) | ( x32 & n32874 ) | ( n6918 & n32874 ) ;
  assign n32879 = ( n19328 & n32877 ) | ( n19328 & n32878 ) | ( n32877 & n32878 ) ;
  assign n32880 = x32 & ~n6918 ;
  assign n32881 = ~n32874 & n32880 ;
  assign n32882 = x32 & ~n32874 ;
  assign n32883 = ( ~n19328 & n32881 ) | ( ~n19328 & n32882 ) | ( n32881 & n32882 ) ;
  assign n32884 = ( n32876 & ~n32879 ) | ( n32876 & n32883 ) | ( ~n32879 & n32883 ) ;
  assign n32885 = n32789 & n32884 ;
  assign n32886 = ~n32772 & n32885 ;
  assign n32887 = ( n32797 & n32884 ) | ( n32797 & n32886 ) | ( n32884 & n32886 ) ;
  assign n32888 = n32789 | n32884 ;
  assign n32889 = ( ~n32772 & n32884 ) | ( ~n32772 & n32888 ) | ( n32884 & n32888 ) ;
  assign n32890 = n32797 | n32889 ;
  assign n32891 = ~n32887 & n32890 ;
  assign n32892 = n32763 | n32769 ;
  assign n32893 = n32738 | n32743 ;
  assign n33057 = n32690 | n32696 ;
  assign n33058 = ( n32690 & ~n32693 ) | ( n32690 & n33057 ) | ( ~n32693 & n33057 ) ;
  assign n32894 = ( ~n32619 & n32636 ) | ( ~n32619 & n32639 ) | ( n32636 & n32639 ) ;
  assign n32980 = n32581 | n32589 ;
  assign n32981 = ( n32581 & ~n32586 ) | ( n32581 & n32980 ) | ( ~n32586 & n32980 ) ;
  assign n32895 = n32532 & ~n32557 ;
  assign n32896 = ( n32532 & n32552 ) | ( n32532 & n32895 ) | ( n32552 & n32895 ) ;
  assign n32897 = n32551 | n32896 ;
  assign n32898 = x95 & n18290 ;
  assign n32899 = x63 & x94 ;
  assign n32900 = ~n18290 & n32899 ;
  assign n32901 = n32898 | n32900 ;
  assign n32902 = n32196 | n32540 ;
  assign n32903 = ( n32540 & ~n32542 ) | ( n32540 & n32902 ) | ( ~n32542 & n32902 ) ;
  assign n32904 = n32901 & ~n32903 ;
  assign n32905 = ~n32901 & n32903 ;
  assign n32906 = n32904 | n32905 ;
  assign n32907 = n5834 & ~n5850 ;
  assign n32908 = x97 & n17141 ;
  assign n32909 = x96 & ~n17140 ;
  assign n32910 = n17724 & n32909 ;
  assign n32911 = n32908 | n32910 ;
  assign n32912 = x98 & n17146 ;
  assign n32913 = n17149 | n32912 ;
  assign n32914 = n32911 | n32913 ;
  assign n32915 = x62 & ~n32914 ;
  assign n32916 = ~n32906 & n32915 ;
  assign n32917 = x62 & x98 ;
  assign n32918 = n17146 & n32917 ;
  assign n32919 = x62 & ~n32918 ;
  assign n32920 = ~n32911 & n32919 ;
  assign n32921 = ~n32906 & n32920 ;
  assign n32922 = ( ~n32907 & n32916 ) | ( ~n32907 & n32921 ) | ( n32916 & n32921 ) ;
  assign n32923 = ~x62 & n32914 ;
  assign n32924 = ~x62 & n32912 ;
  assign n32925 = ( ~x62 & n32911 ) | ( ~x62 & n32924 ) | ( n32911 & n32924 ) ;
  assign n32926 = ( ~n5850 & n32923 ) | ( ~n5850 & n32925 ) | ( n32923 & n32925 ) ;
  assign n32927 = n32923 & n32925 ;
  assign n32928 = ( n5834 & n32926 ) | ( n5834 & n32927 ) | ( n32926 & n32927 ) ;
  assign n32929 = ( ~n32906 & n32922 ) | ( ~n32906 & n32928 ) | ( n32922 & n32928 ) ;
  assign n32930 = n32906 & ~n32915 ;
  assign n32931 = n32906 & ~n32920 ;
  assign n32932 = ( n32907 & n32930 ) | ( n32907 & n32931 ) | ( n32930 & n32931 ) ;
  assign n32933 = ~n32928 & n32932 ;
  assign n32934 = n32929 | n32933 ;
  assign n32935 = n32551 & ~n32934 ;
  assign n32936 = ( n32896 & ~n32934 ) | ( n32896 & n32935 ) | ( ~n32934 & n32935 ) ;
  assign n32937 = n32897 & ~n32936 ;
  assign n32938 = n32934 | n32935 ;
  assign n32939 = x101 & n15552 ;
  assign n32940 = x100 & n15547 ;
  assign n32941 = x99 & ~n15546 ;
  assign n32942 = n16123 & n32941 ;
  assign n32943 = n32940 | n32942 ;
  assign n32944 = n32939 | n32943 ;
  assign n32945 = n15555 | n32939 ;
  assign n32946 = n32943 | n32945 ;
  assign n32947 = ( n6844 & n32944 ) | ( n6844 & n32946 ) | ( n32944 & n32946 ) ;
  assign n32948 = x59 & n32946 ;
  assign n32949 = x59 & n32939 ;
  assign n32950 = ( x59 & n32943 ) | ( x59 & n32949 ) | ( n32943 & n32949 ) ;
  assign n32951 = ( n6844 & n32948 ) | ( n6844 & n32950 ) | ( n32948 & n32950 ) ;
  assign n32952 = x59 & ~n32950 ;
  assign n32953 = x59 & ~n32946 ;
  assign n32954 = ( ~n6844 & n32952 ) | ( ~n6844 & n32953 ) | ( n32952 & n32953 ) ;
  assign n32955 = ( n32947 & ~n32951 ) | ( n32947 & n32954 ) | ( ~n32951 & n32954 ) ;
  assign n32956 = n32896 & ~n32955 ;
  assign n32957 = ( n32938 & ~n32955 ) | ( n32938 & n32956 ) | ( ~n32955 & n32956 ) ;
  assign n32958 = ~n32937 & n32957 ;
  assign n32959 = ~n32896 & n32955 ;
  assign n32960 = ~n32938 & n32959 ;
  assign n32961 = ( n32937 & n32955 ) | ( n32937 & n32960 ) | ( n32955 & n32960 ) ;
  assign n32962 = n32958 | n32961 ;
  assign n32963 = x104 & n14045 ;
  assign n32964 = x103 & n14040 ;
  assign n32965 = x102 & ~n14039 ;
  assign n32966 = n14552 & n32965 ;
  assign n32967 = n32964 | n32966 ;
  assign n32968 = n32963 | n32967 ;
  assign n32969 = n14048 | n32963 ;
  assign n32970 = n32967 | n32969 ;
  assign n32971 = ( n7911 & n32968 ) | ( n7911 & n32970 ) | ( n32968 & n32970 ) ;
  assign n32972 = x56 & n32970 ;
  assign n32973 = x56 & n32963 ;
  assign n32974 = ( x56 & n32967 ) | ( x56 & n32973 ) | ( n32967 & n32973 ) ;
  assign n32975 = ( n7911 & n32972 ) | ( n7911 & n32974 ) | ( n32972 & n32974 ) ;
  assign n32976 = x56 & ~n32974 ;
  assign n32977 = x56 & ~n32970 ;
  assign n32978 = ( ~n7911 & n32976 ) | ( ~n7911 & n32977 ) | ( n32976 & n32977 ) ;
  assign n32979 = ( n32971 & ~n32975 ) | ( n32971 & n32978 ) | ( ~n32975 & n32978 ) ;
  assign n32982 = ( ~n32962 & n32979 ) | ( ~n32962 & n32981 ) | ( n32979 & n32981 ) ;
  assign n32983 = ( n32962 & ~n32979 ) | ( n32962 & n32982 ) | ( ~n32979 & n32982 ) ;
  assign n32984 = ( ~n32981 & n32982 ) | ( ~n32981 & n32983 ) | ( n32982 & n32983 ) ;
  assign n32985 = n32610 & ~n32984 ;
  assign n32986 = ( n32616 & ~n32984 ) | ( n32616 & n32985 ) | ( ~n32984 & n32985 ) ;
  assign n32987 = ~n32610 & n32984 ;
  assign n32988 = ~n32616 & n32987 ;
  assign n32989 = n32986 | n32988 ;
  assign n32990 = x107 & n12574 ;
  assign n32991 = x106 & n12569 ;
  assign n32992 = x105 & ~n12568 ;
  assign n32993 = n13076 & n32992 ;
  assign n32994 = n32991 | n32993 ;
  assign n32995 = n32990 | n32994 ;
  assign n32996 = n12577 | n32990 ;
  assign n32997 = n32994 | n32996 ;
  assign n32998 = ( n9084 & n32995 ) | ( n9084 & n32997 ) | ( n32995 & n32997 ) ;
  assign n32999 = x53 & n32997 ;
  assign n33000 = x53 & n32990 ;
  assign n33001 = ( x53 & n32994 ) | ( x53 & n33000 ) | ( n32994 & n33000 ) ;
  assign n33002 = ( n9084 & n32999 ) | ( n9084 & n33001 ) | ( n32999 & n33001 ) ;
  assign n33003 = x53 & ~n33001 ;
  assign n33004 = x53 & ~n32997 ;
  assign n33005 = ( ~n9084 & n33003 ) | ( ~n9084 & n33004 ) | ( n33003 & n33004 ) ;
  assign n33006 = ( n32998 & ~n33002 ) | ( n32998 & n33005 ) | ( ~n33002 & n33005 ) ;
  assign n33007 = n32989 | n33006 ;
  assign n33008 = n32989 & ~n33006 ;
  assign n33009 = ( ~n32989 & n33007 ) | ( ~n32989 & n33008 ) | ( n33007 & n33008 ) ;
  assign n33010 = ~n32894 & n33009 ;
  assign n33011 = n32894 & ~n33009 ;
  assign n33012 = n33010 | n33011 ;
  assign n33013 = x110 & n11205 ;
  assign n33014 = x109 & n11200 ;
  assign n33015 = x108 & ~n11199 ;
  assign n33016 = n11679 & n33015 ;
  assign n33017 = n33014 | n33016 ;
  assign n33018 = n33013 | n33017 ;
  assign n33019 = n11208 | n33013 ;
  assign n33020 = n33017 | n33019 ;
  assign n33021 = ( n10330 & n33018 ) | ( n10330 & n33020 ) | ( n33018 & n33020 ) ;
  assign n33022 = x50 & n33020 ;
  assign n33023 = x50 & n33013 ;
  assign n33024 = ( x50 & n33017 ) | ( x50 & n33023 ) | ( n33017 & n33023 ) ;
  assign n33025 = ( n10330 & n33022 ) | ( n10330 & n33024 ) | ( n33022 & n33024 ) ;
  assign n33026 = x50 & ~n33024 ;
  assign n33027 = x50 & ~n33020 ;
  assign n33028 = ( ~n10330 & n33026 ) | ( ~n10330 & n33027 ) | ( n33026 & n33027 ) ;
  assign n33029 = ( n33021 & ~n33025 ) | ( n33021 & n33028 ) | ( ~n33025 & n33028 ) ;
  assign n33030 = n33012 & n33029 ;
  assign n33031 = n32639 | n33029 ;
  assign n33032 = n32636 | n33029 ;
  assign n33033 = ( ~n32619 & n33031 ) | ( ~n32619 & n33032 ) | ( n33031 & n33032 ) ;
  assign n33034 = ( ~n33009 & n33029 ) | ( ~n33009 & n33033 ) | ( n33029 & n33033 ) ;
  assign n33035 = n33010 | n33034 ;
  assign n33036 = ~n33030 & n33035 ;
  assign n33037 = ~n32664 & n32666 ;
  assign n33038 = ( n32664 & n32669 ) | ( n32664 & ~n33037 ) | ( n32669 & ~n33037 ) ;
  assign n33039 = n33036 & ~n33038 ;
  assign n33040 = ~n33036 & n33038 ;
  assign n33041 = n33039 | n33040 ;
  assign n33042 = x113 & n9933 ;
  assign n33043 = x112 & n9928 ;
  assign n33044 = x111 & ~n9927 ;
  assign n33045 = n10379 & n33044 ;
  assign n33046 = n33043 | n33045 ;
  assign n33047 = n33042 | n33046 ;
  assign n33048 = n9936 | n33042 ;
  assign n33049 = n33046 | n33048 ;
  assign n33050 = ( ~n11642 & n33047 ) | ( ~n11642 & n33049 ) | ( n33047 & n33049 ) ;
  assign n33051 = n33047 & n33049 ;
  assign n33052 = ( n11626 & n33050 ) | ( n11626 & n33051 ) | ( n33050 & n33051 ) ;
  assign n33053 = x47 & n33052 ;
  assign n33054 = x47 & ~n33052 ;
  assign n33055 = ( n33052 & ~n33053 ) | ( n33052 & n33054 ) | ( ~n33053 & n33054 ) ;
  assign n33056 = n33041 & n33055 ;
  assign n33059 = n33056 & n33058 ;
  assign n33060 = n33035 & ~n33055 ;
  assign n33061 = ~n33030 & n33060 ;
  assign n33062 = ( n33038 & n33055 ) | ( n33038 & ~n33061 ) | ( n33055 & ~n33061 ) ;
  assign n33063 = n33039 | n33062 ;
  assign n33064 = ( n33058 & n33059 ) | ( n33058 & ~n33063 ) | ( n33059 & ~n33063 ) ;
  assign n33065 = ~n33056 & n33063 ;
  assign n33066 = ~n33058 & n33065 ;
  assign n33067 = n33064 | n33066 ;
  assign n33068 = x116 & n8724 ;
  assign n33069 = x115 & n8719 ;
  assign n33070 = x114 & ~n8718 ;
  assign n33071 = n9149 & n33070 ;
  assign n33072 = n33069 | n33071 ;
  assign n33073 = n33068 | n33072 ;
  assign n33074 = n8727 | n33068 ;
  assign n33075 = n33072 | n33074 ;
  assign n33076 = ( ~n13040 & n33073 ) | ( ~n13040 & n33075 ) | ( n33073 & n33075 ) ;
  assign n33077 = n33073 & n33075 ;
  assign n33078 = ( n13022 & n33076 ) | ( n13022 & n33077 ) | ( n33076 & n33077 ) ;
  assign n33079 = x44 & n33078 ;
  assign n33080 = x44 & ~n33078 ;
  assign n33081 = ( n33078 & ~n33079 ) | ( n33078 & n33080 ) | ( ~n33079 & n33080 ) ;
  assign n33082 = n33066 | n33081 ;
  assign n33083 = n33064 | n33082 ;
  assign n33084 = ~n33081 & n33083 ;
  assign n33085 = ( ~n33067 & n33083 ) | ( ~n33067 & n33084 ) | ( n33083 & n33084 ) ;
  assign n33086 = n32714 | n32719 ;
  assign n33087 = ( n32714 & ~n32716 ) | ( n32714 & n33086 ) | ( ~n32716 & n33086 ) ;
  assign n33088 = n33085 & n33087 ;
  assign n33089 = n33085 | n33087 ;
  assign n33090 = ~n33088 & n33089 ;
  assign n33091 = x119 & n7566 ;
  assign n33092 = x118 & n7561 ;
  assign n33093 = x117 & ~n7560 ;
  assign n33094 = n7953 & n33093 ;
  assign n33095 = n33092 | n33094 ;
  assign n33096 = n33091 | n33095 ;
  assign n33097 = n7569 | n33091 ;
  assign n33098 = n33095 | n33097 ;
  assign n33099 = ( n14496 & n33096 ) | ( n14496 & n33098 ) | ( n33096 & n33098 ) ;
  assign n33100 = x41 & n33098 ;
  assign n33101 = x41 & n33091 ;
  assign n33102 = ( x41 & n33095 ) | ( x41 & n33101 ) | ( n33095 & n33101 ) ;
  assign n33103 = ( n14496 & n33100 ) | ( n14496 & n33102 ) | ( n33100 & n33102 ) ;
  assign n33104 = x41 & ~n33102 ;
  assign n33105 = x41 & ~n33098 ;
  assign n33106 = ( ~n14496 & n33104 ) | ( ~n14496 & n33105 ) | ( n33104 & n33105 ) ;
  assign n33107 = ( n33099 & ~n33103 ) | ( n33099 & n33106 ) | ( ~n33103 & n33106 ) ;
  assign n33108 = ~n33090 & n33107 ;
  assign n33109 = n33090 & ~n33107 ;
  assign n33110 = n33108 | n33109 ;
  assign n33111 = n32893 & ~n33110 ;
  assign n33112 = ~n32893 & n33110 ;
  assign n33113 = n33111 | n33112 ;
  assign n33114 = x122 & n6536 ;
  assign n33115 = x121 & n6531 ;
  assign n33116 = x120 & ~n6530 ;
  assign n33117 = n6871 & n33116 ;
  assign n33118 = n33115 | n33117 ;
  assign n33119 = n33114 | n33118 ;
  assign n33120 = n6539 | n33114 ;
  assign n33121 = n33118 | n33120 ;
  assign n33122 = ( n16043 & n33119 ) | ( n16043 & n33121 ) | ( n33119 & n33121 ) ;
  assign n33123 = x38 & n33121 ;
  assign n33124 = x38 & n33114 ;
  assign n33125 = ( x38 & n33118 ) | ( x38 & n33124 ) | ( n33118 & n33124 ) ;
  assign n33126 = ( n16043 & n33123 ) | ( n16043 & n33125 ) | ( n33123 & n33125 ) ;
  assign n33127 = x38 & ~n33125 ;
  assign n33128 = x38 & ~n33121 ;
  assign n33129 = ( ~n16043 & n33127 ) | ( ~n16043 & n33128 ) | ( n33127 & n33128 ) ;
  assign n33130 = ( n33122 & ~n33126 ) | ( n33122 & n33129 ) | ( ~n33126 & n33129 ) ;
  assign n33131 = n33113 | n33130 ;
  assign n33132 = n33113 & ~n33130 ;
  assign n33133 = ( ~n33113 & n33131 ) | ( ~n33113 & n33132 ) | ( n33131 & n33132 ) ;
  assign n33134 = ~n32892 & n33133 ;
  assign n33135 = n32892 & ~n33133 ;
  assign n33136 = n33134 | n33135 ;
  assign n33137 = ( n32870 & n32891 ) | ( n32870 & ~n33136 ) | ( n32891 & ~n33136 ) ;
  assign n33138 = ( ~n32891 & n33136 ) | ( ~n32891 & n33137 ) | ( n33136 & n33137 ) ;
  assign n33139 = ( ~n32870 & n33137 ) | ( ~n32870 & n33138 ) | ( n33137 & n33138 ) ;
  assign n33143 = ~n33139 & n33142 ;
  assign n33144 = n33142 & ~n33143 ;
  assign n33145 = n33139 | n33142 ;
  assign n33146 = ~n33144 & n33145 ;
  assign n33147 = ~n32832 & n32834 ;
  assign n33148 = ( ~n32832 & n32844 ) | ( ~n32832 & n33147 ) | ( n32844 & n33147 ) ;
  assign n33149 = n32832 | n32848 ;
  assign n33150 = ( n32511 & n33147 ) | ( n32511 & ~n33149 ) | ( n33147 & ~n33149 ) ;
  assign n33151 = ( n32507 & ~n33147 ) | ( n32507 & n33149 ) | ( ~n33147 & n33149 ) ;
  assign n33152 = ( n32151 & n33150 ) | ( n32151 & ~n33151 ) | ( n33150 & ~n33151 ) ;
  assign n33153 = ( ~n30754 & n33148 ) | ( ~n30754 & n33152 ) | ( n33148 & n33152 ) ;
  assign n33154 = n33146 & n33153 ;
  assign n33155 = n33146 | n33147 ;
  assign n33156 = n32832 & ~n33146 ;
  assign n33157 = ( n32844 & n33155 ) | ( n32844 & ~n33156 ) | ( n33155 & ~n33156 ) ;
  assign n33158 = ~n33146 & n33151 ;
  assign n33159 = ~n33146 & n33149 ;
  assign n33160 = ( n32511 & n33155 ) | ( n32511 & ~n33159 ) | ( n33155 & ~n33159 ) ;
  assign n33161 = ( n32151 & ~n33158 ) | ( n32151 & n33160 ) | ( ~n33158 & n33160 ) ;
  assign n33162 = ( ~n30754 & n33157 ) | ( ~n30754 & n33161 ) | ( n33157 & n33161 ) ;
  assign n33163 = ~n33154 & n33162 ;
  assign n33325 = ( n33040 & ~n33041 ) | ( n33040 & n33062 ) | ( ~n33041 & n33062 ) ;
  assign n33164 = n32936 | n32961 ;
  assign n33165 = n32905 | n32928 ;
  assign n33166 = ~n32905 & n32906 ;
  assign n33167 = ( n32922 & n33165 ) | ( n32922 & ~n33166 ) | ( n33165 & ~n33166 ) ;
  assign n33168 = x96 & n18290 ;
  assign n33169 = x63 & x95 ;
  assign n33170 = ~n18290 & n33169 ;
  assign n33171 = n33168 | n33170 ;
  assign n33172 = n32901 & ~n33171 ;
  assign n33173 = ~n32901 & n33171 ;
  assign n33174 = n33172 | n33173 ;
  assign n33175 = n32901 | n33174 ;
  assign n33176 = n32903 & ~n33175 ;
  assign n33177 = ( n32928 & ~n33174 ) | ( n32928 & n33176 ) | ( ~n33174 & n33176 ) ;
  assign n33178 = ( n32906 & n33174 ) | ( n32906 & ~n33176 ) | ( n33174 & ~n33176 ) ;
  assign n33179 = ( n32922 & n33177 ) | ( n32922 & ~n33178 ) | ( n33177 & ~n33178 ) ;
  assign n33180 = n33167 & ~n33179 ;
  assign n33181 = x99 & n17146 ;
  assign n33182 = x98 & n17141 ;
  assign n33183 = x97 & ~n17140 ;
  assign n33184 = n17724 & n33183 ;
  assign n33185 = n33182 | n33184 ;
  assign n33186 = n33181 | n33185 ;
  assign n33187 = n17149 | n33181 ;
  assign n33188 = n33185 | n33187 ;
  assign n33189 = ( n6164 & n33186 ) | ( n6164 & n33188 ) | ( n33186 & n33188 ) ;
  assign n33190 = x62 & n33188 ;
  assign n33191 = x62 & n33181 ;
  assign n33192 = ( x62 & n33185 ) | ( x62 & n33191 ) | ( n33185 & n33191 ) ;
  assign n33193 = ( n6164 & n33190 ) | ( n6164 & n33192 ) | ( n33190 & n33192 ) ;
  assign n33194 = x62 & ~n33192 ;
  assign n33195 = x62 & ~n33188 ;
  assign n33196 = ( ~n6164 & n33194 ) | ( ~n6164 & n33195 ) | ( n33194 & n33195 ) ;
  assign n33197 = ( n33189 & ~n33193 ) | ( n33189 & n33196 ) | ( ~n33193 & n33196 ) ;
  assign n33198 = n33174 | n33176 ;
  assign n33199 = n32928 | n33198 ;
  assign n33200 = n32906 & ~n33198 ;
  assign n33201 = ( n32922 & n33199 ) | ( n32922 & ~n33200 ) | ( n33199 & ~n33200 ) ;
  assign n33202 = n33197 & ~n33201 ;
  assign n33203 = ( n33180 & n33197 ) | ( n33180 & n33202 ) | ( n33197 & n33202 ) ;
  assign n33204 = ~n33197 & n33201 ;
  assign n33205 = ~n33180 & n33204 ;
  assign n33206 = n33203 | n33205 ;
  assign n33207 = x102 & n15552 ;
  assign n33208 = x101 & n15547 ;
  assign n33209 = x100 & ~n15546 ;
  assign n33210 = n16123 & n33209 ;
  assign n33211 = n33208 | n33210 ;
  assign n33212 = n33207 | n33211 ;
  assign n33213 = n15555 | n33207 ;
  assign n33214 = n33211 | n33213 ;
  assign n33215 = ( n7178 & n33212 ) | ( n7178 & n33214 ) | ( n33212 & n33214 ) ;
  assign n33216 = x59 & n33214 ;
  assign n33217 = x59 & n33207 ;
  assign n33218 = ( x59 & n33211 ) | ( x59 & n33217 ) | ( n33211 & n33217 ) ;
  assign n33219 = ( n7178 & n33216 ) | ( n7178 & n33218 ) | ( n33216 & n33218 ) ;
  assign n33220 = x59 & ~n33218 ;
  assign n33221 = x59 & ~n33214 ;
  assign n33222 = ( ~n7178 & n33220 ) | ( ~n7178 & n33221 ) | ( n33220 & n33221 ) ;
  assign n33223 = ( n33215 & ~n33219 ) | ( n33215 & n33222 ) | ( ~n33219 & n33222 ) ;
  assign n33224 = n33206 | n33223 ;
  assign n33225 = n33206 & n33223 ;
  assign n33226 = n33224 & ~n33225 ;
  assign n33227 = n33164 & ~n33226 ;
  assign n33228 = ~n33164 & n33226 ;
  assign n33229 = n33227 | n33228 ;
  assign n33230 = x105 & n14045 ;
  assign n33231 = x104 & n14040 ;
  assign n33232 = x103 & ~n14039 ;
  assign n33233 = n14552 & n33232 ;
  assign n33234 = n33231 | n33233 ;
  assign n33235 = n33230 | n33234 ;
  assign n33236 = n14048 | n33230 ;
  assign n33237 = n33234 | n33236 ;
  assign n33238 = ( n8273 & n33235 ) | ( n8273 & n33237 ) | ( n33235 & n33237 ) ;
  assign n33239 = x56 & n33237 ;
  assign n33240 = x56 & n33230 ;
  assign n33241 = ( x56 & n33234 ) | ( x56 & n33240 ) | ( n33234 & n33240 ) ;
  assign n33242 = ( n8273 & n33239 ) | ( n8273 & n33241 ) | ( n33239 & n33241 ) ;
  assign n33243 = x56 & ~n33241 ;
  assign n33244 = x56 & ~n33237 ;
  assign n33245 = ( ~n8273 & n33243 ) | ( ~n8273 & n33244 ) | ( n33243 & n33244 ) ;
  assign n33246 = ( n33238 & ~n33242 ) | ( n33238 & n33245 ) | ( ~n33242 & n33245 ) ;
  assign n33247 = ~n33229 & n33246 ;
  assign n33248 = n33229 & ~n33246 ;
  assign n33249 = n33247 | n33248 ;
  assign n33250 = ~n32962 & n32981 ;
  assign n33251 = n32981 & ~n33250 ;
  assign n33252 = n32962 | n33250 ;
  assign n33253 = ~n33251 & n33252 ;
  assign n33254 = n32979 | n33250 ;
  assign n33255 = ( n33250 & ~n33253 ) | ( n33250 & n33254 ) | ( ~n33253 & n33254 ) ;
  assign n33256 = ~n33249 & n33255 ;
  assign n33257 = n33249 & ~n33255 ;
  assign n33258 = n33256 | n33257 ;
  assign n33259 = x108 & n12574 ;
  assign n33260 = x107 & n12569 ;
  assign n33261 = x106 & ~n12568 ;
  assign n33262 = n13076 & n33261 ;
  assign n33263 = n33260 | n33262 ;
  assign n33264 = n33259 | n33263 ;
  assign n33265 = n12577 | n33259 ;
  assign n33266 = n33263 | n33265 ;
  assign n33267 = ( n9479 & n33264 ) | ( n9479 & n33266 ) | ( n33264 & n33266 ) ;
  assign n33268 = x53 & n33266 ;
  assign n33269 = x53 & n33259 ;
  assign n33270 = ( x53 & n33263 ) | ( x53 & n33269 ) | ( n33263 & n33269 ) ;
  assign n33271 = ( n9479 & n33268 ) | ( n9479 & n33270 ) | ( n33268 & n33270 ) ;
  assign n33272 = x53 & ~n33270 ;
  assign n33273 = x53 & ~n33266 ;
  assign n33274 = ( ~n9479 & n33272 ) | ( ~n9479 & n33273 ) | ( n33272 & n33273 ) ;
  assign n33275 = ( n33267 & ~n33271 ) | ( n33267 & n33274 ) | ( ~n33271 & n33274 ) ;
  assign n33276 = ~n33258 & n33275 ;
  assign n33277 = n33258 & ~n33275 ;
  assign n33278 = n33276 | n33277 ;
  assign n33279 = n32986 | n33006 ;
  assign n33280 = ( n32986 & ~n32989 ) | ( n32986 & n33279 ) | ( ~n32989 & n33279 ) ;
  assign n33281 = ~n33278 & n33280 ;
  assign n33282 = n33278 & ~n33280 ;
  assign n33283 = n33281 | n33282 ;
  assign n33284 = x111 & n11205 ;
  assign n33285 = x110 & n11200 ;
  assign n33286 = x109 & ~n11199 ;
  assign n33287 = n11679 & n33286 ;
  assign n33288 = n33285 | n33287 ;
  assign n33289 = n33284 | n33288 ;
  assign n33290 = n11208 | n33284 ;
  assign n33291 = n33288 | n33290 ;
  assign n33292 = ( n10749 & n33289 ) | ( n10749 & n33291 ) | ( n33289 & n33291 ) ;
  assign n33293 = x50 & n33291 ;
  assign n33294 = x50 & n33284 ;
  assign n33295 = ( x50 & n33288 ) | ( x50 & n33294 ) | ( n33288 & n33294 ) ;
  assign n33296 = ( n10749 & n33293 ) | ( n10749 & n33295 ) | ( n33293 & n33295 ) ;
  assign n33297 = x50 & ~n33295 ;
  assign n33298 = x50 & ~n33291 ;
  assign n33299 = ( ~n10749 & n33297 ) | ( ~n10749 & n33298 ) | ( n33297 & n33298 ) ;
  assign n33300 = ( n33292 & ~n33296 ) | ( n33292 & n33299 ) | ( ~n33296 & n33299 ) ;
  assign n33301 = n33283 | n33300 ;
  assign n33302 = n33283 & ~n33300 ;
  assign n33303 = ( ~n33283 & n33301 ) | ( ~n33283 & n33302 ) | ( n33301 & n33302 ) ;
  assign n33304 = ( n33011 & ~n33012 ) | ( n33011 & n33034 ) | ( ~n33012 & n33034 ) ;
  assign n33305 = n33303 & ~n33304 ;
  assign n33306 = ~n33303 & n33304 ;
  assign n33307 = n33305 | n33306 ;
  assign n33308 = x114 & n9933 ;
  assign n33309 = x113 & n9928 ;
  assign n33310 = x112 & ~n9927 ;
  assign n33311 = n10379 & n33310 ;
  assign n33312 = n33309 | n33311 ;
  assign n33313 = n33308 | n33312 ;
  assign n33314 = n9936 | n33308 ;
  assign n33315 = n33312 | n33314 ;
  assign n33316 = ( ~n12095 & n33313 ) | ( ~n12095 & n33315 ) | ( n33313 & n33315 ) ;
  assign n33317 = n33313 & n33315 ;
  assign n33318 = ( n12079 & n33316 ) | ( n12079 & n33317 ) | ( n33316 & n33317 ) ;
  assign n33319 = x47 & n33318 ;
  assign n33320 = x47 & ~n33318 ;
  assign n33321 = ( n33318 & ~n33319 ) | ( n33318 & n33320 ) | ( ~n33319 & n33320 ) ;
  assign n33322 = n33307 & ~n33321 ;
  assign n33323 = ~n33307 & n33321 ;
  assign n33324 = n33322 | n33323 ;
  assign n33326 = ~n33324 & n33325 ;
  assign n33327 = n33325 & ~n33326 ;
  assign n33328 = n33324 | n33325 ;
  assign n33329 = x117 & n8724 ;
  assign n33330 = x116 & n8719 ;
  assign n33331 = x115 & ~n8718 ;
  assign n33332 = n9149 & n33331 ;
  assign n33333 = n33330 | n33332 ;
  assign n33334 = n33329 | n33333 ;
  assign n33335 = n8727 | n33329 ;
  assign n33336 = n33333 | n33335 ;
  assign n33337 = ( ~n13522 & n33334 ) | ( ~n13522 & n33336 ) | ( n33334 & n33336 ) ;
  assign n33338 = n33334 & n33336 ;
  assign n33339 = ( n13503 & n33337 ) | ( n13503 & n33338 ) | ( n33337 & n33338 ) ;
  assign n33340 = x44 & n33339 ;
  assign n33341 = x44 & ~n33339 ;
  assign n33342 = ( n33339 & ~n33340 ) | ( n33339 & n33341 ) | ( ~n33340 & n33341 ) ;
  assign n33343 = n33328 & ~n33342 ;
  assign n33344 = ~n33327 & n33343 ;
  assign n33345 = ~n33328 & n33342 ;
  assign n33346 = ( n33327 & n33342 ) | ( n33327 & n33345 ) | ( n33342 & n33345 ) ;
  assign n33347 = n33344 | n33346 ;
  assign n33348 = ~n33066 & n33081 ;
  assign n33349 = ~n33064 & n33348 ;
  assign n33350 = n33064 & ~n33347 ;
  assign n33351 = ( ~n33347 & n33349 ) | ( ~n33347 & n33350 ) | ( n33349 & n33350 ) ;
  assign n33352 = ~n33064 & n33347 ;
  assign n33353 = ~n33349 & n33352 ;
  assign n33354 = n33351 | n33353 ;
  assign n33355 = x120 & n7566 ;
  assign n33356 = x119 & n7561 ;
  assign n33357 = x118 & ~n7560 ;
  assign n33358 = n7953 & n33357 ;
  assign n33359 = n33356 | n33358 ;
  assign n33360 = n33355 | n33359 ;
  assign n33361 = n7569 | n33355 ;
  assign n33362 = n33359 | n33361 ;
  assign n33363 = ( n14991 & n33360 ) | ( n14991 & n33362 ) | ( n33360 & n33362 ) ;
  assign n33364 = x41 & n33362 ;
  assign n33365 = x41 & n33355 ;
  assign n33366 = ( x41 & n33359 ) | ( x41 & n33365 ) | ( n33359 & n33365 ) ;
  assign n33367 = ( n14991 & n33364 ) | ( n14991 & n33366 ) | ( n33364 & n33366 ) ;
  assign n33368 = x41 & ~n33366 ;
  assign n33369 = x41 & ~n33362 ;
  assign n33370 = ( ~n14991 & n33368 ) | ( ~n14991 & n33369 ) | ( n33368 & n33369 ) ;
  assign n33371 = ( n33363 & ~n33367 ) | ( n33363 & n33370 ) | ( ~n33367 & n33370 ) ;
  assign n33372 = ~n33354 & n33371 ;
  assign n33373 = n33354 & ~n33371 ;
  assign n33374 = n33372 | n33373 ;
  assign n33375 = ( ~n33085 & n33087 ) | ( ~n33085 & n33107 ) | ( n33087 & n33107 ) ;
  assign n33376 = ~n33374 & n33375 ;
  assign n33377 = n33374 & ~n33375 ;
  assign n33378 = n33376 | n33377 ;
  assign n33379 = x123 & n6536 ;
  assign n33380 = x122 & n6531 ;
  assign n33381 = x121 & ~n6530 ;
  assign n33382 = n6871 & n33381 ;
  assign n33383 = n33380 | n33382 ;
  assign n33384 = n33379 | n33383 ;
  assign n33385 = n6539 | n33379 ;
  assign n33386 = n33383 | n33385 ;
  assign n33387 = ( n16086 & n33384 ) | ( n16086 & n33386 ) | ( n33384 & n33386 ) ;
  assign n33388 = x38 & n33386 ;
  assign n33389 = x38 & n33379 ;
  assign n33390 = ( x38 & n33383 ) | ( x38 & n33389 ) | ( n33383 & n33389 ) ;
  assign n33391 = ( n16086 & n33388 ) | ( n16086 & n33390 ) | ( n33388 & n33390 ) ;
  assign n33392 = x38 & ~n33390 ;
  assign n33393 = x38 & ~n33386 ;
  assign n33394 = ( ~n16086 & n33392 ) | ( ~n16086 & n33393 ) | ( n33392 & n33393 ) ;
  assign n33395 = ( n33387 & ~n33391 ) | ( n33387 & n33394 ) | ( ~n33391 & n33394 ) ;
  assign n33396 = n33378 | n33395 ;
  assign n33397 = n33378 & ~n33395 ;
  assign n33398 = ( ~n33378 & n33396 ) | ( ~n33378 & n33397 ) | ( n33396 & n33397 ) ;
  assign n33399 = n33111 | n33130 ;
  assign n33400 = ( n33111 & ~n33113 ) | ( n33111 & n33399 ) | ( ~n33113 & n33399 ) ;
  assign n33401 = n33398 & ~n33400 ;
  assign n33402 = ~n33398 & n33400 ;
  assign n33403 = n33401 | n33402 ;
  assign n33404 = x126 & n5554 ;
  assign n33405 = x125 & n5549 ;
  assign n33406 = x124 & ~n5548 ;
  assign n33407 = n5893 & n33406 ;
  assign n33408 = n33405 | n33407 ;
  assign n33409 = n33404 | n33408 ;
  assign n33410 = n5557 | n33404 ;
  assign n33411 = n33408 | n33410 ;
  assign n33412 = ( n18220 & n33409 ) | ( n18220 & n33411 ) | ( n33409 & n33411 ) ;
  assign n33413 = x35 & n33411 ;
  assign n33414 = x35 & n33404 ;
  assign n33415 = ( x35 & n33408 ) | ( x35 & n33414 ) | ( n33408 & n33414 ) ;
  assign n33416 = ( n18220 & n33413 ) | ( n18220 & n33415 ) | ( n33413 & n33415 ) ;
  assign n33417 = x35 & ~n33415 ;
  assign n33418 = x35 & ~n33411 ;
  assign n33419 = ( ~n18220 & n33417 ) | ( ~n18220 & n33418 ) | ( n33417 & n33418 ) ;
  assign n33420 = ( n33412 & ~n33416 ) | ( n33412 & n33419 ) | ( ~n33416 & n33419 ) ;
  assign n33421 = n33403 & n33420 ;
  assign n33422 = n33398 & ~n33420 ;
  assign n33423 = ( n33400 & n33420 ) | ( n33400 & ~n33422 ) | ( n33420 & ~n33422 ) ;
  assign n33424 = n33401 | n33423 ;
  assign n33425 = ~n33421 & n33424 ;
  assign n33426 = x127 & ~n4625 ;
  assign n33427 = n4943 & n33426 ;
  assign n33428 = n4634 & n19877 ;
  assign n33429 = n33427 | n33428 ;
  assign n33430 = n4634 & n19880 ;
  assign n33431 = n33427 | n33430 ;
  assign n33432 = ( n18202 & n33429 ) | ( n18202 & n33431 ) | ( n33429 & n33431 ) ;
  assign n33433 = n33429 & n33431 ;
  assign n33434 = ( n18212 & n33432 ) | ( n18212 & n33433 ) | ( n33432 & n33433 ) ;
  assign n33435 = ( n18214 & n33432 ) | ( n18214 & n33433 ) | ( n33432 & n33433 ) ;
  assign n33436 = ( n14002 & n33434 ) | ( n14002 & n33435 ) | ( n33434 & n33435 ) ;
  assign n33437 = x32 & n33434 ;
  assign n33438 = x32 & n33435 ;
  assign n33439 = ( n14002 & n33437 ) | ( n14002 & n33438 ) | ( n33437 & n33438 ) ;
  assign n33440 = x32 & ~n33438 ;
  assign n33441 = x32 & ~n33437 ;
  assign n33442 = ( ~n14002 & n33440 ) | ( ~n14002 & n33441 ) | ( n33440 & n33441 ) ;
  assign n33443 = ( n33436 & ~n33439 ) | ( n33436 & n33442 ) | ( ~n33439 & n33442 ) ;
  assign n33444 = n32870 | n33135 ;
  assign n33445 = ( n33135 & ~n33136 ) | ( n33135 & n33444 ) | ( ~n33136 & n33444 ) ;
  assign n33446 = ( n33425 & n33443 ) | ( n33425 & ~n33445 ) | ( n33443 & ~n33445 ) ;
  assign n33447 = ( ~n33443 & n33445 ) | ( ~n33443 & n33446 ) | ( n33445 & n33446 ) ;
  assign n33448 = ( ~n33425 & n33446 ) | ( ~n33425 & n33447 ) | ( n33446 & n33447 ) ;
  assign n33449 = n32870 & ~n33136 ;
  assign n33450 = ~n32870 & n33136 ;
  assign n33451 = n33449 | n33450 ;
  assign n33452 = ~n32887 & n33451 ;
  assign n33453 = ( n32887 & n32891 ) | ( n32887 & ~n33452 ) | ( n32891 & ~n33452 ) ;
  assign n33454 = n33448 & n33453 ;
  assign n33455 = ~n33448 & n33453 ;
  assign n33456 = n33448 | n33455 ;
  assign n33457 = ~n33454 & n33456 ;
  assign n33458 = ~n33143 & n33146 ;
  assign n33459 = ( ~n33143 & n33147 ) | ( ~n33143 & n33458 ) | ( n33147 & n33458 ) ;
  assign n33460 = n33457 | n33459 ;
  assign n33461 = n32832 | n33143 ;
  assign n33462 = ( n33143 & ~n33146 ) | ( n33143 & n33461 ) | ( ~n33146 & n33461 ) ;
  assign n33463 = ~n33457 & n33462 ;
  assign n33464 = ( n32844 & n33460 ) | ( n32844 & ~n33463 ) | ( n33460 & ~n33463 ) ;
  assign n33465 = n33143 | n33159 ;
  assign n33466 = ~n33143 & n33155 ;
  assign n33467 = ( n32511 & ~n33465 ) | ( n32511 & n33466 ) | ( ~n33465 & n33466 ) ;
  assign n33468 = n33457 | n33467 ;
  assign n33469 = n33457 | n33458 ;
  assign n33470 = n33143 & ~n33457 ;
  assign n33471 = ( n33151 & ~n33469 ) | ( n33151 & n33470 ) | ( ~n33469 & n33470 ) ;
  assign n33472 = ( n32151 & n33468 ) | ( n32151 & ~n33471 ) | ( n33468 & ~n33471 ) ;
  assign n33473 = ( ~n30754 & n33464 ) | ( ~n30754 & n33472 ) | ( n33464 & n33472 ) ;
  assign n33474 = ( n32844 & n33459 ) | ( n32844 & ~n33462 ) | ( n33459 & ~n33462 ) ;
  assign n33475 = ( n33143 & n33151 ) | ( n33143 & ~n33458 ) | ( n33151 & ~n33458 ) ;
  assign n33476 = ( n32151 & n33467 ) | ( n32151 & ~n33475 ) | ( n33467 & ~n33475 ) ;
  assign n33477 = ( ~n30754 & n33474 ) | ( ~n30754 & n33476 ) | ( n33474 & n33476 ) ;
  assign n33478 = ( n33448 & n33453 ) | ( n33448 & n33477 ) | ( n33453 & n33477 ) ;
  assign n33479 = ( n33454 & n33473 ) | ( n33454 & ~n33478 ) | ( n33473 & ~n33478 ) ;
  assign n33480 = n33326 | n33346 ;
  assign n33481 = x100 & n17146 ;
  assign n33482 = x99 & n17141 ;
  assign n33483 = x98 & ~n17140 ;
  assign n33484 = n17724 & n33483 ;
  assign n33485 = n33482 | n33484 ;
  assign n33486 = n33481 | n33485 ;
  assign n33487 = n17149 | n33481 ;
  assign n33488 = n33485 | n33487 ;
  assign n33489 = ( n6483 & n33486 ) | ( n6483 & n33488 ) | ( n33486 & n33488 ) ;
  assign n33490 = x62 & n33488 ;
  assign n33491 = x62 & n33481 ;
  assign n33492 = ( x62 & n33485 ) | ( x62 & n33491 ) | ( n33485 & n33491 ) ;
  assign n33493 = ( n6483 & n33490 ) | ( n6483 & n33492 ) | ( n33490 & n33492 ) ;
  assign n33494 = x62 & ~n33492 ;
  assign n33495 = x62 & ~n33488 ;
  assign n33496 = ( ~n6483 & n33494 ) | ( ~n6483 & n33495 ) | ( n33494 & n33495 ) ;
  assign n33497 = ( n33489 & ~n33493 ) | ( n33489 & n33496 ) | ( ~n33493 & n33496 ) ;
  assign n33498 = n33172 | n33176 ;
  assign n33499 = ~n33172 & n33174 ;
  assign n33500 = ( n32928 & n33498 ) | ( n32928 & ~n33499 ) | ( n33498 & ~n33499 ) ;
  assign n33501 = ( n32906 & ~n33498 ) | ( n32906 & n33499 ) | ( ~n33498 & n33499 ) ;
  assign n33502 = ( n32922 & n33500 ) | ( n32922 & ~n33501 ) | ( n33500 & ~n33501 ) ;
  assign n33503 = x97 & n18290 ;
  assign n33504 = x63 & x96 ;
  assign n33505 = ~n18290 & n33504 ;
  assign n33506 = n33503 | n33505 ;
  assign n33507 = ~x32 & n33506 ;
  assign n33508 = x32 & ~n33506 ;
  assign n33509 = n33507 | n33508 ;
  assign n33510 = n33171 | n33509 ;
  assign n33511 = ~n33509 & n33510 ;
  assign n33512 = ( ~n33171 & n33510 ) | ( ~n33171 & n33511 ) | ( n33510 & n33511 ) ;
  assign n33513 = n33498 & ~n33512 ;
  assign n33514 = n33499 | n33510 ;
  assign n33515 = n33171 & n33172 ;
  assign n33516 = ( n33171 & ~n33174 ) | ( n33171 & n33515 ) | ( ~n33174 & n33515 ) ;
  assign n33517 = ( n33511 & n33514 ) | ( n33511 & ~n33516 ) | ( n33514 & ~n33516 ) ;
  assign n33518 = ( n32928 & n33513 ) | ( n32928 & ~n33517 ) | ( n33513 & ~n33517 ) ;
  assign n33519 = ( n32906 & ~n33513 ) | ( n32906 & n33517 ) | ( ~n33513 & n33517 ) ;
  assign n33520 = ( n32922 & n33518 ) | ( n32922 & ~n33519 ) | ( n33518 & ~n33519 ) ;
  assign n33521 = n33502 & ~n33520 ;
  assign n33522 = n33498 | n33512 ;
  assign n33523 = n33499 & ~n33510 ;
  assign n33524 = n33171 & n33499 ;
  assign n33525 = ( ~n33511 & n33523 ) | ( ~n33511 & n33524 ) | ( n33523 & n33524 ) ;
  assign n33526 = ( n32928 & n33522 ) | ( n32928 & ~n33525 ) | ( n33522 & ~n33525 ) ;
  assign n33527 = ( n32906 & ~n33522 ) | ( n32906 & n33525 ) | ( ~n33522 & n33525 ) ;
  assign n33528 = ( n32922 & n33526 ) | ( n32922 & ~n33527 ) | ( n33526 & ~n33527 ) ;
  assign n33529 = n33497 & n33528 ;
  assign n33530 = ~n33521 & n33529 ;
  assign n33531 = n33497 & ~n33530 ;
  assign n33532 = x103 & n15552 ;
  assign n33533 = x102 & n15547 ;
  assign n33534 = x101 & ~n15546 ;
  assign n33535 = n16123 & n33534 ;
  assign n33536 = n33533 | n33535 ;
  assign n33537 = n33532 | n33536 ;
  assign n33538 = n15555 | n33532 ;
  assign n33539 = n33536 | n33538 ;
  assign n33540 = ( n7529 & n33537 ) | ( n7529 & n33539 ) | ( n33537 & n33539 ) ;
  assign n33541 = x59 & n33539 ;
  assign n33542 = x59 & n33532 ;
  assign n33543 = ( x59 & n33536 ) | ( x59 & n33542 ) | ( n33536 & n33542 ) ;
  assign n33544 = ( n7529 & n33541 ) | ( n7529 & n33543 ) | ( n33541 & n33543 ) ;
  assign n33545 = x59 & ~n33543 ;
  assign n33546 = x59 & ~n33539 ;
  assign n33547 = ( ~n7529 & n33545 ) | ( ~n7529 & n33546 ) | ( n33545 & n33546 ) ;
  assign n33548 = ( n33540 & ~n33544 ) | ( n33540 & n33547 ) | ( ~n33544 & n33547 ) ;
  assign n33549 = n33530 & n33548 ;
  assign n33550 = ~n33528 & n33548 ;
  assign n33551 = ( n33521 & n33548 ) | ( n33521 & n33550 ) | ( n33548 & n33550 ) ;
  assign n33552 = ( ~n33531 & n33549 ) | ( ~n33531 & n33551 ) | ( n33549 & n33551 ) ;
  assign n33553 = n33530 | n33548 ;
  assign n33554 = n33528 & ~n33548 ;
  assign n33555 = ~n33521 & n33554 ;
  assign n33556 = ( n33531 & ~n33553 ) | ( n33531 & n33555 ) | ( ~n33553 & n33555 ) ;
  assign n33557 = n33552 | n33556 ;
  assign n33558 = n33203 | n33223 ;
  assign n33559 = ( n33203 & ~n33206 ) | ( n33203 & n33558 ) | ( ~n33206 & n33558 ) ;
  assign n33560 = ~n33557 & n33559 ;
  assign n33561 = n33557 & ~n33559 ;
  assign n33562 = n33560 | n33561 ;
  assign n33563 = x106 & n14045 ;
  assign n33564 = x105 & n14040 ;
  assign n33565 = x104 & ~n14039 ;
  assign n33566 = n14552 & n33565 ;
  assign n33567 = n33564 | n33566 ;
  assign n33568 = n33563 | n33567 ;
  assign n33569 = n14048 | n33563 ;
  assign n33570 = n33567 | n33569 ;
  assign n33571 = ( n8656 & n33568 ) | ( n8656 & n33570 ) | ( n33568 & n33570 ) ;
  assign n33572 = x56 & n33570 ;
  assign n33573 = x56 & n33563 ;
  assign n33574 = ( x56 & n33567 ) | ( x56 & n33573 ) | ( n33567 & n33573 ) ;
  assign n33575 = ( n8656 & n33572 ) | ( n8656 & n33574 ) | ( n33572 & n33574 ) ;
  assign n33576 = x56 & ~n33574 ;
  assign n33577 = x56 & ~n33570 ;
  assign n33578 = ( ~n8656 & n33576 ) | ( ~n8656 & n33577 ) | ( n33576 & n33577 ) ;
  assign n33579 = ( n33571 & ~n33575 ) | ( n33571 & n33578 ) | ( ~n33575 & n33578 ) ;
  assign n33580 = ~n33562 & n33579 ;
  assign n33581 = n33562 | n33580 ;
  assign n33582 = n33562 & n33579 ;
  assign n33583 = n33581 & ~n33582 ;
  assign n33584 = n33226 & ~n33246 ;
  assign n33585 = ( n33164 & n33246 ) | ( n33164 & ~n33584 ) | ( n33246 & ~n33584 ) ;
  assign n33586 = ( n33227 & ~n33229 ) | ( n33227 & n33585 ) | ( ~n33229 & n33585 ) ;
  assign n33587 = n33583 & ~n33586 ;
  assign n33588 = ~n33583 & n33586 ;
  assign n33589 = n33587 | n33588 ;
  assign n33590 = x109 & n12574 ;
  assign n33591 = x108 & n12569 ;
  assign n33592 = x107 & ~n12568 ;
  assign n33593 = n13076 & n33592 ;
  assign n33594 = n33591 | n33593 ;
  assign n33595 = n33590 | n33594 ;
  assign n33596 = n12577 | n33590 ;
  assign n33597 = n33594 | n33596 ;
  assign n33598 = ( n9878 & n33595 ) | ( n9878 & n33597 ) | ( n33595 & n33597 ) ;
  assign n33599 = x53 & n33597 ;
  assign n33600 = x53 & n33590 ;
  assign n33601 = ( x53 & n33594 ) | ( x53 & n33600 ) | ( n33594 & n33600 ) ;
  assign n33602 = ( n9878 & n33599 ) | ( n9878 & n33601 ) | ( n33599 & n33601 ) ;
  assign n33603 = x53 & ~n33601 ;
  assign n33604 = x53 & ~n33597 ;
  assign n33605 = ( ~n9878 & n33603 ) | ( ~n9878 & n33604 ) | ( n33603 & n33604 ) ;
  assign n33606 = ( n33598 & ~n33602 ) | ( n33598 & n33605 ) | ( ~n33602 & n33605 ) ;
  assign n33607 = ~n33589 & n33606 ;
  assign n33608 = n33589 | n33607 ;
  assign n33610 = n33256 | n33275 ;
  assign n33611 = ( n33256 & ~n33258 ) | ( n33256 & n33610 ) | ( ~n33258 & n33610 ) ;
  assign n33609 = n33589 & n33606 ;
  assign n33612 = n33609 & n33611 ;
  assign n33613 = ( ~n33608 & n33611 ) | ( ~n33608 & n33612 ) | ( n33611 & n33612 ) ;
  assign n33614 = n33609 | n33611 ;
  assign n33615 = n33608 & ~n33614 ;
  assign n33616 = n33613 | n33615 ;
  assign n33617 = x112 & n11205 ;
  assign n33618 = x111 & n11200 ;
  assign n33619 = x110 & ~n11199 ;
  assign n33620 = n11679 & n33619 ;
  assign n33621 = n33618 | n33620 ;
  assign n33622 = n33617 | n33621 ;
  assign n33623 = n11208 | n33617 ;
  assign n33624 = n33621 | n33623 ;
  assign n33625 = ( n11172 & n33622 ) | ( n11172 & n33624 ) | ( n33622 & n33624 ) ;
  assign n33626 = x50 & n33624 ;
  assign n33627 = x50 & n33617 ;
  assign n33628 = ( x50 & n33621 ) | ( x50 & n33627 ) | ( n33621 & n33627 ) ;
  assign n33629 = ( n11172 & n33626 ) | ( n11172 & n33628 ) | ( n33626 & n33628 ) ;
  assign n33630 = x50 & ~n33628 ;
  assign n33631 = x50 & ~n33624 ;
  assign n33632 = ( ~n11172 & n33630 ) | ( ~n11172 & n33631 ) | ( n33630 & n33631 ) ;
  assign n33633 = ( n33625 & ~n33629 ) | ( n33625 & n33632 ) | ( ~n33629 & n33632 ) ;
  assign n33634 = ~n33616 & n33633 ;
  assign n33635 = n33616 | n33634 ;
  assign n33637 = n33280 | n33300 ;
  assign n33638 = ( ~n33278 & n33300 ) | ( ~n33278 & n33637 ) | ( n33300 & n33637 ) ;
  assign n33639 = ( n33281 & ~n33283 ) | ( n33281 & n33638 ) | ( ~n33283 & n33638 ) ;
  assign n33636 = n33616 & n33633 ;
  assign n33640 = n33636 & n33639 ;
  assign n33641 = ( ~n33635 & n33639 ) | ( ~n33635 & n33640 ) | ( n33639 & n33640 ) ;
  assign n33642 = n33636 | n33639 ;
  assign n33643 = n33635 & ~n33642 ;
  assign n33644 = n33641 | n33643 ;
  assign n33645 = x115 & n9933 ;
  assign n33646 = x114 & n9928 ;
  assign n33647 = x113 & ~n9927 ;
  assign n33648 = n10379 & n33647 ;
  assign n33649 = n33646 | n33648 ;
  assign n33650 = n33645 | n33649 ;
  assign n33651 = n9936 | n33645 ;
  assign n33652 = n33649 | n33651 ;
  assign n33653 = ( ~n12550 & n33650 ) | ( ~n12550 & n33652 ) | ( n33650 & n33652 ) ;
  assign n33654 = n33650 & n33652 ;
  assign n33655 = ( n12532 & n33653 ) | ( n12532 & n33654 ) | ( n33653 & n33654 ) ;
  assign n33656 = x47 & n33655 ;
  assign n33657 = x47 & ~n33655 ;
  assign n33658 = ( n33655 & ~n33656 ) | ( n33655 & n33657 ) | ( ~n33656 & n33657 ) ;
  assign n33659 = ~n33644 & n33658 ;
  assign n33660 = n33644 & ~n33658 ;
  assign n33661 = n33659 | n33660 ;
  assign n33662 = n33304 | n33321 ;
  assign n33663 = ( ~n33303 & n33321 ) | ( ~n33303 & n33662 ) | ( n33321 & n33662 ) ;
  assign n33664 = ( n33306 & ~n33307 ) | ( n33306 & n33663 ) | ( ~n33307 & n33663 ) ;
  assign n33665 = ~n33661 & n33664 ;
  assign n33666 = n33661 | n33665 ;
  assign n33667 = x118 & n8724 ;
  assign n33668 = x117 & n8719 ;
  assign n33669 = x116 & ~n8718 ;
  assign n33670 = n9149 & n33669 ;
  assign n33671 = n33668 | n33670 ;
  assign n33672 = n33667 | n33671 ;
  assign n33673 = n8727 | n33667 ;
  assign n33674 = n33671 | n33673 ;
  assign n33675 = ( ~n14002 & n33672 ) | ( ~n14002 & n33674 ) | ( n33672 & n33674 ) ;
  assign n33676 = n33672 & n33674 ;
  assign n33677 = ( n13981 & n33675 ) | ( n13981 & n33676 ) | ( n33675 & n33676 ) ;
  assign n33678 = x44 & n33677 ;
  assign n33679 = x44 & ~n33677 ;
  assign n33680 = ( n33677 & ~n33678 ) | ( n33677 & n33679 ) | ( ~n33678 & n33679 ) ;
  assign n33681 = n33664 & n33680 ;
  assign n33682 = n33661 & n33681 ;
  assign n33683 = ( ~n33666 & n33680 ) | ( ~n33666 & n33682 ) | ( n33680 & n33682 ) ;
  assign n33684 = n33664 | n33680 ;
  assign n33685 = ( n33661 & n33680 ) | ( n33661 & n33684 ) | ( n33680 & n33684 ) ;
  assign n33686 = n33666 & ~n33685 ;
  assign n33687 = n33683 | n33686 ;
  assign n33688 = n33480 & ~n33687 ;
  assign n33689 = ~n33480 & n33687 ;
  assign n33690 = n33688 | n33689 ;
  assign n33691 = x121 & n7566 ;
  assign n33692 = x120 & n7561 ;
  assign n33693 = x119 & ~n7560 ;
  assign n33694 = n7953 & n33693 ;
  assign n33695 = n33692 | n33694 ;
  assign n33696 = n33691 | n33695 ;
  assign n33697 = n7569 | n33691 ;
  assign n33698 = n33695 | n33697 ;
  assign n33699 = ( n15501 & n33696 ) | ( n15501 & n33698 ) | ( n33696 & n33698 ) ;
  assign n33700 = x41 & n33698 ;
  assign n33701 = x41 & n33691 ;
  assign n33702 = ( x41 & n33695 ) | ( x41 & n33701 ) | ( n33695 & n33701 ) ;
  assign n33703 = ( n15501 & n33700 ) | ( n15501 & n33702 ) | ( n33700 & n33702 ) ;
  assign n33704 = x41 & ~n33702 ;
  assign n33705 = x41 & ~n33698 ;
  assign n33706 = ( ~n15501 & n33704 ) | ( ~n15501 & n33705 ) | ( n33704 & n33705 ) ;
  assign n33707 = ( n33699 & ~n33703 ) | ( n33699 & n33706 ) | ( ~n33703 & n33706 ) ;
  assign n33708 = ~n33690 & n33707 ;
  assign n33709 = n33690 | n33708 ;
  assign n33711 = n33349 | n33371 ;
  assign n33712 = n33347 & ~n33371 ;
  assign n33713 = ( n33350 & n33711 ) | ( n33350 & ~n33712 ) | ( n33711 & ~n33712 ) ;
  assign n33714 = ( n33351 & ~n33354 ) | ( n33351 & n33713 ) | ( ~n33354 & n33713 ) ;
  assign n33710 = n33690 & n33707 ;
  assign n33715 = n33710 & n33714 ;
  assign n33716 = ( ~n33709 & n33714 ) | ( ~n33709 & n33715 ) | ( n33714 & n33715 ) ;
  assign n33717 = n33710 | n33714 ;
  assign n33718 = n33709 & ~n33717 ;
  assign n33719 = n33716 | n33718 ;
  assign n33720 = x124 & n6536 ;
  assign n33721 = x123 & n6531 ;
  assign n33722 = x122 & ~n6530 ;
  assign n33723 = n6871 & n33722 ;
  assign n33724 = n33721 | n33723 ;
  assign n33725 = n33720 | n33724 ;
  assign n33726 = n6539 | n33720 ;
  assign n33727 = n33724 | n33726 ;
  assign n33728 = ( n17084 & n33725 ) | ( n17084 & n33727 ) | ( n33725 & n33727 ) ;
  assign n33729 = x38 & n33727 ;
  assign n33730 = x38 & n33720 ;
  assign n33731 = ( x38 & n33724 ) | ( x38 & n33730 ) | ( n33724 & n33730 ) ;
  assign n33732 = ( n17084 & n33729 ) | ( n17084 & n33731 ) | ( n33729 & n33731 ) ;
  assign n33733 = x38 & ~n33731 ;
  assign n33734 = x38 & ~n33727 ;
  assign n33735 = ( ~n17084 & n33733 ) | ( ~n17084 & n33734 ) | ( n33733 & n33734 ) ;
  assign n33736 = ( n33728 & ~n33732 ) | ( n33728 & n33735 ) | ( ~n33732 & n33735 ) ;
  assign n33737 = ~n33719 & n33736 ;
  assign n33738 = n33719 | n33737 ;
  assign n33739 = n33375 | n33395 ;
  assign n33740 = ( ~n33374 & n33395 ) | ( ~n33374 & n33739 ) | ( n33395 & n33739 ) ;
  assign n33741 = ( n33376 & ~n33378 ) | ( n33376 & n33740 ) | ( ~n33378 & n33740 ) ;
  assign n33742 = n33719 & n33736 ;
  assign n33743 = n33741 & n33742 ;
  assign n33744 = ( ~n33738 & n33741 ) | ( ~n33738 & n33743 ) | ( n33741 & n33743 ) ;
  assign n33745 = n33741 | n33742 ;
  assign n33746 = n33738 & ~n33745 ;
  assign n33747 = n33744 | n33746 ;
  assign n33765 = ( n33402 & ~n33403 ) | ( n33402 & n33423 ) | ( ~n33403 & n33423 ) ;
  assign n33748 = x127 & n5554 ;
  assign n33749 = x126 & n5549 ;
  assign n33750 = x125 & ~n5548 ;
  assign n33751 = n5893 & n33750 ;
  assign n33752 = n33749 | n33751 ;
  assign n33753 = n33748 | n33752 ;
  assign n33754 = n5557 | n33748 ;
  assign n33755 = n33752 | n33754 ;
  assign n33756 = ( n18763 & n33753 ) | ( n18763 & n33755 ) | ( n33753 & n33755 ) ;
  assign n33757 = x35 & n33755 ;
  assign n33758 = x35 & n33748 ;
  assign n33759 = ( x35 & n33752 ) | ( x35 & n33758 ) | ( n33752 & n33758 ) ;
  assign n33760 = ( n18763 & n33757 ) | ( n18763 & n33759 ) | ( n33757 & n33759 ) ;
  assign n33761 = x35 & ~n33759 ;
  assign n33762 = x35 & ~n33755 ;
  assign n33763 = ( ~n18763 & n33761 ) | ( ~n18763 & n33762 ) | ( n33761 & n33762 ) ;
  assign n33764 = ( n33756 & ~n33760 ) | ( n33756 & n33763 ) | ( ~n33760 & n33763 ) ;
  assign n33766 = n33764 & n33765 ;
  assign n33767 = n33765 & ~n33766 ;
  assign n33768 = ~n33747 & n33764 ;
  assign n33769 = ~n33765 & n33768 ;
  assign n33770 = ( ~n33747 & n33767 ) | ( ~n33747 & n33769 ) | ( n33767 & n33769 ) ;
  assign n33771 = n33747 & ~n33764 ;
  assign n33772 = ( n33747 & n33765 ) | ( n33747 & n33771 ) | ( n33765 & n33771 ) ;
  assign n33773 = ~n33767 & n33772 ;
  assign n33774 = n33770 | n33773 ;
  assign n33775 = n33443 & n33445 ;
  assign n33776 = n33445 & ~n33775 ;
  assign n33777 = n33443 & ~n33445 ;
  assign n33778 = n33425 | n33777 ;
  assign n33779 = n33776 | n33778 ;
  assign n33780 = ( ~n33425 & n33775 ) | ( ~n33425 & n33779 ) | ( n33775 & n33779 ) ;
  assign n33781 = ~n33774 & n33780 ;
  assign n33782 = n33774 & ~n33780 ;
  assign n33783 = n33781 | n33782 ;
  assign n33784 = ~n33455 & n33472 ;
  assign n33785 = ~n33455 & n33457 ;
  assign n33786 = ( ~n33455 & n33459 ) | ( ~n33455 & n33785 ) | ( n33459 & n33785 ) ;
  assign n33787 = ( n33455 & n33462 ) | ( n33455 & ~n33785 ) | ( n33462 & ~n33785 ) ;
  assign n33788 = ( n32844 & n33786 ) | ( n32844 & ~n33787 ) | ( n33786 & ~n33787 ) ;
  assign n33789 = ( ~n30754 & n33784 ) | ( ~n30754 & n33788 ) | ( n33784 & n33788 ) ;
  assign n33790 = n33783 & n33789 ;
  assign n33791 = n33455 & ~n33783 ;
  assign n33792 = n33783 | n33785 ;
  assign n33793 = ( n33459 & ~n33791 ) | ( n33459 & n33792 ) | ( ~n33791 & n33792 ) ;
  assign n33794 = ( n33462 & n33791 ) | ( n33462 & ~n33792 ) | ( n33791 & ~n33792 ) ;
  assign n33795 = ( n32844 & n33793 ) | ( n32844 & ~n33794 ) | ( n33793 & ~n33794 ) ;
  assign n33796 = ( n33472 & n33783 ) | ( n33472 & ~n33791 ) | ( n33783 & ~n33791 ) ;
  assign n33797 = ( ~n30754 & n33795 ) | ( ~n30754 & n33796 ) | ( n33795 & n33796 ) ;
  assign n33798 = ~n33790 & n33797 ;
  assign n33799 = ~n33781 & n33792 ;
  assign n33800 = n33455 | n33781 ;
  assign n33801 = ( n33781 & ~n33783 ) | ( n33781 & n33800 ) | ( ~n33783 & n33800 ) ;
  assign n33802 = ( n33459 & n33799 ) | ( n33459 & ~n33801 ) | ( n33799 & ~n33801 ) ;
  assign n33803 = ( n33462 & ~n33799 ) | ( n33462 & n33801 ) | ( ~n33799 & n33801 ) ;
  assign n33804 = ( n32844 & n33802 ) | ( n32844 & ~n33803 ) | ( n33802 & ~n33803 ) ;
  assign n33805 = ~n33781 & n33783 ;
  assign n33806 = ( n33472 & ~n33801 ) | ( n33472 & n33805 ) | ( ~n33801 & n33805 ) ;
  assign n33807 = ( ~n30754 & n33804 ) | ( ~n30754 & n33806 ) | ( n33804 & n33806 ) ;
  assign n33808 = x125 & n6536 ;
  assign n33809 = x124 & n6531 ;
  assign n33810 = x123 & ~n6530 ;
  assign n33811 = n6871 & n33810 ;
  assign n33812 = n33809 | n33811 ;
  assign n33813 = n33808 | n33812 ;
  assign n33814 = n6539 | n33808 ;
  assign n33815 = n33812 | n33814 ;
  assign n33816 = ( n17670 & n33813 ) | ( n17670 & n33815 ) | ( n33813 & n33815 ) ;
  assign n33817 = x38 & n33815 ;
  assign n33818 = x38 & n33808 ;
  assign n33819 = ( x38 & n33812 ) | ( x38 & n33818 ) | ( n33812 & n33818 ) ;
  assign n33820 = ( n17670 & n33817 ) | ( n17670 & n33819 ) | ( n33817 & n33819 ) ;
  assign n33821 = x38 & ~n33819 ;
  assign n33822 = x38 & ~n33815 ;
  assign n33823 = ( ~n17670 & n33821 ) | ( ~n17670 & n33822 ) | ( n33821 & n33822 ) ;
  assign n33824 = ( n33816 & ~n33820 ) | ( n33816 & n33823 ) | ( ~n33820 & n33823 ) ;
  assign n33825 = x127 & n5549 ;
  assign n33826 = x126 & ~n5548 ;
  assign n33827 = n5893 & n33826 ;
  assign n33828 = n33825 | n33827 ;
  assign n33829 = n5557 | n33828 ;
  assign n33830 = ( n19328 & n33828 ) | ( n19328 & n33829 ) | ( n33828 & n33829 ) ;
  assign n33831 = x35 & n33828 ;
  assign n33832 = ( x35 & n8000 ) | ( x35 & n33828 ) | ( n8000 & n33828 ) ;
  assign n33833 = ( n19328 & n33831 ) | ( n19328 & n33832 ) | ( n33831 & n33832 ) ;
  assign n33834 = x35 & ~n8000 ;
  assign n33835 = ~n33828 & n33834 ;
  assign n33836 = x35 & ~n33828 ;
  assign n33837 = ( ~n19328 & n33835 ) | ( ~n19328 & n33836 ) | ( n33835 & n33836 ) ;
  assign n33838 = ( n33830 & ~n33833 ) | ( n33830 & n33837 ) | ( ~n33833 & n33837 ) ;
  assign n33839 = n33736 & n33838 ;
  assign n33840 = ~n33719 & n33839 ;
  assign n33841 = ( n33744 & n33838 ) | ( n33744 & n33840 ) | ( n33838 & n33840 ) ;
  assign n33842 = n33736 | n33838 ;
  assign n33843 = ( ~n33719 & n33838 ) | ( ~n33719 & n33842 ) | ( n33838 & n33842 ) ;
  assign n33844 = n33744 | n33843 ;
  assign n33845 = ~n33841 & n33844 ;
  assign n33846 = n33634 | n33641 ;
  assign n33847 = x98 & n18290 ;
  assign n33848 = x63 & x97 ;
  assign n33849 = ~n18290 & n33848 ;
  assign n33850 = n33847 | n33849 ;
  assign n33851 = n33171 | n33507 ;
  assign n33852 = ( n33507 & ~n33509 ) | ( n33507 & n33851 ) | ( ~n33509 & n33851 ) ;
  assign n33853 = n33850 & ~n33852 ;
  assign n33854 = ~n33850 & n33852 ;
  assign n33855 = n33853 | n33854 ;
  assign n33856 = x100 & n17141 ;
  assign n33857 = x99 & ~n17140 ;
  assign n33858 = n17724 & n33857 ;
  assign n33859 = n33856 | n33858 ;
  assign n33860 = x101 & n17146 ;
  assign n33861 = n17149 | n33860 ;
  assign n33862 = n33859 | n33861 ;
  assign n33863 = x62 & ~n33862 ;
  assign n33864 = ~n33855 & n33863 ;
  assign n33865 = x62 & x101 ;
  assign n33866 = n17146 & n33865 ;
  assign n33867 = x62 & ~n33866 ;
  assign n33868 = ~n33859 & n33867 ;
  assign n33869 = ~n33855 & n33868 ;
  assign n33870 = ( ~n6844 & n33864 ) | ( ~n6844 & n33869 ) | ( n33864 & n33869 ) ;
  assign n33871 = ~x62 & n33862 ;
  assign n33872 = ~x62 & n33860 ;
  assign n33873 = ( ~x62 & n33859 ) | ( ~x62 & n33872 ) | ( n33859 & n33872 ) ;
  assign n33874 = ( n6844 & n33871 ) | ( n6844 & n33873 ) | ( n33871 & n33873 ) ;
  assign n33875 = ( ~n33855 & n33870 ) | ( ~n33855 & n33874 ) | ( n33870 & n33874 ) ;
  assign n33876 = n33855 & ~n33863 ;
  assign n33877 = n33855 & ~n33868 ;
  assign n33878 = ( n6844 & n33876 ) | ( n6844 & n33877 ) | ( n33876 & n33877 ) ;
  assign n33879 = ~n33874 & n33878 ;
  assign n33880 = n33875 | n33879 ;
  assign n33881 = n33497 & ~n33528 ;
  assign n33882 = ( n33497 & n33521 ) | ( n33497 & n33881 ) | ( n33521 & n33881 ) ;
  assign n33884 = x104 & n15552 ;
  assign n33885 = x103 & n15547 ;
  assign n33886 = x102 & ~n15546 ;
  assign n33887 = n16123 & n33886 ;
  assign n33888 = n33885 | n33887 ;
  assign n33889 = n33884 | n33888 ;
  assign n33890 = n15555 | n33884 ;
  assign n33891 = n33888 | n33890 ;
  assign n33892 = ( n7911 & n33889 ) | ( n7911 & n33891 ) | ( n33889 & n33891 ) ;
  assign n33893 = x59 & n33891 ;
  assign n33894 = x59 & n33884 ;
  assign n33895 = ( x59 & n33888 ) | ( x59 & n33894 ) | ( n33888 & n33894 ) ;
  assign n33896 = ( n7911 & n33893 ) | ( n7911 & n33895 ) | ( n33893 & n33895 ) ;
  assign n33897 = x59 & ~n33895 ;
  assign n33898 = x59 & ~n33891 ;
  assign n33899 = ( ~n7911 & n33897 ) | ( ~n7911 & n33898 ) | ( n33897 & n33898 ) ;
  assign n33900 = ( n33892 & ~n33896 ) | ( n33892 & n33899 ) | ( ~n33896 & n33899 ) ;
  assign n33901 = ( ~n33520 & n33880 ) | ( ~n33520 & n33900 ) | ( n33880 & n33900 ) ;
  assign n33902 = n33880 & n33900 ;
  assign n33903 = ( ~n33882 & n33901 ) | ( ~n33882 & n33902 ) | ( n33901 & n33902 ) ;
  assign n33883 = n33520 | n33882 ;
  assign n33904 = ( n33883 & ~n33900 ) | ( n33883 & n33903 ) | ( ~n33900 & n33903 ) ;
  assign n33905 = ( ~n33880 & n33903 ) | ( ~n33880 & n33904 ) | ( n33903 & n33904 ) ;
  assign n33906 = n33552 | n33559 ;
  assign n33907 = ( n33552 & ~n33557 ) | ( n33552 & n33906 ) | ( ~n33557 & n33906 ) ;
  assign n33908 = ~n33905 & n33907 ;
  assign n33909 = n33905 & ~n33907 ;
  assign n33910 = n33908 | n33909 ;
  assign n33911 = x107 & n14045 ;
  assign n33912 = x106 & n14040 ;
  assign n33913 = x105 & ~n14039 ;
  assign n33914 = n14552 & n33913 ;
  assign n33915 = n33912 | n33914 ;
  assign n33916 = n33911 | n33915 ;
  assign n33917 = n14048 | n33911 ;
  assign n33918 = n33915 | n33917 ;
  assign n33919 = ( n9084 & n33916 ) | ( n9084 & n33918 ) | ( n33916 & n33918 ) ;
  assign n33920 = x56 & n33918 ;
  assign n33921 = x56 & n33911 ;
  assign n33922 = ( x56 & n33915 ) | ( x56 & n33921 ) | ( n33915 & n33921 ) ;
  assign n33923 = ( n9084 & n33920 ) | ( n9084 & n33922 ) | ( n33920 & n33922 ) ;
  assign n33924 = x56 & ~n33922 ;
  assign n33925 = x56 & ~n33918 ;
  assign n33926 = ( ~n9084 & n33924 ) | ( ~n9084 & n33925 ) | ( n33924 & n33925 ) ;
  assign n33927 = ( n33919 & ~n33923 ) | ( n33919 & n33926 ) | ( ~n33923 & n33926 ) ;
  assign n33928 = n33910 | n33927 ;
  assign n33929 = n33910 & ~n33927 ;
  assign n33930 = ( ~n33910 & n33928 ) | ( ~n33910 & n33929 ) | ( n33928 & n33929 ) ;
  assign n33931 = n33580 | n33586 ;
  assign n33932 = ( n33580 & ~n33583 ) | ( n33580 & n33931 ) | ( ~n33583 & n33931 ) ;
  assign n33933 = n33930 & ~n33932 ;
  assign n33934 = ~n33930 & n33932 ;
  assign n33935 = n33933 | n33934 ;
  assign n33936 = x110 & n12574 ;
  assign n33937 = x109 & n12569 ;
  assign n33938 = x108 & ~n12568 ;
  assign n33939 = n13076 & n33938 ;
  assign n33940 = n33937 | n33939 ;
  assign n33941 = n33936 | n33940 ;
  assign n33942 = n12577 | n33936 ;
  assign n33943 = n33940 | n33942 ;
  assign n33944 = ( n10330 & n33941 ) | ( n10330 & n33943 ) | ( n33941 & n33943 ) ;
  assign n33945 = x53 & n33943 ;
  assign n33946 = x53 & n33936 ;
  assign n33947 = ( x53 & n33940 ) | ( x53 & n33946 ) | ( n33940 & n33946 ) ;
  assign n33948 = ( n10330 & n33945 ) | ( n10330 & n33947 ) | ( n33945 & n33947 ) ;
  assign n33949 = x53 & ~n33947 ;
  assign n33950 = x53 & ~n33943 ;
  assign n33951 = ( ~n10330 & n33949 ) | ( ~n10330 & n33950 ) | ( n33949 & n33950 ) ;
  assign n33952 = ( n33944 & ~n33948 ) | ( n33944 & n33951 ) | ( ~n33948 & n33951 ) ;
  assign n33953 = n33935 & n33952 ;
  assign n33954 = n33930 & ~n33952 ;
  assign n33955 = ( n33932 & n33952 ) | ( n33932 & ~n33954 ) | ( n33952 & ~n33954 ) ;
  assign n33956 = n33933 | n33955 ;
  assign n33957 = ~n33953 & n33956 ;
  assign n33958 = n33607 | n33613 ;
  assign n33959 = n33957 & ~n33958 ;
  assign n33960 = ~n33957 & n33958 ;
  assign n33961 = n33959 | n33960 ;
  assign n33962 = x113 & n11205 ;
  assign n33963 = x112 & n11200 ;
  assign n33964 = x111 & ~n11199 ;
  assign n33965 = n11679 & n33964 ;
  assign n33966 = n33963 | n33965 ;
  assign n33967 = n33962 | n33966 ;
  assign n33968 = n11208 | n33962 ;
  assign n33969 = n33966 | n33968 ;
  assign n33970 = ( ~n11642 & n33967 ) | ( ~n11642 & n33969 ) | ( n33967 & n33969 ) ;
  assign n33971 = n33967 & n33969 ;
  assign n33972 = ( n11626 & n33970 ) | ( n11626 & n33971 ) | ( n33970 & n33971 ) ;
  assign n33973 = x50 & n33972 ;
  assign n33974 = x50 & ~n33972 ;
  assign n33975 = ( n33972 & ~n33973 ) | ( n33972 & n33974 ) | ( ~n33973 & n33974 ) ;
  assign n33976 = n33961 & n33975 ;
  assign n33977 = n33846 & n33976 ;
  assign n33978 = n33956 & ~n33975 ;
  assign n33979 = ~n33953 & n33978 ;
  assign n33980 = ( n33958 & n33975 ) | ( n33958 & ~n33979 ) | ( n33975 & ~n33979 ) ;
  assign n33981 = n33959 | n33980 ;
  assign n33982 = ( n33846 & n33977 ) | ( n33846 & ~n33981 ) | ( n33977 & ~n33981 ) ;
  assign n33983 = ~n33976 & n33981 ;
  assign n33984 = ~n33846 & n33983 ;
  assign n33985 = n33982 | n33984 ;
  assign n33986 = x116 & n9933 ;
  assign n33987 = x115 & n9928 ;
  assign n33988 = x114 & ~n9927 ;
  assign n33989 = n10379 & n33988 ;
  assign n33990 = n33987 | n33989 ;
  assign n33991 = n33986 | n33990 ;
  assign n33992 = n9936 | n33986 ;
  assign n33993 = n33990 | n33992 ;
  assign n33994 = ( ~n13040 & n33991 ) | ( ~n13040 & n33993 ) | ( n33991 & n33993 ) ;
  assign n33995 = n33991 & n33993 ;
  assign n33996 = ( n13022 & n33994 ) | ( n13022 & n33995 ) | ( n33994 & n33995 ) ;
  assign n33997 = x47 & n33996 ;
  assign n33998 = x47 & ~n33996 ;
  assign n33999 = ( n33996 & ~n33997 ) | ( n33996 & n33998 ) | ( ~n33997 & n33998 ) ;
  assign n34000 = n33659 | n33664 ;
  assign n34001 = ( n33659 & ~n33661 ) | ( n33659 & n34000 ) | ( ~n33661 & n34000 ) ;
  assign n34002 = ( n33985 & ~n33999 ) | ( n33985 & n34001 ) | ( ~n33999 & n34001 ) ;
  assign n34003 = ( ~n33985 & n33999 ) | ( ~n33985 & n34002 ) | ( n33999 & n34002 ) ;
  assign n34004 = x119 & n8724 ;
  assign n34005 = x118 & n8719 ;
  assign n34006 = x117 & ~n8718 ;
  assign n34007 = n9149 & n34006 ;
  assign n34008 = n34005 | n34007 ;
  assign n34009 = n34004 | n34008 ;
  assign n34010 = n8727 | n34004 ;
  assign n34011 = n34008 | n34010 ;
  assign n34012 = ( n14496 & n34009 ) | ( n14496 & n34011 ) | ( n34009 & n34011 ) ;
  assign n34013 = x44 & n34011 ;
  assign n34014 = x44 & n34004 ;
  assign n34015 = ( x44 & n34008 ) | ( x44 & n34014 ) | ( n34008 & n34014 ) ;
  assign n34016 = ( n14496 & n34013 ) | ( n14496 & n34015 ) | ( n34013 & n34015 ) ;
  assign n34017 = x44 & ~n34015 ;
  assign n34018 = x44 & ~n34011 ;
  assign n34019 = ( ~n14496 & n34017 ) | ( ~n14496 & n34018 ) | ( n34017 & n34018 ) ;
  assign n34020 = ( n34012 & ~n34016 ) | ( n34012 & n34019 ) | ( ~n34016 & n34019 ) ;
  assign n34021 = ~n34002 & n34020 ;
  assign n34022 = n34001 & n34020 ;
  assign n34023 = ( ~n34003 & n34021 ) | ( ~n34003 & n34022 ) | ( n34021 & n34022 ) ;
  assign n34024 = n34002 & ~n34020 ;
  assign n34025 = n34001 | n34020 ;
  assign n34026 = ( n34003 & n34024 ) | ( n34003 & ~n34025 ) | ( n34024 & ~n34025 ) ;
  assign n34027 = n34023 | n34026 ;
  assign n34028 = n33683 | n33688 ;
  assign n34029 = ~n34027 & n34028 ;
  assign n34030 = n34027 & ~n34028 ;
  assign n34031 = n34029 | n34030 ;
  assign n34032 = x122 & n7566 ;
  assign n34033 = x121 & n7561 ;
  assign n34034 = x120 & ~n7560 ;
  assign n34035 = n7953 & n34034 ;
  assign n34036 = n34033 | n34035 ;
  assign n34037 = n34032 | n34036 ;
  assign n34038 = n7569 | n34032 ;
  assign n34039 = n34036 | n34038 ;
  assign n34040 = ( n16043 & n34037 ) | ( n16043 & n34039 ) | ( n34037 & n34039 ) ;
  assign n34041 = x41 & n34039 ;
  assign n34042 = x41 & n34032 ;
  assign n34043 = ( x41 & n34036 ) | ( x41 & n34042 ) | ( n34036 & n34042 ) ;
  assign n34044 = ( n16043 & n34041 ) | ( n16043 & n34043 ) | ( n34041 & n34043 ) ;
  assign n34045 = x41 & ~n34043 ;
  assign n34046 = x41 & ~n34039 ;
  assign n34047 = ( ~n16043 & n34045 ) | ( ~n16043 & n34046 ) | ( n34045 & n34046 ) ;
  assign n34048 = ( n34040 & ~n34044 ) | ( n34040 & n34047 ) | ( ~n34044 & n34047 ) ;
  assign n34049 = n34031 | n34048 ;
  assign n34050 = n34031 & ~n34048 ;
  assign n34051 = ( ~n34031 & n34049 ) | ( ~n34031 & n34050 ) | ( n34049 & n34050 ) ;
  assign n34052 = n33708 | n33714 ;
  assign n34053 = ~n33708 & n33709 ;
  assign n34054 = ( n33715 & n34052 ) | ( n33715 & ~n34053 ) | ( n34052 & ~n34053 ) ;
  assign n34055 = n34051 & ~n34054 ;
  assign n34056 = ~n34051 & n34054 ;
  assign n34057 = n34055 | n34056 ;
  assign n34058 = ( n33824 & n33845 ) | ( n33824 & ~n34057 ) | ( n33845 & ~n34057 ) ;
  assign n34059 = ( ~n33845 & n34057 ) | ( ~n33845 & n34058 ) | ( n34057 & n34058 ) ;
  assign n34060 = ( ~n33824 & n34058 ) | ( ~n33824 & n34059 ) | ( n34058 & n34059 ) ;
  assign n34061 = n33766 | n33769 ;
  assign n34062 = ( n33747 & ~n33765 ) | ( n33747 & n33771 ) | ( ~n33765 & n33771 ) ;
  assign n34063 = ( n33767 & n34061 ) | ( n33767 & ~n34062 ) | ( n34061 & ~n34062 ) ;
  assign n34064 = ~n34060 & n34063 ;
  assign n34065 = n34060 & ~n34063 ;
  assign n34066 = n34064 | n34065 ;
  assign n34067 = n33807 & n34066 ;
  assign n34068 = n33803 & ~n34066 ;
  assign n34069 = n33801 & ~n34066 ;
  assign n34070 = n33799 | n34066 ;
  assign n34071 = ( n33459 & ~n34069 ) | ( n33459 & n34070 ) | ( ~n34069 & n34070 ) ;
  assign n34072 = ( n32844 & ~n34068 ) | ( n32844 & n34071 ) | ( ~n34068 & n34071 ) ;
  assign n34073 = n33781 & ~n34066 ;
  assign n34074 = ( n33783 & n34066 ) | ( n33783 & ~n34073 ) | ( n34066 & ~n34073 ) ;
  assign n34075 = ( n33472 & ~n34069 ) | ( n33472 & n34074 ) | ( ~n34069 & n34074 ) ;
  assign n34076 = ( ~n30754 & n34072 ) | ( ~n30754 & n34075 ) | ( n34072 & n34075 ) ;
  assign n34077 = ~n34067 & n34076 ;
  assign n34225 = ( n33960 & ~n33961 ) | ( n33960 & n33980 ) | ( ~n33961 & n33980 ) ;
  assign n34078 = n33854 | n33875 ;
  assign n34079 = x99 & n18290 ;
  assign n34080 = x63 & x98 ;
  assign n34081 = ~n18290 & n34080 ;
  assign n34082 = n34079 | n34081 ;
  assign n34083 = n33850 & ~n34082 ;
  assign n34084 = ~n33850 & n34082 ;
  assign n34085 = n34083 | n34084 ;
  assign n34086 = n33850 | n34085 ;
  assign n34087 = n33852 & ~n34086 ;
  assign n34088 = ( n33875 & ~n34085 ) | ( n33875 & n34087 ) | ( ~n34085 & n34087 ) ;
  assign n34089 = n34078 & ~n34088 ;
  assign n34090 = x102 & n17146 ;
  assign n34091 = x101 & n17141 ;
  assign n34092 = x100 & ~n17140 ;
  assign n34093 = n17724 & n34092 ;
  assign n34094 = n34091 | n34093 ;
  assign n34095 = n34090 | n34094 ;
  assign n34096 = n17149 | n34090 ;
  assign n34097 = n34094 | n34096 ;
  assign n34098 = ( n7178 & n34095 ) | ( n7178 & n34097 ) | ( n34095 & n34097 ) ;
  assign n34099 = x62 & n34097 ;
  assign n34100 = x62 & n34090 ;
  assign n34101 = ( x62 & n34094 ) | ( x62 & n34100 ) | ( n34094 & n34100 ) ;
  assign n34102 = ( n7178 & n34099 ) | ( n7178 & n34101 ) | ( n34099 & n34101 ) ;
  assign n34103 = x62 & ~n34101 ;
  assign n34104 = x62 & ~n34097 ;
  assign n34105 = ( ~n7178 & n34103 ) | ( ~n7178 & n34104 ) | ( n34103 & n34104 ) ;
  assign n34106 = ( n34098 & ~n34102 ) | ( n34098 & n34105 ) | ( ~n34102 & n34105 ) ;
  assign n34107 = n34085 | n34087 ;
  assign n34108 = n33875 | n34107 ;
  assign n34109 = n34106 & ~n34108 ;
  assign n34110 = ( n34089 & n34106 ) | ( n34089 & n34109 ) | ( n34106 & n34109 ) ;
  assign n34111 = ~n34106 & n34108 ;
  assign n34112 = ~n34089 & n34111 ;
  assign n34113 = n34110 | n34112 ;
  assign n34114 = x105 & n15552 ;
  assign n34115 = x104 & n15547 ;
  assign n34116 = x103 & ~n15546 ;
  assign n34117 = n16123 & n34116 ;
  assign n34118 = n34115 | n34117 ;
  assign n34119 = n34114 | n34118 ;
  assign n34120 = n15555 | n34114 ;
  assign n34121 = n34118 | n34120 ;
  assign n34122 = ( n8273 & n34119 ) | ( n8273 & n34121 ) | ( n34119 & n34121 ) ;
  assign n34123 = x59 & n34121 ;
  assign n34124 = x59 & n34114 ;
  assign n34125 = ( x59 & n34118 ) | ( x59 & n34124 ) | ( n34118 & n34124 ) ;
  assign n34126 = ( n8273 & n34123 ) | ( n8273 & n34125 ) | ( n34123 & n34125 ) ;
  assign n34127 = x59 & ~n34125 ;
  assign n34128 = x59 & ~n34121 ;
  assign n34129 = ( ~n8273 & n34127 ) | ( ~n8273 & n34128 ) | ( n34127 & n34128 ) ;
  assign n34130 = ( n34122 & ~n34126 ) | ( n34122 & n34129 ) | ( ~n34126 & n34129 ) ;
  assign n34131 = n34113 | n34130 ;
  assign n34132 = n34113 & n34130 ;
  assign n34133 = n34131 & ~n34132 ;
  assign n34134 = n33520 & ~n33880 ;
  assign n34135 = ( ~n33880 & n33882 ) | ( ~n33880 & n34134 ) | ( n33882 & n34134 ) ;
  assign n34136 = n33883 & ~n34135 ;
  assign n34137 = n33880 | n34135 ;
  assign n34138 = ~n34136 & n34137 ;
  assign n34139 = n33900 | n34135 ;
  assign n34140 = ( n34135 & ~n34138 ) | ( n34135 & n34139 ) | ( ~n34138 & n34139 ) ;
  assign n34141 = ~n34133 & n34140 ;
  assign n34142 = n34133 & ~n34140 ;
  assign n34143 = n34141 | n34142 ;
  assign n34144 = x108 & n14045 ;
  assign n34145 = x107 & n14040 ;
  assign n34146 = x106 & ~n14039 ;
  assign n34147 = n14552 & n34146 ;
  assign n34148 = n34145 | n34147 ;
  assign n34149 = n34144 | n34148 ;
  assign n34150 = n14048 | n34144 ;
  assign n34151 = n34148 | n34150 ;
  assign n34152 = ( n9479 & n34149 ) | ( n9479 & n34151 ) | ( n34149 & n34151 ) ;
  assign n34153 = x56 & n34151 ;
  assign n34154 = x56 & n34144 ;
  assign n34155 = ( x56 & n34148 ) | ( x56 & n34154 ) | ( n34148 & n34154 ) ;
  assign n34156 = ( n9479 & n34153 ) | ( n9479 & n34155 ) | ( n34153 & n34155 ) ;
  assign n34157 = x56 & ~n34155 ;
  assign n34158 = x56 & ~n34151 ;
  assign n34159 = ( ~n9479 & n34157 ) | ( ~n9479 & n34158 ) | ( n34157 & n34158 ) ;
  assign n34160 = ( n34152 & ~n34156 ) | ( n34152 & n34159 ) | ( ~n34156 & n34159 ) ;
  assign n34161 = ~n34143 & n34160 ;
  assign n34162 = n34143 & ~n34160 ;
  assign n34163 = n34161 | n34162 ;
  assign n34164 = n33905 & ~n33927 ;
  assign n34165 = ( n33907 & n33927 ) | ( n33907 & ~n34164 ) | ( n33927 & ~n34164 ) ;
  assign n34166 = ( n33908 & ~n33910 ) | ( n33908 & n34165 ) | ( ~n33910 & n34165 ) ;
  assign n34167 = ~n34163 & n34166 ;
  assign n34168 = n34163 & ~n34166 ;
  assign n34169 = n34167 | n34168 ;
  assign n34170 = x111 & n12574 ;
  assign n34171 = x110 & n12569 ;
  assign n34172 = x109 & ~n12568 ;
  assign n34173 = n13076 & n34172 ;
  assign n34174 = n34171 | n34173 ;
  assign n34175 = n34170 | n34174 ;
  assign n34176 = n12577 | n34170 ;
  assign n34177 = n34174 | n34176 ;
  assign n34178 = ( n10749 & n34175 ) | ( n10749 & n34177 ) | ( n34175 & n34177 ) ;
  assign n34179 = x53 & n34177 ;
  assign n34180 = x53 & n34170 ;
  assign n34181 = ( x53 & n34174 ) | ( x53 & n34180 ) | ( n34174 & n34180 ) ;
  assign n34182 = ( n10749 & n34179 ) | ( n10749 & n34181 ) | ( n34179 & n34181 ) ;
  assign n34183 = x53 & ~n34181 ;
  assign n34184 = x53 & ~n34177 ;
  assign n34185 = ( ~n10749 & n34183 ) | ( ~n10749 & n34184 ) | ( n34183 & n34184 ) ;
  assign n34186 = ( n34178 & ~n34182 ) | ( n34178 & n34185 ) | ( ~n34182 & n34185 ) ;
  assign n34187 = n34169 | n34186 ;
  assign n34188 = n34169 & ~n34186 ;
  assign n34189 = ( ~n34169 & n34187 ) | ( ~n34169 & n34188 ) | ( n34187 & n34188 ) ;
  assign n34190 = ( n33934 & ~n33935 ) | ( n33934 & n33955 ) | ( ~n33935 & n33955 ) ;
  assign n34191 = n34189 & ~n34190 ;
  assign n34192 = ~n34189 & n34190 ;
  assign n34193 = n34191 | n34192 ;
  assign n34194 = x114 & n11205 ;
  assign n34195 = x113 & n11200 ;
  assign n34196 = x112 & ~n11199 ;
  assign n34197 = n11679 & n34196 ;
  assign n34198 = n34195 | n34197 ;
  assign n34199 = n34194 | n34198 ;
  assign n34200 = n11208 | n34194 ;
  assign n34201 = n34198 | n34200 ;
  assign n34202 = ( ~n12095 & n34199 ) | ( ~n12095 & n34201 ) | ( n34199 & n34201 ) ;
  assign n34203 = n34199 & n34201 ;
  assign n34204 = ( n12079 & n34202 ) | ( n12079 & n34203 ) | ( n34202 & n34203 ) ;
  assign n34205 = x50 & n34204 ;
  assign n34206 = x50 & ~n34204 ;
  assign n34207 = ( n34204 & ~n34205 ) | ( n34204 & n34206 ) | ( ~n34205 & n34206 ) ;
  assign n34208 = n34193 & ~n34207 ;
  assign n34209 = ~n34193 & n34207 ;
  assign n34210 = n34208 | n34209 ;
  assign n34211 = x117 & n9933 ;
  assign n34212 = x116 & n9928 ;
  assign n34213 = x115 & ~n9927 ;
  assign n34214 = n10379 & n34213 ;
  assign n34215 = n34212 | n34214 ;
  assign n34216 = n34211 | n34215 ;
  assign n34217 = n9936 | n34211 ;
  assign n34218 = n34215 | n34217 ;
  assign n34219 = ( ~n13522 & n34216 ) | ( ~n13522 & n34218 ) | ( n34216 & n34218 ) ;
  assign n34220 = n34216 & n34218 ;
  assign n34221 = ( n13503 & n34219 ) | ( n13503 & n34220 ) | ( n34219 & n34220 ) ;
  assign n34222 = x47 & n34221 ;
  assign n34223 = x47 & ~n34221 ;
  assign n34224 = ( n34221 & ~n34222 ) | ( n34221 & n34223 ) | ( ~n34222 & n34223 ) ;
  assign n34226 = ( ~n34210 & n34224 ) | ( ~n34210 & n34225 ) | ( n34224 & n34225 ) ;
  assign n34227 = ( n34210 & ~n34224 ) | ( n34210 & n34225 ) | ( ~n34224 & n34225 ) ;
  assign n34228 = ( ~n34225 & n34226 ) | ( ~n34225 & n34227 ) | ( n34226 & n34227 ) ;
  assign n34229 = ~n33984 & n33999 ;
  assign n34230 = ~n33982 & n34229 ;
  assign n34231 = n33982 & ~n34228 ;
  assign n34232 = ( ~n34228 & n34230 ) | ( ~n34228 & n34231 ) | ( n34230 & n34231 ) ;
  assign n34233 = ~n33982 & n34228 ;
  assign n34234 = ~n34230 & n34233 ;
  assign n34235 = n34232 | n34234 ;
  assign n34236 = x120 & n8724 ;
  assign n34237 = x119 & n8719 ;
  assign n34238 = x118 & ~n8718 ;
  assign n34239 = n9149 & n34238 ;
  assign n34240 = n34237 | n34239 ;
  assign n34241 = n34236 | n34240 ;
  assign n34242 = n8727 | n34236 ;
  assign n34243 = n34240 | n34242 ;
  assign n34244 = ( n14991 & n34241 ) | ( n14991 & n34243 ) | ( n34241 & n34243 ) ;
  assign n34245 = x44 & n34243 ;
  assign n34246 = x44 & n34236 ;
  assign n34247 = ( x44 & n34240 ) | ( x44 & n34246 ) | ( n34240 & n34246 ) ;
  assign n34248 = ( n14991 & n34245 ) | ( n14991 & n34247 ) | ( n34245 & n34247 ) ;
  assign n34249 = x44 & ~n34247 ;
  assign n34250 = x44 & ~n34243 ;
  assign n34251 = ( ~n14991 & n34249 ) | ( ~n14991 & n34250 ) | ( n34249 & n34250 ) ;
  assign n34252 = ( n34244 & ~n34248 ) | ( n34244 & n34251 ) | ( ~n34248 & n34251 ) ;
  assign n34253 = ~n34235 & n34252 ;
  assign n34254 = n34235 & ~n34252 ;
  assign n34255 = n34253 | n34254 ;
  assign n34256 = n33985 | n34230 ;
  assign n34257 = n33984 & n33999 ;
  assign n34258 = ( n33982 & n33999 ) | ( n33982 & n34257 ) | ( n33999 & n34257 ) ;
  assign n34259 = n34001 & n34258 ;
  assign n34260 = ( n34001 & ~n34256 ) | ( n34001 & n34259 ) | ( ~n34256 & n34259 ) ;
  assign n34261 = n34023 | n34260 ;
  assign n34262 = ~n34255 & n34261 ;
  assign n34263 = n34255 & ~n34261 ;
  assign n34264 = n34262 | n34263 ;
  assign n34265 = x123 & n7566 ;
  assign n34266 = x122 & n7561 ;
  assign n34267 = x121 & ~n7560 ;
  assign n34268 = n7953 & n34267 ;
  assign n34269 = n34266 | n34268 ;
  assign n34270 = n34265 | n34269 ;
  assign n34271 = n7569 | n34265 ;
  assign n34272 = n34269 | n34271 ;
  assign n34273 = ( n16086 & n34270 ) | ( n16086 & n34272 ) | ( n34270 & n34272 ) ;
  assign n34274 = x41 & n34272 ;
  assign n34275 = x41 & n34265 ;
  assign n34276 = ( x41 & n34269 ) | ( x41 & n34275 ) | ( n34269 & n34275 ) ;
  assign n34277 = ( n16086 & n34274 ) | ( n16086 & n34276 ) | ( n34274 & n34276 ) ;
  assign n34278 = x41 & ~n34276 ;
  assign n34279 = x41 & ~n34272 ;
  assign n34280 = ( ~n16086 & n34278 ) | ( ~n16086 & n34279 ) | ( n34278 & n34279 ) ;
  assign n34281 = ( n34273 & ~n34277 ) | ( n34273 & n34280 ) | ( ~n34277 & n34280 ) ;
  assign n34282 = ~n34264 & n34281 ;
  assign n34283 = n34264 | n34282 ;
  assign n34285 = n34027 & ~n34048 ;
  assign n34286 = ( n34028 & n34048 ) | ( n34028 & ~n34285 ) | ( n34048 & ~n34285 ) ;
  assign n34287 = ( n34029 & ~n34031 ) | ( n34029 & n34286 ) | ( ~n34031 & n34286 ) ;
  assign n34284 = n34264 & n34281 ;
  assign n34288 = n34284 & n34287 ;
  assign n34289 = ( ~n34283 & n34287 ) | ( ~n34283 & n34288 ) | ( n34287 & n34288 ) ;
  assign n34290 = n34284 | n34287 ;
  assign n34291 = n34283 & ~n34290 ;
  assign n34292 = n34289 | n34291 ;
  assign n34293 = x126 & n6536 ;
  assign n34294 = x125 & n6531 ;
  assign n34295 = x124 & ~n6530 ;
  assign n34296 = n6871 & n34295 ;
  assign n34297 = n34294 | n34296 ;
  assign n34298 = n34293 | n34297 ;
  assign n34299 = n6539 | n34293 ;
  assign n34300 = n34297 | n34299 ;
  assign n34301 = ( n18220 & n34298 ) | ( n18220 & n34300 ) | ( n34298 & n34300 ) ;
  assign n34302 = x38 & n34300 ;
  assign n34303 = x38 & n34293 ;
  assign n34304 = ( x38 & n34297 ) | ( x38 & n34303 ) | ( n34297 & n34303 ) ;
  assign n34305 = ( n18220 & n34302 ) | ( n18220 & n34304 ) | ( n34302 & n34304 ) ;
  assign n34306 = x38 & ~n34304 ;
  assign n34307 = x38 & ~n34300 ;
  assign n34308 = ( ~n18220 & n34306 ) | ( ~n18220 & n34307 ) | ( n34306 & n34307 ) ;
  assign n34309 = ( n34301 & ~n34305 ) | ( n34301 & n34308 ) | ( ~n34305 & n34308 ) ;
  assign n34310 = n34292 | n34309 ;
  assign n34311 = n34292 & ~n34309 ;
  assign n34312 = ( ~n34292 & n34310 ) | ( ~n34292 & n34311 ) | ( n34310 & n34311 ) ;
  assign n34313 = x127 & ~n5548 ;
  assign n34314 = n5893 & n34313 ;
  assign n34315 = n5557 & n19877 ;
  assign n34316 = n34314 | n34315 ;
  assign n34317 = n5557 & n19880 ;
  assign n34318 = n34314 | n34317 ;
  assign n34319 = ( n18202 & n34316 ) | ( n18202 & n34318 ) | ( n34316 & n34318 ) ;
  assign n34320 = n34316 & n34318 ;
  assign n34321 = ( n18212 & n34319 ) | ( n18212 & n34320 ) | ( n34319 & n34320 ) ;
  assign n34322 = ( n18214 & n34319 ) | ( n18214 & n34320 ) | ( n34319 & n34320 ) ;
  assign n34323 = ( n14002 & n34321 ) | ( n14002 & n34322 ) | ( n34321 & n34322 ) ;
  assign n34324 = x35 & n34321 ;
  assign n34325 = x35 & n34322 ;
  assign n34326 = ( n14002 & n34324 ) | ( n14002 & n34325 ) | ( n34324 & n34325 ) ;
  assign n34327 = x35 & ~n34325 ;
  assign n34328 = x35 & ~n34324 ;
  assign n34329 = ( ~n14002 & n34327 ) | ( ~n14002 & n34328 ) | ( n34327 & n34328 ) ;
  assign n34330 = ( n34323 & ~n34326 ) | ( n34323 & n34329 ) | ( ~n34326 & n34329 ) ;
  assign n34331 = n33824 | n34056 ;
  assign n34332 = ( n34056 & ~n34057 ) | ( n34056 & n34331 ) | ( ~n34057 & n34331 ) ;
  assign n34333 = ( n34312 & n34330 ) | ( n34312 & ~n34332 ) | ( n34330 & ~n34332 ) ;
  assign n34334 = ( n34312 & ~n34330 ) | ( n34312 & n34332 ) | ( ~n34330 & n34332 ) ;
  assign n34335 = ( ~n34312 & n34333 ) | ( ~n34312 & n34334 ) | ( n34333 & n34334 ) ;
  assign n34336 = n33824 & ~n34057 ;
  assign n34337 = ~n33824 & n34057 ;
  assign n34338 = n34336 | n34337 ;
  assign n34339 = ~n33841 & n34338 ;
  assign n34340 = ( n33841 & n33845 ) | ( n33841 & ~n34339 ) | ( n33845 & ~n34339 ) ;
  assign n34341 = ~n34335 & n34340 ;
  assign n34342 = n34335 & ~n34340 ;
  assign n34343 = n34341 | n34342 ;
  assign n34344 = ~n34064 & n34071 ;
  assign n34345 = ~n34064 & n34066 ;
  assign n34346 = ( n33803 & n34064 ) | ( n33803 & ~n34345 ) | ( n34064 & ~n34345 ) ;
  assign n34347 = ( n32844 & n34344 ) | ( n32844 & ~n34346 ) | ( n34344 & ~n34346 ) ;
  assign n34348 = ~n34064 & n34074 ;
  assign n34349 = ( n33801 & n34064 ) | ( n33801 & ~n34345 ) | ( n34064 & ~n34345 ) ;
  assign n34350 = ( n33472 & n34348 ) | ( n33472 & ~n34349 ) | ( n34348 & ~n34349 ) ;
  assign n34351 = ( ~n30754 & n34347 ) | ( ~n30754 & n34350 ) | ( n34347 & n34350 ) ;
  assign n34352 = n34343 & n34351 ;
  assign n34353 = n34064 & ~n34343 ;
  assign n34354 = ( n34071 & n34343 ) | ( n34071 & ~n34353 ) | ( n34343 & ~n34353 ) ;
  assign n34355 = n34343 | n34345 ;
  assign n34356 = ( n33803 & n34353 ) | ( n33803 & ~n34355 ) | ( n34353 & ~n34355 ) ;
  assign n34357 = ( n32844 & n34354 ) | ( n32844 & ~n34356 ) | ( n34354 & ~n34356 ) ;
  assign n34358 = ( n33801 & n34353 ) | ( n33801 & ~n34355 ) | ( n34353 & ~n34355 ) ;
  assign n34359 = ( n34074 & n34343 ) | ( n34074 & ~n34353 ) | ( n34343 & ~n34353 ) ;
  assign n34360 = ( n33472 & ~n34358 ) | ( n33472 & n34359 ) | ( ~n34358 & n34359 ) ;
  assign n34361 = ( ~n30754 & n34357 ) | ( ~n30754 & n34360 ) | ( n34357 & n34360 ) ;
  assign n34362 = ~n34352 & n34361 ;
  assign n34363 = n34083 | n34087 ;
  assign n34364 = x100 & n18290 ;
  assign n34365 = x63 & x99 ;
  assign n34366 = ~n18290 & n34365 ;
  assign n34367 = n34364 | n34366 ;
  assign n34368 = x35 & n34082 ;
  assign n34369 = x35 | n34082 ;
  assign n34370 = ~n34368 & n34369 ;
  assign n34371 = n34367 & ~n34370 ;
  assign n34372 = ~n34367 & n34370 ;
  assign n34373 = n34371 | n34372 ;
  assign n34374 = n34363 & ~n34373 ;
  assign n34375 = ~n34083 & n34085 ;
  assign n34376 = n34373 | n34375 ;
  assign n34377 = ( n33875 & n34374 ) | ( n33875 & ~n34376 ) | ( n34374 & ~n34376 ) ;
  assign n34378 = ~n34363 & n34373 ;
  assign n34379 = n34373 & n34375 ;
  assign n34380 = ( ~n33875 & n34378 ) | ( ~n33875 & n34379 ) | ( n34378 & n34379 ) ;
  assign n34381 = n34377 | n34380 ;
  assign n34382 = x103 & n17146 ;
  assign n34383 = x102 & n17141 ;
  assign n34384 = x101 & ~n17140 ;
  assign n34385 = n17724 & n34384 ;
  assign n34386 = n34383 | n34385 ;
  assign n34387 = n34382 | n34386 ;
  assign n34388 = n17149 | n34382 ;
  assign n34389 = n34386 | n34388 ;
  assign n34390 = ( n7529 & n34387 ) | ( n7529 & n34389 ) | ( n34387 & n34389 ) ;
  assign n34391 = x62 & n34389 ;
  assign n34392 = x62 & n34382 ;
  assign n34393 = ( x62 & n34386 ) | ( x62 & n34392 ) | ( n34386 & n34392 ) ;
  assign n34394 = ( n7529 & n34391 ) | ( n7529 & n34393 ) | ( n34391 & n34393 ) ;
  assign n34395 = x62 & ~n34393 ;
  assign n34396 = x62 & ~n34389 ;
  assign n34397 = ( ~n7529 & n34395 ) | ( ~n7529 & n34396 ) | ( n34395 & n34396 ) ;
  assign n34398 = ( n34390 & ~n34394 ) | ( n34390 & n34397 ) | ( ~n34394 & n34397 ) ;
  assign n34399 = n34381 & ~n34398 ;
  assign n34400 = ~n34381 & n34398 ;
  assign n34401 = n34399 | n34400 ;
  assign n34402 = x106 & n15552 ;
  assign n34403 = x105 & n15547 ;
  assign n34404 = x104 & ~n15546 ;
  assign n34405 = n16123 & n34404 ;
  assign n34406 = n34403 | n34405 ;
  assign n34407 = n34402 | n34406 ;
  assign n34408 = n15555 | n34402 ;
  assign n34409 = n34406 | n34408 ;
  assign n34410 = ( n8656 & n34407 ) | ( n8656 & n34409 ) | ( n34407 & n34409 ) ;
  assign n34411 = x59 & n34409 ;
  assign n34412 = x59 & n34402 ;
  assign n34413 = ( x59 & n34406 ) | ( x59 & n34412 ) | ( n34406 & n34412 ) ;
  assign n34414 = ( n8656 & n34411 ) | ( n8656 & n34413 ) | ( n34411 & n34413 ) ;
  assign n34415 = x59 & ~n34413 ;
  assign n34416 = x59 & ~n34409 ;
  assign n34417 = ( ~n8656 & n34415 ) | ( ~n8656 & n34416 ) | ( n34415 & n34416 ) ;
  assign n34418 = ( n34410 & ~n34414 ) | ( n34410 & n34417 ) | ( ~n34414 & n34417 ) ;
  assign n34419 = ~n34401 & n34418 ;
  assign n34420 = n34401 | n34419 ;
  assign n34421 = n34401 & n34418 ;
  assign n34422 = n34110 | n34130 ;
  assign n34423 = ( n34110 & ~n34113 ) | ( n34110 & n34422 ) | ( ~n34113 & n34422 ) ;
  assign n34424 = ~n34421 & n34423 ;
  assign n34425 = n34420 & n34424 ;
  assign n34426 = n34421 & ~n34423 ;
  assign n34427 = ( n34420 & n34423 ) | ( n34420 & ~n34426 ) | ( n34423 & ~n34426 ) ;
  assign n34428 = ~n34425 & n34427 ;
  assign n34429 = x109 & n14045 ;
  assign n34430 = x108 & n14040 ;
  assign n34431 = x107 & ~n14039 ;
  assign n34432 = n14552 & n34431 ;
  assign n34433 = n34430 | n34432 ;
  assign n34434 = n34429 | n34433 ;
  assign n34435 = n14048 | n34429 ;
  assign n34436 = n34433 | n34435 ;
  assign n34437 = ( n9878 & n34434 ) | ( n9878 & n34436 ) | ( n34434 & n34436 ) ;
  assign n34438 = x56 & n34436 ;
  assign n34439 = x56 & n34429 ;
  assign n34440 = ( x56 & n34433 ) | ( x56 & n34439 ) | ( n34433 & n34439 ) ;
  assign n34441 = ( n9878 & n34438 ) | ( n9878 & n34440 ) | ( n34438 & n34440 ) ;
  assign n34442 = x56 & ~n34440 ;
  assign n34443 = x56 & ~n34436 ;
  assign n34444 = ( ~n9878 & n34442 ) | ( ~n9878 & n34443 ) | ( n34442 & n34443 ) ;
  assign n34445 = ( n34437 & ~n34441 ) | ( n34437 & n34444 ) | ( ~n34441 & n34444 ) ;
  assign n34446 = ~n34428 & n34445 ;
  assign n34447 = n34428 & ~n34445 ;
  assign n34448 = n34446 | n34447 ;
  assign n34449 = n34141 | n34160 ;
  assign n34450 = ( n34141 & ~n34143 ) | ( n34141 & n34449 ) | ( ~n34143 & n34449 ) ;
  assign n34451 = n34448 & ~n34450 ;
  assign n34452 = ~n34448 & n34450 ;
  assign n34453 = n34451 | n34452 ;
  assign n34454 = x112 & n12574 ;
  assign n34455 = x111 & n12569 ;
  assign n34456 = x110 & ~n12568 ;
  assign n34457 = n13076 & n34456 ;
  assign n34458 = n34455 | n34457 ;
  assign n34459 = n34454 | n34458 ;
  assign n34460 = n12577 | n34454 ;
  assign n34461 = n34458 | n34460 ;
  assign n34462 = ( n11172 & n34459 ) | ( n11172 & n34461 ) | ( n34459 & n34461 ) ;
  assign n34463 = x53 & n34461 ;
  assign n34464 = x53 & n34454 ;
  assign n34465 = ( x53 & n34458 ) | ( x53 & n34464 ) | ( n34458 & n34464 ) ;
  assign n34466 = ( n11172 & n34463 ) | ( n11172 & n34465 ) | ( n34463 & n34465 ) ;
  assign n34467 = x53 & ~n34465 ;
  assign n34468 = x53 & ~n34461 ;
  assign n34469 = ( ~n11172 & n34467 ) | ( ~n11172 & n34468 ) | ( n34467 & n34468 ) ;
  assign n34470 = ( n34462 & ~n34466 ) | ( n34462 & n34469 ) | ( ~n34466 & n34469 ) ;
  assign n34471 = ~n34453 & n34470 ;
  assign n34472 = n34453 | n34471 ;
  assign n34474 = n34166 | n34186 ;
  assign n34475 = ( ~n34163 & n34186 ) | ( ~n34163 & n34474 ) | ( n34186 & n34474 ) ;
  assign n34476 = ( n34167 & ~n34169 ) | ( n34167 & n34475 ) | ( ~n34169 & n34475 ) ;
  assign n34473 = n34453 & n34470 ;
  assign n34477 = n34473 & n34476 ;
  assign n34478 = ( ~n34472 & n34476 ) | ( ~n34472 & n34477 ) | ( n34476 & n34477 ) ;
  assign n34479 = n34473 | n34476 ;
  assign n34480 = n34472 & ~n34479 ;
  assign n34481 = n34478 | n34480 ;
  assign n34482 = x115 & n11205 ;
  assign n34483 = x114 & n11200 ;
  assign n34484 = x113 & ~n11199 ;
  assign n34485 = n11679 & n34484 ;
  assign n34486 = n34483 | n34485 ;
  assign n34487 = n34482 | n34486 ;
  assign n34488 = n11208 | n34482 ;
  assign n34489 = n34486 | n34488 ;
  assign n34490 = ( ~n12550 & n34487 ) | ( ~n12550 & n34489 ) | ( n34487 & n34489 ) ;
  assign n34491 = n34487 & n34489 ;
  assign n34492 = ( n12532 & n34490 ) | ( n12532 & n34491 ) | ( n34490 & n34491 ) ;
  assign n34493 = x50 & n34492 ;
  assign n34494 = x50 & ~n34492 ;
  assign n34495 = ( n34492 & ~n34493 ) | ( n34492 & n34494 ) | ( ~n34493 & n34494 ) ;
  assign n34496 = n34481 & ~n34495 ;
  assign n34497 = ~n34481 & n34495 ;
  assign n34498 = n34496 | n34497 ;
  assign n34499 = n34192 | n34207 ;
  assign n34500 = ( n34192 & ~n34193 ) | ( n34192 & n34499 ) | ( ~n34193 & n34499 ) ;
  assign n34501 = ~n34498 & n34500 ;
  assign n34502 = n34498 & ~n34500 ;
  assign n34503 = n34501 | n34502 ;
  assign n34504 = x118 & n9933 ;
  assign n34505 = x117 & n9928 ;
  assign n34506 = x116 & ~n9927 ;
  assign n34507 = n10379 & n34506 ;
  assign n34508 = n34505 | n34507 ;
  assign n34509 = n34504 | n34508 ;
  assign n34510 = n9936 | n34504 ;
  assign n34511 = n34508 | n34510 ;
  assign n34512 = ( ~n14002 & n34509 ) | ( ~n14002 & n34511 ) | ( n34509 & n34511 ) ;
  assign n34513 = n34509 & n34511 ;
  assign n34514 = ( n13981 & n34512 ) | ( n13981 & n34513 ) | ( n34512 & n34513 ) ;
  assign n34515 = x47 & n34514 ;
  assign n34516 = x47 & ~n34514 ;
  assign n34517 = ( n34514 & ~n34515 ) | ( n34514 & n34516 ) | ( ~n34515 & n34516 ) ;
  assign n34518 = ~n34503 & n34517 ;
  assign n34519 = n34503 & ~n34517 ;
  assign n34520 = n34518 | n34519 ;
  assign n34521 = ~n34210 & n34225 ;
  assign n34522 = n34225 & ~n34521 ;
  assign n34523 = ~n34210 & n34224 ;
  assign n34524 = ~n34225 & n34523 ;
  assign n34525 = n34521 | n34524 ;
  assign n34526 = n34224 | n34521 ;
  assign n34527 = ( n34522 & n34525 ) | ( n34522 & n34526 ) | ( n34525 & n34526 ) ;
  assign n34528 = ~n34520 & n34527 ;
  assign n34529 = n34520 & ~n34527 ;
  assign n34530 = n34528 | n34529 ;
  assign n34531 = x121 & n8724 ;
  assign n34532 = x120 & n8719 ;
  assign n34533 = x119 & ~n8718 ;
  assign n34534 = n9149 & n34533 ;
  assign n34535 = n34532 | n34534 ;
  assign n34536 = n34531 | n34535 ;
  assign n34537 = n8727 | n34531 ;
  assign n34538 = n34535 | n34537 ;
  assign n34539 = ( n15501 & n34536 ) | ( n15501 & n34538 ) | ( n34536 & n34538 ) ;
  assign n34540 = x44 & n34538 ;
  assign n34541 = x44 & n34531 ;
  assign n34542 = ( x44 & n34535 ) | ( x44 & n34541 ) | ( n34535 & n34541 ) ;
  assign n34543 = ( n15501 & n34540 ) | ( n15501 & n34542 ) | ( n34540 & n34542 ) ;
  assign n34544 = x44 & ~n34542 ;
  assign n34545 = x44 & ~n34538 ;
  assign n34546 = ( ~n15501 & n34544 ) | ( ~n15501 & n34545 ) | ( n34544 & n34545 ) ;
  assign n34547 = ( n34539 & ~n34543 ) | ( n34539 & n34546 ) | ( ~n34543 & n34546 ) ;
  assign n34548 = ~n34530 & n34547 ;
  assign n34549 = n34530 | n34548 ;
  assign n34550 = n34232 | n34252 ;
  assign n34551 = ( n34232 & ~n34235 ) | ( n34232 & n34550 ) | ( ~n34235 & n34550 ) ;
  assign n34552 = n34530 & n34547 ;
  assign n34553 = n34551 & n34552 ;
  assign n34554 = ( ~n34549 & n34551 ) | ( ~n34549 & n34553 ) | ( n34551 & n34553 ) ;
  assign n34555 = n34551 | n34552 ;
  assign n34556 = n34549 & ~n34555 ;
  assign n34557 = n34554 | n34556 ;
  assign n34558 = x124 & n7566 ;
  assign n34559 = x123 & n7561 ;
  assign n34560 = x122 & ~n7560 ;
  assign n34561 = n7953 & n34560 ;
  assign n34562 = n34559 | n34561 ;
  assign n34563 = n34558 | n34562 ;
  assign n34564 = n7569 | n34558 ;
  assign n34565 = n34562 | n34564 ;
  assign n34566 = ( n17084 & n34563 ) | ( n17084 & n34565 ) | ( n34563 & n34565 ) ;
  assign n34567 = x41 & n34565 ;
  assign n34568 = x41 & n34558 ;
  assign n34569 = ( x41 & n34562 ) | ( x41 & n34568 ) | ( n34562 & n34568 ) ;
  assign n34570 = ( n17084 & n34567 ) | ( n17084 & n34569 ) | ( n34567 & n34569 ) ;
  assign n34571 = x41 & ~n34569 ;
  assign n34572 = x41 & ~n34565 ;
  assign n34573 = ( ~n17084 & n34571 ) | ( ~n17084 & n34572 ) | ( n34571 & n34572 ) ;
  assign n34574 = ( n34566 & ~n34570 ) | ( n34566 & n34573 ) | ( ~n34570 & n34573 ) ;
  assign n34575 = ~n34557 & n34574 ;
  assign n34576 = n34557 | n34575 ;
  assign n34578 = n34262 | n34281 ;
  assign n34579 = ( n34262 & ~n34264 ) | ( n34262 & n34578 ) | ( ~n34264 & n34578 ) ;
  assign n34577 = n34557 & n34574 ;
  assign n34580 = n34577 & n34579 ;
  assign n34581 = ( ~n34576 & n34579 ) | ( ~n34576 & n34580 ) | ( n34579 & n34580 ) ;
  assign n34582 = n34577 | n34579 ;
  assign n34583 = n34576 & ~n34582 ;
  assign n34584 = n34581 | n34583 ;
  assign n34585 = x127 & n6536 ;
  assign n34586 = x126 & n6531 ;
  assign n34587 = x125 & ~n6530 ;
  assign n34588 = n6871 & n34587 ;
  assign n34589 = n34586 | n34588 ;
  assign n34590 = n34585 | n34589 ;
  assign n34591 = n6539 | n34585 ;
  assign n34592 = n34589 | n34591 ;
  assign n34593 = ( n18763 & n34590 ) | ( n18763 & n34592 ) | ( n34590 & n34592 ) ;
  assign n34594 = x38 & n34592 ;
  assign n34595 = x38 & n34585 ;
  assign n34596 = ( x38 & n34589 ) | ( x38 & n34595 ) | ( n34589 & n34595 ) ;
  assign n34597 = ( n18763 & n34594 ) | ( n18763 & n34596 ) | ( n34594 & n34596 ) ;
  assign n34598 = x38 & ~n34596 ;
  assign n34599 = x38 & ~n34592 ;
  assign n34600 = ( ~n18763 & n34598 ) | ( ~n18763 & n34599 ) | ( n34598 & n34599 ) ;
  assign n34601 = ( n34593 & ~n34597 ) | ( n34593 & n34600 ) | ( ~n34597 & n34600 ) ;
  assign n34602 = ~n34584 & n34601 ;
  assign n34603 = n34584 | n34602 ;
  assign n34605 = n34287 | n34309 ;
  assign n34606 = n34283 & ~n34309 ;
  assign n34607 = ( n34288 & n34605 ) | ( n34288 & ~n34606 ) | ( n34605 & ~n34606 ) ;
  assign n34608 = ( n34289 & ~n34292 ) | ( n34289 & n34607 ) | ( ~n34292 & n34607 ) ;
  assign n34604 = n34584 & n34601 ;
  assign n34609 = n34604 & n34608 ;
  assign n34610 = ( ~n34603 & n34608 ) | ( ~n34603 & n34609 ) | ( n34608 & n34609 ) ;
  assign n34611 = n34604 | n34608 ;
  assign n34612 = n34603 & ~n34611 ;
  assign n34613 = n34610 | n34612 ;
  assign n34614 = n34330 & n34332 ;
  assign n34615 = n34332 & ~n34614 ;
  assign n34616 = n34330 & ~n34332 ;
  assign n34617 = ~n34312 & n34616 ;
  assign n34618 = ( ~n34312 & n34615 ) | ( ~n34312 & n34617 ) | ( n34615 & n34617 ) ;
  assign n34619 = ~n34613 & n34614 ;
  assign n34620 = ( ~n34613 & n34618 ) | ( ~n34613 & n34619 ) | ( n34618 & n34619 ) ;
  assign n34621 = n34613 & ~n34614 ;
  assign n34622 = ~n34618 & n34621 ;
  assign n34623 = n34620 | n34622 ;
  assign n34624 = ~n34341 & n34357 ;
  assign n34625 = ~n34341 & n34355 ;
  assign n34626 = n34341 | n34353 ;
  assign n34627 = ( n33801 & ~n34625 ) | ( n33801 & n34626 ) | ( ~n34625 & n34626 ) ;
  assign n34628 = ~n34341 & n34343 ;
  assign n34629 = ( n34074 & ~n34626 ) | ( n34074 & n34628 ) | ( ~n34626 & n34628 ) ;
  assign n34630 = ( n33472 & ~n34627 ) | ( n33472 & n34629 ) | ( ~n34627 & n34629 ) ;
  assign n34631 = ( ~n30754 & n34624 ) | ( ~n30754 & n34630 ) | ( n34624 & n34630 ) ;
  assign n34632 = n34623 & n34631 ;
  assign n34633 = n34341 & ~n34623 ;
  assign n34634 = ( n34357 & n34623 ) | ( n34357 & ~n34633 ) | ( n34623 & ~n34633 ) ;
  assign n34635 = ~n34623 & n34627 ;
  assign n34636 = ~n34623 & n34626 ;
  assign n34637 = n34623 | n34628 ;
  assign n34638 = ( n34074 & ~n34636 ) | ( n34074 & n34637 ) | ( ~n34636 & n34637 ) ;
  assign n34639 = ( n33472 & ~n34635 ) | ( n33472 & n34638 ) | ( ~n34635 & n34638 ) ;
  assign n34640 = ( ~n30754 & n34634 ) | ( ~n30754 & n34639 ) | ( n34634 & n34639 ) ;
  assign n34641 = ~n34632 & n34640 ;
  assign n34642 = x125 & n7566 ;
  assign n34643 = x124 & n7561 ;
  assign n34644 = x123 & ~n7560 ;
  assign n34645 = n7953 & n34644 ;
  assign n34646 = n34643 | n34645 ;
  assign n34647 = n34642 | n34646 ;
  assign n34648 = n7569 | n34642 ;
  assign n34649 = n34646 | n34648 ;
  assign n34650 = ( n17670 & n34647 ) | ( n17670 & n34649 ) | ( n34647 & n34649 ) ;
  assign n34651 = x41 & n34649 ;
  assign n34652 = x41 & n34642 ;
  assign n34653 = ( x41 & n34646 ) | ( x41 & n34652 ) | ( n34646 & n34652 ) ;
  assign n34654 = ( n17670 & n34651 ) | ( n17670 & n34653 ) | ( n34651 & n34653 ) ;
  assign n34655 = x41 & ~n34653 ;
  assign n34656 = x41 & ~n34649 ;
  assign n34657 = ( ~n17670 & n34655 ) | ( ~n17670 & n34656 ) | ( n34655 & n34656 ) ;
  assign n34658 = ( n34650 & ~n34654 ) | ( n34650 & n34657 ) | ( ~n34654 & n34657 ) ;
  assign n34659 = x127 & n6531 ;
  assign n34660 = x126 & ~n6530 ;
  assign n34661 = n6871 & n34660 ;
  assign n34662 = n34659 | n34661 ;
  assign n34663 = n6539 | n34662 ;
  assign n34664 = ( n19328 & n34662 ) | ( n19328 & n34663 ) | ( n34662 & n34663 ) ;
  assign n34665 = x38 & n34662 ;
  assign n34666 = ( x38 & n9196 ) | ( x38 & n34662 ) | ( n9196 & n34662 ) ;
  assign n34667 = ( n19328 & n34665 ) | ( n19328 & n34666 ) | ( n34665 & n34666 ) ;
  assign n34668 = x38 & ~n9196 ;
  assign n34669 = ~n34662 & n34668 ;
  assign n34670 = x38 & ~n34662 ;
  assign n34671 = ( ~n19328 & n34669 ) | ( ~n19328 & n34670 ) | ( n34669 & n34670 ) ;
  assign n34672 = ( n34664 & ~n34667 ) | ( n34664 & n34671 ) | ( ~n34667 & n34671 ) ;
  assign n34673 = n34574 & n34672 ;
  assign n34674 = ~n34557 & n34673 ;
  assign n34675 = ( n34581 & n34672 ) | ( n34581 & n34674 ) | ( n34672 & n34674 ) ;
  assign n34676 = n34574 | n34672 ;
  assign n34677 = ( ~n34557 & n34672 ) | ( ~n34557 & n34676 ) | ( n34672 & n34676 ) ;
  assign n34678 = n34581 | n34677 ;
  assign n34679 = ~n34675 & n34678 ;
  assign n34680 = x103 & n17141 ;
  assign n34681 = x102 & ~n17140 ;
  assign n34682 = n17724 & n34681 ;
  assign n34683 = n34680 | n34682 ;
  assign n34684 = x104 & n17146 ;
  assign n34685 = n17149 | n34684 ;
  assign n34686 = n34683 | n34685 ;
  assign n34687 = ~x62 & n34686 ;
  assign n34688 = ~x62 & n34684 ;
  assign n34689 = ( ~x62 & n34683 ) | ( ~x62 & n34688 ) | ( n34683 & n34688 ) ;
  assign n34690 = ( n7911 & n34687 ) | ( n7911 & n34689 ) | ( n34687 & n34689 ) ;
  assign n34691 = x62 & ~n34686 ;
  assign n34692 = x62 & x104 ;
  assign n34693 = n17146 & n34692 ;
  assign n34694 = x62 & ~n34693 ;
  assign n34695 = ~n34683 & n34694 ;
  assign n34696 = ( ~n7911 & n34691 ) | ( ~n7911 & n34695 ) | ( n34691 & n34695 ) ;
  assign n34697 = n34690 | n34696 ;
  assign n34698 = ( ~x35 & n34082 ) | ( ~x35 & n34367 ) | ( n34082 & n34367 ) ;
  assign n34699 = x101 & n18290 ;
  assign n34700 = x63 & x100 ;
  assign n34701 = ~n18290 & n34700 ;
  assign n34702 = n34699 | n34701 ;
  assign n34703 = n34698 & ~n34702 ;
  assign n34704 = n34698 & ~n34703 ;
  assign n34705 = n34698 | n34702 ;
  assign n34706 = ~n34704 & n34705 ;
  assign n34707 = n34697 & ~n34706 ;
  assign n34708 = ~n34697 & n34706 ;
  assign n34709 = n34707 | n34708 ;
  assign n34710 = n34377 | n34398 ;
  assign n34711 = ( n34377 & ~n34381 ) | ( n34377 & n34710 ) | ( ~n34381 & n34710 ) ;
  assign n34712 = n34709 & ~n34711 ;
  assign n34713 = ~n34709 & n34711 ;
  assign n34714 = n34712 | n34713 ;
  assign n34715 = x107 & n15552 ;
  assign n34716 = x106 & n15547 ;
  assign n34717 = x105 & ~n15546 ;
  assign n34718 = n16123 & n34717 ;
  assign n34719 = n34716 | n34718 ;
  assign n34720 = n34715 | n34719 ;
  assign n34721 = n15555 | n34715 ;
  assign n34722 = n34719 | n34721 ;
  assign n34723 = ( n9084 & n34720 ) | ( n9084 & n34722 ) | ( n34720 & n34722 ) ;
  assign n34724 = x59 & n34722 ;
  assign n34725 = x59 & n34715 ;
  assign n34726 = ( x59 & n34719 ) | ( x59 & n34725 ) | ( n34719 & n34725 ) ;
  assign n34727 = ( n9084 & n34724 ) | ( n9084 & n34726 ) | ( n34724 & n34726 ) ;
  assign n34728 = x59 & ~n34726 ;
  assign n34729 = x59 & ~n34722 ;
  assign n34730 = ( ~n9084 & n34728 ) | ( ~n9084 & n34729 ) | ( n34728 & n34729 ) ;
  assign n34731 = ( n34723 & ~n34727 ) | ( n34723 & n34730 ) | ( ~n34727 & n34730 ) ;
  assign n34732 = n34714 & n34731 ;
  assign n34733 = n34709 & ~n34731 ;
  assign n34734 = ( n34711 & n34731 ) | ( n34711 & ~n34733 ) | ( n34731 & ~n34733 ) ;
  assign n34735 = n34712 | n34734 ;
  assign n34736 = ~n34732 & n34735 ;
  assign n34737 = n34421 & n34423 ;
  assign n34738 = ( ~n34420 & n34423 ) | ( ~n34420 & n34737 ) | ( n34423 & n34737 ) ;
  assign n34739 = n34419 | n34738 ;
  assign n34740 = n34736 & ~n34739 ;
  assign n34741 = ~n34736 & n34739 ;
  assign n34742 = n34740 | n34741 ;
  assign n34743 = x110 & n14045 ;
  assign n34744 = x109 & n14040 ;
  assign n34745 = x108 & ~n14039 ;
  assign n34746 = n14552 & n34745 ;
  assign n34747 = n34744 | n34746 ;
  assign n34748 = n34743 | n34747 ;
  assign n34749 = n14048 | n34743 ;
  assign n34750 = n34747 | n34749 ;
  assign n34751 = ( n10330 & n34748 ) | ( n10330 & n34750 ) | ( n34748 & n34750 ) ;
  assign n34752 = x56 & n34750 ;
  assign n34753 = x56 & n34743 ;
  assign n34754 = ( x56 & n34747 ) | ( x56 & n34753 ) | ( n34747 & n34753 ) ;
  assign n34755 = ( n10330 & n34752 ) | ( n10330 & n34754 ) | ( n34752 & n34754 ) ;
  assign n34756 = x56 & ~n34754 ;
  assign n34757 = x56 & ~n34750 ;
  assign n34758 = ( ~n10330 & n34756 ) | ( ~n10330 & n34757 ) | ( n34756 & n34757 ) ;
  assign n34759 = ( n34751 & ~n34755 ) | ( n34751 & n34758 ) | ( ~n34755 & n34758 ) ;
  assign n34760 = n34742 & n34759 ;
  assign n34761 = n34735 & ~n34759 ;
  assign n34762 = ~n34732 & n34761 ;
  assign n34763 = ( n34739 & n34759 ) | ( n34739 & ~n34762 ) | ( n34759 & ~n34762 ) ;
  assign n34764 = n34740 | n34763 ;
  assign n34765 = ~n34760 & n34764 ;
  assign n34766 = n34446 | n34450 ;
  assign n34767 = ( n34446 & ~n34448 ) | ( n34446 & n34766 ) | ( ~n34448 & n34766 ) ;
  assign n34768 = n34765 & ~n34767 ;
  assign n34769 = ~n34765 & n34767 ;
  assign n34770 = n34768 | n34769 ;
  assign n34771 = x113 & n12574 ;
  assign n34772 = x112 & n12569 ;
  assign n34773 = x111 & ~n12568 ;
  assign n34774 = n13076 & n34773 ;
  assign n34775 = n34772 | n34774 ;
  assign n34776 = n34771 | n34775 ;
  assign n34777 = n12577 | n34771 ;
  assign n34778 = n34775 | n34777 ;
  assign n34779 = ( ~n11642 & n34776 ) | ( ~n11642 & n34778 ) | ( n34776 & n34778 ) ;
  assign n34780 = n34776 & n34778 ;
  assign n34781 = ( n11626 & n34779 ) | ( n11626 & n34780 ) | ( n34779 & n34780 ) ;
  assign n34782 = x53 & n34781 ;
  assign n34783 = x53 & ~n34781 ;
  assign n34784 = ( n34781 & ~n34782 ) | ( n34781 & n34783 ) | ( ~n34782 & n34783 ) ;
  assign n34785 = n34770 & n34784 ;
  assign n34786 = n34767 | n34784 ;
  assign n34787 = ( ~n34765 & n34784 ) | ( ~n34765 & n34786 ) | ( n34784 & n34786 ) ;
  assign n34788 = n34768 | n34787 ;
  assign n34789 = ~n34785 & n34788 ;
  assign n34790 = n34471 | n34478 ;
  assign n34791 = n34789 & ~n34790 ;
  assign n34792 = ~n34789 & n34790 ;
  assign n34793 = n34791 | n34792 ;
  assign n34794 = x116 & n11205 ;
  assign n34795 = x115 & n11200 ;
  assign n34796 = x114 & ~n11199 ;
  assign n34797 = n11679 & n34796 ;
  assign n34798 = n34795 | n34797 ;
  assign n34799 = n34794 | n34798 ;
  assign n34800 = n11208 | n34794 ;
  assign n34801 = n34798 | n34800 ;
  assign n34802 = ( ~n13040 & n34799 ) | ( ~n13040 & n34801 ) | ( n34799 & n34801 ) ;
  assign n34803 = n34799 & n34801 ;
  assign n34804 = ( n13022 & n34802 ) | ( n13022 & n34803 ) | ( n34802 & n34803 ) ;
  assign n34805 = x50 & n34804 ;
  assign n34806 = x50 & ~n34804 ;
  assign n34807 = ( n34804 & ~n34805 ) | ( n34804 & n34806 ) | ( ~n34805 & n34806 ) ;
  assign n34808 = n34793 & n34807 ;
  assign n34809 = n34792 | n34807 ;
  assign n34810 = n34791 | n34809 ;
  assign n34811 = ~n34808 & n34810 ;
  assign n34812 = n34497 | n34500 ;
  assign n34813 = ( n34497 & ~n34498 ) | ( n34497 & n34812 ) | ( ~n34498 & n34812 ) ;
  assign n34814 = ~n34811 & n34813 ;
  assign n34815 = n34811 & ~n34813 ;
  assign n34816 = n34814 | n34815 ;
  assign n34817 = x119 & n9933 ;
  assign n34818 = x118 & n9928 ;
  assign n34819 = x117 & ~n9927 ;
  assign n34820 = n10379 & n34819 ;
  assign n34821 = n34818 | n34820 ;
  assign n34822 = n34817 | n34821 ;
  assign n34823 = n9936 | n34817 ;
  assign n34824 = n34821 | n34823 ;
  assign n34825 = ( n14496 & n34822 ) | ( n14496 & n34824 ) | ( n34822 & n34824 ) ;
  assign n34826 = x47 & n34824 ;
  assign n34827 = x47 & n34817 ;
  assign n34828 = ( x47 & n34821 ) | ( x47 & n34827 ) | ( n34821 & n34827 ) ;
  assign n34829 = ( n14496 & n34826 ) | ( n14496 & n34828 ) | ( n34826 & n34828 ) ;
  assign n34830 = x47 & ~n34828 ;
  assign n34831 = x47 & ~n34824 ;
  assign n34832 = ( ~n14496 & n34830 ) | ( ~n14496 & n34831 ) | ( n34830 & n34831 ) ;
  assign n34833 = ( n34825 & ~n34829 ) | ( n34825 & n34832 ) | ( ~n34829 & n34832 ) ;
  assign n34834 = ~n34816 & n34833 ;
  assign n34835 = n34816 | n34834 ;
  assign n34837 = ~n34518 & n34520 ;
  assign n34838 = ( n34518 & n34527 ) | ( n34518 & ~n34837 ) | ( n34527 & ~n34837 ) ;
  assign n34836 = n34816 & n34833 ;
  assign n34839 = n34836 & n34838 ;
  assign n34840 = ( ~n34835 & n34838 ) | ( ~n34835 & n34839 ) | ( n34838 & n34839 ) ;
  assign n34841 = n34836 | n34838 ;
  assign n34842 = n34835 & ~n34841 ;
  assign n34843 = n34840 | n34842 ;
  assign n34844 = x122 & n8724 ;
  assign n34845 = x121 & n8719 ;
  assign n34846 = x120 & ~n8718 ;
  assign n34847 = n9149 & n34846 ;
  assign n34848 = n34845 | n34847 ;
  assign n34849 = n34844 | n34848 ;
  assign n34850 = n8727 | n34844 ;
  assign n34851 = n34848 | n34850 ;
  assign n34852 = ( n16043 & n34849 ) | ( n16043 & n34851 ) | ( n34849 & n34851 ) ;
  assign n34853 = x44 & n34851 ;
  assign n34854 = x44 & n34844 ;
  assign n34855 = ( x44 & n34848 ) | ( x44 & n34854 ) | ( n34848 & n34854 ) ;
  assign n34856 = ( n16043 & n34853 ) | ( n16043 & n34855 ) | ( n34853 & n34855 ) ;
  assign n34857 = x44 & ~n34855 ;
  assign n34858 = x44 & ~n34851 ;
  assign n34859 = ( ~n16043 & n34857 ) | ( ~n16043 & n34858 ) | ( n34857 & n34858 ) ;
  assign n34860 = ( n34852 & ~n34856 ) | ( n34852 & n34859 ) | ( ~n34856 & n34859 ) ;
  assign n34861 = ~n34843 & n34860 ;
  assign n34862 = n34843 | n34861 ;
  assign n34864 = n34548 | n34551 ;
  assign n34865 = ~n34548 & n34549 ;
  assign n34866 = ( n34553 & n34864 ) | ( n34553 & ~n34865 ) | ( n34864 & ~n34865 ) ;
  assign n34863 = n34843 & n34860 ;
  assign n34867 = n34863 & n34866 ;
  assign n34868 = ( ~n34862 & n34866 ) | ( ~n34862 & n34867 ) | ( n34866 & n34867 ) ;
  assign n34869 = n34863 | n34866 ;
  assign n34870 = n34862 & ~n34869 ;
  assign n34871 = n34868 | n34870 ;
  assign n34872 = ( n34658 & n34679 ) | ( n34658 & ~n34871 ) | ( n34679 & ~n34871 ) ;
  assign n34873 = ( ~n34679 & n34871 ) | ( ~n34679 & n34872 ) | ( n34871 & n34872 ) ;
  assign n34874 = ( ~n34658 & n34872 ) | ( ~n34658 & n34873 ) | ( n34872 & n34873 ) ;
  assign n34875 = n34602 | n34608 ;
  assign n34876 = ~n34602 & n34603 ;
  assign n34877 = ( n34609 & n34875 ) | ( n34609 & ~n34876 ) | ( n34875 & ~n34876 ) ;
  assign n34878 = n34874 & ~n34877 ;
  assign n34879 = ~n34874 & n34877 ;
  assign n34880 = n34878 | n34879 ;
  assign n34881 = ~n34620 & n34623 ;
  assign n34882 = n34341 | n34620 ;
  assign n34883 = ( n34620 & ~n34623 ) | ( n34620 & n34882 ) | ( ~n34623 & n34882 ) ;
  assign n34884 = ( n34357 & n34881 ) | ( n34357 & ~n34883 ) | ( n34881 & ~n34883 ) ;
  assign n34885 = ( n34620 & n34627 ) | ( n34620 & ~n34881 ) | ( n34627 & ~n34881 ) ;
  assign n34886 = n34620 | n34636 ;
  assign n34887 = ~n34620 & n34637 ;
  assign n34888 = ( n34074 & ~n34886 ) | ( n34074 & n34887 ) | ( ~n34886 & n34887 ) ;
  assign n34889 = ( n33472 & ~n34885 ) | ( n33472 & n34888 ) | ( ~n34885 & n34888 ) ;
  assign n34890 = ( ~n30754 & n34884 ) | ( ~n30754 & n34889 ) | ( n34884 & n34889 ) ;
  assign n34891 = n34880 & n34890 ;
  assign n34892 = ~n34880 & n34883 ;
  assign n34893 = n34620 & ~n34880 ;
  assign n34894 = ( n34623 & n34880 ) | ( n34623 & ~n34893 ) | ( n34880 & ~n34893 ) ;
  assign n34895 = ( n34357 & ~n34892 ) | ( n34357 & n34894 ) | ( ~n34892 & n34894 ) ;
  assign n34896 = n34880 | n34888 ;
  assign n34897 = n34880 | n34881 ;
  assign n34898 = ( n34627 & n34893 ) | ( n34627 & ~n34897 ) | ( n34893 & ~n34897 ) ;
  assign n34899 = ( n33472 & n34896 ) | ( n33472 & ~n34898 ) | ( n34896 & ~n34898 ) ;
  assign n34900 = ( ~n30754 & n34895 ) | ( ~n30754 & n34899 ) | ( n34895 & n34899 ) ;
  assign n34901 = ~n34891 & n34900 ;
  assign n34920 = n34658 | n34868 ;
  assign n34921 = ( n34868 & ~n34871 ) | ( n34868 & n34920 ) | ( ~n34871 & n34920 ) ;
  assign n34902 = x127 & ~n6530 ;
  assign n34903 = n6871 & n34902 ;
  assign n34904 = n6539 & n19877 ;
  assign n34905 = n34903 | n34904 ;
  assign n34906 = n6539 & n19880 ;
  assign n34907 = n34903 | n34906 ;
  assign n34908 = ( n18202 & n34905 ) | ( n18202 & n34907 ) | ( n34905 & n34907 ) ;
  assign n34909 = n34905 & n34907 ;
  assign n34910 = ( n18212 & n34908 ) | ( n18212 & n34909 ) | ( n34908 & n34909 ) ;
  assign n34911 = ( n18214 & n34908 ) | ( n18214 & n34909 ) | ( n34908 & n34909 ) ;
  assign n34912 = ( n14002 & n34910 ) | ( n14002 & n34911 ) | ( n34910 & n34911 ) ;
  assign n34913 = x38 & n34910 ;
  assign n34914 = x38 & n34911 ;
  assign n34915 = ( n14002 & n34913 ) | ( n14002 & n34914 ) | ( n34913 & n34914 ) ;
  assign n34916 = x38 & ~n34914 ;
  assign n34917 = x38 & ~n34913 ;
  assign n34918 = ( ~n14002 & n34916 ) | ( ~n14002 & n34917 ) | ( n34916 & n34917 ) ;
  assign n34919 = ( n34912 & ~n34915 ) | ( n34912 & n34918 ) | ( ~n34915 & n34918 ) ;
  assign n34922 = n34919 & n34921 ;
  assign n34923 = n34921 & ~n34922 ;
  assign n35042 = ( n34769 & ~n34770 ) | ( n34769 & n34787 ) | ( ~n34770 & n34787 ) ;
  assign n34924 = x102 & n18290 ;
  assign n34925 = x63 & x101 ;
  assign n34926 = ~n18290 & n34925 ;
  assign n34927 = n34924 | n34926 ;
  assign n34928 = ~n34702 & n34927 ;
  assign n34929 = n34702 | n34928 ;
  assign n34930 = n34927 & ~n34928 ;
  assign n34931 = n34929 & ~n34930 ;
  assign n34932 = n34703 & ~n34931 ;
  assign n34933 = n34931 | n34932 ;
  assign n34934 = n34706 & ~n34933 ;
  assign n34935 = ( n34697 & n34933 ) | ( n34697 & ~n34934 ) | ( n34933 & ~n34934 ) ;
  assign n34936 = ~n34703 & n34705 ;
  assign n34937 = ~n34704 & n34936 ;
  assign n34938 = n34931 & ~n34937 ;
  assign n34939 = n34703 & n34931 ;
  assign n34940 = ( n34697 & n34938 ) | ( n34697 & n34939 ) | ( n34938 & n34939 ) ;
  assign n34941 = n34935 & ~n34940 ;
  assign n34942 = x105 & n17146 ;
  assign n34943 = x104 & n17141 ;
  assign n34944 = x103 & ~n17140 ;
  assign n34945 = n17724 & n34944 ;
  assign n34946 = n34943 | n34945 ;
  assign n34947 = n34942 | n34946 ;
  assign n34948 = n17149 | n34942 ;
  assign n34949 = n34946 | n34948 ;
  assign n34950 = ( n8273 & n34947 ) | ( n8273 & n34949 ) | ( n34947 & n34949 ) ;
  assign n34951 = x62 & n34949 ;
  assign n34952 = x62 & n34942 ;
  assign n34953 = ( x62 & n34946 ) | ( x62 & n34952 ) | ( n34946 & n34952 ) ;
  assign n34954 = ( n8273 & n34951 ) | ( n8273 & n34953 ) | ( n34951 & n34953 ) ;
  assign n34955 = x62 & ~n34953 ;
  assign n34956 = x62 & ~n34949 ;
  assign n34957 = ( ~n8273 & n34955 ) | ( ~n8273 & n34956 ) | ( n34955 & n34956 ) ;
  assign n34958 = ( n34950 & ~n34954 ) | ( n34950 & n34957 ) | ( ~n34954 & n34957 ) ;
  assign n34959 = ~n34941 & n34958 ;
  assign n34960 = n34941 & ~n34958 ;
  assign n34961 = n34959 | n34960 ;
  assign n34962 = x108 & n15552 ;
  assign n34963 = x107 & n15547 ;
  assign n34964 = x106 & ~n15546 ;
  assign n34965 = n16123 & n34964 ;
  assign n34966 = n34963 | n34965 ;
  assign n34967 = n34962 | n34966 ;
  assign n34968 = n15555 | n34962 ;
  assign n34969 = n34966 | n34968 ;
  assign n34970 = ( n9479 & n34967 ) | ( n9479 & n34969 ) | ( n34967 & n34969 ) ;
  assign n34971 = x59 & n34969 ;
  assign n34972 = x59 & n34962 ;
  assign n34973 = ( x59 & n34966 ) | ( x59 & n34972 ) | ( n34966 & n34972 ) ;
  assign n34974 = ( n9479 & n34971 ) | ( n9479 & n34973 ) | ( n34971 & n34973 ) ;
  assign n34975 = x59 & ~n34973 ;
  assign n34976 = x59 & ~n34969 ;
  assign n34977 = ( ~n9479 & n34975 ) | ( ~n9479 & n34976 ) | ( n34975 & n34976 ) ;
  assign n34978 = ( n34970 & ~n34974 ) | ( n34970 & n34977 ) | ( ~n34974 & n34977 ) ;
  assign n34979 = n34961 | n34978 ;
  assign n34980 = n34961 & n34978 ;
  assign n34981 = n34979 & ~n34980 ;
  assign n34982 = ( n34713 & ~n34714 ) | ( n34713 & n34734 ) | ( ~n34714 & n34734 ) ;
  assign n34983 = n34981 & ~n34982 ;
  assign n34984 = ~n34981 & n34982 ;
  assign n34985 = n34983 | n34984 ;
  assign n34986 = x111 & n14045 ;
  assign n34987 = x110 & n14040 ;
  assign n34988 = x109 & ~n14039 ;
  assign n34989 = n14552 & n34988 ;
  assign n34990 = n34987 | n34989 ;
  assign n34991 = n34986 | n34990 ;
  assign n34992 = n14048 | n34986 ;
  assign n34993 = n34990 | n34992 ;
  assign n34994 = ( n10749 & n34991 ) | ( n10749 & n34993 ) | ( n34991 & n34993 ) ;
  assign n34995 = x56 & n34993 ;
  assign n34996 = x56 & n34986 ;
  assign n34997 = ( x56 & n34990 ) | ( x56 & n34996 ) | ( n34990 & n34996 ) ;
  assign n34998 = ( n10749 & n34995 ) | ( n10749 & n34997 ) | ( n34995 & n34997 ) ;
  assign n34999 = x56 & ~n34997 ;
  assign n35000 = x56 & ~n34993 ;
  assign n35001 = ( ~n10749 & n34999 ) | ( ~n10749 & n35000 ) | ( n34999 & n35000 ) ;
  assign n35002 = ( n34994 & ~n34998 ) | ( n34994 & n35001 ) | ( ~n34998 & n35001 ) ;
  assign n35003 = n34985 & n35002 ;
  assign n35004 = n34984 | n35002 ;
  assign n35005 = n34983 | n35004 ;
  assign n35006 = ~n35003 & n35005 ;
  assign n35007 = ( n34741 & ~n34742 ) | ( n34741 & n34763 ) | ( ~n34742 & n34763 ) ;
  assign n35008 = n35006 & ~n35007 ;
  assign n35009 = ~n35006 & n35007 ;
  assign n35010 = n35008 | n35009 ;
  assign n35011 = x114 & n12574 ;
  assign n35012 = x113 & n12569 ;
  assign n35013 = x112 & ~n12568 ;
  assign n35014 = n13076 & n35013 ;
  assign n35015 = n35012 | n35014 ;
  assign n35016 = n35011 | n35015 ;
  assign n35017 = n12577 | n35011 ;
  assign n35018 = n35015 | n35017 ;
  assign n35019 = ( ~n12095 & n35016 ) | ( ~n12095 & n35018 ) | ( n35016 & n35018 ) ;
  assign n35020 = n35016 & n35018 ;
  assign n35021 = ( n12079 & n35019 ) | ( n12079 & n35020 ) | ( n35019 & n35020 ) ;
  assign n35022 = x53 & n35021 ;
  assign n35023 = x53 & ~n35021 ;
  assign n35024 = ( n35021 & ~n35022 ) | ( n35021 & n35023 ) | ( ~n35022 & n35023 ) ;
  assign n35025 = n35010 & ~n35024 ;
  assign n35026 = ~n35010 & n35024 ;
  assign n35027 = n35025 | n35026 ;
  assign n35028 = x117 & n11205 ;
  assign n35029 = x116 & n11200 ;
  assign n35030 = x115 & ~n11199 ;
  assign n35031 = n11679 & n35030 ;
  assign n35032 = n35029 | n35031 ;
  assign n35033 = n35028 | n35032 ;
  assign n35034 = n11208 | n35028 ;
  assign n35035 = n35032 | n35034 ;
  assign n35036 = ( ~n13522 & n35033 ) | ( ~n13522 & n35035 ) | ( n35033 & n35035 ) ;
  assign n35037 = n35033 & n35035 ;
  assign n35038 = ( n13503 & n35036 ) | ( n13503 & n35037 ) | ( n35036 & n35037 ) ;
  assign n35039 = x50 & n35038 ;
  assign n35040 = x50 & ~n35038 ;
  assign n35041 = ( n35038 & ~n35039 ) | ( n35038 & n35040 ) | ( ~n35039 & n35040 ) ;
  assign n35043 = ( ~n35027 & n35041 ) | ( ~n35027 & n35042 ) | ( n35041 & n35042 ) ;
  assign n35044 = ( n35027 & ~n35041 ) | ( n35027 & n35043 ) | ( ~n35041 & n35043 ) ;
  assign n35045 = ( ~n35042 & n35043 ) | ( ~n35042 & n35044 ) | ( n35043 & n35044 ) ;
  assign n35046 = ( n34792 & ~n34793 ) | ( n34792 & n34809 ) | ( ~n34793 & n34809 ) ;
  assign n35047 = ~n35045 & n35046 ;
  assign n35048 = n35045 & ~n35046 ;
  assign n35049 = n35047 | n35048 ;
  assign n35050 = x120 & n9933 ;
  assign n35051 = x119 & n9928 ;
  assign n35052 = x118 & ~n9927 ;
  assign n35053 = n10379 & n35052 ;
  assign n35054 = n35051 | n35053 ;
  assign n35055 = n35050 | n35054 ;
  assign n35056 = n9936 | n35050 ;
  assign n35057 = n35054 | n35056 ;
  assign n35058 = ( n14991 & n35055 ) | ( n14991 & n35057 ) | ( n35055 & n35057 ) ;
  assign n35059 = x47 & n35057 ;
  assign n35060 = x47 & n35050 ;
  assign n35061 = ( x47 & n35054 ) | ( x47 & n35060 ) | ( n35054 & n35060 ) ;
  assign n35062 = ( n14991 & n35059 ) | ( n14991 & n35061 ) | ( n35059 & n35061 ) ;
  assign n35063 = x47 & ~n35061 ;
  assign n35064 = x47 & ~n35057 ;
  assign n35065 = ( ~n14991 & n35063 ) | ( ~n14991 & n35064 ) | ( n35063 & n35064 ) ;
  assign n35066 = ( n35058 & ~n35062 ) | ( n35058 & n35065 ) | ( ~n35062 & n35065 ) ;
  assign n35067 = ~n35049 & n35066 ;
  assign n35068 = n35049 & ~n35066 ;
  assign n35069 = n35067 | n35068 ;
  assign n35070 = n34813 | n34833 ;
  assign n35071 = ( ~n34811 & n34833 ) | ( ~n34811 & n35070 ) | ( n34833 & n35070 ) ;
  assign n35072 = ( n34814 & ~n34816 ) | ( n34814 & n35071 ) | ( ~n34816 & n35071 ) ;
  assign n35073 = ~n35069 & n35072 ;
  assign n35074 = n35069 & ~n35072 ;
  assign n35075 = n35073 | n35074 ;
  assign n35076 = x123 & n8724 ;
  assign n35077 = x122 & n8719 ;
  assign n35078 = x121 & ~n8718 ;
  assign n35079 = n9149 & n35078 ;
  assign n35080 = n35077 | n35079 ;
  assign n35081 = n35076 | n35080 ;
  assign n35082 = n8727 | n35076 ;
  assign n35083 = n35080 | n35082 ;
  assign n35084 = ( n16086 & n35081 ) | ( n16086 & n35083 ) | ( n35081 & n35083 ) ;
  assign n35085 = x44 & n35083 ;
  assign n35086 = x44 & n35076 ;
  assign n35087 = ( x44 & n35080 ) | ( x44 & n35086 ) | ( n35080 & n35086 ) ;
  assign n35088 = ( n16086 & n35085 ) | ( n16086 & n35087 ) | ( n35085 & n35087 ) ;
  assign n35089 = x44 & ~n35087 ;
  assign n35090 = x44 & ~n35083 ;
  assign n35091 = ( ~n16086 & n35089 ) | ( ~n16086 & n35090 ) | ( n35089 & n35090 ) ;
  assign n35092 = ( n35084 & ~n35088 ) | ( n35084 & n35091 ) | ( ~n35088 & n35091 ) ;
  assign n35093 = n35075 | n35092 ;
  assign n35094 = n35075 & ~n35092 ;
  assign n35095 = ( ~n35075 & n35093 ) | ( ~n35075 & n35094 ) | ( n35093 & n35094 ) ;
  assign n35096 = n34838 | n34860 ;
  assign n35097 = n34835 & ~n34860 ;
  assign n35098 = ( n34839 & n35096 ) | ( n34839 & ~n35097 ) | ( n35096 & ~n35097 ) ;
  assign n35099 = ( n34840 & ~n34843 ) | ( n34840 & n35098 ) | ( ~n34843 & n35098 ) ;
  assign n35100 = n35095 & ~n35099 ;
  assign n35101 = ~n35095 & n35099 ;
  assign n35102 = n35100 | n35101 ;
  assign n35103 = x126 & n7566 ;
  assign n35104 = x125 & n7561 ;
  assign n35105 = x124 & ~n7560 ;
  assign n35106 = n7953 & n35105 ;
  assign n35107 = n35104 | n35106 ;
  assign n35108 = n35103 | n35107 ;
  assign n35109 = n7569 | n35103 ;
  assign n35110 = n35107 | n35109 ;
  assign n35111 = ( n18220 & n35108 ) | ( n18220 & n35110 ) | ( n35108 & n35110 ) ;
  assign n35112 = x41 & n35110 ;
  assign n35113 = x41 & n35103 ;
  assign n35114 = ( x41 & n35107 ) | ( x41 & n35113 ) | ( n35107 & n35113 ) ;
  assign n35115 = ( n18220 & n35112 ) | ( n18220 & n35114 ) | ( n35112 & n35114 ) ;
  assign n35116 = x41 & ~n35114 ;
  assign n35117 = x41 & ~n35110 ;
  assign n35118 = ( ~n18220 & n35116 ) | ( ~n18220 & n35117 ) | ( n35116 & n35117 ) ;
  assign n35119 = ( n35111 & ~n35115 ) | ( n35111 & n35118 ) | ( ~n35115 & n35118 ) ;
  assign n35120 = n35102 & n35119 ;
  assign n35121 = n35095 & ~n35119 ;
  assign n35122 = ( n35099 & n35119 ) | ( n35099 & ~n35121 ) | ( n35119 & ~n35121 ) ;
  assign n35123 = n35100 | n35122 ;
  assign n35124 = ~n35120 & n35123 ;
  assign n35125 = n34919 & ~n34921 ;
  assign n35126 = n35124 & n35125 ;
  assign n35127 = ( n34923 & n35124 ) | ( n34923 & n35126 ) | ( n35124 & n35126 ) ;
  assign n35128 = n35124 | n35125 ;
  assign n35129 = n34923 | n35128 ;
  assign n35130 = ~n35127 & n35129 ;
  assign n35131 = n34658 & ~n34871 ;
  assign n35132 = ~n34658 & n34871 ;
  assign n35133 = n35131 | n35132 ;
  assign n35134 = ~n34675 & n35133 ;
  assign n35135 = ( n34675 & n34679 ) | ( n34675 & ~n35134 ) | ( n34679 & ~n35134 ) ;
  assign n35136 = ~n35130 & n35135 ;
  assign n35137 = n35130 & ~n35135 ;
  assign n35138 = n35136 | n35137 ;
  assign n35139 = ~n34879 & n34894 ;
  assign n35140 = ~n34879 & n34880 ;
  assign n35141 = ( n34879 & n34883 ) | ( n34879 & ~n35140 ) | ( n34883 & ~n35140 ) ;
  assign n35142 = ( n34357 & n35139 ) | ( n34357 & ~n35141 ) | ( n35139 & ~n35141 ) ;
  assign n35143 = ~n34879 & n34897 ;
  assign n35144 = n34879 | n34893 ;
  assign n35145 = ( n34627 & ~n35143 ) | ( n34627 & n35144 ) | ( ~n35143 & n35144 ) ;
  assign n35146 = ( ~n34879 & n34888 ) | ( ~n34879 & n35140 ) | ( n34888 & n35140 ) ;
  assign n35147 = ( n33472 & ~n35145 ) | ( n33472 & n35146 ) | ( ~n35145 & n35146 ) ;
  assign n35148 = ( ~n30754 & n35142 ) | ( ~n30754 & n35147 ) | ( n35142 & n35147 ) ;
  assign n35149 = n35138 & n35148 ;
  assign n35150 = n35138 | n35140 ;
  assign n35151 = n34879 & ~n35138 ;
  assign n35152 = ( n34883 & ~n35150 ) | ( n34883 & n35151 ) | ( ~n35150 & n35151 ) ;
  assign n35153 = ( n34894 & n35138 ) | ( n34894 & ~n35151 ) | ( n35138 & ~n35151 ) ;
  assign n35154 = ( n34357 & ~n35152 ) | ( n34357 & n35153 ) | ( ~n35152 & n35153 ) ;
  assign n35155 = n35138 | n35143 ;
  assign n35156 = ~n35138 & n35144 ;
  assign n35157 = ( n34627 & ~n35155 ) | ( n34627 & n35156 ) | ( ~n35155 & n35156 ) ;
  assign n35158 = ( n34888 & n35150 ) | ( n34888 & ~n35151 ) | ( n35150 & ~n35151 ) ;
  assign n35159 = ( n33472 & ~n35157 ) | ( n33472 & n35158 ) | ( ~n35157 & n35158 ) ;
  assign n35160 = ( ~n30754 & n35154 ) | ( ~n30754 & n35159 ) | ( n35154 & n35159 ) ;
  assign n35161 = ~n35149 & n35160 ;
  assign n35162 = n34958 | n34978 ;
  assign n35163 = ( ~n34941 & n34978 ) | ( ~n34941 & n35162 ) | ( n34978 & n35162 ) ;
  assign n35164 = ( n34959 & ~n34961 ) | ( n34959 & n35163 ) | ( ~n34961 & n35163 ) ;
  assign n35165 = x103 & n18290 ;
  assign n35166 = x63 & x102 ;
  assign n35167 = ~n18290 & n35166 ;
  assign n35168 = n35165 | n35167 ;
  assign n35169 = x38 & n34702 ;
  assign n35170 = x38 | n34702 ;
  assign n35171 = ~n35169 & n35170 ;
  assign n35172 = n35168 & ~n35171 ;
  assign n35173 = ~n35168 & n35171 ;
  assign n35174 = n35172 | n35173 ;
  assign n35175 = ~n34928 & n34931 ;
  assign n35176 = n34703 | n34928 ;
  assign n35177 = ( n34928 & ~n34931 ) | ( n34928 & n35176 ) | ( ~n34931 & n35176 ) ;
  assign n35178 = ~n35175 & n35177 ;
  assign n35179 = ~n35174 & n35178 ;
  assign n35180 = ( n34706 & n35175 ) | ( n34706 & ~n35177 ) | ( n35175 & ~n35177 ) ;
  assign n35181 = n35174 | n35180 ;
  assign n35182 = ( n34697 & n35179 ) | ( n34697 & ~n35181 ) | ( n35179 & ~n35181 ) ;
  assign n35183 = n35174 & ~n35178 ;
  assign n35184 = n35174 & n35180 ;
  assign n35185 = ( ~n34697 & n35183 ) | ( ~n34697 & n35184 ) | ( n35183 & n35184 ) ;
  assign n35186 = n35182 | n35185 ;
  assign n35187 = x106 & n17146 ;
  assign n35188 = x105 & n17141 ;
  assign n35189 = x104 & ~n17140 ;
  assign n35190 = n17724 & n35189 ;
  assign n35191 = n35188 | n35190 ;
  assign n35192 = n35187 | n35191 ;
  assign n35193 = n17149 | n35187 ;
  assign n35194 = n35191 | n35193 ;
  assign n35195 = ( n8656 & n35192 ) | ( n8656 & n35194 ) | ( n35192 & n35194 ) ;
  assign n35196 = x62 & n35194 ;
  assign n35197 = x62 & n35187 ;
  assign n35198 = ( x62 & n35191 ) | ( x62 & n35197 ) | ( n35191 & n35197 ) ;
  assign n35199 = ( n8656 & n35196 ) | ( n8656 & n35198 ) | ( n35196 & n35198 ) ;
  assign n35200 = x62 & ~n35198 ;
  assign n35201 = x62 & ~n35194 ;
  assign n35202 = ( ~n8656 & n35200 ) | ( ~n8656 & n35201 ) | ( n35200 & n35201 ) ;
  assign n35203 = ( n35195 & ~n35199 ) | ( n35195 & n35202 ) | ( ~n35199 & n35202 ) ;
  assign n35204 = ~n35186 & n35203 ;
  assign n35205 = n35186 | n35204 ;
  assign n35206 = x109 & n15552 ;
  assign n35207 = x108 & n15547 ;
  assign n35208 = x107 & ~n15546 ;
  assign n35209 = n16123 & n35208 ;
  assign n35210 = n35207 | n35209 ;
  assign n35211 = n35206 | n35210 ;
  assign n35212 = n15555 | n35206 ;
  assign n35213 = n35210 | n35212 ;
  assign n35214 = ( n9878 & n35211 ) | ( n9878 & n35213 ) | ( n35211 & n35213 ) ;
  assign n35215 = x59 & n35213 ;
  assign n35216 = x59 & n35206 ;
  assign n35217 = ( x59 & n35210 ) | ( x59 & n35216 ) | ( n35210 & n35216 ) ;
  assign n35218 = ( n9878 & n35215 ) | ( n9878 & n35217 ) | ( n35215 & n35217 ) ;
  assign n35219 = x59 & ~n35217 ;
  assign n35220 = x59 & ~n35213 ;
  assign n35221 = ( ~n9878 & n35219 ) | ( ~n9878 & n35220 ) | ( n35219 & n35220 ) ;
  assign n35222 = ( n35214 & ~n35218 ) | ( n35214 & n35221 ) | ( ~n35218 & n35221 ) ;
  assign n35223 = n35203 & n35222 ;
  assign n35224 = n35186 & n35223 ;
  assign n35225 = ( ~n35205 & n35222 ) | ( ~n35205 & n35224 ) | ( n35222 & n35224 ) ;
  assign n35226 = n35203 | n35222 ;
  assign n35227 = ( n35186 & n35222 ) | ( n35186 & n35226 ) | ( n35222 & n35226 ) ;
  assign n35228 = n35205 & ~n35227 ;
  assign n35229 = n35225 | n35228 ;
  assign n35230 = n35164 & n35229 ;
  assign n35231 = n35164 | n35229 ;
  assign n35232 = ~n35230 & n35231 ;
  assign n35233 = x112 & n14045 ;
  assign n35234 = x111 & n14040 ;
  assign n35235 = x110 & ~n14039 ;
  assign n35236 = n14552 & n35235 ;
  assign n35237 = n35234 | n35236 ;
  assign n35238 = n35233 | n35237 ;
  assign n35239 = n14048 | n35233 ;
  assign n35240 = n35237 | n35239 ;
  assign n35241 = ( n11172 & n35238 ) | ( n11172 & n35240 ) | ( n35238 & n35240 ) ;
  assign n35242 = x56 & n35240 ;
  assign n35243 = x56 & n35233 ;
  assign n35244 = ( x56 & n35237 ) | ( x56 & n35243 ) | ( n35237 & n35243 ) ;
  assign n35245 = ( n11172 & n35242 ) | ( n11172 & n35244 ) | ( n35242 & n35244 ) ;
  assign n35246 = x56 & ~n35244 ;
  assign n35247 = x56 & ~n35240 ;
  assign n35248 = ( ~n11172 & n35246 ) | ( ~n11172 & n35247 ) | ( n35246 & n35247 ) ;
  assign n35249 = ( n35241 & ~n35245 ) | ( n35241 & n35248 ) | ( ~n35245 & n35248 ) ;
  assign n35250 = ~n35232 & n35249 ;
  assign n35251 = n35232 & ~n35249 ;
  assign n35252 = n35250 | n35251 ;
  assign n35253 = ( n34984 & ~n34985 ) | ( n34984 & n35004 ) | ( ~n34985 & n35004 ) ;
  assign n35254 = n35252 & ~n35253 ;
  assign n35255 = ~n35252 & n35253 ;
  assign n35256 = n35254 | n35255 ;
  assign n35257 = x115 & n12574 ;
  assign n35258 = x114 & n12569 ;
  assign n35259 = x113 & ~n12568 ;
  assign n35260 = n13076 & n35259 ;
  assign n35261 = n35258 | n35260 ;
  assign n35262 = n35257 | n35261 ;
  assign n35263 = n12577 | n35257 ;
  assign n35264 = n35261 | n35263 ;
  assign n35265 = ( ~n12550 & n35262 ) | ( ~n12550 & n35264 ) | ( n35262 & n35264 ) ;
  assign n35266 = n35262 & n35264 ;
  assign n35267 = ( n12532 & n35265 ) | ( n12532 & n35266 ) | ( n35265 & n35266 ) ;
  assign n35268 = x53 & n35267 ;
  assign n35269 = x53 & ~n35267 ;
  assign n35270 = ( n35267 & ~n35268 ) | ( n35267 & n35269 ) | ( ~n35268 & n35269 ) ;
  assign n35271 = n35256 & ~n35270 ;
  assign n35272 = ~n35256 & n35270 ;
  assign n35273 = n35271 | n35272 ;
  assign n35274 = n35006 & ~n35024 ;
  assign n35275 = ( n35007 & n35024 ) | ( n35007 & ~n35274 ) | ( n35024 & ~n35274 ) ;
  assign n35276 = ( n35009 & ~n35010 ) | ( n35009 & n35275 ) | ( ~n35010 & n35275 ) ;
  assign n35277 = ~n35273 & n35276 ;
  assign n35278 = n35273 & ~n35276 ;
  assign n35279 = n35277 | n35278 ;
  assign n35280 = x118 & n11205 ;
  assign n35281 = x117 & n11200 ;
  assign n35282 = x116 & ~n11199 ;
  assign n35283 = n11679 & n35282 ;
  assign n35284 = n35281 | n35283 ;
  assign n35285 = n35280 | n35284 ;
  assign n35286 = n11208 | n35280 ;
  assign n35287 = n35284 | n35286 ;
  assign n35288 = ( ~n14002 & n35285 ) | ( ~n14002 & n35287 ) | ( n35285 & n35287 ) ;
  assign n35289 = n35285 & n35287 ;
  assign n35290 = ( n13981 & n35288 ) | ( n13981 & n35289 ) | ( n35288 & n35289 ) ;
  assign n35291 = x50 & n35290 ;
  assign n35292 = x50 & ~n35290 ;
  assign n35293 = ( n35290 & ~n35291 ) | ( n35290 & n35292 ) | ( ~n35291 & n35292 ) ;
  assign n35294 = ~n35279 & n35293 ;
  assign n35295 = n35279 & ~n35293 ;
  assign n35296 = n35294 | n35295 ;
  assign n35297 = ~n35027 & n35042 ;
  assign n35298 = n35042 & ~n35297 ;
  assign n35299 = n35027 | n35297 ;
  assign n35300 = ~n35298 & n35299 ;
  assign n35301 = n35041 | n35297 ;
  assign n35302 = ( n35297 & ~n35300 ) | ( n35297 & n35301 ) | ( ~n35300 & n35301 ) ;
  assign n35303 = ~n35296 & n35302 ;
  assign n35304 = n35296 & ~n35302 ;
  assign n35305 = n35303 | n35304 ;
  assign n35306 = x121 & n9933 ;
  assign n35307 = x120 & n9928 ;
  assign n35308 = x119 & ~n9927 ;
  assign n35309 = n10379 & n35308 ;
  assign n35310 = n35307 | n35309 ;
  assign n35311 = n35306 | n35310 ;
  assign n35312 = n9936 | n35306 ;
  assign n35313 = n35310 | n35312 ;
  assign n35314 = ( n15501 & n35311 ) | ( n15501 & n35313 ) | ( n35311 & n35313 ) ;
  assign n35315 = x47 & n35313 ;
  assign n35316 = x47 & n35306 ;
  assign n35317 = ( x47 & n35310 ) | ( x47 & n35316 ) | ( n35310 & n35316 ) ;
  assign n35318 = ( n15501 & n35315 ) | ( n15501 & n35317 ) | ( n35315 & n35317 ) ;
  assign n35319 = x47 & ~n35317 ;
  assign n35320 = x47 & ~n35313 ;
  assign n35321 = ( ~n15501 & n35319 ) | ( ~n15501 & n35320 ) | ( n35319 & n35320 ) ;
  assign n35322 = ( n35314 & ~n35318 ) | ( n35314 & n35321 ) | ( ~n35318 & n35321 ) ;
  assign n35323 = ~n35305 & n35322 ;
  assign n35324 = n35305 | n35323 ;
  assign n35325 = n35045 & ~n35066 ;
  assign n35326 = ( n35046 & n35066 ) | ( n35046 & ~n35325 ) | ( n35066 & ~n35325 ) ;
  assign n35327 = ( n35047 & ~n35049 ) | ( n35047 & n35326 ) | ( ~n35049 & n35326 ) ;
  assign n35328 = n35305 & n35322 ;
  assign n35329 = n35327 & n35328 ;
  assign n35330 = ( ~n35324 & n35327 ) | ( ~n35324 & n35329 ) | ( n35327 & n35329 ) ;
  assign n35331 = n35327 | n35328 ;
  assign n35332 = n35324 & ~n35331 ;
  assign n35333 = n35330 | n35332 ;
  assign n35334 = x124 & n8724 ;
  assign n35335 = x123 & n8719 ;
  assign n35336 = x122 & ~n8718 ;
  assign n35337 = n9149 & n35336 ;
  assign n35338 = n35335 | n35337 ;
  assign n35339 = n35334 | n35338 ;
  assign n35340 = n8727 | n35334 ;
  assign n35341 = n35338 | n35340 ;
  assign n35342 = ( n17084 & n35339 ) | ( n17084 & n35341 ) | ( n35339 & n35341 ) ;
  assign n35343 = x44 & n35341 ;
  assign n35344 = x44 & n35334 ;
  assign n35345 = ( x44 & n35338 ) | ( x44 & n35344 ) | ( n35338 & n35344 ) ;
  assign n35346 = ( n17084 & n35343 ) | ( n17084 & n35345 ) | ( n35343 & n35345 ) ;
  assign n35347 = x44 & ~n35345 ;
  assign n35348 = x44 & ~n35341 ;
  assign n35349 = ( ~n17084 & n35347 ) | ( ~n17084 & n35348 ) | ( n35347 & n35348 ) ;
  assign n35350 = ( n35342 & ~n35346 ) | ( n35342 & n35349 ) | ( ~n35346 & n35349 ) ;
  assign n35351 = ~n35333 & n35350 ;
  assign n35352 = n35333 | n35351 ;
  assign n35353 = n35073 | n35092 ;
  assign n35354 = ( n35073 & ~n35075 ) | ( n35073 & n35353 ) | ( ~n35075 & n35353 ) ;
  assign n35355 = n35333 & n35350 ;
  assign n35356 = n35354 & n35355 ;
  assign n35357 = ( ~n35352 & n35354 ) | ( ~n35352 & n35356 ) | ( n35354 & n35356 ) ;
  assign n35358 = n35354 | n35355 ;
  assign n35359 = n35352 & ~n35358 ;
  assign n35360 = n35357 | n35359 ;
  assign n35361 = x127 & n7566 ;
  assign n35362 = x126 & n7561 ;
  assign n35363 = x125 & ~n7560 ;
  assign n35364 = n7953 & n35363 ;
  assign n35365 = n35362 | n35364 ;
  assign n35366 = n35361 | n35365 ;
  assign n35367 = n7569 | n35361 ;
  assign n35368 = n35365 | n35367 ;
  assign n35369 = ( n18763 & n35366 ) | ( n18763 & n35368 ) | ( n35366 & n35368 ) ;
  assign n35370 = x41 & n35368 ;
  assign n35371 = x41 & n35361 ;
  assign n35372 = ( x41 & n35365 ) | ( x41 & n35371 ) | ( n35365 & n35371 ) ;
  assign n35373 = ( n18763 & n35370 ) | ( n18763 & n35372 ) | ( n35370 & n35372 ) ;
  assign n35374 = x41 & ~n35372 ;
  assign n35375 = x41 & ~n35368 ;
  assign n35376 = ( ~n18763 & n35374 ) | ( ~n18763 & n35375 ) | ( n35374 & n35375 ) ;
  assign n35377 = ( n35369 & ~n35373 ) | ( n35369 & n35376 ) | ( ~n35373 & n35376 ) ;
  assign n35378 = ~n35360 & n35377 ;
  assign n35379 = n35360 | n35378 ;
  assign n35380 = n35360 & n35377 ;
  assign n35381 = n35379 & ~n35380 ;
  assign n35382 = ( n35101 & ~n35102 ) | ( n35101 & n35122 ) | ( ~n35102 & n35122 ) ;
  assign n35383 = n35381 & ~n35382 ;
  assign n35384 = ~n35381 & n35382 ;
  assign n35385 = n35383 | n35384 ;
  assign n35386 = ( n34919 & n34921 ) | ( n34919 & ~n35124 ) | ( n34921 & ~n35124 ) ;
  assign n35387 = ~n35385 & n35386 ;
  assign n35388 = n35385 & ~n35386 ;
  assign n35389 = n35387 | n35388 ;
  assign n35390 = ~n35136 & n35150 ;
  assign n35391 = n35136 | n35151 ;
  assign n35392 = ( n34883 & ~n35390 ) | ( n34883 & n35391 ) | ( ~n35390 & n35391 ) ;
  assign n35393 = ~n35136 & n35138 ;
  assign n35394 = ( n34894 & ~n35391 ) | ( n34894 & n35393 ) | ( ~n35391 & n35393 ) ;
  assign n35395 = ( n34357 & ~n35392 ) | ( n34357 & n35394 ) | ( ~n35392 & n35394 ) ;
  assign n35396 = ~n35136 & n35155 ;
  assign n35397 = n35136 | n35156 ;
  assign n35398 = ( n34627 & ~n35396 ) | ( n34627 & n35397 ) | ( ~n35396 & n35397 ) ;
  assign n35399 = ( n34888 & n35390 ) | ( n34888 & ~n35391 ) | ( n35390 & ~n35391 ) ;
  assign n35400 = ( n33472 & ~n35398 ) | ( n33472 & n35399 ) | ( ~n35398 & n35399 ) ;
  assign n35401 = ( ~n30754 & n35395 ) | ( ~n30754 & n35400 ) | ( n35395 & n35400 ) ;
  assign n35402 = n35389 & n35401 ;
  assign n35403 = ~n35389 & n35392 ;
  assign n35404 = ~n35389 & n35391 ;
  assign n35405 = n35389 | n35393 ;
  assign n35406 = ( n34894 & ~n35404 ) | ( n34894 & n35405 ) | ( ~n35404 & n35405 ) ;
  assign n35407 = ( n34357 & ~n35403 ) | ( n34357 & n35406 ) | ( ~n35403 & n35406 ) ;
  assign n35408 = n35389 | n35396 ;
  assign n35409 = ~n35389 & n35397 ;
  assign n35410 = ( n34627 & ~n35408 ) | ( n34627 & n35409 ) | ( ~n35408 & n35409 ) ;
  assign n35411 = n35389 | n35390 ;
  assign n35412 = ( n34888 & ~n35404 ) | ( n34888 & n35411 ) | ( ~n35404 & n35411 ) ;
  assign n35413 = ( n33468 & ~n35410 ) | ( n33468 & n35412 ) | ( ~n35410 & n35412 ) ;
  assign n35414 = ( n33471 & n35410 ) | ( n33471 & ~n35412 ) | ( n35410 & ~n35412 ) ;
  assign n35415 = ( n32151 & n35413 ) | ( n32151 & ~n35414 ) | ( n35413 & ~n35414 ) ;
  assign n35416 = ( ~n30754 & n35407 ) | ( ~n30754 & n35415 ) | ( n35407 & n35415 ) ;
  assign n35417 = ~n35402 & n35416 ;
  assign n35418 = x125 & n8724 ;
  assign n35419 = x124 & n8719 ;
  assign n35420 = x123 & ~n8718 ;
  assign n35421 = n9149 & n35420 ;
  assign n35422 = n35419 | n35421 ;
  assign n35423 = n35418 | n35422 ;
  assign n35424 = n8727 | n35418 ;
  assign n35425 = n35422 | n35424 ;
  assign n35426 = ( n17670 & n35423 ) | ( n17670 & n35425 ) | ( n35423 & n35425 ) ;
  assign n35427 = x44 & n35425 ;
  assign n35428 = x44 & n35418 ;
  assign n35429 = ( x44 & n35422 ) | ( x44 & n35428 ) | ( n35422 & n35428 ) ;
  assign n35430 = ( n17670 & n35427 ) | ( n17670 & n35429 ) | ( n35427 & n35429 ) ;
  assign n35431 = x44 & ~n35429 ;
  assign n35432 = x44 & ~n35425 ;
  assign n35433 = ( ~n17670 & n35431 ) | ( ~n17670 & n35432 ) | ( n35431 & n35432 ) ;
  assign n35434 = ( n35426 & ~n35430 ) | ( n35426 & n35433 ) | ( ~n35430 & n35433 ) ;
  assign n35435 = x127 & n7561 ;
  assign n35436 = x126 & ~n7560 ;
  assign n35437 = n7953 & n35436 ;
  assign n35438 = n35435 | n35437 ;
  assign n35439 = n7569 | n35438 ;
  assign n35440 = ( n19328 & n35438 ) | ( n19328 & n35439 ) | ( n35438 & n35439 ) ;
  assign n35441 = x41 & n35438 ;
  assign n35442 = ( x41 & n10426 ) | ( x41 & n35438 ) | ( n10426 & n35438 ) ;
  assign n35443 = ( n19328 & n35441 ) | ( n19328 & n35442 ) | ( n35441 & n35442 ) ;
  assign n35444 = x41 & ~n10426 ;
  assign n35445 = ~n35438 & n35444 ;
  assign n35446 = x41 & ~n35438 ;
  assign n35447 = ( ~n19328 & n35445 ) | ( ~n19328 & n35446 ) | ( n35445 & n35446 ) ;
  assign n35448 = ( n35440 & ~n35443 ) | ( n35440 & n35447 ) | ( ~n35443 & n35447 ) ;
  assign n35449 = n35350 & n35448 ;
  assign n35450 = ~n35333 & n35449 ;
  assign n35451 = ( n35357 & n35448 ) | ( n35357 & n35450 ) | ( n35448 & n35450 ) ;
  assign n35452 = n35350 | n35448 ;
  assign n35453 = ( ~n35333 & n35448 ) | ( ~n35333 & n35452 ) | ( n35448 & n35452 ) ;
  assign n35454 = n35357 | n35453 ;
  assign n35455 = ~n35451 & n35454 ;
  assign n35456 = n35323 | n35330 ;
  assign n35457 = x104 & n18290 ;
  assign n35458 = x63 & x103 ;
  assign n35459 = ~n18290 & n35458 ;
  assign n35460 = n35457 | n35459 ;
  assign n35461 = ( ~x38 & n34702 ) | ( ~x38 & n35168 ) | ( n34702 & n35168 ) ;
  assign n35462 = ~n35460 & n35461 ;
  assign n35463 = n35460 & ~n35461 ;
  assign n35464 = n35462 | n35463 ;
  assign n35466 = x106 & n17141 ;
  assign n35467 = x105 & ~n17140 ;
  assign n35468 = n17724 & n35467 ;
  assign n35469 = n35466 | n35468 ;
  assign n35465 = x107 & n17146 ;
  assign n35471 = n17149 | n35465 ;
  assign n35472 = n35469 | n35471 ;
  assign n35470 = n35465 | n35469 ;
  assign n35473 = n35470 & n35472 ;
  assign n35474 = ( n9084 & n35472 ) | ( n9084 & n35473 ) | ( n35472 & n35473 ) ;
  assign n35475 = x62 & n35473 ;
  assign n35476 = x62 & n35472 ;
  assign n35477 = ( n9084 & n35475 ) | ( n9084 & n35476 ) | ( n35475 & n35476 ) ;
  assign n35478 = x62 & ~n35473 ;
  assign n35479 = x62 & ~n35472 ;
  assign n35480 = ( ~n9084 & n35478 ) | ( ~n9084 & n35479 ) | ( n35478 & n35479 ) ;
  assign n35481 = ( n35474 & ~n35477 ) | ( n35474 & n35480 ) | ( ~n35477 & n35480 ) ;
  assign n35482 = ~n35464 & n35481 ;
  assign n35483 = n35464 & ~n35481 ;
  assign n35484 = n35482 | n35483 ;
  assign n35485 = n35182 | n35203 ;
  assign n35486 = ( n35182 & ~n35186 ) | ( n35182 & n35485 ) | ( ~n35186 & n35485 ) ;
  assign n35487 = ~n35484 & n35486 ;
  assign n35488 = n35484 & ~n35486 ;
  assign n35489 = n35487 | n35488 ;
  assign n35490 = x110 & n15552 ;
  assign n35491 = x109 & n15547 ;
  assign n35492 = x108 & ~n15546 ;
  assign n35493 = n16123 & n35492 ;
  assign n35494 = n35491 | n35493 ;
  assign n35495 = n35490 | n35494 ;
  assign n35496 = n15555 | n35490 ;
  assign n35497 = n35494 | n35496 ;
  assign n35498 = ( n10330 & n35495 ) | ( n10330 & n35497 ) | ( n35495 & n35497 ) ;
  assign n35499 = x59 & n35497 ;
  assign n35500 = x59 & n35490 ;
  assign n35501 = ( x59 & n35494 ) | ( x59 & n35500 ) | ( n35494 & n35500 ) ;
  assign n35502 = ( n10330 & n35499 ) | ( n10330 & n35501 ) | ( n35499 & n35501 ) ;
  assign n35503 = x59 & ~n35501 ;
  assign n35504 = x59 & ~n35497 ;
  assign n35505 = ( ~n10330 & n35503 ) | ( ~n10330 & n35504 ) | ( n35503 & n35504 ) ;
  assign n35506 = ( n35498 & ~n35502 ) | ( n35498 & n35505 ) | ( ~n35502 & n35505 ) ;
  assign n35507 = n35489 | n35506 ;
  assign n35508 = n35489 & ~n35506 ;
  assign n35509 = ( ~n35489 & n35507 ) | ( ~n35489 & n35508 ) | ( n35507 & n35508 ) ;
  assign n35510 = n35164 | n35225 ;
  assign n35511 = ( n35225 & ~n35229 ) | ( n35225 & n35510 ) | ( ~n35229 & n35510 ) ;
  assign n35512 = n35509 & ~n35511 ;
  assign n35513 = ~n35509 & n35511 ;
  assign n35514 = n35512 | n35513 ;
  assign n35515 = x113 & n14045 ;
  assign n35516 = x112 & n14040 ;
  assign n35517 = x111 & ~n14039 ;
  assign n35518 = n14552 & n35517 ;
  assign n35519 = n35516 | n35518 ;
  assign n35520 = n35515 | n35519 ;
  assign n35521 = n14048 | n35515 ;
  assign n35522 = n35519 | n35521 ;
  assign n35523 = ( ~n11642 & n35520 ) | ( ~n11642 & n35522 ) | ( n35520 & n35522 ) ;
  assign n35524 = n35520 & n35522 ;
  assign n35525 = ( n11626 & n35523 ) | ( n11626 & n35524 ) | ( n35523 & n35524 ) ;
  assign n35526 = x56 & n35525 ;
  assign n35527 = x56 & ~n35525 ;
  assign n35528 = ( n35525 & ~n35526 ) | ( n35525 & n35527 ) | ( ~n35526 & n35527 ) ;
  assign n35529 = n35514 & n35528 ;
  assign n35530 = n35513 | n35528 ;
  assign n35531 = n35512 | n35530 ;
  assign n35532 = ~n35529 & n35531 ;
  assign n35533 = n35250 | n35253 ;
  assign n35534 = ( n35250 & ~n35252 ) | ( n35250 & n35533 ) | ( ~n35252 & n35533 ) ;
  assign n35535 = n35532 & ~n35534 ;
  assign n35536 = ~n35532 & n35534 ;
  assign n35537 = n35535 | n35536 ;
  assign n35538 = x116 & n12574 ;
  assign n35539 = x115 & n12569 ;
  assign n35540 = x114 & ~n12568 ;
  assign n35541 = n13076 & n35540 ;
  assign n35542 = n35539 | n35541 ;
  assign n35543 = n35538 | n35542 ;
  assign n35544 = n12577 | n35538 ;
  assign n35545 = n35542 | n35544 ;
  assign n35546 = ( ~n13040 & n35543 ) | ( ~n13040 & n35545 ) | ( n35543 & n35545 ) ;
  assign n35547 = n35543 & n35545 ;
  assign n35548 = ( n13022 & n35546 ) | ( n13022 & n35547 ) | ( n35546 & n35547 ) ;
  assign n35549 = x53 & n35548 ;
  assign n35550 = x53 & ~n35548 ;
  assign n35551 = ( n35548 & ~n35549 ) | ( n35548 & n35550 ) | ( ~n35549 & n35550 ) ;
  assign n35552 = n35537 & n35551 ;
  assign n35553 = n35536 | n35551 ;
  assign n35554 = n35535 | n35553 ;
  assign n35555 = ~n35552 & n35554 ;
  assign n35556 = n35272 | n35277 ;
  assign n35557 = n35555 & n35556 ;
  assign n35558 = n35555 | n35556 ;
  assign n35559 = ~n35557 & n35558 ;
  assign n35560 = x119 & n11205 ;
  assign n35561 = x118 & n11200 ;
  assign n35562 = x117 & ~n11199 ;
  assign n35563 = n11679 & n35562 ;
  assign n35564 = n35561 | n35563 ;
  assign n35565 = n35560 | n35564 ;
  assign n35566 = n11208 | n35560 ;
  assign n35567 = n35564 | n35566 ;
  assign n35568 = ( n14496 & n35565 ) | ( n14496 & n35567 ) | ( n35565 & n35567 ) ;
  assign n35569 = x50 & n35567 ;
  assign n35570 = x50 & n35560 ;
  assign n35571 = ( x50 & n35564 ) | ( x50 & n35570 ) | ( n35564 & n35570 ) ;
  assign n35572 = ( n14496 & n35569 ) | ( n14496 & n35571 ) | ( n35569 & n35571 ) ;
  assign n35573 = x50 & ~n35571 ;
  assign n35574 = x50 & ~n35567 ;
  assign n35575 = ( ~n14496 & n35573 ) | ( ~n14496 & n35574 ) | ( n35573 & n35574 ) ;
  assign n35576 = ( n35568 & ~n35572 ) | ( n35568 & n35575 ) | ( ~n35572 & n35575 ) ;
  assign n35577 = ~n35559 & n35576 ;
  assign n35578 = n35559 & ~n35576 ;
  assign n35579 = n35577 | n35578 ;
  assign n35580 = ~n35294 & n35296 ;
  assign n35581 = ( n35294 & n35302 ) | ( n35294 & ~n35580 ) | ( n35302 & ~n35580 ) ;
  assign n35582 = n35579 & ~n35581 ;
  assign n35583 = ~n35579 & n35581 ;
  assign n35584 = x122 & n9933 ;
  assign n35585 = x121 & n9928 ;
  assign n35586 = x120 & ~n9927 ;
  assign n35587 = n10379 & n35586 ;
  assign n35588 = n35585 | n35587 ;
  assign n35589 = n35584 | n35588 ;
  assign n35590 = n9936 | n35584 ;
  assign n35591 = n35588 | n35590 ;
  assign n35592 = ( n16043 & n35589 ) | ( n16043 & n35591 ) | ( n35589 & n35591 ) ;
  assign n35593 = x47 & n35591 ;
  assign n35594 = x47 & n35584 ;
  assign n35595 = ( x47 & n35588 ) | ( x47 & n35594 ) | ( n35588 & n35594 ) ;
  assign n35596 = ( n16043 & n35593 ) | ( n16043 & n35595 ) | ( n35593 & n35595 ) ;
  assign n35597 = x47 & ~n35595 ;
  assign n35598 = x47 & ~n35591 ;
  assign n35599 = ( ~n16043 & n35597 ) | ( ~n16043 & n35598 ) | ( n35597 & n35598 ) ;
  assign n35600 = ( n35592 & ~n35596 ) | ( n35592 & n35599 ) | ( ~n35596 & n35599 ) ;
  assign n35601 = n35583 | n35600 ;
  assign n35602 = n35582 | n35601 ;
  assign n35603 = n35582 | n35583 ;
  assign n35604 = n35600 & n35603 ;
  assign n35605 = n35323 & n35604 ;
  assign n35606 = ( n35330 & n35604 ) | ( n35330 & n35605 ) | ( n35604 & n35605 ) ;
  assign n35607 = ( n35456 & ~n35602 ) | ( n35456 & n35606 ) | ( ~n35602 & n35606 ) ;
  assign n35608 = n35323 | n35604 ;
  assign n35609 = n35330 | n35608 ;
  assign n35610 = n35602 & ~n35609 ;
  assign n35611 = n35607 | n35610 ;
  assign n35612 = ( n35434 & n35455 ) | ( n35434 & ~n35611 ) | ( n35455 & ~n35611 ) ;
  assign n35613 = ( ~n35455 & n35611 ) | ( ~n35455 & n35612 ) | ( n35611 & n35612 ) ;
  assign n35614 = ( ~n35434 & n35612 ) | ( ~n35434 & n35613 ) | ( n35612 & n35613 ) ;
  assign n35615 = n35378 | n35382 ;
  assign n35616 = ( n35378 & ~n35381 ) | ( n35378 & n35615 ) | ( ~n35381 & n35615 ) ;
  assign n35617 = n35614 & ~n35616 ;
  assign n35618 = ~n35614 & n35616 ;
  assign n35619 = n35617 | n35618 ;
  assign n35620 = ~n35387 & n35415 ;
  assign n35621 = ~n35387 & n35389 ;
  assign n35622 = ( n35387 & n35392 ) | ( n35387 & ~n35621 ) | ( n35392 & ~n35621 ) ;
  assign n35623 = n35387 | n35404 ;
  assign n35624 = ~n35387 & n35405 ;
  assign n35625 = ( n34894 & ~n35623 ) | ( n34894 & n35624 ) | ( ~n35623 & n35624 ) ;
  assign n35626 = ( n34357 & ~n35622 ) | ( n34357 & n35625 ) | ( ~n35622 & n35625 ) ;
  assign n35627 = ( ~n30754 & n35620 ) | ( ~n30754 & n35626 ) | ( n35620 & n35626 ) ;
  assign n35628 = n35619 & n35627 ;
  assign n35629 = n35619 | n35625 ;
  assign n35630 = n35387 & ~n35619 ;
  assign n35631 = n35619 | n35621 ;
  assign n35632 = ( n35392 & n35630 ) | ( n35392 & ~n35631 ) | ( n35630 & ~n35631 ) ;
  assign n35633 = ( n34357 & n35629 ) | ( n34357 & ~n35632 ) | ( n35629 & ~n35632 ) ;
  assign n35634 = ( n35415 & n35619 ) | ( n35415 & ~n35630 ) | ( n35619 & ~n35630 ) ;
  assign n35635 = ( ~n30754 & n35633 ) | ( ~n30754 & n35634 ) | ( n35633 & n35634 ) ;
  assign n35636 = ~n35628 & n35635 ;
  assign n35741 = ( n35536 & ~n35537 ) | ( n35536 & n35553 ) | ( ~n35537 & n35553 ) ;
  assign n35718 = ( n35513 & ~n35514 ) | ( n35513 & n35530 ) | ( ~n35514 & n35530 ) ;
  assign n35637 = x108 & n17146 ;
  assign n35638 = x107 & n17141 ;
  assign n35639 = x106 & ~n17140 ;
  assign n35640 = n17724 & n35639 ;
  assign n35641 = n35638 | n35640 ;
  assign n35642 = n35637 | n35641 ;
  assign n35643 = n17149 | n35637 ;
  assign n35644 = n35641 | n35643 ;
  assign n35645 = ( n9479 & n35642 ) | ( n9479 & n35644 ) | ( n35642 & n35644 ) ;
  assign n35646 = x62 & n35644 ;
  assign n35647 = x62 & n35637 ;
  assign n35648 = ( x62 & n35641 ) | ( x62 & n35647 ) | ( n35641 & n35647 ) ;
  assign n35649 = ( n9479 & n35646 ) | ( n9479 & n35648 ) | ( n35646 & n35648 ) ;
  assign n35650 = x62 & ~n35648 ;
  assign n35651 = x62 & ~n35644 ;
  assign n35652 = ( ~n9479 & n35650 ) | ( ~n9479 & n35651 ) | ( n35650 & n35651 ) ;
  assign n35653 = ( n35645 & ~n35649 ) | ( n35645 & n35652 ) | ( ~n35649 & n35652 ) ;
  assign n35654 = ~n35462 & n35464 ;
  assign n35655 = x105 & n18290 ;
  assign n35656 = x63 & x104 ;
  assign n35657 = ~n18290 & n35656 ;
  assign n35658 = n35655 | n35657 ;
  assign n35659 = ~n35460 & n35658 ;
  assign n35660 = n35460 | n35659 ;
  assign n35661 = n35658 & ~n35659 ;
  assign n35662 = n35660 & ~n35661 ;
  assign n35663 = n35654 & ~n35662 ;
  assign n35664 = n35462 | n35662 ;
  assign n35665 = ( n35481 & ~n35663 ) | ( n35481 & n35664 ) | ( ~n35663 & n35664 ) ;
  assign n35666 = n35653 | n35665 ;
  assign n35667 = n35654 | n35662 ;
  assign n35668 = n35462 & ~n35662 ;
  assign n35669 = ( n35481 & ~n35667 ) | ( n35481 & n35668 ) | ( ~n35667 & n35668 ) ;
  assign n35670 = ( n35462 & n35482 ) | ( n35462 & ~n35669 ) | ( n35482 & ~n35669 ) ;
  assign n35671 = ( n35653 & n35666 ) | ( n35653 & ~n35670 ) | ( n35666 & ~n35670 ) ;
  assign n35672 = n35653 & n35665 ;
  assign n35673 = ~n35670 & n35672 ;
  assign n35674 = n35671 & ~n35673 ;
  assign n35675 = x111 & n15552 ;
  assign n35676 = x110 & n15547 ;
  assign n35677 = x109 & ~n15546 ;
  assign n35678 = n16123 & n35677 ;
  assign n35679 = n35676 | n35678 ;
  assign n35680 = n35675 | n35679 ;
  assign n35681 = n15555 | n35675 ;
  assign n35682 = n35679 | n35681 ;
  assign n35683 = ( n10749 & n35680 ) | ( n10749 & n35682 ) | ( n35680 & n35682 ) ;
  assign n35684 = x59 & n35682 ;
  assign n35685 = x59 & n35675 ;
  assign n35686 = ( x59 & n35679 ) | ( x59 & n35685 ) | ( n35679 & n35685 ) ;
  assign n35687 = ( n10749 & n35684 ) | ( n10749 & n35686 ) | ( n35684 & n35686 ) ;
  assign n35688 = x59 & ~n35686 ;
  assign n35689 = x59 & ~n35682 ;
  assign n35690 = ( ~n10749 & n35688 ) | ( ~n10749 & n35689 ) | ( n35688 & n35689 ) ;
  assign n35691 = ( n35683 & ~n35687 ) | ( n35683 & n35690 ) | ( ~n35687 & n35690 ) ;
  assign n35692 = ~n35674 & n35691 ;
  assign n35693 = n35674 & ~n35691 ;
  assign n35694 = n35692 | n35693 ;
  assign n35695 = n35484 & ~n35506 ;
  assign n35696 = ( n35486 & n35506 ) | ( n35486 & ~n35695 ) | ( n35506 & ~n35695 ) ;
  assign n35697 = ( n35487 & ~n35489 ) | ( n35487 & n35696 ) | ( ~n35489 & n35696 ) ;
  assign n35698 = n35694 & ~n35697 ;
  assign n35699 = ~n35694 & n35697 ;
  assign n35700 = n35698 | n35699 ;
  assign n35701 = x114 & n14045 ;
  assign n35702 = x113 & n14040 ;
  assign n35703 = x112 & ~n14039 ;
  assign n35704 = n14552 & n35703 ;
  assign n35705 = n35702 | n35704 ;
  assign n35706 = n35701 | n35705 ;
  assign n35707 = n14048 | n35701 ;
  assign n35708 = n35705 | n35707 ;
  assign n35709 = ( ~n12095 & n35706 ) | ( ~n12095 & n35708 ) | ( n35706 & n35708 ) ;
  assign n35710 = n35706 & n35708 ;
  assign n35711 = ( n12079 & n35709 ) | ( n12079 & n35710 ) | ( n35709 & n35710 ) ;
  assign n35712 = x56 & n35711 ;
  assign n35713 = x56 & ~n35711 ;
  assign n35714 = ( n35711 & ~n35712 ) | ( n35711 & n35713 ) | ( ~n35712 & n35713 ) ;
  assign n35715 = n35700 & ~n35714 ;
  assign n35716 = ~n35700 & n35714 ;
  assign n35717 = n35715 | n35716 ;
  assign n35719 = ~n35717 & n35718 ;
  assign n35720 = n35718 & ~n35719 ;
  assign n35721 = n35717 | n35718 ;
  assign n35722 = x117 & n12574 ;
  assign n35723 = x116 & n12569 ;
  assign n35724 = x115 & ~n12568 ;
  assign n35725 = n13076 & n35724 ;
  assign n35726 = n35723 | n35725 ;
  assign n35727 = n35722 | n35726 ;
  assign n35728 = n12577 | n35722 ;
  assign n35729 = n35726 | n35728 ;
  assign n35730 = ( ~n13522 & n35727 ) | ( ~n13522 & n35729 ) | ( n35727 & n35729 ) ;
  assign n35731 = n35727 & n35729 ;
  assign n35732 = ( n13503 & n35730 ) | ( n13503 & n35731 ) | ( n35730 & n35731 ) ;
  assign n35733 = x53 & n35732 ;
  assign n35734 = x53 & ~n35732 ;
  assign n35735 = ( n35732 & ~n35733 ) | ( n35732 & n35734 ) | ( ~n35733 & n35734 ) ;
  assign n35736 = n35721 & ~n35735 ;
  assign n35737 = ~n35720 & n35736 ;
  assign n35738 = ~n35721 & n35735 ;
  assign n35739 = ( n35720 & n35735 ) | ( n35720 & n35738 ) | ( n35735 & n35738 ) ;
  assign n35740 = n35737 | n35739 ;
  assign n35742 = ~n35740 & n35741 ;
  assign n35743 = n35741 & ~n35742 ;
  assign n35744 = n35740 | n35741 ;
  assign n35745 = x120 & n11205 ;
  assign n35746 = x119 & n11200 ;
  assign n35747 = x118 & ~n11199 ;
  assign n35748 = n11679 & n35747 ;
  assign n35749 = n35746 | n35748 ;
  assign n35750 = n35745 | n35749 ;
  assign n35751 = n11208 | n35745 ;
  assign n35752 = n35749 | n35751 ;
  assign n35753 = ( n14991 & n35750 ) | ( n14991 & n35752 ) | ( n35750 & n35752 ) ;
  assign n35754 = x50 & n35752 ;
  assign n35755 = x50 & n35745 ;
  assign n35756 = ( x50 & n35749 ) | ( x50 & n35755 ) | ( n35749 & n35755 ) ;
  assign n35757 = ( n14991 & n35754 ) | ( n14991 & n35756 ) | ( n35754 & n35756 ) ;
  assign n35758 = x50 & ~n35756 ;
  assign n35759 = x50 & ~n35752 ;
  assign n35760 = ( ~n14991 & n35758 ) | ( ~n14991 & n35759 ) | ( n35758 & n35759 ) ;
  assign n35761 = ( n35753 & ~n35757 ) | ( n35753 & n35760 ) | ( ~n35757 & n35760 ) ;
  assign n35762 = n35744 & ~n35761 ;
  assign n35763 = ~n35743 & n35762 ;
  assign n35764 = ~n35744 & n35761 ;
  assign n35765 = ( n35743 & n35761 ) | ( n35743 & n35764 ) | ( n35761 & n35764 ) ;
  assign n35766 = n35763 | n35765 ;
  assign n35767 = ~n35555 & n35556 ;
  assign n35768 = ~n35766 & n35767 ;
  assign n35769 = ( n35577 & ~n35766 ) | ( n35577 & n35768 ) | ( ~n35766 & n35768 ) ;
  assign n35770 = n35766 & ~n35767 ;
  assign n35771 = ~n35577 & n35770 ;
  assign n35772 = n35769 | n35771 ;
  assign n35773 = x123 & n9933 ;
  assign n35774 = x122 & n9928 ;
  assign n35775 = x121 & ~n9927 ;
  assign n35776 = n10379 & n35775 ;
  assign n35777 = n35774 | n35776 ;
  assign n35778 = n35773 | n35777 ;
  assign n35779 = n9936 | n35773 ;
  assign n35780 = n35777 | n35779 ;
  assign n35781 = ( n16086 & n35778 ) | ( n16086 & n35780 ) | ( n35778 & n35780 ) ;
  assign n35782 = x47 & n35780 ;
  assign n35783 = x47 & n35773 ;
  assign n35784 = ( x47 & n35777 ) | ( x47 & n35783 ) | ( n35777 & n35783 ) ;
  assign n35785 = ( n16086 & n35782 ) | ( n16086 & n35784 ) | ( n35782 & n35784 ) ;
  assign n35786 = x47 & ~n35784 ;
  assign n35787 = x47 & ~n35780 ;
  assign n35788 = ( ~n16086 & n35786 ) | ( ~n16086 & n35787 ) | ( n35786 & n35787 ) ;
  assign n35789 = ( n35781 & ~n35785 ) | ( n35781 & n35788 ) | ( ~n35785 & n35788 ) ;
  assign n35790 = n35772 | n35789 ;
  assign n35791 = n35772 & ~n35789 ;
  assign n35792 = ( ~n35772 & n35790 ) | ( ~n35772 & n35791 ) | ( n35790 & n35791 ) ;
  assign n35793 = ( n35583 & n35601 ) | ( n35583 & ~n35603 ) | ( n35601 & ~n35603 ) ;
  assign n35794 = n35792 & ~n35793 ;
  assign n35795 = ~n35792 & n35793 ;
  assign n35796 = n35794 | n35795 ;
  assign n35797 = x126 & n8724 ;
  assign n35798 = x125 & n8719 ;
  assign n35799 = x124 & ~n8718 ;
  assign n35800 = n9149 & n35799 ;
  assign n35801 = n35798 | n35800 ;
  assign n35802 = n35797 | n35801 ;
  assign n35803 = n8727 | n35797 ;
  assign n35804 = n35801 | n35803 ;
  assign n35805 = ( n18220 & n35802 ) | ( n18220 & n35804 ) | ( n35802 & n35804 ) ;
  assign n35806 = x44 & n35804 ;
  assign n35807 = x44 & n35797 ;
  assign n35808 = ( x44 & n35801 ) | ( x44 & n35807 ) | ( n35801 & n35807 ) ;
  assign n35809 = ( n18220 & n35806 ) | ( n18220 & n35808 ) | ( n35806 & n35808 ) ;
  assign n35810 = x44 & ~n35808 ;
  assign n35811 = x44 & ~n35804 ;
  assign n35812 = ( ~n18220 & n35810 ) | ( ~n18220 & n35811 ) | ( n35810 & n35811 ) ;
  assign n35813 = ( n35805 & ~n35809 ) | ( n35805 & n35812 ) | ( ~n35809 & n35812 ) ;
  assign n35814 = n35796 & n35813 ;
  assign n35815 = n35795 | n35813 ;
  assign n35816 = n35794 | n35815 ;
  assign n35817 = ~n35814 & n35816 ;
  assign n35818 = x127 & ~n7560 ;
  assign n35819 = n7953 & n35818 ;
  assign n35820 = n7569 & n19877 ;
  assign n35821 = n35819 | n35820 ;
  assign n35822 = n7569 & n19880 ;
  assign n35823 = n35819 | n35822 ;
  assign n35824 = ( n18202 & n35821 ) | ( n18202 & n35823 ) | ( n35821 & n35823 ) ;
  assign n35825 = n35821 & n35823 ;
  assign n35826 = ( n18212 & n35824 ) | ( n18212 & n35825 ) | ( n35824 & n35825 ) ;
  assign n35827 = ( n18214 & n35824 ) | ( n18214 & n35825 ) | ( n35824 & n35825 ) ;
  assign n35828 = ( n14002 & n35826 ) | ( n14002 & n35827 ) | ( n35826 & n35827 ) ;
  assign n35829 = x41 & n35826 ;
  assign n35830 = x41 & n35827 ;
  assign n35831 = ( n14002 & n35829 ) | ( n14002 & n35830 ) | ( n35829 & n35830 ) ;
  assign n35832 = x41 & ~n35830 ;
  assign n35833 = x41 & ~n35829 ;
  assign n35834 = ( ~n14002 & n35832 ) | ( ~n14002 & n35833 ) | ( n35832 & n35833 ) ;
  assign n35835 = ( n35828 & ~n35831 ) | ( n35828 & n35834 ) | ( ~n35831 & n35834 ) ;
  assign n35836 = n35434 | n35607 ;
  assign n35837 = ( n35607 & ~n35611 ) | ( n35607 & n35836 ) | ( ~n35611 & n35836 ) ;
  assign n35838 = ( n35817 & n35835 ) | ( n35817 & ~n35837 ) | ( n35835 & ~n35837 ) ;
  assign n35839 = ( ~n35835 & n35837 ) | ( ~n35835 & n35838 ) | ( n35837 & n35838 ) ;
  assign n35840 = ( ~n35817 & n35838 ) | ( ~n35817 & n35839 ) | ( n35838 & n35839 ) ;
  assign n35841 = n35434 & ~n35611 ;
  assign n35842 = ~n35434 & n35611 ;
  assign n35843 = n35841 | n35842 ;
  assign n35844 = ~n35451 & n35843 ;
  assign n35845 = ( n35451 & n35455 ) | ( n35451 & ~n35844 ) | ( n35455 & ~n35844 ) ;
  assign n35846 = ~n35840 & n35845 ;
  assign n35847 = n35840 & ~n35845 ;
  assign n35848 = n35846 | n35847 ;
  assign n35849 = n35618 | n35630 ;
  assign n35850 = ~n35618 & n35631 ;
  assign n35851 = ( n35392 & n35849 ) | ( n35392 & ~n35850 ) | ( n35849 & ~n35850 ) ;
  assign n35852 = ~n35618 & n35619 ;
  assign n35853 = ( ~n35618 & n35625 ) | ( ~n35618 & n35852 ) | ( n35625 & n35852 ) ;
  assign n35854 = ( n34357 & ~n35851 ) | ( n34357 & n35853 ) | ( ~n35851 & n35853 ) ;
  assign n35855 = ( n35415 & ~n35849 ) | ( n35415 & n35852 ) | ( ~n35849 & n35852 ) ;
  assign n35856 = ( ~n30754 & n35854 ) | ( ~n30754 & n35855 ) | ( n35854 & n35855 ) ;
  assign n35857 = n35848 & n35856 ;
  assign n35858 = n35848 | n35850 ;
  assign n35859 = n35618 & ~n35848 ;
  assign n35860 = ( n35630 & ~n35848 ) | ( n35630 & n35859 ) | ( ~n35848 & n35859 ) ;
  assign n35861 = ( n35392 & ~n35858 ) | ( n35392 & n35860 ) | ( ~n35858 & n35860 ) ;
  assign n35862 = ( n35619 & n35848 ) | ( n35619 & ~n35859 ) | ( n35848 & ~n35859 ) ;
  assign n35863 = ( n35625 & ~n35859 ) | ( n35625 & n35862 ) | ( ~n35859 & n35862 ) ;
  assign n35864 = ( n34357 & ~n35861 ) | ( n34357 & n35863 ) | ( ~n35861 & n35863 ) ;
  assign n35865 = ( n35415 & ~n35860 ) | ( n35415 & n35862 ) | ( ~n35860 & n35862 ) ;
  assign n35866 = ( ~n30754 & n35864 ) | ( ~n30754 & n35865 ) | ( n35864 & n35865 ) ;
  assign n35867 = ~n35857 & n35866 ;
  assign n35868 = n35742 | n35765 ;
  assign n35869 = n35719 | n35739 ;
  assign n35870 = x41 & n35460 ;
  assign n35871 = x41 | n35460 ;
  assign n35872 = ~n35870 & n35871 ;
  assign n35873 = x106 & n18290 ;
  assign n35874 = x63 & x105 ;
  assign n35875 = ~n18290 & n35874 ;
  assign n35876 = n35873 | n35875 ;
  assign n35877 = n35872 & ~n35876 ;
  assign n35878 = ~n35872 & n35876 ;
  assign n35879 = n35877 | n35878 ;
  assign n35880 = x108 & n17141 ;
  assign n35881 = x107 & ~n17140 ;
  assign n35882 = n17724 & n35881 ;
  assign n35883 = n35880 | n35882 ;
  assign n35884 = x109 & n17146 ;
  assign n35885 = n17149 | n35884 ;
  assign n35886 = n35883 | n35885 ;
  assign n35887 = ~x62 & n35886 ;
  assign n35888 = ~x62 & n35884 ;
  assign n35889 = ( ~x62 & n35883 ) | ( ~x62 & n35888 ) | ( n35883 & n35888 ) ;
  assign n35890 = ( n9878 & n35887 ) | ( n9878 & n35889 ) | ( n35887 & n35889 ) ;
  assign n35891 = x62 & ~n35886 ;
  assign n35892 = x62 & x109 ;
  assign n35893 = n17146 & n35892 ;
  assign n35894 = x62 & ~n35893 ;
  assign n35895 = ~n35883 & n35894 ;
  assign n35896 = ( ~n9878 & n35891 ) | ( ~n9878 & n35895 ) | ( n35891 & n35895 ) ;
  assign n35897 = n35890 | n35896 ;
  assign n35898 = ~n35879 & n35897 ;
  assign n35899 = n35879 & ~n35897 ;
  assign n35900 = n35898 | n35899 ;
  assign n35901 = ~n35659 & n35662 ;
  assign n35902 = ( n35654 & ~n35659 ) | ( n35654 & n35901 ) | ( ~n35659 & n35901 ) ;
  assign n35903 = n35462 | n35659 ;
  assign n35904 = ( n35659 & ~n35662 ) | ( n35659 & n35903 ) | ( ~n35662 & n35903 ) ;
  assign n35905 = ( n35481 & ~n35902 ) | ( n35481 & n35904 ) | ( ~n35902 & n35904 ) ;
  assign n35906 = n35900 & ~n35905 ;
  assign n35907 = ~n35900 & n35905 ;
  assign n35908 = n35906 | n35907 ;
  assign n35909 = x112 & n15552 ;
  assign n35910 = x111 & n15547 ;
  assign n35911 = x110 & ~n15546 ;
  assign n35912 = n16123 & n35911 ;
  assign n35913 = n35910 | n35912 ;
  assign n35914 = n35909 | n35913 ;
  assign n35915 = n15555 | n35909 ;
  assign n35916 = n35913 | n35915 ;
  assign n35917 = ( n11172 & n35914 ) | ( n11172 & n35916 ) | ( n35914 & n35916 ) ;
  assign n35918 = x59 & n35916 ;
  assign n35919 = x59 & n35909 ;
  assign n35920 = ( x59 & n35913 ) | ( x59 & n35919 ) | ( n35913 & n35919 ) ;
  assign n35921 = ( n11172 & n35918 ) | ( n11172 & n35920 ) | ( n35918 & n35920 ) ;
  assign n35922 = x59 & ~n35920 ;
  assign n35923 = x59 & ~n35916 ;
  assign n35924 = ( ~n11172 & n35922 ) | ( ~n11172 & n35923 ) | ( n35922 & n35923 ) ;
  assign n35925 = ( n35917 & ~n35921 ) | ( n35917 & n35924 ) | ( ~n35921 & n35924 ) ;
  assign n35926 = ~n35908 & n35925 ;
  assign n35927 = n35908 | n35926 ;
  assign n35928 = ( n35653 & ~n35665 ) | ( n35653 & n35691 ) | ( ~n35665 & n35691 ) ;
  assign n35929 = n35653 | n35691 ;
  assign n35930 = ( n35670 & n35928 ) | ( n35670 & n35929 ) | ( n35928 & n35929 ) ;
  assign n35931 = n35925 & n35930 ;
  assign n35932 = n35908 & n35931 ;
  assign n35933 = ( ~n35927 & n35930 ) | ( ~n35927 & n35932 ) | ( n35930 & n35932 ) ;
  assign n35934 = n35925 | n35930 ;
  assign n35935 = ( n35908 & n35930 ) | ( n35908 & n35934 ) | ( n35930 & n35934 ) ;
  assign n35936 = n35927 & ~n35935 ;
  assign n35937 = n35933 | n35936 ;
  assign n35938 = x115 & n14045 ;
  assign n35939 = x114 & n14040 ;
  assign n35940 = x113 & ~n14039 ;
  assign n35941 = n14552 & n35940 ;
  assign n35942 = n35939 | n35941 ;
  assign n35943 = n35938 | n35942 ;
  assign n35944 = n14048 | n35938 ;
  assign n35945 = n35942 | n35944 ;
  assign n35946 = ( ~n12550 & n35943 ) | ( ~n12550 & n35945 ) | ( n35943 & n35945 ) ;
  assign n35947 = n35943 & n35945 ;
  assign n35948 = ( n12532 & n35946 ) | ( n12532 & n35947 ) | ( n35946 & n35947 ) ;
  assign n35949 = x56 & n35948 ;
  assign n35950 = x56 & ~n35948 ;
  assign n35951 = ( n35948 & ~n35949 ) | ( n35948 & n35950 ) | ( ~n35949 & n35950 ) ;
  assign n35952 = ~n35937 & n35951 ;
  assign n35953 = n35937 | n35952 ;
  assign n35954 = n35699 | n35714 ;
  assign n35955 = ( n35699 & ~n35700 ) | ( n35699 & n35954 ) | ( ~n35700 & n35954 ) ;
  assign n35956 = n35937 & n35951 ;
  assign n35957 = n35955 & n35956 ;
  assign n35958 = ( ~n35953 & n35955 ) | ( ~n35953 & n35957 ) | ( n35955 & n35957 ) ;
  assign n35959 = n35955 | n35956 ;
  assign n35960 = n35953 & ~n35959 ;
  assign n35961 = n35958 | n35960 ;
  assign n35962 = x118 & n12574 ;
  assign n35963 = x117 & n12569 ;
  assign n35964 = x116 & ~n12568 ;
  assign n35965 = n13076 & n35964 ;
  assign n35966 = n35963 | n35965 ;
  assign n35967 = n35962 | n35966 ;
  assign n35968 = n12577 | n35962 ;
  assign n35969 = n35966 | n35968 ;
  assign n35970 = ( ~n14002 & n35967 ) | ( ~n14002 & n35969 ) | ( n35967 & n35969 ) ;
  assign n35971 = n35967 & n35969 ;
  assign n35972 = ( n13981 & n35970 ) | ( n13981 & n35971 ) | ( n35970 & n35971 ) ;
  assign n35973 = x53 & n35972 ;
  assign n35974 = x53 & ~n35972 ;
  assign n35975 = ( n35972 & ~n35973 ) | ( n35972 & n35974 ) | ( ~n35973 & n35974 ) ;
  assign n35976 = n35961 & ~n35975 ;
  assign n35977 = ~n35961 & n35975 ;
  assign n35978 = n35976 | n35977 ;
  assign n35979 = n35869 & ~n35978 ;
  assign n35980 = ~n35869 & n35978 ;
  assign n35981 = n35979 | n35980 ;
  assign n35982 = x121 & n11205 ;
  assign n35983 = x120 & n11200 ;
  assign n35984 = x119 & ~n11199 ;
  assign n35985 = n11679 & n35984 ;
  assign n35986 = n35983 | n35985 ;
  assign n35987 = n35982 | n35986 ;
  assign n35988 = n11208 | n35982 ;
  assign n35989 = n35986 | n35988 ;
  assign n35990 = ( n15501 & n35987 ) | ( n15501 & n35989 ) | ( n35987 & n35989 ) ;
  assign n35991 = x50 & n35989 ;
  assign n35992 = x50 & n35982 ;
  assign n35993 = ( x50 & n35986 ) | ( x50 & n35992 ) | ( n35986 & n35992 ) ;
  assign n35994 = ( n15501 & n35991 ) | ( n15501 & n35993 ) | ( n35991 & n35993 ) ;
  assign n35995 = x50 & ~n35993 ;
  assign n35996 = x50 & ~n35989 ;
  assign n35997 = ( ~n15501 & n35995 ) | ( ~n15501 & n35996 ) | ( n35995 & n35996 ) ;
  assign n35998 = ( n35990 & ~n35994 ) | ( n35990 & n35997 ) | ( ~n35994 & n35997 ) ;
  assign n35999 = n35981 & ~n35998 ;
  assign n36000 = ~n35981 & n35998 ;
  assign n36001 = n35999 | n36000 ;
  assign n36002 = n35868 & ~n36001 ;
  assign n36003 = ~n35868 & n36001 ;
  assign n36004 = n36002 | n36003 ;
  assign n36005 = x124 & n9933 ;
  assign n36006 = x123 & n9928 ;
  assign n36007 = x122 & ~n9927 ;
  assign n36008 = n10379 & n36007 ;
  assign n36009 = n36006 | n36008 ;
  assign n36010 = n36005 | n36009 ;
  assign n36011 = n9936 | n36005 ;
  assign n36012 = n36009 | n36011 ;
  assign n36013 = ( n17084 & n36010 ) | ( n17084 & n36012 ) | ( n36010 & n36012 ) ;
  assign n36014 = x47 & n36012 ;
  assign n36015 = x47 & n36005 ;
  assign n36016 = ( x47 & n36009 ) | ( x47 & n36015 ) | ( n36009 & n36015 ) ;
  assign n36017 = ( n17084 & n36014 ) | ( n17084 & n36016 ) | ( n36014 & n36016 ) ;
  assign n36018 = x47 & ~n36016 ;
  assign n36019 = x47 & ~n36012 ;
  assign n36020 = ( ~n17084 & n36018 ) | ( ~n17084 & n36019 ) | ( n36018 & n36019 ) ;
  assign n36021 = ( n36013 & ~n36017 ) | ( n36013 & n36020 ) | ( ~n36017 & n36020 ) ;
  assign n36022 = ~n36004 & n36021 ;
  assign n36023 = n36004 | n36022 ;
  assign n36024 = n36004 & n36021 ;
  assign n36025 = n36023 & ~n36024 ;
  assign n36026 = n35769 | n35789 ;
  assign n36027 = ( n35769 & ~n35772 ) | ( n35769 & n36026 ) | ( ~n35772 & n36026 ) ;
  assign n36028 = n36025 & ~n36027 ;
  assign n36029 = ~n36025 & n36027 ;
  assign n36030 = n36028 | n36029 ;
  assign n36031 = x127 & n8724 ;
  assign n36032 = x126 & n8719 ;
  assign n36033 = x125 & ~n8718 ;
  assign n36034 = n9149 & n36033 ;
  assign n36035 = n36032 | n36034 ;
  assign n36036 = n36031 | n36035 ;
  assign n36037 = n8727 | n36031 ;
  assign n36038 = n36035 | n36037 ;
  assign n36039 = ( n18763 & n36036 ) | ( n18763 & n36038 ) | ( n36036 & n36038 ) ;
  assign n36040 = x44 & n36038 ;
  assign n36041 = x44 & n36031 ;
  assign n36042 = ( x44 & n36035 ) | ( x44 & n36041 ) | ( n36035 & n36041 ) ;
  assign n36043 = ( n18763 & n36040 ) | ( n18763 & n36042 ) | ( n36040 & n36042 ) ;
  assign n36044 = x44 & ~n36042 ;
  assign n36045 = x44 & ~n36038 ;
  assign n36046 = ( ~n18763 & n36044 ) | ( ~n18763 & n36045 ) | ( n36044 & n36045 ) ;
  assign n36047 = ( n36039 & ~n36043 ) | ( n36039 & n36046 ) | ( ~n36043 & n36046 ) ;
  assign n36048 = ~n36030 & n36047 ;
  assign n36049 = n36030 | n36048 ;
  assign n36050 = ( n35795 & ~n35796 ) | ( n35795 & n35815 ) | ( ~n35796 & n35815 ) ;
  assign n36051 = n36030 & n36047 ;
  assign n36052 = n36050 & n36051 ;
  assign n36053 = ( ~n36049 & n36050 ) | ( ~n36049 & n36052 ) | ( n36050 & n36052 ) ;
  assign n36054 = n36050 | n36051 ;
  assign n36055 = n36049 & ~n36054 ;
  assign n36056 = n36053 | n36055 ;
  assign n36057 = n35835 & n35837 ;
  assign n36058 = n35837 & ~n36057 ;
  assign n36059 = ~n35817 & n35835 ;
  assign n36060 = ~n35837 & n36059 ;
  assign n36061 = ( ~n35817 & n36058 ) | ( ~n35817 & n36060 ) | ( n36058 & n36060 ) ;
  assign n36062 = ~n36056 & n36057 ;
  assign n36063 = ( ~n36056 & n36061 ) | ( ~n36056 & n36062 ) | ( n36061 & n36062 ) ;
  assign n36064 = n36056 & ~n36057 ;
  assign n36065 = ~n36061 & n36064 ;
  assign n36066 = n36063 | n36065 ;
  assign n36067 = ~n35846 & n35858 ;
  assign n36068 = n35846 | n35859 ;
  assign n36069 = ~n35846 & n35848 ;
  assign n36070 = ( n35630 & n36068 ) | ( n35630 & ~n36069 ) | ( n36068 & ~n36069 ) ;
  assign n36071 = ( n35392 & ~n36067 ) | ( n35392 & n36070 ) | ( ~n36067 & n36070 ) ;
  assign n36072 = ~n35846 & n35862 ;
  assign n36073 = ( n35625 & ~n36068 ) | ( n35625 & n36072 ) | ( ~n36068 & n36072 ) ;
  assign n36074 = ( n34357 & ~n36071 ) | ( n34357 & n36073 ) | ( ~n36071 & n36073 ) ;
  assign n36075 = ( n35415 & ~n36070 ) | ( n35415 & n36072 ) | ( ~n36070 & n36072 ) ;
  assign n36076 = ( ~n30754 & n36074 ) | ( ~n30754 & n36075 ) | ( n36074 & n36075 ) ;
  assign n36077 = n36066 & n36076 ;
  assign n36078 = ~n36066 & n36070 ;
  assign n36079 = n36066 | n36067 ;
  assign n36080 = ( n35392 & n36078 ) | ( n35392 & ~n36079 ) | ( n36078 & ~n36079 ) ;
  assign n36081 = ~n36066 & n36068 ;
  assign n36082 = n35846 & ~n36066 ;
  assign n36083 = ( n35862 & n36066 ) | ( n35862 & ~n36082 ) | ( n36066 & ~n36082 ) ;
  assign n36084 = ( n35625 & ~n36081 ) | ( n35625 & n36083 ) | ( ~n36081 & n36083 ) ;
  assign n36085 = ( n34357 & ~n36080 ) | ( n34357 & n36084 ) | ( ~n36080 & n36084 ) ;
  assign n36086 = ( n35415 & ~n36078 ) | ( n35415 & n36083 ) | ( ~n36078 & n36083 ) ;
  assign n36087 = ( ~n30754 & n36085 ) | ( ~n30754 & n36086 ) | ( n36085 & n36086 ) ;
  assign n36088 = ~n36077 & n36087 ;
  assign n36089 = x127 & n8719 ;
  assign n36090 = x126 & ~n8718 ;
  assign n36091 = n9149 & n36090 ;
  assign n36092 = n36089 | n36091 ;
  assign n36093 = n8727 | n36092 ;
  assign n36094 = ( n19328 & n36092 ) | ( n19328 & n36093 ) | ( n36092 & n36093 ) ;
  assign n36095 = x44 & n36092 ;
  assign n36096 = ( x44 & n11726 ) | ( x44 & n36092 ) | ( n11726 & n36092 ) ;
  assign n36097 = ( n19328 & n36095 ) | ( n19328 & n36096 ) | ( n36095 & n36096 ) ;
  assign n36098 = x44 & ~n11726 ;
  assign n36099 = ~n36092 & n36098 ;
  assign n36100 = x44 & ~n36092 ;
  assign n36101 = ( ~n19328 & n36099 ) | ( ~n19328 & n36100 ) | ( n36099 & n36100 ) ;
  assign n36102 = ( n36094 & ~n36097 ) | ( n36094 & n36101 ) | ( ~n36097 & n36101 ) ;
  assign n36103 = n36022 | n36027 ;
  assign n36104 = ( n36022 & ~n36025 ) | ( n36022 & n36103 ) | ( ~n36025 & n36103 ) ;
  assign n36105 = n36102 & n36104 ;
  assign n36106 = n36102 | n36104 ;
  assign n36107 = ~n36105 & n36106 ;
  assign n36108 = n36000 | n36002 ;
  assign n36109 = n35977 | n35979 ;
  assign n36110 = ( ~x41 & n35460 ) | ( ~x41 & n35876 ) | ( n35460 & n35876 ) ;
  assign n36111 = x107 & n18290 ;
  assign n36112 = x63 & x106 ;
  assign n36113 = ~n18290 & n36112 ;
  assign n36114 = n36111 | n36113 ;
  assign n36115 = n36110 & ~n36114 ;
  assign n36116 = n36110 & ~n36115 ;
  assign n36117 = n36110 | n36114 ;
  assign n36118 = ~n36116 & n36117 ;
  assign n36120 = x109 & n17141 ;
  assign n36121 = x108 & ~n17140 ;
  assign n36122 = n17724 & n36121 ;
  assign n36123 = n36120 | n36122 ;
  assign n36119 = x110 & n17146 ;
  assign n36125 = n17149 | n36119 ;
  assign n36126 = n36123 | n36125 ;
  assign n36124 = n36119 | n36123 ;
  assign n36127 = n36124 & n36126 ;
  assign n36128 = ( n10330 & n36126 ) | ( n10330 & n36127 ) | ( n36126 & n36127 ) ;
  assign n36129 = x62 & n36127 ;
  assign n36130 = x62 & n36126 ;
  assign n36131 = ( n10330 & n36129 ) | ( n10330 & n36130 ) | ( n36129 & n36130 ) ;
  assign n36132 = x62 & ~n36127 ;
  assign n36133 = x62 & ~n36126 ;
  assign n36134 = ( ~n10330 & n36132 ) | ( ~n10330 & n36133 ) | ( n36132 & n36133 ) ;
  assign n36135 = ( n36128 & ~n36131 ) | ( n36128 & n36134 ) | ( ~n36131 & n36134 ) ;
  assign n36136 = ~n36118 & n36135 ;
  assign n36137 = n36118 & ~n36135 ;
  assign n36138 = n36136 | n36137 ;
  assign n36139 = n35898 | n35905 ;
  assign n36140 = ( n35898 & ~n35900 ) | ( n35898 & n36139 ) | ( ~n35900 & n36139 ) ;
  assign n36141 = ~n36138 & n36140 ;
  assign n36142 = n36138 & ~n36140 ;
  assign n36143 = n36141 | n36142 ;
  assign n36144 = x113 & n15552 ;
  assign n36145 = x112 & n15547 ;
  assign n36146 = x111 & ~n15546 ;
  assign n36147 = n16123 & n36146 ;
  assign n36148 = n36145 | n36147 ;
  assign n36149 = n36144 | n36148 ;
  assign n36150 = n15555 | n36144 ;
  assign n36151 = n36148 | n36150 ;
  assign n36152 = ( ~n11642 & n36149 ) | ( ~n11642 & n36151 ) | ( n36149 & n36151 ) ;
  assign n36153 = n36149 & n36151 ;
  assign n36154 = ( n11626 & n36152 ) | ( n11626 & n36153 ) | ( n36152 & n36153 ) ;
  assign n36155 = x59 & n36154 ;
  assign n36156 = x59 & ~n36154 ;
  assign n36157 = ( n36154 & ~n36155 ) | ( n36154 & n36156 ) | ( ~n36155 & n36156 ) ;
  assign n36158 = n36143 | n36157 ;
  assign n36159 = n36143 & ~n36157 ;
  assign n36160 = ( ~n36143 & n36158 ) | ( ~n36143 & n36159 ) | ( n36158 & n36159 ) ;
  assign n36161 = n35926 | n35932 ;
  assign n36162 = ( ~n35908 & n35930 ) | ( ~n35908 & n35934 ) | ( n35930 & n35934 ) ;
  assign n36163 = ( ~n35927 & n36161 ) | ( ~n35927 & n36162 ) | ( n36161 & n36162 ) ;
  assign n36164 = n36160 & ~n36163 ;
  assign n36165 = ~n36160 & n36163 ;
  assign n36166 = n36164 | n36165 ;
  assign n36167 = x116 & n14045 ;
  assign n36168 = x115 & n14040 ;
  assign n36169 = x114 & ~n14039 ;
  assign n36170 = n14552 & n36169 ;
  assign n36171 = n36168 | n36170 ;
  assign n36172 = n36167 | n36171 ;
  assign n36173 = n14048 | n36167 ;
  assign n36174 = n36171 | n36173 ;
  assign n36175 = ( ~n13040 & n36172 ) | ( ~n13040 & n36174 ) | ( n36172 & n36174 ) ;
  assign n36176 = n36172 & n36174 ;
  assign n36177 = ( n13022 & n36175 ) | ( n13022 & n36176 ) | ( n36175 & n36176 ) ;
  assign n36178 = x56 & n36177 ;
  assign n36179 = x56 & ~n36177 ;
  assign n36180 = ( n36177 & ~n36178 ) | ( n36177 & n36179 ) | ( ~n36178 & n36179 ) ;
  assign n36181 = n36166 & n36180 ;
  assign n36182 = n36165 | n36180 ;
  assign n36183 = n36164 | n36182 ;
  assign n36184 = ~n36181 & n36183 ;
  assign n36185 = n35952 | n35958 ;
  assign n36186 = n36184 & ~n36185 ;
  assign n36187 = x119 & n12574 ;
  assign n36188 = x118 & n12569 ;
  assign n36189 = x117 & ~n12568 ;
  assign n36190 = n13076 & n36189 ;
  assign n36191 = n36188 | n36190 ;
  assign n36192 = n36187 | n36191 ;
  assign n36193 = n12577 | n36187 ;
  assign n36194 = n36191 | n36193 ;
  assign n36195 = ( n14496 & n36192 ) | ( n14496 & n36194 ) | ( n36192 & n36194 ) ;
  assign n36196 = x53 & n36194 ;
  assign n36197 = x53 & n36187 ;
  assign n36198 = ( x53 & n36191 ) | ( x53 & n36197 ) | ( n36191 & n36197 ) ;
  assign n36199 = ( n14496 & n36196 ) | ( n14496 & n36198 ) | ( n36196 & n36198 ) ;
  assign n36200 = x53 & ~n36198 ;
  assign n36201 = x53 & ~n36194 ;
  assign n36202 = ( ~n14496 & n36200 ) | ( ~n14496 & n36201 ) | ( n36200 & n36201 ) ;
  assign n36203 = ( n36195 & ~n36199 ) | ( n36195 & n36202 ) | ( ~n36199 & n36202 ) ;
  assign n36204 = n36184 & ~n36203 ;
  assign n36205 = ( n36185 & n36203 ) | ( n36185 & ~n36204 ) | ( n36203 & ~n36204 ) ;
  assign n36206 = n36186 | n36205 ;
  assign n36207 = ~n36184 & n36185 ;
  assign n36208 = n36186 | n36207 ;
  assign n36209 = n36203 & n36208 ;
  assign n36210 = ~n36109 & n36209 ;
  assign n36211 = ( n36109 & n36206 ) | ( n36109 & ~n36210 ) | ( n36206 & ~n36210 ) ;
  assign n36212 = x122 & n11205 ;
  assign n36213 = x121 & n11200 ;
  assign n36214 = x120 & ~n11199 ;
  assign n36215 = n11679 & n36214 ;
  assign n36216 = n36213 | n36215 ;
  assign n36217 = n36212 | n36216 ;
  assign n36218 = n11208 | n36212 ;
  assign n36219 = n36216 | n36218 ;
  assign n36220 = ( n16043 & n36217 ) | ( n16043 & n36219 ) | ( n36217 & n36219 ) ;
  assign n36221 = x50 & n36219 ;
  assign n36222 = x50 & n36212 ;
  assign n36223 = ( x50 & n36216 ) | ( x50 & n36222 ) | ( n36216 & n36222 ) ;
  assign n36224 = ( n16043 & n36221 ) | ( n16043 & n36223 ) | ( n36221 & n36223 ) ;
  assign n36225 = x50 & ~n36223 ;
  assign n36226 = x50 & ~n36219 ;
  assign n36227 = ( ~n16043 & n36225 ) | ( ~n16043 & n36226 ) | ( n36225 & n36226 ) ;
  assign n36228 = ( n36220 & ~n36224 ) | ( n36220 & n36227 ) | ( ~n36224 & n36227 ) ;
  assign n36229 = n36206 & ~n36209 ;
  assign n36230 = n36109 & n36229 ;
  assign n36231 = n36228 | n36230 ;
  assign n36232 = n36211 & ~n36231 ;
  assign n36233 = n36228 & n36230 ;
  assign n36234 = ( ~n36211 & n36228 ) | ( ~n36211 & n36233 ) | ( n36228 & n36233 ) ;
  assign n36235 = n36232 | n36234 ;
  assign n36236 = n36108 & ~n36235 ;
  assign n36237 = n36108 & ~n36236 ;
  assign n36238 = n36235 | n36236 ;
  assign n36239 = ~n36237 & n36238 ;
  assign n36240 = x125 & n9933 ;
  assign n36241 = x124 & n9928 ;
  assign n36242 = x123 & ~n9927 ;
  assign n36243 = n10379 & n36242 ;
  assign n36244 = n36241 | n36243 ;
  assign n36245 = n36240 | n36244 ;
  assign n36246 = n9936 | n36240 ;
  assign n36247 = n36244 | n36246 ;
  assign n36248 = ( n17670 & n36245 ) | ( n17670 & n36247 ) | ( n36245 & n36247 ) ;
  assign n36249 = x47 & n36247 ;
  assign n36250 = x47 & n36240 ;
  assign n36251 = ( x47 & n36244 ) | ( x47 & n36250 ) | ( n36244 & n36250 ) ;
  assign n36252 = ( n17670 & n36249 ) | ( n17670 & n36251 ) | ( n36249 & n36251 ) ;
  assign n36253 = x47 & ~n36251 ;
  assign n36254 = x47 & ~n36247 ;
  assign n36255 = ( ~n17670 & n36253 ) | ( ~n17670 & n36254 ) | ( n36253 & n36254 ) ;
  assign n36256 = ( n36248 & ~n36252 ) | ( n36248 & n36255 ) | ( ~n36252 & n36255 ) ;
  assign n36257 = n36239 & n36256 ;
  assign n36258 = n36239 | n36256 ;
  assign n36259 = ~n36257 & n36258 ;
  assign n36260 = n36107 & ~n36259 ;
  assign n36261 = n36107 | n36259 ;
  assign n36262 = ( ~n36107 & n36260 ) | ( ~n36107 & n36261 ) | ( n36260 & n36261 ) ;
  assign n36263 = n36048 | n36053 ;
  assign n36264 = n36262 & ~n36263 ;
  assign n36265 = ~n36262 & n36263 ;
  assign n36266 = n36264 | n36265 ;
  assign n36267 = ~n36063 & n36079 ;
  assign n36268 = ~n36063 & n36066 ;
  assign n36269 = ( n36063 & n36070 ) | ( n36063 & ~n36268 ) | ( n36070 & ~n36268 ) ;
  assign n36270 = ( n35392 & ~n36267 ) | ( n35392 & n36269 ) | ( ~n36267 & n36269 ) ;
  assign n36271 = n36063 | n36081 ;
  assign n36272 = n36063 | n36082 ;
  assign n36273 = ( n35862 & n36268 ) | ( n35862 & ~n36272 ) | ( n36268 & ~n36272 ) ;
  assign n36274 = ( n35625 & ~n36271 ) | ( n35625 & n36273 ) | ( ~n36271 & n36273 ) ;
  assign n36275 = ( n34357 & ~n36270 ) | ( n34357 & n36274 ) | ( ~n36270 & n36274 ) ;
  assign n36276 = ( n35415 & ~n36269 ) | ( n35415 & n36273 ) | ( ~n36269 & n36273 ) ;
  assign n36277 = ( ~n30754 & n36275 ) | ( ~n30754 & n36276 ) | ( n36275 & n36276 ) ;
  assign n36278 = n36266 & n36277 ;
  assign n36279 = ~n36266 & n36270 ;
  assign n36280 = ~n36266 & n36271 ;
  assign n36281 = n36266 | n36268 ;
  assign n36282 = ~n36266 & n36272 ;
  assign n36283 = ( n35862 & n36281 ) | ( n35862 & ~n36282 ) | ( n36281 & ~n36282 ) ;
  assign n36284 = ( n35625 & ~n36280 ) | ( n35625 & n36283 ) | ( ~n36280 & n36283 ) ;
  assign n36285 = ( n34357 & ~n36279 ) | ( n34357 & n36284 ) | ( ~n36279 & n36284 ) ;
  assign n36286 = n36063 & ~n36266 ;
  assign n36287 = ( n36070 & ~n36281 ) | ( n36070 & n36286 ) | ( ~n36281 & n36286 ) ;
  assign n36288 = ( n35415 & n36283 ) | ( n35415 & ~n36287 ) | ( n36283 & ~n36287 ) ;
  assign n36289 = ( ~n30754 & n36285 ) | ( ~n30754 & n36288 ) | ( n36285 & n36288 ) ;
  assign n36290 = ~n36278 & n36289 ;
  assign n36291 = x127 & ~n8718 ;
  assign n36292 = n9149 & n36291 ;
  assign n36293 = n8727 & n19877 ;
  assign n36294 = n36292 | n36293 ;
  assign n36295 = n8727 & n19880 ;
  assign n36296 = n36292 | n36295 ;
  assign n36297 = ( n18202 & n36294 ) | ( n18202 & n36296 ) | ( n36294 & n36296 ) ;
  assign n36298 = n36294 & n36296 ;
  assign n36299 = ( n18212 & n36297 ) | ( n18212 & n36298 ) | ( n36297 & n36298 ) ;
  assign n36300 = ( n18214 & n36297 ) | ( n18214 & n36298 ) | ( n36297 & n36298 ) ;
  assign n36301 = ( n14002 & n36299 ) | ( n14002 & n36300 ) | ( n36299 & n36300 ) ;
  assign n36302 = x44 & n36299 ;
  assign n36303 = x44 & n36300 ;
  assign n36304 = ( n14002 & n36302 ) | ( n14002 & n36303 ) | ( n36302 & n36303 ) ;
  assign n36305 = x44 & ~n36303 ;
  assign n36306 = x44 & ~n36302 ;
  assign n36307 = ( ~n14002 & n36305 ) | ( ~n14002 & n36306 ) | ( n36305 & n36306 ) ;
  assign n36308 = ( n36301 & ~n36304 ) | ( n36301 & n36307 ) | ( ~n36304 & n36307 ) ;
  assign n36309 = n36236 & n36308 ;
  assign n36310 = n36256 & n36308 ;
  assign n36311 = ( n36236 & n36308 ) | ( n36236 & n36310 ) | ( n36308 & n36310 ) ;
  assign n36312 = ( ~n36239 & n36309 ) | ( ~n36239 & n36311 ) | ( n36309 & n36311 ) ;
  assign n36313 = n36236 | n36308 ;
  assign n36314 = n36256 | n36308 ;
  assign n36315 = n36236 | n36314 ;
  assign n36316 = ( ~n36239 & n36313 ) | ( ~n36239 & n36315 ) | ( n36313 & n36315 ) ;
  assign n36317 = ~n36312 & n36316 ;
  assign n36392 = ( n36165 & ~n36166 ) | ( n36165 & n36182 ) | ( ~n36166 & n36182 ) ;
  assign n36386 = n36138 & ~n36157 ;
  assign n36387 = ( n36140 & n36157 ) | ( n36140 & ~n36386 ) | ( n36157 & ~n36386 ) ;
  assign n36388 = ( n36141 & ~n36143 ) | ( n36141 & n36387 ) | ( ~n36143 & n36387 ) ;
  assign n36318 = x108 & n18290 ;
  assign n36319 = x63 & x107 ;
  assign n36320 = ~n18290 & n36319 ;
  assign n36321 = n36318 | n36320 ;
  assign n36322 = ~n36114 & n36321 ;
  assign n36323 = n36114 & ~n36321 ;
  assign n36324 = n36322 | n36323 ;
  assign n36326 = x110 & n17141 ;
  assign n36327 = x109 & ~n17140 ;
  assign n36328 = n17724 & n36327 ;
  assign n36329 = n36326 | n36328 ;
  assign n36325 = x111 & n17146 ;
  assign n36331 = n17149 | n36325 ;
  assign n36332 = n36329 | n36331 ;
  assign n36330 = n36325 | n36329 ;
  assign n36333 = n36330 & n36332 ;
  assign n36334 = ( n10749 & n36332 ) | ( n10749 & n36333 ) | ( n36332 & n36333 ) ;
  assign n36335 = x62 & n36333 ;
  assign n36336 = x62 & n36332 ;
  assign n36337 = ( n10749 & n36335 ) | ( n10749 & n36336 ) | ( n36335 & n36336 ) ;
  assign n36338 = x62 & ~n36333 ;
  assign n36339 = x62 & ~n36332 ;
  assign n36340 = ( ~n10749 & n36338 ) | ( ~n10749 & n36339 ) | ( n36338 & n36339 ) ;
  assign n36341 = ( n36334 & ~n36337 ) | ( n36334 & n36340 ) | ( ~n36337 & n36340 ) ;
  assign n36342 = ~n36324 & n36341 ;
  assign n36343 = n36324 & ~n36341 ;
  assign n36344 = n36342 | n36343 ;
  assign n36345 = ~n36115 & n36117 ;
  assign n36346 = ~n36116 & n36345 ;
  assign n36347 = ( n36115 & n36135 ) | ( n36115 & ~n36346 ) | ( n36135 & ~n36346 ) ;
  assign n36348 = n36344 & n36347 ;
  assign n36349 = ~n36344 & n36347 ;
  assign n36350 = x114 & n15552 ;
  assign n36351 = x113 & n15547 ;
  assign n36352 = x112 & ~n15546 ;
  assign n36353 = n16123 & n36352 ;
  assign n36354 = n36351 | n36353 ;
  assign n36355 = n36350 | n36354 ;
  assign n36356 = n15555 | n36350 ;
  assign n36357 = n36354 | n36356 ;
  assign n36358 = ( ~n12095 & n36355 ) | ( ~n12095 & n36357 ) | ( n36355 & n36357 ) ;
  assign n36359 = n36355 & n36357 ;
  assign n36360 = ( n12079 & n36358 ) | ( n12079 & n36359 ) | ( n36358 & n36359 ) ;
  assign n36361 = x59 & n36360 ;
  assign n36362 = x59 & ~n36360 ;
  assign n36363 = ( n36360 & ~n36361 ) | ( n36360 & n36362 ) | ( ~n36361 & n36362 ) ;
  assign n36364 = n36344 & ~n36363 ;
  assign n36365 = ( n36349 & ~n36363 ) | ( n36349 & n36364 ) | ( ~n36363 & n36364 ) ;
  assign n36366 = ~n36348 & n36365 ;
  assign n36367 = n36344 | n36349 ;
  assign n36368 = n36347 & n36363 ;
  assign n36369 = n36344 & n36368 ;
  assign n36370 = ( n36363 & ~n36367 ) | ( n36363 & n36369 ) | ( ~n36367 & n36369 ) ;
  assign n36371 = n36366 | n36370 ;
  assign n36372 = x117 & n14045 ;
  assign n36373 = x116 & n14040 ;
  assign n36374 = x115 & ~n14039 ;
  assign n36375 = n14552 & n36374 ;
  assign n36376 = n36373 | n36375 ;
  assign n36377 = n36372 | n36376 ;
  assign n36378 = n14048 | n36372 ;
  assign n36379 = n36376 | n36378 ;
  assign n36380 = ( ~n13522 & n36377 ) | ( ~n13522 & n36379 ) | ( n36377 & n36379 ) ;
  assign n36381 = n36377 & n36379 ;
  assign n36382 = ( n13503 & n36380 ) | ( n13503 & n36381 ) | ( n36380 & n36381 ) ;
  assign n36383 = x56 & n36382 ;
  assign n36384 = x56 & ~n36382 ;
  assign n36385 = ( n36382 & ~n36383 ) | ( n36382 & n36384 ) | ( ~n36383 & n36384 ) ;
  assign n36389 = ( ~n36371 & n36385 ) | ( ~n36371 & n36388 ) | ( n36385 & n36388 ) ;
  assign n36390 = ( n36371 & ~n36385 ) | ( n36371 & n36389 ) | ( ~n36385 & n36389 ) ;
  assign n36391 = ( ~n36388 & n36389 ) | ( ~n36388 & n36390 ) | ( n36389 & n36390 ) ;
  assign n36393 = ~n36391 & n36392 ;
  assign n36394 = n36392 & ~n36393 ;
  assign n36395 = x120 & n12574 ;
  assign n36396 = x119 & n12569 ;
  assign n36397 = x118 & ~n12568 ;
  assign n36398 = n13076 & n36397 ;
  assign n36399 = n36396 | n36398 ;
  assign n36400 = n36395 | n36399 ;
  assign n36401 = n12577 | n36395 ;
  assign n36402 = n36399 | n36401 ;
  assign n36403 = ( n14991 & n36400 ) | ( n14991 & n36402 ) | ( n36400 & n36402 ) ;
  assign n36404 = x53 & n36402 ;
  assign n36405 = x53 & n36395 ;
  assign n36406 = ( x53 & n36399 ) | ( x53 & n36405 ) | ( n36399 & n36405 ) ;
  assign n36407 = ( n14991 & n36404 ) | ( n14991 & n36406 ) | ( n36404 & n36406 ) ;
  assign n36408 = x53 & ~n36406 ;
  assign n36409 = x53 & ~n36402 ;
  assign n36410 = ( ~n14991 & n36408 ) | ( ~n14991 & n36409 ) | ( n36408 & n36409 ) ;
  assign n36411 = ( n36403 & ~n36407 ) | ( n36403 & n36410 ) | ( ~n36407 & n36410 ) ;
  assign n36412 = n36389 & ~n36411 ;
  assign n36413 = n36388 | n36411 ;
  assign n36414 = ( n36390 & n36412 ) | ( n36390 & ~n36413 ) | ( n36412 & ~n36413 ) ;
  assign n36415 = ( n36392 & ~n36411 ) | ( n36392 & n36414 ) | ( ~n36411 & n36414 ) ;
  assign n36416 = ~n36394 & n36415 ;
  assign n36417 = ~n36389 & n36411 ;
  assign n36418 = n36388 & n36411 ;
  assign n36419 = ( ~n36390 & n36417 ) | ( ~n36390 & n36418 ) | ( n36417 & n36418 ) ;
  assign n36420 = ~n36392 & n36419 ;
  assign n36421 = ( n36394 & n36411 ) | ( n36394 & n36420 ) | ( n36411 & n36420 ) ;
  assign n36422 = n36416 | n36421 ;
  assign n36423 = ( n36205 & n36207 ) | ( n36205 & ~n36208 ) | ( n36207 & ~n36208 ) ;
  assign n36424 = ~n36422 & n36423 ;
  assign n36425 = n36422 & ~n36423 ;
  assign n36426 = n36424 | n36425 ;
  assign n36427 = x123 & n11205 ;
  assign n36428 = x122 & n11200 ;
  assign n36429 = x121 & ~n11199 ;
  assign n36430 = n11679 & n36429 ;
  assign n36431 = n36428 | n36430 ;
  assign n36432 = n36427 | n36431 ;
  assign n36433 = n11208 | n36427 ;
  assign n36434 = n36431 | n36433 ;
  assign n36435 = ( n16086 & n36432 ) | ( n16086 & n36434 ) | ( n36432 & n36434 ) ;
  assign n36436 = x50 & n36434 ;
  assign n36437 = x50 & n36427 ;
  assign n36438 = ( x50 & n36431 ) | ( x50 & n36437 ) | ( n36431 & n36437 ) ;
  assign n36439 = ( n16086 & n36436 ) | ( n16086 & n36438 ) | ( n36436 & n36438 ) ;
  assign n36440 = x50 & ~n36438 ;
  assign n36441 = x50 & ~n36434 ;
  assign n36442 = ( ~n16086 & n36440 ) | ( ~n16086 & n36441 ) | ( n36440 & n36441 ) ;
  assign n36443 = ( n36435 & ~n36439 ) | ( n36435 & n36442 ) | ( ~n36439 & n36442 ) ;
  assign n36444 = n36426 | n36443 ;
  assign n36445 = n36426 & ~n36443 ;
  assign n36446 = ( ~n36426 & n36444 ) | ( ~n36426 & n36445 ) | ( n36444 & n36445 ) ;
  assign n36447 = ( n36109 & n36228 ) | ( n36109 & ~n36229 ) | ( n36228 & ~n36229 ) ;
  assign n36448 = ~n36446 & n36447 ;
  assign n36449 = n36446 | n36448 ;
  assign n36450 = x126 & n9933 ;
  assign n36451 = x125 & n9928 ;
  assign n36452 = x124 & ~n9927 ;
  assign n36453 = n10379 & n36452 ;
  assign n36454 = n36451 | n36453 ;
  assign n36455 = n36450 | n36454 ;
  assign n36456 = n9936 | n36450 ;
  assign n36457 = n36454 | n36456 ;
  assign n36458 = ( n18220 & n36455 ) | ( n18220 & n36457 ) | ( n36455 & n36457 ) ;
  assign n36459 = x47 & n36457 ;
  assign n36460 = x47 & n36450 ;
  assign n36461 = ( x47 & n36454 ) | ( x47 & n36460 ) | ( n36454 & n36460 ) ;
  assign n36462 = ( n18220 & n36459 ) | ( n18220 & n36461 ) | ( n36459 & n36461 ) ;
  assign n36463 = x47 & ~n36461 ;
  assign n36464 = x47 & ~n36457 ;
  assign n36465 = ( ~n18220 & n36463 ) | ( ~n18220 & n36464 ) | ( n36463 & n36464 ) ;
  assign n36466 = ( n36458 & ~n36462 ) | ( n36458 & n36465 ) | ( ~n36462 & n36465 ) ;
  assign n36467 = n36447 & n36466 ;
  assign n36468 = n36446 & n36467 ;
  assign n36469 = ( ~n36449 & n36466 ) | ( ~n36449 & n36468 ) | ( n36466 & n36468 ) ;
  assign n36470 = n36447 | n36466 ;
  assign n36471 = ( n36446 & n36466 ) | ( n36446 & n36470 ) | ( n36466 & n36470 ) ;
  assign n36472 = n36449 & ~n36471 ;
  assign n36473 = n36469 | n36472 ;
  assign n36474 = n36317 & n36473 ;
  assign n36475 = n36317 | n36473 ;
  assign n36476 = ~n36474 & n36475 ;
  assign n36477 = ~n36105 & n36259 ;
  assign n36478 = ( n36105 & n36107 ) | ( n36105 & ~n36477 ) | ( n36107 & ~n36477 ) ;
  assign n36479 = ~n36476 & n36478 ;
  assign n36480 = n36476 & ~n36478 ;
  assign n36481 = n36479 | n36480 ;
  assign n36482 = ~n36265 & n36266 ;
  assign n36483 = ( n36265 & n36270 ) | ( n36265 & ~n36482 ) | ( n36270 & ~n36482 ) ;
  assign n36484 = ~n36265 & n36283 ;
  assign n36485 = n36265 | n36280 ;
  assign n36486 = ( n35625 & n36484 ) | ( n35625 & ~n36485 ) | ( n36484 & ~n36485 ) ;
  assign n36487 = ( n34357 & ~n36483 ) | ( n34357 & n36486 ) | ( ~n36483 & n36486 ) ;
  assign n36488 = ~n36265 & n36281 ;
  assign n36489 = n36265 | n36286 ;
  assign n36490 = ( n36070 & ~n36488 ) | ( n36070 & n36489 ) | ( ~n36488 & n36489 ) ;
  assign n36491 = ( n35415 & n36484 ) | ( n35415 & ~n36490 ) | ( n36484 & ~n36490 ) ;
  assign n36492 = ( ~n30754 & n36487 ) | ( ~n30754 & n36491 ) | ( n36487 & n36491 ) ;
  assign n36493 = n36481 & n36492 ;
  assign n36494 = n36481 | n36482 ;
  assign n36495 = n36265 & ~n36481 ;
  assign n36496 = ( n36270 & ~n36494 ) | ( n36270 & n36495 ) | ( ~n36494 & n36495 ) ;
  assign n36497 = ~n36481 & n36485 ;
  assign n36498 = ( n36283 & n36481 ) | ( n36283 & ~n36495 ) | ( n36481 & ~n36495 ) ;
  assign n36499 = ( n35625 & ~n36497 ) | ( n35625 & n36498 ) | ( ~n36497 & n36498 ) ;
  assign n36500 = ( n34357 & ~n36496 ) | ( n34357 & n36499 ) | ( ~n36496 & n36499 ) ;
  assign n36501 = n36481 | n36488 ;
  assign n36502 = ~n36481 & n36489 ;
  assign n36503 = ( n36070 & ~n36501 ) | ( n36070 & n36502 ) | ( ~n36501 & n36502 ) ;
  assign n36504 = ( n35415 & n36498 ) | ( n35415 & ~n36503 ) | ( n36498 & ~n36503 ) ;
  assign n36505 = ( ~n30754 & n36500 ) | ( ~n30754 & n36504 ) | ( n36500 & n36504 ) ;
  assign n36506 = ~n36493 & n36505 ;
  assign n36507 = x115 & n15552 ;
  assign n36508 = x114 & n15547 ;
  assign n36509 = x113 & ~n15546 ;
  assign n36510 = n16123 & n36509 ;
  assign n36511 = n36508 | n36510 ;
  assign n36512 = n36507 | n36511 ;
  assign n36513 = n15555 | n36507 ;
  assign n36514 = n36511 | n36513 ;
  assign n36515 = ( ~n12550 & n36512 ) | ( ~n12550 & n36514 ) | ( n36512 & n36514 ) ;
  assign n36516 = n36512 & n36514 ;
  assign n36517 = ( n12532 & n36515 ) | ( n12532 & n36516 ) | ( n36515 & n36516 ) ;
  assign n36518 = x59 & n36517 ;
  assign n36519 = x59 & ~n36517 ;
  assign n36520 = ( n36517 & ~n36518 ) | ( n36517 & n36519 ) | ( ~n36518 & n36519 ) ;
  assign n36521 = x109 & n18290 ;
  assign n36522 = x63 & x108 ;
  assign n36523 = ~n18290 & n36522 ;
  assign n36524 = n36521 | n36523 ;
  assign n36525 = ~x44 & n36524 ;
  assign n36526 = x44 & ~n36524 ;
  assign n36527 = n36525 | n36526 ;
  assign n36528 = n36114 | n36527 ;
  assign n36529 = ~n36527 & n36528 ;
  assign n36530 = ~n36322 & n36324 ;
  assign n36531 = n36528 | n36530 ;
  assign n36532 = n36114 & n36322 ;
  assign n36533 = ( n36114 & ~n36324 ) | ( n36114 & n36532 ) | ( ~n36324 & n36532 ) ;
  assign n36534 = ( n36529 & n36531 ) | ( n36529 & ~n36533 ) | ( n36531 & ~n36533 ) ;
  assign n36535 = ~n36114 & n36322 ;
  assign n36536 = ~n36527 & n36535 ;
  assign n36537 = ( ~n36529 & n36532 ) | ( ~n36529 & n36536 ) | ( n36532 & n36536 ) ;
  assign n36538 = ( n36341 & ~n36534 ) | ( n36341 & n36537 ) | ( ~n36534 & n36537 ) ;
  assign n36539 = ( n36322 & n36342 ) | ( n36322 & ~n36538 ) | ( n36342 & ~n36538 ) ;
  assign n36540 = x112 & n17146 ;
  assign n36541 = x111 & n17141 ;
  assign n36542 = x110 & ~n17140 ;
  assign n36543 = n17724 & n36542 ;
  assign n36544 = n36541 | n36543 ;
  assign n36545 = n36540 | n36544 ;
  assign n36546 = n17149 | n36540 ;
  assign n36547 = n36544 | n36546 ;
  assign n36548 = ( n11172 & n36545 ) | ( n11172 & n36547 ) | ( n36545 & n36547 ) ;
  assign n36549 = x62 & n36547 ;
  assign n36550 = x62 & n36540 ;
  assign n36551 = ( x62 & n36544 ) | ( x62 & n36550 ) | ( n36544 & n36550 ) ;
  assign n36552 = ( n11172 & n36549 ) | ( n11172 & n36551 ) | ( n36549 & n36551 ) ;
  assign n36553 = x62 & ~n36551 ;
  assign n36554 = x62 & ~n36547 ;
  assign n36555 = ( ~n11172 & n36553 ) | ( ~n11172 & n36554 ) | ( n36553 & n36554 ) ;
  assign n36556 = ( n36548 & ~n36552 ) | ( n36548 & n36555 ) | ( ~n36552 & n36555 ) ;
  assign n36557 = ~n36528 & n36530 ;
  assign n36558 = n36114 & n36530 ;
  assign n36559 = ( ~n36529 & n36557 ) | ( ~n36529 & n36558 ) | ( n36557 & n36558 ) ;
  assign n36560 = n36322 | n36528 ;
  assign n36561 = n36114 & ~n36322 ;
  assign n36562 = ( n36529 & n36560 ) | ( n36529 & ~n36561 ) | ( n36560 & ~n36561 ) ;
  assign n36563 = ( n36341 & ~n36559 ) | ( n36341 & n36562 ) | ( ~n36559 & n36562 ) ;
  assign n36564 = n36556 & n36563 ;
  assign n36565 = ~n36539 & n36564 ;
  assign n36566 = n36520 & n36565 ;
  assign n36567 = n36556 | n36563 ;
  assign n36568 = ( ~n36539 & n36556 ) | ( ~n36539 & n36567 ) | ( n36556 & n36567 ) ;
  assign n36569 = ( n36520 & n36566 ) | ( n36520 & ~n36568 ) | ( n36566 & ~n36568 ) ;
  assign n36570 = n36520 | n36565 ;
  assign n36571 = n36568 & ~n36570 ;
  assign n36572 = n36569 | n36571 ;
  assign n36573 = n36349 | n36369 ;
  assign n36574 = n36347 | n36363 ;
  assign n36575 = ( ~n36344 & n36363 ) | ( ~n36344 & n36574 ) | ( n36363 & n36574 ) ;
  assign n36576 = ( ~n36367 & n36573 ) | ( ~n36367 & n36575 ) | ( n36573 & n36575 ) ;
  assign n36577 = ~n36572 & n36576 ;
  assign n36578 = n36572 & ~n36576 ;
  assign n36579 = n36577 | n36578 ;
  assign n36580 = x118 & n14045 ;
  assign n36581 = x117 & n14040 ;
  assign n36582 = x116 & ~n14039 ;
  assign n36583 = n14552 & n36582 ;
  assign n36584 = n36581 | n36583 ;
  assign n36585 = n36580 | n36584 ;
  assign n36586 = n14048 | n36580 ;
  assign n36587 = n36584 | n36586 ;
  assign n36588 = ( ~n14002 & n36585 ) | ( ~n14002 & n36587 ) | ( n36585 & n36587 ) ;
  assign n36589 = n36585 & n36587 ;
  assign n36590 = ( n13981 & n36588 ) | ( n13981 & n36589 ) | ( n36588 & n36589 ) ;
  assign n36591 = x56 & n36590 ;
  assign n36592 = x56 & ~n36590 ;
  assign n36593 = ( n36590 & ~n36591 ) | ( n36590 & n36592 ) | ( ~n36591 & n36592 ) ;
  assign n36594 = n36579 & ~n36593 ;
  assign n36595 = ~n36579 & n36593 ;
  assign n36596 = n36594 | n36595 ;
  assign n36597 = ~n36371 & n36388 ;
  assign n36598 = n36388 & ~n36597 ;
  assign n36599 = n36371 | n36597 ;
  assign n36600 = ~n36598 & n36599 ;
  assign n36601 = n36385 | n36597 ;
  assign n36602 = ( n36597 & ~n36600 ) | ( n36597 & n36601 ) | ( ~n36600 & n36601 ) ;
  assign n36603 = ~n36596 & n36602 ;
  assign n36604 = n36596 & ~n36602 ;
  assign n36605 = n36603 | n36604 ;
  assign n36606 = x121 & n12574 ;
  assign n36607 = x120 & n12569 ;
  assign n36608 = x119 & ~n12568 ;
  assign n36609 = n13076 & n36608 ;
  assign n36610 = n36607 | n36609 ;
  assign n36611 = n36606 | n36610 ;
  assign n36612 = n12577 | n36606 ;
  assign n36613 = n36610 | n36612 ;
  assign n36614 = ( n15501 & n36611 ) | ( n15501 & n36613 ) | ( n36611 & n36613 ) ;
  assign n36615 = x53 & n36613 ;
  assign n36616 = x53 & n36606 ;
  assign n36617 = ( x53 & n36610 ) | ( x53 & n36616 ) | ( n36610 & n36616 ) ;
  assign n36618 = ( n15501 & n36615 ) | ( n15501 & n36617 ) | ( n36615 & n36617 ) ;
  assign n36619 = x53 & ~n36617 ;
  assign n36620 = x53 & ~n36613 ;
  assign n36621 = ( ~n15501 & n36619 ) | ( ~n15501 & n36620 ) | ( n36619 & n36620 ) ;
  assign n36622 = ( n36614 & ~n36618 ) | ( n36614 & n36621 ) | ( ~n36618 & n36621 ) ;
  assign n36623 = n36605 & ~n36622 ;
  assign n36624 = ~n36605 & n36622 ;
  assign n36625 = n36623 | n36624 ;
  assign n36626 = n36393 | n36420 ;
  assign n36627 = ( n36392 & n36411 ) | ( n36392 & ~n36414 ) | ( n36411 & ~n36414 ) ;
  assign n36628 = ( n36394 & n36626 ) | ( n36394 & n36627 ) | ( n36626 & n36627 ) ;
  assign n36629 = ~n36625 & n36628 ;
  assign n36630 = n36625 & ~n36628 ;
  assign n36631 = n36629 | n36630 ;
  assign n36632 = x124 & n11205 ;
  assign n36633 = x123 & n11200 ;
  assign n36634 = x122 & ~n11199 ;
  assign n36635 = n11679 & n36634 ;
  assign n36636 = n36633 | n36635 ;
  assign n36637 = n36632 | n36636 ;
  assign n36638 = n11208 | n36632 ;
  assign n36639 = n36636 | n36638 ;
  assign n36640 = ( n17084 & n36637 ) | ( n17084 & n36639 ) | ( n36637 & n36639 ) ;
  assign n36641 = x50 & n36639 ;
  assign n36642 = x50 & n36632 ;
  assign n36643 = ( x50 & n36636 ) | ( x50 & n36642 ) | ( n36636 & n36642 ) ;
  assign n36644 = ( n17084 & n36641 ) | ( n17084 & n36643 ) | ( n36641 & n36643 ) ;
  assign n36645 = x50 & ~n36643 ;
  assign n36646 = x50 & ~n36639 ;
  assign n36647 = ( ~n17084 & n36645 ) | ( ~n17084 & n36646 ) | ( n36645 & n36646 ) ;
  assign n36648 = ( n36640 & ~n36644 ) | ( n36640 & n36647 ) | ( ~n36644 & n36647 ) ;
  assign n36649 = n36631 & ~n36648 ;
  assign n36650 = ~n36631 & n36648 ;
  assign n36651 = n36649 | n36650 ;
  assign n36652 = n36422 & ~n36443 ;
  assign n36653 = ( n36423 & n36443 ) | ( n36423 & ~n36652 ) | ( n36443 & ~n36652 ) ;
  assign n36654 = ( n36424 & ~n36426 ) | ( n36424 & n36653 ) | ( ~n36426 & n36653 ) ;
  assign n36655 = ~n36651 & n36654 ;
  assign n36656 = n36651 & ~n36654 ;
  assign n36657 = n36655 | n36656 ;
  assign n36658 = x127 & n9933 ;
  assign n36659 = x126 & n9928 ;
  assign n36660 = x125 & ~n9927 ;
  assign n36661 = n10379 & n36660 ;
  assign n36662 = n36659 | n36661 ;
  assign n36663 = n36658 | n36662 ;
  assign n36664 = n9936 | n36658 ;
  assign n36665 = n36662 | n36664 ;
  assign n36666 = ( n18763 & n36663 ) | ( n18763 & n36665 ) | ( n36663 & n36665 ) ;
  assign n36667 = x47 & n36665 ;
  assign n36668 = x47 & n36658 ;
  assign n36669 = ( x47 & n36662 ) | ( x47 & n36668 ) | ( n36662 & n36668 ) ;
  assign n36670 = ( n18763 & n36667 ) | ( n18763 & n36669 ) | ( n36667 & n36669 ) ;
  assign n36671 = x47 & ~n36669 ;
  assign n36672 = x47 & ~n36665 ;
  assign n36673 = ( ~n18763 & n36671 ) | ( ~n18763 & n36672 ) | ( n36671 & n36672 ) ;
  assign n36674 = ( n36666 & ~n36670 ) | ( n36666 & n36673 ) | ( ~n36670 & n36673 ) ;
  assign n36675 = ~n36657 & n36674 ;
  assign n36676 = n36657 | n36675 ;
  assign n36677 = n36657 & n36674 ;
  assign n36678 = n36676 & ~n36677 ;
  assign n36679 = n36448 | n36468 ;
  assign n36680 = n36448 | n36466 ;
  assign n36681 = ( ~n36449 & n36679 ) | ( ~n36449 & n36680 ) | ( n36679 & n36680 ) ;
  assign n36682 = n36678 & ~n36681 ;
  assign n36683 = ~n36678 & n36681 ;
  assign n36684 = n36682 | n36683 ;
  assign n36685 = ~n36312 & n36473 ;
  assign n36686 = ( n36312 & n36317 ) | ( n36312 & ~n36685 ) | ( n36317 & ~n36685 ) ;
  assign n36687 = ~n36684 & n36686 ;
  assign n36688 = n36684 & ~n36686 ;
  assign n36689 = n36687 | n36688 ;
  assign n36690 = ~n36479 & n36499 ;
  assign n36691 = ~n36479 & n36494 ;
  assign n36692 = n36479 | n36495 ;
  assign n36693 = ( n36270 & ~n36691 ) | ( n36270 & n36692 ) | ( ~n36691 & n36692 ) ;
  assign n36694 = ( n34354 & n36690 ) | ( n34354 & ~n36693 ) | ( n36690 & ~n36693 ) ;
  assign n36695 = ( n34356 & ~n36690 ) | ( n34356 & n36693 ) | ( ~n36690 & n36693 ) ;
  assign n36696 = ( n32844 & n36694 ) | ( n32844 & ~n36695 ) | ( n36694 & ~n36695 ) ;
  assign n36697 = n36479 | n36503 ;
  assign n36698 = ~n36479 & n36481 ;
  assign n36699 = ( n36283 & ~n36692 ) | ( n36283 & n36698 ) | ( ~n36692 & n36698 ) ;
  assign n36700 = ( n35413 & ~n36697 ) | ( n35413 & n36699 ) | ( ~n36697 & n36699 ) ;
  assign n36701 = ( n35414 & n36697 ) | ( n35414 & ~n36699 ) | ( n36697 & ~n36699 ) ;
  assign n36702 = ( n32151 & n36700 ) | ( n32151 & ~n36701 ) | ( n36700 & ~n36701 ) ;
  assign n36703 = ( ~n30751 & n36696 ) | ( ~n30751 & n36702 ) | ( n36696 & n36702 ) ;
  assign n36704 = ( ~n30750 & n36696 ) | ( ~n30750 & n36702 ) | ( n36696 & n36702 ) ;
  assign n36705 = ( ~n25522 & n36703 ) | ( ~n25522 & n36704 ) | ( n36703 & n36704 ) ;
  assign n36706 = ( ~n25519 & n36703 ) | ( ~n25519 & n36704 ) | ( n36703 & n36704 ) ;
  assign n36707 = ( ~n22794 & n36705 ) | ( ~n22794 & n36706 ) | ( n36705 & n36706 ) ;
  assign n36708 = n36689 & n36707 ;
  assign n36709 = n36689 | n36704 ;
  assign n36710 = n36689 | n36703 ;
  assign n36711 = ( ~n25522 & n36709 ) | ( ~n25522 & n36710 ) | ( n36709 & n36710 ) ;
  assign n36712 = ( ~n25519 & n36709 ) | ( ~n25519 & n36710 ) | ( n36709 & n36710 ) ;
  assign n36713 = ( ~n22790 & n36711 ) | ( ~n22790 & n36712 ) | ( n36711 & n36712 ) ;
  assign n36714 = ( ~n22793 & n36711 ) | ( ~n22793 & n36712 ) | ( n36711 & n36712 ) ;
  assign n36715 = ( ~n21078 & n36713 ) | ( ~n21078 & n36714 ) | ( n36713 & n36714 ) ;
  assign n36716 = ~n36708 & n36715 ;
  assign n36717 = x127 & n9928 ;
  assign n36718 = x126 & ~n9927 ;
  assign n36719 = n10379 & n36718 ;
  assign n36720 = n36717 | n36719 ;
  assign n36721 = n9936 | n36720 ;
  assign n36722 = ( n19328 & n36720 ) | ( n19328 & n36721 ) | ( n36720 & n36721 ) ;
  assign n36723 = x47 & n36720 ;
  assign n36724 = ( x47 & n13065 ) | ( x47 & n36720 ) | ( n13065 & n36720 ) ;
  assign n36725 = ( n19328 & n36723 ) | ( n19328 & n36724 ) | ( n36723 & n36724 ) ;
  assign n36726 = x47 & ~n13065 ;
  assign n36727 = ~n36720 & n36726 ;
  assign n36728 = x47 & ~n36720 ;
  assign n36729 = ( ~n19328 & n36727 ) | ( ~n19328 & n36728 ) | ( n36727 & n36728 ) ;
  assign n36730 = ( n36722 & ~n36725 ) | ( n36722 & n36729 ) | ( ~n36725 & n36729 ) ;
  assign n36731 = n36648 & n36730 ;
  assign n36732 = ~n36631 & n36731 ;
  assign n36733 = ( n36655 & n36730 ) | ( n36655 & n36732 ) | ( n36730 & n36732 ) ;
  assign n36734 = n36648 | n36730 ;
  assign n36735 = ( ~n36631 & n36730 ) | ( ~n36631 & n36734 ) | ( n36730 & n36734 ) ;
  assign n36736 = n36655 | n36735 ;
  assign n36737 = ~n36733 & n36736 ;
  assign n36738 = n36556 & ~n36563 ;
  assign n36739 = ( n36539 & n36556 ) | ( n36539 & n36738 ) | ( n36556 & n36738 ) ;
  assign n36740 = n36538 | n36739 ;
  assign n36741 = x110 & n18290 ;
  assign n36742 = x63 & x109 ;
  assign n36743 = ~n18290 & n36742 ;
  assign n36744 = n36741 | n36743 ;
  assign n36745 = n36114 | n36525 ;
  assign n36746 = ( n36525 & ~n36527 ) | ( n36525 & n36745 ) | ( ~n36527 & n36745 ) ;
  assign n36747 = n36744 & ~n36746 ;
  assign n36748 = ~n36744 & n36746 ;
  assign n36749 = n36747 | n36748 ;
  assign n36750 = x113 & n17146 ;
  assign n36751 = x112 & n17141 ;
  assign n36752 = x111 & ~n17140 ;
  assign n36753 = n17724 & n36752 ;
  assign n36754 = n36751 | n36753 ;
  assign n36755 = n36750 | n36754 ;
  assign n36756 = n17149 | n36750 ;
  assign n36757 = n36754 | n36756 ;
  assign n36758 = ( ~n11642 & n36755 ) | ( ~n11642 & n36757 ) | ( n36755 & n36757 ) ;
  assign n36759 = n36755 & n36757 ;
  assign n36760 = ( n11626 & n36758 ) | ( n11626 & n36759 ) | ( n36758 & n36759 ) ;
  assign n36761 = ~x62 & n36760 ;
  assign n36762 = x62 & n36757 ;
  assign n36763 = x62 & x113 ;
  assign n36764 = n17146 & n36763 ;
  assign n36765 = ( x62 & n36754 ) | ( x62 & n36764 ) | ( n36754 & n36764 ) ;
  assign n36766 = ( ~n11642 & n36762 ) | ( ~n11642 & n36765 ) | ( n36762 & n36765 ) ;
  assign n36767 = n36762 & n36765 ;
  assign n36768 = ( n11626 & n36766 ) | ( n11626 & n36767 ) | ( n36766 & n36767 ) ;
  assign n36769 = x62 & ~n36749 ;
  assign n36770 = ~n36768 & n36769 ;
  assign n36771 = ( ~n36749 & n36761 ) | ( ~n36749 & n36770 ) | ( n36761 & n36770 ) ;
  assign n36772 = ~x62 & n36749 ;
  assign n36773 = ( n36749 & n36768 ) | ( n36749 & n36772 ) | ( n36768 & n36772 ) ;
  assign n36774 = ~n36761 & n36773 ;
  assign n36775 = n36771 | n36774 ;
  assign n36776 = n36538 & ~n36775 ;
  assign n36777 = ( n36739 & ~n36775 ) | ( n36739 & n36776 ) | ( ~n36775 & n36776 ) ;
  assign n36778 = n36740 & ~n36777 ;
  assign n36779 = x116 & n15552 ;
  assign n36780 = x115 & n15547 ;
  assign n36781 = x114 & ~n15546 ;
  assign n36782 = n16123 & n36781 ;
  assign n36783 = n36780 | n36782 ;
  assign n36784 = n36779 | n36783 ;
  assign n36785 = n15555 | n36779 ;
  assign n36786 = n36783 | n36785 ;
  assign n36787 = ( ~n13040 & n36784 ) | ( ~n13040 & n36786 ) | ( n36784 & n36786 ) ;
  assign n36788 = n36784 & n36786 ;
  assign n36789 = ( n13022 & n36787 ) | ( n13022 & n36788 ) | ( n36787 & n36788 ) ;
  assign n36790 = x59 & n36789 ;
  assign n36791 = x59 & ~n36789 ;
  assign n36792 = ( n36789 & ~n36790 ) | ( n36789 & n36791 ) | ( ~n36790 & n36791 ) ;
  assign n36793 = n36538 | n36775 ;
  assign n36794 = n36739 | n36793 ;
  assign n36795 = ~n36792 & n36794 ;
  assign n36796 = ~n36778 & n36795 ;
  assign n36797 = n36792 & ~n36794 ;
  assign n36798 = ( n36778 & n36792 ) | ( n36778 & n36797 ) | ( n36792 & n36797 ) ;
  assign n36799 = n36796 | n36798 ;
  assign n36800 = n36569 | n36576 ;
  assign n36801 = ( n36569 & ~n36572 ) | ( n36569 & n36800 ) | ( ~n36572 & n36800 ) ;
  assign n36802 = ~n36799 & n36801 ;
  assign n36803 = n36799 & ~n36801 ;
  assign n36804 = n36802 | n36803 ;
  assign n36805 = x119 & n14045 ;
  assign n36806 = x118 & n14040 ;
  assign n36807 = x117 & ~n14039 ;
  assign n36808 = n14552 & n36807 ;
  assign n36809 = n36806 | n36808 ;
  assign n36810 = n36805 | n36809 ;
  assign n36811 = n14048 | n36805 ;
  assign n36812 = n36809 | n36811 ;
  assign n36813 = ( n14496 & n36810 ) | ( n14496 & n36812 ) | ( n36810 & n36812 ) ;
  assign n36814 = x56 & n36812 ;
  assign n36815 = x56 & n36805 ;
  assign n36816 = ( x56 & n36809 ) | ( x56 & n36815 ) | ( n36809 & n36815 ) ;
  assign n36817 = ( n14496 & n36814 ) | ( n14496 & n36816 ) | ( n36814 & n36816 ) ;
  assign n36818 = x56 & ~n36816 ;
  assign n36819 = x56 & ~n36812 ;
  assign n36820 = ( ~n14496 & n36818 ) | ( ~n14496 & n36819 ) | ( n36818 & n36819 ) ;
  assign n36821 = ( n36813 & ~n36817 ) | ( n36813 & n36820 ) | ( ~n36817 & n36820 ) ;
  assign n36822 = n36804 | n36821 ;
  assign n36823 = n36804 & ~n36821 ;
  assign n36824 = ( ~n36804 & n36822 ) | ( ~n36804 & n36823 ) | ( n36822 & n36823 ) ;
  assign n36825 = n36595 | n36603 ;
  assign n36826 = n36824 & n36825 ;
  assign n36827 = n36824 | n36825 ;
  assign n36828 = ~n36826 & n36827 ;
  assign n36829 = x122 & n12574 ;
  assign n36830 = x121 & n12569 ;
  assign n36831 = x120 & ~n12568 ;
  assign n36832 = n13076 & n36831 ;
  assign n36833 = n36830 | n36832 ;
  assign n36834 = n36829 | n36833 ;
  assign n36835 = n12577 | n36829 ;
  assign n36836 = n36833 | n36835 ;
  assign n36837 = ( n16043 & n36834 ) | ( n16043 & n36836 ) | ( n36834 & n36836 ) ;
  assign n36838 = x53 & n36836 ;
  assign n36839 = x53 & n36829 ;
  assign n36840 = ( x53 & n36833 ) | ( x53 & n36839 ) | ( n36833 & n36839 ) ;
  assign n36841 = ( n16043 & n36838 ) | ( n16043 & n36840 ) | ( n36838 & n36840 ) ;
  assign n36842 = x53 & ~n36840 ;
  assign n36843 = x53 & ~n36836 ;
  assign n36844 = ( ~n16043 & n36842 ) | ( ~n16043 & n36843 ) | ( n36842 & n36843 ) ;
  assign n36845 = ( n36837 & ~n36841 ) | ( n36837 & n36844 ) | ( ~n36841 & n36844 ) ;
  assign n36846 = n36828 & ~n36845 ;
  assign n36847 = ~n36828 & n36845 ;
  assign n36848 = n36846 | n36847 ;
  assign n36849 = n36624 | n36628 ;
  assign n36850 = ( n36624 & ~n36625 ) | ( n36624 & n36849 ) | ( ~n36625 & n36849 ) ;
  assign n36851 = ~n36848 & n36850 ;
  assign n36852 = n36848 | n36851 ;
  assign n36853 = x125 & n11205 ;
  assign n36854 = x124 & n11200 ;
  assign n36855 = x123 & ~n11199 ;
  assign n36856 = n11679 & n36855 ;
  assign n36857 = n36854 | n36856 ;
  assign n36858 = n36853 | n36857 ;
  assign n36859 = n11208 | n36853 ;
  assign n36860 = n36857 | n36859 ;
  assign n36861 = ( n17670 & n36858 ) | ( n17670 & n36860 ) | ( n36858 & n36860 ) ;
  assign n36862 = x50 & n36860 ;
  assign n36863 = x50 & n36853 ;
  assign n36864 = ( x50 & n36857 ) | ( x50 & n36863 ) | ( n36857 & n36863 ) ;
  assign n36865 = ( n17670 & n36862 ) | ( n17670 & n36864 ) | ( n36862 & n36864 ) ;
  assign n36866 = x50 & ~n36864 ;
  assign n36867 = x50 & ~n36860 ;
  assign n36868 = ( ~n17670 & n36866 ) | ( ~n17670 & n36867 ) | ( n36866 & n36867 ) ;
  assign n36869 = ( n36861 & ~n36865 ) | ( n36861 & n36868 ) | ( ~n36865 & n36868 ) ;
  assign n36870 = ~n36850 & n36869 ;
  assign n36871 = ( ~n36848 & n36869 ) | ( ~n36848 & n36870 ) | ( n36869 & n36870 ) ;
  assign n36872 = n36852 & n36871 ;
  assign n36873 = n36850 & ~n36869 ;
  assign n36874 = n36848 & n36873 ;
  assign n36875 = ( n36852 & n36869 ) | ( n36852 & ~n36874 ) | ( n36869 & ~n36874 ) ;
  assign n36876 = ~n36872 & n36875 ;
  assign n36877 = n36737 & ~n36876 ;
  assign n36878 = n36737 | n36876 ;
  assign n36879 = ( ~n36737 & n36877 ) | ( ~n36737 & n36878 ) | ( n36877 & n36878 ) ;
  assign n36880 = n36675 & ~n36879 ;
  assign n36881 = ( n36683 & ~n36879 ) | ( n36683 & n36880 ) | ( ~n36879 & n36880 ) ;
  assign n36882 = ~n36675 & n36879 ;
  assign n36883 = ~n36683 & n36882 ;
  assign n36884 = n36881 | n36883 ;
  assign n36885 = ~n36687 & n36715 ;
  assign n36886 = n36884 & n36885 ;
  assign n36887 = n36687 & ~n36884 ;
  assign n36888 = ( n36715 & n36884 ) | ( n36715 & ~n36887 ) | ( n36884 & ~n36887 ) ;
  assign n36889 = ~n36886 & n36888 ;
  assign n36890 = x127 & ~n9927 ;
  assign n36891 = n10379 & n36890 ;
  assign n36892 = n9936 | n36891 ;
  assign n36893 = n19877 | n36891 ;
  assign n36894 = n36892 & n36893 ;
  assign n36895 = n19880 | n36891 ;
  assign n36896 = n36892 & n36895 ;
  assign n36897 = ( n18202 & n36894 ) | ( n18202 & n36896 ) | ( n36894 & n36896 ) ;
  assign n36898 = n36894 & n36896 ;
  assign n36899 = ( n18212 & n36897 ) | ( n18212 & n36898 ) | ( n36897 & n36898 ) ;
  assign n36900 = ( n18214 & n36897 ) | ( n18214 & n36898 ) | ( n36897 & n36898 ) ;
  assign n36901 = ( n14002 & n36899 ) | ( n14002 & n36900 ) | ( n36899 & n36900 ) ;
  assign n36902 = x47 & n36899 ;
  assign n36903 = x47 & n36900 ;
  assign n36904 = ( n14002 & n36902 ) | ( n14002 & n36903 ) | ( n36902 & n36903 ) ;
  assign n36905 = x47 & ~n36903 ;
  assign n36906 = x47 & ~n36902 ;
  assign n36907 = ( ~n14002 & n36905 ) | ( ~n14002 & n36906 ) | ( n36905 & n36906 ) ;
  assign n36908 = ( n36901 & ~n36904 ) | ( n36901 & n36907 ) | ( ~n36904 & n36907 ) ;
  assign n36909 = n36848 & n36850 ;
  assign n36910 = n36850 | n36869 ;
  assign n36911 = ( ~n36848 & n36869 ) | ( ~n36848 & n36910 ) | ( n36869 & n36910 ) ;
  assign n36912 = ( n36851 & n36909 ) | ( n36851 & n36911 ) | ( n36909 & n36911 ) ;
  assign n36913 = n36851 | n36911 ;
  assign n36914 = ( ~n36852 & n36912 ) | ( ~n36852 & n36913 ) | ( n36912 & n36913 ) ;
  assign n36915 = n36908 & n36914 ;
  assign n36916 = n36908 | n36914 ;
  assign n36917 = ~n36915 & n36916 ;
  assign n36918 = n36777 | n36798 ;
  assign n36919 = n36748 | n36771 ;
  assign n36920 = x111 & n18290 ;
  assign n36921 = x63 & x110 ;
  assign n36922 = ~n18290 & n36921 ;
  assign n36923 = n36920 | n36922 ;
  assign n36924 = ~n36744 & n36923 ;
  assign n36925 = n36744 & ~n36923 ;
  assign n36926 = n36924 | n36925 ;
  assign n36927 = n36744 | n36926 ;
  assign n36928 = n36746 & ~n36927 ;
  assign n36929 = ( n36771 & ~n36926 ) | ( n36771 & n36928 ) | ( ~n36926 & n36928 ) ;
  assign n36930 = n36919 & ~n36929 ;
  assign n36931 = x114 & n17146 ;
  assign n36932 = x113 & n17141 ;
  assign n36933 = x112 & ~n17140 ;
  assign n36934 = n17724 & n36933 ;
  assign n36935 = n36932 | n36934 ;
  assign n36936 = n36931 | n36935 ;
  assign n36937 = n17149 | n36931 ;
  assign n36938 = n36935 | n36937 ;
  assign n36939 = ( ~n12095 & n36936 ) | ( ~n12095 & n36938 ) | ( n36936 & n36938 ) ;
  assign n36940 = n36936 & n36938 ;
  assign n36941 = ( n12079 & n36939 ) | ( n12079 & n36940 ) | ( n36939 & n36940 ) ;
  assign n36942 = x62 & n36941 ;
  assign n36943 = x62 & ~n36941 ;
  assign n36944 = ( n36941 & ~n36942 ) | ( n36941 & n36943 ) | ( ~n36942 & n36943 ) ;
  assign n36945 = n36926 | n36928 ;
  assign n36946 = n36771 | n36945 ;
  assign n36947 = n36944 | n36946 ;
  assign n36948 = ( ~n36930 & n36944 ) | ( ~n36930 & n36947 ) | ( n36944 & n36947 ) ;
  assign n36949 = n36944 & n36946 ;
  assign n36950 = ~n36930 & n36949 ;
  assign n36951 = n36948 & ~n36950 ;
  assign n36952 = x117 & n15552 ;
  assign n36953 = x116 & n15547 ;
  assign n36954 = x115 & ~n15546 ;
  assign n36955 = n16123 & n36954 ;
  assign n36956 = n36953 | n36955 ;
  assign n36957 = n36952 | n36956 ;
  assign n36958 = n15555 | n36952 ;
  assign n36959 = n36956 | n36958 ;
  assign n36960 = ( ~n13522 & n36957 ) | ( ~n13522 & n36959 ) | ( n36957 & n36959 ) ;
  assign n36961 = n36957 & n36959 ;
  assign n36962 = ( n13503 & n36960 ) | ( n13503 & n36961 ) | ( n36960 & n36961 ) ;
  assign n36963 = x59 & n36962 ;
  assign n36964 = x59 & ~n36962 ;
  assign n36965 = ( n36962 & ~n36963 ) | ( n36962 & n36964 ) | ( ~n36963 & n36964 ) ;
  assign n36966 = ~n36951 & n36965 ;
  assign n36967 = n36951 & ~n36965 ;
  assign n36968 = n36966 | n36967 ;
  assign n36969 = n36918 & ~n36968 ;
  assign n36970 = n36918 & ~n36969 ;
  assign n36971 = n36968 | n36969 ;
  assign n36972 = ~n36970 & n36971 ;
  assign n36973 = x120 & n14045 ;
  assign n36974 = x119 & n14040 ;
  assign n36975 = x118 & ~n14039 ;
  assign n36976 = n14552 & n36975 ;
  assign n36977 = n36974 | n36976 ;
  assign n36978 = n36973 | n36977 ;
  assign n36979 = n14048 | n36973 ;
  assign n36980 = n36977 | n36979 ;
  assign n36981 = ( n14991 & n36978 ) | ( n14991 & n36980 ) | ( n36978 & n36980 ) ;
  assign n36982 = x56 & n36980 ;
  assign n36983 = x56 & n36973 ;
  assign n36984 = ( x56 & n36977 ) | ( x56 & n36983 ) | ( n36977 & n36983 ) ;
  assign n36985 = ( n14991 & n36982 ) | ( n14991 & n36984 ) | ( n36982 & n36984 ) ;
  assign n36986 = x56 & ~n36984 ;
  assign n36987 = x56 & ~n36980 ;
  assign n36988 = ( ~n14991 & n36986 ) | ( ~n14991 & n36987 ) | ( n36986 & n36987 ) ;
  assign n36989 = ( n36981 & ~n36985 ) | ( n36981 & n36988 ) | ( ~n36985 & n36988 ) ;
  assign n36990 = ~n36972 & n36989 ;
  assign n36991 = n36968 & ~n36989 ;
  assign n36992 = ( n36969 & ~n36989 ) | ( n36969 & n36991 ) | ( ~n36989 & n36991 ) ;
  assign n36993 = ~n36970 & n36992 ;
  assign n36994 = n36802 | n36821 ;
  assign n36995 = ( n36802 & ~n36804 ) | ( n36802 & n36994 ) | ( ~n36804 & n36994 ) ;
  assign n36996 = ~n36993 & n36995 ;
  assign n36997 = ~n36990 & n36996 ;
  assign n36998 = n36993 & ~n36995 ;
  assign n36999 = ( n36990 & ~n36995 ) | ( n36990 & n36998 ) | ( ~n36995 & n36998 ) ;
  assign n37000 = n36997 | n36999 ;
  assign n37001 = x123 & n12574 ;
  assign n37002 = x122 & n12569 ;
  assign n37003 = x121 & ~n12568 ;
  assign n37004 = n13076 & n37003 ;
  assign n37005 = n37002 | n37004 ;
  assign n37006 = n37001 | n37005 ;
  assign n37007 = n12577 | n37001 ;
  assign n37008 = n37005 | n37007 ;
  assign n37009 = ( n16086 & n37006 ) | ( n16086 & n37008 ) | ( n37006 & n37008 ) ;
  assign n37010 = x53 & n37008 ;
  assign n37011 = x53 & n37001 ;
  assign n37012 = ( x53 & n37005 ) | ( x53 & n37011 ) | ( n37005 & n37011 ) ;
  assign n37013 = ( n16086 & n37010 ) | ( n16086 & n37012 ) | ( n37010 & n37012 ) ;
  assign n37014 = x53 & ~n37012 ;
  assign n37015 = x53 & ~n37008 ;
  assign n37016 = ( ~n16086 & n37014 ) | ( ~n16086 & n37015 ) | ( n37014 & n37015 ) ;
  assign n37017 = ( n37009 & ~n37013 ) | ( n37009 & n37016 ) | ( ~n37013 & n37016 ) ;
  assign n37018 = n37000 | n37017 ;
  assign n37019 = n37000 & ~n37017 ;
  assign n37020 = ( ~n37000 & n37018 ) | ( ~n37000 & n37019 ) | ( n37018 & n37019 ) ;
  assign n37021 = ( ~n36824 & n36825 ) | ( ~n36824 & n36845 ) | ( n36825 & n36845 ) ;
  assign n37022 = ~n37020 & n37021 ;
  assign n37023 = n37020 | n37022 ;
  assign n37024 = x126 & n11205 ;
  assign n37025 = x125 & n11200 ;
  assign n37026 = x124 & ~n11199 ;
  assign n37027 = n11679 & n37026 ;
  assign n37028 = n37025 | n37027 ;
  assign n37029 = n37024 | n37028 ;
  assign n37030 = n11208 | n37024 ;
  assign n37031 = n37028 | n37030 ;
  assign n37032 = ( n18220 & n37029 ) | ( n18220 & n37031 ) | ( n37029 & n37031 ) ;
  assign n37033 = x50 & n37031 ;
  assign n37034 = x50 & n37024 ;
  assign n37035 = ( x50 & n37028 ) | ( x50 & n37034 ) | ( n37028 & n37034 ) ;
  assign n37036 = ( n18220 & n37033 ) | ( n18220 & n37035 ) | ( n37033 & n37035 ) ;
  assign n37037 = x50 & ~n37035 ;
  assign n37038 = x50 & ~n37031 ;
  assign n37039 = ( ~n18220 & n37037 ) | ( ~n18220 & n37038 ) | ( n37037 & n37038 ) ;
  assign n37040 = ( n37032 & ~n37036 ) | ( n37032 & n37039 ) | ( ~n37036 & n37039 ) ;
  assign n37041 = n37021 & n37040 ;
  assign n37042 = n37020 & n37041 ;
  assign n37043 = ( ~n37023 & n37040 ) | ( ~n37023 & n37042 ) | ( n37040 & n37042 ) ;
  assign n37044 = n37021 | n37040 ;
  assign n37045 = ( n37020 & n37040 ) | ( n37020 & n37044 ) | ( n37040 & n37044 ) ;
  assign n37046 = n37023 & ~n37045 ;
  assign n37047 = n37043 | n37046 ;
  assign n37048 = n36917 & ~n37047 ;
  assign n37049 = n36917 & ~n37048 ;
  assign n37050 = ~n36733 & n36876 ;
  assign n37051 = ( n36733 & n36737 ) | ( n36733 & ~n37050 ) | ( n36737 & ~n37050 ) ;
  assign n37052 = n36917 | n37047 ;
  assign n37053 = n37051 & ~n37052 ;
  assign n37054 = ( n37049 & n37051 ) | ( n37049 & n37053 ) | ( n37051 & n37053 ) ;
  assign n37055 = ~n37051 & n37052 ;
  assign n37056 = ~n37049 & n37055 ;
  assign n37057 = n37054 | n37056 ;
  assign n37058 = ~n36881 & n36884 ;
  assign n37059 = ( n36687 & n36881 ) | ( n36687 & ~n37058 ) | ( n36881 & ~n37058 ) ;
  assign n37060 = ( n36715 & n37058 ) | ( n36715 & ~n37059 ) | ( n37058 & ~n37059 ) ;
  assign n37061 = n37057 & n37060 ;
  assign n37062 = ~n37057 & n37059 ;
  assign n37063 = n36881 & ~n37057 ;
  assign n37064 = ( n36884 & n37057 ) | ( n36884 & ~n37063 ) | ( n37057 & ~n37063 ) ;
  assign n37065 = ( n36715 & ~n37062 ) | ( n36715 & n37064 ) | ( ~n37062 & n37064 ) ;
  assign n37066 = ~n37061 & n37065 ;
  assign n37067 = x118 & n15552 ;
  assign n37068 = x117 & n15547 ;
  assign n37069 = x116 & ~n15546 ;
  assign n37070 = n16123 & n37069 ;
  assign n37071 = n37068 | n37070 ;
  assign n37072 = n37067 | n37071 ;
  assign n37073 = n15555 | n37067 ;
  assign n37074 = n37071 | n37073 ;
  assign n37075 = ( ~n14002 & n37072 ) | ( ~n14002 & n37074 ) | ( n37072 & n37074 ) ;
  assign n37076 = n37072 & n37074 ;
  assign n37077 = ( n13981 & n37075 ) | ( n13981 & n37076 ) | ( n37075 & n37076 ) ;
  assign n37078 = x59 & n37077 ;
  assign n37079 = x59 & ~n37077 ;
  assign n37080 = ( n37077 & ~n37078 ) | ( n37077 & n37079 ) | ( ~n37078 & n37079 ) ;
  assign n37081 = n36925 | n36928 ;
  assign n37082 = ~n36925 & n36926 ;
  assign n37083 = ( n36771 & n37081 ) | ( n36771 & ~n37082 ) | ( n37081 & ~n37082 ) ;
  assign n37084 = x115 & n17146 ;
  assign n37085 = x114 & n17141 ;
  assign n37086 = x113 & ~n17140 ;
  assign n37087 = n17724 & n37086 ;
  assign n37088 = n37085 | n37087 ;
  assign n37089 = n37084 | n37088 ;
  assign n37090 = n17149 | n37084 ;
  assign n37091 = n37088 | n37090 ;
  assign n37092 = ( ~n12550 & n37089 ) | ( ~n12550 & n37091 ) | ( n37089 & n37091 ) ;
  assign n37093 = n37089 & n37091 ;
  assign n37094 = ( n12532 & n37092 ) | ( n12532 & n37093 ) | ( n37092 & n37093 ) ;
  assign n37095 = ~x62 & n37094 ;
  assign n37096 = x62 & n37091 ;
  assign n37097 = x62 & x115 ;
  assign n37098 = n17146 & n37097 ;
  assign n37099 = ( x62 & n37088 ) | ( x62 & n37098 ) | ( n37088 & n37098 ) ;
  assign n37100 = ( ~n12550 & n37096 ) | ( ~n12550 & n37099 ) | ( n37096 & n37099 ) ;
  assign n37101 = n37096 & n37099 ;
  assign n37102 = ( n12532 & n37100 ) | ( n12532 & n37101 ) | ( n37100 & n37101 ) ;
  assign n37103 = x62 & ~n37102 ;
  assign n37104 = n37095 | n37103 ;
  assign n37105 = x112 & n18290 ;
  assign n37106 = x63 & x111 ;
  assign n37107 = ~n18290 & n37106 ;
  assign n37108 = n37105 | n37107 ;
  assign n37109 = x47 & n36923 ;
  assign n37110 = x47 | n36923 ;
  assign n37111 = ~n37109 & n37110 ;
  assign n37112 = n37108 & ~n37111 ;
  assign n37113 = ~n37108 & n37111 ;
  assign n37114 = n37112 | n37113 ;
  assign n37115 = n37104 & ~n37114 ;
  assign n37116 = ~n37104 & n37114 ;
  assign n37117 = n37115 | n37116 ;
  assign n37118 = n37083 | n37117 ;
  assign n37119 = n37080 & n37083 ;
  assign n37120 = n37117 & n37119 ;
  assign n37121 = ( n37080 & ~n37118 ) | ( n37080 & n37120 ) | ( ~n37118 & n37120 ) ;
  assign n37122 = n37080 | n37083 ;
  assign n37123 = ( n37080 & n37117 ) | ( n37080 & n37122 ) | ( n37117 & n37122 ) ;
  assign n37124 = n37118 & ~n37123 ;
  assign n37125 = n37121 | n37124 ;
  assign n37126 = ( n36944 & ~n36946 ) | ( n36944 & n36965 ) | ( ~n36946 & n36965 ) ;
  assign n37127 = n36944 | n36965 ;
  assign n37128 = ( n36930 & n37126 ) | ( n36930 & n37127 ) | ( n37126 & n37127 ) ;
  assign n37129 = ~n37125 & n37128 ;
  assign n37130 = n37125 & ~n37128 ;
  assign n37131 = n37129 | n37130 ;
  assign n37132 = x121 & n14045 ;
  assign n37133 = x120 & n14040 ;
  assign n37134 = x119 & ~n14039 ;
  assign n37135 = n14552 & n37134 ;
  assign n37136 = n37133 | n37135 ;
  assign n37137 = n37132 | n37136 ;
  assign n37138 = n14048 | n37132 ;
  assign n37139 = n37136 | n37138 ;
  assign n37140 = ( n15501 & n37137 ) | ( n15501 & n37139 ) | ( n37137 & n37139 ) ;
  assign n37141 = x56 & n37139 ;
  assign n37142 = x56 & n37132 ;
  assign n37143 = ( x56 & n37136 ) | ( x56 & n37142 ) | ( n37136 & n37142 ) ;
  assign n37144 = ( n15501 & n37141 ) | ( n15501 & n37143 ) | ( n37141 & n37143 ) ;
  assign n37145 = x56 & ~n37143 ;
  assign n37146 = x56 & ~n37139 ;
  assign n37147 = ( ~n15501 & n37145 ) | ( ~n15501 & n37146 ) | ( n37145 & n37146 ) ;
  assign n37148 = ( n37140 & ~n37144 ) | ( n37140 & n37147 ) | ( ~n37144 & n37147 ) ;
  assign n37149 = n37131 & ~n37148 ;
  assign n37150 = ~n37131 & n37148 ;
  assign n37151 = n37149 | n37150 ;
  assign n37152 = n36969 | n36989 ;
  assign n37153 = ( n36969 & ~n36972 ) | ( n36969 & n37152 ) | ( ~n36972 & n37152 ) ;
  assign n37154 = ~n37151 & n37153 ;
  assign n37155 = n37151 & ~n37153 ;
  assign n37156 = n37154 | n37155 ;
  assign n37157 = x124 & n12574 ;
  assign n37158 = x123 & n12569 ;
  assign n37159 = x122 & ~n12568 ;
  assign n37160 = n13076 & n37159 ;
  assign n37161 = n37158 | n37160 ;
  assign n37162 = n37157 | n37161 ;
  assign n37163 = n12577 | n37157 ;
  assign n37164 = n37161 | n37163 ;
  assign n37165 = ( n17084 & n37162 ) | ( n17084 & n37164 ) | ( n37162 & n37164 ) ;
  assign n37166 = x53 & n37164 ;
  assign n37167 = x53 & n37157 ;
  assign n37168 = ( x53 & n37161 ) | ( x53 & n37167 ) | ( n37161 & n37167 ) ;
  assign n37169 = ( n17084 & n37166 ) | ( n17084 & n37168 ) | ( n37166 & n37168 ) ;
  assign n37170 = x53 & ~n37168 ;
  assign n37171 = x53 & ~n37164 ;
  assign n37172 = ( ~n17084 & n37170 ) | ( ~n17084 & n37171 ) | ( n37170 & n37171 ) ;
  assign n37173 = ( n37165 & ~n37169 ) | ( n37165 & n37172 ) | ( ~n37169 & n37172 ) ;
  assign n37174 = n37156 & ~n37173 ;
  assign n37175 = ~n37156 & n37173 ;
  assign n37176 = n37174 | n37175 ;
  assign n37177 = n36997 | n37017 ;
  assign n37178 = ( n36997 & ~n37000 ) | ( n36997 & n37177 ) | ( ~n37000 & n37177 ) ;
  assign n37179 = ~n37176 & n37178 ;
  assign n37180 = n37176 & ~n37178 ;
  assign n37181 = n37179 | n37180 ;
  assign n37182 = x127 & n11205 ;
  assign n37183 = x126 & n11200 ;
  assign n37184 = x125 & ~n11199 ;
  assign n37185 = n11679 & n37184 ;
  assign n37186 = n37183 | n37185 ;
  assign n37187 = n37182 | n37186 ;
  assign n37188 = n11208 | n37182 ;
  assign n37189 = n37186 | n37188 ;
  assign n37190 = ( n18763 & n37187 ) | ( n18763 & n37189 ) | ( n37187 & n37189 ) ;
  assign n37191 = x50 & n37189 ;
  assign n37192 = x50 & n37182 ;
  assign n37193 = ( x50 & n37186 ) | ( x50 & n37192 ) | ( n37186 & n37192 ) ;
  assign n37194 = ( n18763 & n37191 ) | ( n18763 & n37193 ) | ( n37191 & n37193 ) ;
  assign n37195 = x50 & ~n37193 ;
  assign n37196 = x50 & ~n37189 ;
  assign n37197 = ( ~n18763 & n37195 ) | ( ~n18763 & n37196 ) | ( n37195 & n37196 ) ;
  assign n37198 = ( n37190 & ~n37194 ) | ( n37190 & n37197 ) | ( ~n37194 & n37197 ) ;
  assign n37199 = ~n37181 & n37198 ;
  assign n37200 = n37181 | n37199 ;
  assign n37201 = n37181 & n37198 ;
  assign n37202 = n37022 | n37042 ;
  assign n37203 = n37022 | n37040 ;
  assign n37204 = ( ~n37023 & n37202 ) | ( ~n37023 & n37203 ) | ( n37202 & n37203 ) ;
  assign n37205 = n37201 | n37204 ;
  assign n37206 = n37200 & ~n37205 ;
  assign n37207 = n37201 & n37204 ;
  assign n37208 = ( ~n37200 & n37204 ) | ( ~n37200 & n37207 ) | ( n37204 & n37207 ) ;
  assign n37209 = n37206 | n37208 ;
  assign n37210 = ~n36915 & n37047 ;
  assign n37211 = ( n36915 & n36917 ) | ( n36915 & ~n37210 ) | ( n36917 & ~n37210 ) ;
  assign n37212 = n37209 & ~n37211 ;
  assign n37213 = ~n37209 & n37211 ;
  assign n37214 = n37212 | n37213 ;
  assign n37215 = ~n37054 & n37064 ;
  assign n37216 = ~n37054 & n37057 ;
  assign n37217 = ( n37054 & n37059 ) | ( n37054 & ~n37216 ) | ( n37059 & ~n37216 ) ;
  assign n37218 = ( n36715 & n37215 ) | ( n36715 & ~n37217 ) | ( n37215 & ~n37217 ) ;
  assign n37219 = n37214 & n37218 ;
  assign n37220 = n37054 & ~n37214 ;
  assign n37221 = ( n37057 & n37214 ) | ( n37057 & ~n37220 ) | ( n37214 & ~n37220 ) ;
  assign n37222 = ( n37059 & n37220 ) | ( n37059 & ~n37221 ) | ( n37220 & ~n37221 ) ;
  assign n37223 = ( n37064 & n37214 ) | ( n37064 & ~n37220 ) | ( n37214 & ~n37220 ) ;
  assign n37224 = ( n36715 & ~n37222 ) | ( n36715 & n37223 ) | ( ~n37222 & n37223 ) ;
  assign n37225 = ~n37219 & n37224 ;
  assign n37305 = ~n37150 & n37151 ;
  assign n37306 = ( n37150 & n37153 ) | ( n37150 & ~n37305 ) | ( n37153 & ~n37305 ) ;
  assign n37252 = n37083 | n37115 ;
  assign n37253 = ( n37115 & ~n37117 ) | ( n37115 & n37252 ) | ( ~n37117 & n37252 ) ;
  assign n37226 = x113 & n18290 ;
  assign n37227 = x63 & x112 ;
  assign n37228 = ~n18290 & n37227 ;
  assign n37229 = n37226 | n37228 ;
  assign n37230 = ( ~x47 & n36923 ) | ( ~x47 & n37108 ) | ( n36923 & n37108 ) ;
  assign n37231 = ~n37229 & n37230 ;
  assign n37232 = n37229 & ~n37230 ;
  assign n37233 = n37231 | n37232 ;
  assign n37235 = x115 & n17141 ;
  assign n37236 = x114 & ~n17140 ;
  assign n37237 = n17724 & n37236 ;
  assign n37238 = n37235 | n37237 ;
  assign n37234 = x116 & n17146 ;
  assign n37240 = n17149 | n37234 ;
  assign n37241 = n37238 | n37240 ;
  assign n37239 = n37234 | n37238 ;
  assign n37242 = n37239 & n37241 ;
  assign n37243 = ( ~n13040 & n37241 ) | ( ~n13040 & n37242 ) | ( n37241 & n37242 ) ;
  assign n37244 = n37241 & n37242 ;
  assign n37245 = ( n13022 & n37243 ) | ( n13022 & n37244 ) | ( n37243 & n37244 ) ;
  assign n37246 = x62 & n37245 ;
  assign n37247 = x62 & ~n37245 ;
  assign n37248 = ( n37245 & ~n37246 ) | ( n37245 & n37247 ) | ( ~n37246 & n37247 ) ;
  assign n37249 = ~n37233 & n37248 ;
  assign n37250 = n37233 & ~n37248 ;
  assign n37251 = n37249 | n37250 ;
  assign n37254 = ~n37251 & n37253 ;
  assign n37255 = n37253 & ~n37254 ;
  assign n37256 = x119 & n15552 ;
  assign n37257 = x118 & n15547 ;
  assign n37258 = x117 & ~n15546 ;
  assign n37259 = n16123 & n37258 ;
  assign n37260 = n37257 | n37259 ;
  assign n37261 = n37256 | n37260 ;
  assign n37262 = n15555 | n37256 ;
  assign n37263 = n37260 | n37262 ;
  assign n37264 = ( n14496 & n37261 ) | ( n14496 & n37263 ) | ( n37261 & n37263 ) ;
  assign n37265 = x59 & n37263 ;
  assign n37266 = x59 & n37256 ;
  assign n37267 = ( x59 & n37260 ) | ( x59 & n37266 ) | ( n37260 & n37266 ) ;
  assign n37268 = ( n14496 & n37265 ) | ( n14496 & n37267 ) | ( n37265 & n37267 ) ;
  assign n37269 = x59 & ~n37267 ;
  assign n37270 = x59 & ~n37263 ;
  assign n37271 = ( ~n14496 & n37269 ) | ( ~n14496 & n37270 ) | ( n37269 & n37270 ) ;
  assign n37272 = ( n37264 & ~n37268 ) | ( n37264 & n37271 ) | ( ~n37268 & n37271 ) ;
  assign n37273 = n37251 & ~n37272 ;
  assign n37274 = ( n37253 & ~n37272 ) | ( n37253 & n37273 ) | ( ~n37272 & n37273 ) ;
  assign n37275 = ~n37255 & n37274 ;
  assign n37276 = ~n37251 & n37272 ;
  assign n37277 = ~n37253 & n37276 ;
  assign n37278 = ( n37255 & n37272 ) | ( n37255 & n37277 ) | ( n37272 & n37277 ) ;
  assign n37279 = n37275 | n37278 ;
  assign n37280 = n37121 | n37128 ;
  assign n37281 = ( n37121 & ~n37125 ) | ( n37121 & n37280 ) | ( ~n37125 & n37280 ) ;
  assign n37282 = ~n37279 & n37281 ;
  assign n37283 = n37279 & ~n37281 ;
  assign n37284 = n37282 | n37283 ;
  assign n37285 = x122 & n14045 ;
  assign n37286 = x121 & n14040 ;
  assign n37287 = x120 & ~n14039 ;
  assign n37288 = n14552 & n37287 ;
  assign n37289 = n37286 | n37288 ;
  assign n37290 = n37285 | n37289 ;
  assign n37291 = n14048 | n37285 ;
  assign n37292 = n37289 | n37291 ;
  assign n37293 = ( n16043 & n37290 ) | ( n16043 & n37292 ) | ( n37290 & n37292 ) ;
  assign n37294 = x56 & n37292 ;
  assign n37295 = x56 & n37285 ;
  assign n37296 = ( x56 & n37289 ) | ( x56 & n37295 ) | ( n37289 & n37295 ) ;
  assign n37297 = ( n16043 & n37294 ) | ( n16043 & n37296 ) | ( n37294 & n37296 ) ;
  assign n37298 = x56 & ~n37296 ;
  assign n37299 = x56 & ~n37292 ;
  assign n37300 = ( ~n16043 & n37298 ) | ( ~n16043 & n37299 ) | ( n37298 & n37299 ) ;
  assign n37301 = ( n37293 & ~n37297 ) | ( n37293 & n37300 ) | ( ~n37297 & n37300 ) ;
  assign n37302 = ~n37284 & n37301 ;
  assign n37303 = n37284 & ~n37301 ;
  assign n37304 = n37302 | n37303 ;
  assign n37307 = ~n37304 & n37306 ;
  assign n37308 = n37306 & ~n37307 ;
  assign n37309 = n37304 | n37306 ;
  assign n37310 = x125 & n12574 ;
  assign n37311 = x124 & n12569 ;
  assign n37312 = x123 & ~n12568 ;
  assign n37313 = n13076 & n37312 ;
  assign n37314 = n37311 | n37313 ;
  assign n37315 = n37310 | n37314 ;
  assign n37316 = n12577 | n37310 ;
  assign n37317 = n37314 | n37316 ;
  assign n37318 = ( n17670 & n37315 ) | ( n17670 & n37317 ) | ( n37315 & n37317 ) ;
  assign n37319 = x53 & n37317 ;
  assign n37320 = x53 & n37310 ;
  assign n37321 = ( x53 & n37314 ) | ( x53 & n37320 ) | ( n37314 & n37320 ) ;
  assign n37322 = ( n17670 & n37319 ) | ( n17670 & n37321 ) | ( n37319 & n37321 ) ;
  assign n37323 = x53 & ~n37321 ;
  assign n37324 = x53 & ~n37317 ;
  assign n37325 = ( ~n17670 & n37323 ) | ( ~n17670 & n37324 ) | ( n37323 & n37324 ) ;
  assign n37326 = ( n37318 & ~n37322 ) | ( n37318 & n37325 ) | ( ~n37322 & n37325 ) ;
  assign n37327 = n37309 & ~n37326 ;
  assign n37328 = ~n37308 & n37327 ;
  assign n37329 = ( ~n37304 & n37306 ) | ( ~n37304 & n37326 ) | ( n37306 & n37326 ) ;
  assign n37330 = ~n37307 & n37329 ;
  assign n37331 = n37328 | n37330 ;
  assign n37332 = n37175 | n37178 ;
  assign n37333 = ( n37175 & ~n37176 ) | ( n37175 & n37332 ) | ( ~n37176 & n37332 ) ;
  assign n37334 = ~n37331 & n37333 ;
  assign n37335 = n37331 & ~n37333 ;
  assign n37336 = n37334 | n37335 ;
  assign n37337 = x127 & n11200 ;
  assign n37338 = x126 & ~n11199 ;
  assign n37339 = n11679 & n37338 ;
  assign n37340 = n37337 | n37339 ;
  assign n37341 = n11208 | n37340 ;
  assign n37342 = ( n19328 & n37340 ) | ( n19328 & n37341 ) | ( n37340 & n37341 ) ;
  assign n37343 = x50 & n37340 ;
  assign n37344 = ( x50 & n14541 ) | ( x50 & n37340 ) | ( n14541 & n37340 ) ;
  assign n37345 = ( n19328 & n37343 ) | ( n19328 & n37344 ) | ( n37343 & n37344 ) ;
  assign n37346 = x50 & ~n14541 ;
  assign n37347 = ~n37340 & n37346 ;
  assign n37348 = x50 & ~n37340 ;
  assign n37349 = ( ~n19328 & n37347 ) | ( ~n19328 & n37348 ) | ( n37347 & n37348 ) ;
  assign n37350 = ( n37342 & ~n37345 ) | ( n37342 & n37349 ) | ( ~n37345 & n37349 ) ;
  assign n37351 = n37336 | n37350 ;
  assign n37352 = n37336 & ~n37350 ;
  assign n37353 = ( ~n37336 & n37351 ) | ( ~n37336 & n37352 ) | ( n37351 & n37352 ) ;
  assign n37354 = n37200 & ~n37201 ;
  assign n37355 = n37199 | n37204 ;
  assign n37356 = ( n37199 & ~n37354 ) | ( n37199 & n37355 ) | ( ~n37354 & n37355 ) ;
  assign n37357 = n37353 & ~n37356 ;
  assign n37358 = ~n37353 & n37356 ;
  assign n37359 = n37357 | n37358 ;
  assign n37360 = ~n37213 & n37221 ;
  assign n37361 = n37213 | n37220 ;
  assign n37362 = ( n37059 & ~n37360 ) | ( n37059 & n37361 ) | ( ~n37360 & n37361 ) ;
  assign n37363 = ~n37213 & n37214 ;
  assign n37364 = ( n37064 & ~n37361 ) | ( n37064 & n37363 ) | ( ~n37361 & n37363 ) ;
  assign n37365 = ( n36715 & ~n37362 ) | ( n36715 & n37364 ) | ( ~n37362 & n37364 ) ;
  assign n37366 = n37359 & n37365 ;
  assign n37367 = ~n37359 & n37362 ;
  assign n37368 = n37213 & ~n37359 ;
  assign n37369 = ( n37220 & ~n37359 ) | ( n37220 & n37368 ) | ( ~n37359 & n37368 ) ;
  assign n37370 = ( n37214 & n37359 ) | ( n37214 & ~n37368 ) | ( n37359 & ~n37368 ) ;
  assign n37371 = ( n37064 & ~n37369 ) | ( n37064 & n37370 ) | ( ~n37369 & n37370 ) ;
  assign n37372 = ( n36715 & ~n37367 ) | ( n36715 & n37371 ) | ( ~n37367 & n37371 ) ;
  assign n37373 = ~n37366 & n37372 ;
  assign n37374 = x127 & ~n11199 ;
  assign n37375 = n11679 & n37374 ;
  assign n37376 = n11208 | n37375 ;
  assign n37377 = n19877 | n37375 ;
  assign n37378 = n37376 & n37377 ;
  assign n37379 = n19880 | n37375 ;
  assign n37380 = n37376 & n37379 ;
  assign n37381 = ( n18202 & n37378 ) | ( n18202 & n37380 ) | ( n37378 & n37380 ) ;
  assign n37382 = n37378 & n37380 ;
  assign n37383 = ( n18212 & n37381 ) | ( n18212 & n37382 ) | ( n37381 & n37382 ) ;
  assign n37384 = ( n18214 & n37381 ) | ( n18214 & n37382 ) | ( n37381 & n37382 ) ;
  assign n37385 = ( n14002 & n37383 ) | ( n14002 & n37384 ) | ( n37383 & n37384 ) ;
  assign n37386 = x50 & n37383 ;
  assign n37387 = x50 & n37384 ;
  assign n37388 = ( n14002 & n37386 ) | ( n14002 & n37387 ) | ( n37386 & n37387 ) ;
  assign n37389 = x50 & ~n37387 ;
  assign n37390 = x50 & ~n37386 ;
  assign n37391 = ( ~n14002 & n37389 ) | ( ~n14002 & n37390 ) | ( n37389 & n37390 ) ;
  assign n37392 = ( n37385 & ~n37388 ) | ( n37385 & n37391 ) | ( ~n37388 & n37391 ) ;
  assign n37393 = n37307 & n37392 ;
  assign n37394 = ( n37330 & n37392 ) | ( n37330 & n37393 ) | ( n37392 & n37393 ) ;
  assign n37395 = n37307 | n37392 ;
  assign n37396 = n37330 | n37395 ;
  assign n37397 = ~n37394 & n37396 ;
  assign n37398 = x117 & n17146 ;
  assign n37399 = x116 & n17141 ;
  assign n37400 = x115 & ~n17140 ;
  assign n37401 = n17724 & n37400 ;
  assign n37402 = n37399 | n37401 ;
  assign n37403 = n37398 | n37402 ;
  assign n37404 = n17149 | n37398 ;
  assign n37405 = n37402 | n37404 ;
  assign n37406 = ( ~n13522 & n37403 ) | ( ~n13522 & n37405 ) | ( n37403 & n37405 ) ;
  assign n37407 = n37403 & n37405 ;
  assign n37408 = ( n13503 & n37406 ) | ( n13503 & n37407 ) | ( n37406 & n37407 ) ;
  assign n37409 = ~x62 & n37408 ;
  assign n37410 = x62 & n37405 ;
  assign n37411 = x62 & x117 ;
  assign n37412 = n17146 & n37411 ;
  assign n37413 = ( x62 & n37402 ) | ( x62 & n37412 ) | ( n37402 & n37412 ) ;
  assign n37414 = ( ~n13522 & n37410 ) | ( ~n13522 & n37413 ) | ( n37410 & n37413 ) ;
  assign n37415 = n37410 & n37413 ;
  assign n37416 = ( n13503 & n37414 ) | ( n13503 & n37415 ) | ( n37414 & n37415 ) ;
  assign n37417 = x62 & ~n37416 ;
  assign n37418 = n37409 | n37417 ;
  assign n37419 = x114 & n18290 ;
  assign n37420 = x63 & x113 ;
  assign n37421 = ~n18290 & n37420 ;
  assign n37422 = n37419 | n37421 ;
  assign n37423 = ~n37229 & n37422 ;
  assign n37424 = n37229 | n37423 ;
  assign n37425 = n37422 & ~n37423 ;
  assign n37426 = n37424 & ~n37425 ;
  assign n37427 = n37418 & ~n37426 ;
  assign n37428 = ~n37418 & n37426 ;
  assign n37429 = n37427 | n37428 ;
  assign n37430 = ~n37231 & n37233 ;
  assign n37431 = ( n37231 & n37248 ) | ( n37231 & ~n37430 ) | ( n37248 & ~n37430 ) ;
  assign n37432 = n37429 & ~n37431 ;
  assign n37433 = ~n37429 & n37431 ;
  assign n37434 = n37432 | n37433 ;
  assign n37435 = x120 & n15552 ;
  assign n37436 = x119 & n15547 ;
  assign n37437 = x118 & ~n15546 ;
  assign n37438 = n16123 & n37437 ;
  assign n37439 = n37436 | n37438 ;
  assign n37440 = n37435 | n37439 ;
  assign n37441 = n15555 | n37435 ;
  assign n37442 = n37439 | n37441 ;
  assign n37443 = ( n14991 & n37440 ) | ( n14991 & n37442 ) | ( n37440 & n37442 ) ;
  assign n37444 = x59 & n37442 ;
  assign n37445 = x59 & n37435 ;
  assign n37446 = ( x59 & n37439 ) | ( x59 & n37445 ) | ( n37439 & n37445 ) ;
  assign n37447 = ( n14991 & n37444 ) | ( n14991 & n37446 ) | ( n37444 & n37446 ) ;
  assign n37448 = x59 & ~n37446 ;
  assign n37449 = x59 & ~n37442 ;
  assign n37450 = ( ~n14991 & n37448 ) | ( ~n14991 & n37449 ) | ( n37448 & n37449 ) ;
  assign n37451 = ( n37443 & ~n37447 ) | ( n37443 & n37450 ) | ( ~n37447 & n37450 ) ;
  assign n37452 = n37434 & ~n37451 ;
  assign n37453 = ~n37434 & n37451 ;
  assign n37454 = n37452 | n37453 ;
  assign n37455 = n37254 | n37277 ;
  assign n37456 = ( n37253 & n37272 ) | ( n37253 & ~n37273 ) | ( n37272 & ~n37273 ) ;
  assign n37457 = ( n37255 & n37455 ) | ( n37255 & n37456 ) | ( n37455 & n37456 ) ;
  assign n37458 = ~n37454 & n37457 ;
  assign n37459 = n37454 & ~n37457 ;
  assign n37460 = n37458 | n37459 ;
  assign n37461 = x123 & n14045 ;
  assign n37462 = x122 & n14040 ;
  assign n37463 = x121 & ~n14039 ;
  assign n37464 = n14552 & n37463 ;
  assign n37465 = n37462 | n37464 ;
  assign n37466 = n37461 | n37465 ;
  assign n37467 = n14048 | n37461 ;
  assign n37468 = n37465 | n37467 ;
  assign n37469 = ( n16086 & n37466 ) | ( n16086 & n37468 ) | ( n37466 & n37468 ) ;
  assign n37470 = x56 & n37468 ;
  assign n37471 = x56 & n37461 ;
  assign n37472 = ( x56 & n37465 ) | ( x56 & n37471 ) | ( n37465 & n37471 ) ;
  assign n37473 = ( n16086 & n37470 ) | ( n16086 & n37472 ) | ( n37470 & n37472 ) ;
  assign n37474 = x56 & ~n37472 ;
  assign n37475 = x56 & ~n37468 ;
  assign n37476 = ( ~n16086 & n37474 ) | ( ~n16086 & n37475 ) | ( n37474 & n37475 ) ;
  assign n37477 = ( n37469 & ~n37473 ) | ( n37469 & n37476 ) | ( ~n37473 & n37476 ) ;
  assign n37478 = ~n37460 & n37477 ;
  assign n37479 = n37460 | n37478 ;
  assign n37481 = n37281 | n37301 ;
  assign n37482 = ( ~n37279 & n37301 ) | ( ~n37279 & n37481 ) | ( n37301 & n37481 ) ;
  assign n37483 = ( n37282 & ~n37284 ) | ( n37282 & n37482 ) | ( ~n37284 & n37482 ) ;
  assign n37480 = n37460 & n37477 ;
  assign n37484 = n37480 & n37483 ;
  assign n37485 = ( ~n37479 & n37483 ) | ( ~n37479 & n37484 ) | ( n37483 & n37484 ) ;
  assign n37486 = n37480 | n37483 ;
  assign n37487 = n37479 & ~n37486 ;
  assign n37488 = n37485 | n37487 ;
  assign n37489 = x126 & n12574 ;
  assign n37490 = x125 & n12569 ;
  assign n37491 = x124 & ~n12568 ;
  assign n37492 = n13076 & n37491 ;
  assign n37493 = n37490 | n37492 ;
  assign n37494 = n37489 | n37493 ;
  assign n37495 = n12577 | n37489 ;
  assign n37496 = n37493 | n37495 ;
  assign n37497 = ( n18220 & n37494 ) | ( n18220 & n37496 ) | ( n37494 & n37496 ) ;
  assign n37498 = x53 & n37496 ;
  assign n37499 = x53 & n37489 ;
  assign n37500 = ( x53 & n37493 ) | ( x53 & n37499 ) | ( n37493 & n37499 ) ;
  assign n37501 = ( n18220 & n37498 ) | ( n18220 & n37500 ) | ( n37498 & n37500 ) ;
  assign n37502 = x53 & ~n37500 ;
  assign n37503 = x53 & ~n37496 ;
  assign n37504 = ( ~n18220 & n37502 ) | ( ~n18220 & n37503 ) | ( n37502 & n37503 ) ;
  assign n37505 = ( n37497 & ~n37501 ) | ( n37497 & n37504 ) | ( ~n37501 & n37504 ) ;
  assign n37506 = n37488 | n37505 ;
  assign n37507 = n37488 & ~n37505 ;
  assign n37508 = ( ~n37488 & n37506 ) | ( ~n37488 & n37507 ) | ( n37506 & n37507 ) ;
  assign n37509 = n37397 & ~n37508 ;
  assign n37510 = n37508 | n37509 ;
  assign n37511 = ( ~n37397 & n37509 ) | ( ~n37397 & n37510 ) | ( n37509 & n37510 ) ;
  assign n37512 = n37334 | n37350 ;
  assign n37513 = ( n37334 & ~n37336 ) | ( n37334 & n37512 ) | ( ~n37336 & n37512 ) ;
  assign n37514 = n37511 & ~n37513 ;
  assign n37515 = ~n37511 & n37513 ;
  assign n37516 = n37514 | n37515 ;
  assign n37517 = ~n37358 & n37371 ;
  assign n37518 = ~n37358 & n37359 ;
  assign n37519 = ( n37358 & n37362 ) | ( n37358 & ~n37518 ) | ( n37362 & ~n37518 ) ;
  assign n37520 = ( n36715 & n37517 ) | ( n36715 & ~n37519 ) | ( n37517 & ~n37519 ) ;
  assign n37521 = n37516 & n37520 ;
  assign n37522 = n37358 & ~n37516 ;
  assign n37523 = ( n37359 & n37516 ) | ( n37359 & ~n37522 ) | ( n37516 & ~n37522 ) ;
  assign n37524 = ( n37362 & n37522 ) | ( n37362 & ~n37523 ) | ( n37522 & ~n37523 ) ;
  assign n37525 = ( n37371 & n37516 ) | ( n37371 & ~n37522 ) | ( n37516 & ~n37522 ) ;
  assign n37526 = ( n36715 & ~n37524 ) | ( n36715 & n37525 ) | ( ~n37524 & n37525 ) ;
  assign n37527 = ~n37521 & n37526 ;
  assign n37528 = ~n37423 & n37426 ;
  assign n37529 = ( n37418 & n37423 ) | ( n37418 & ~n37528 ) | ( n37423 & ~n37528 ) ;
  assign n37530 = x115 & n18290 ;
  assign n37531 = x63 & x114 ;
  assign n37532 = ~n18290 & n37531 ;
  assign n37533 = n37530 | n37532 ;
  assign n37534 = ~x50 & n37533 ;
  assign n37535 = x50 & ~n37533 ;
  assign n37536 = n37534 | n37535 ;
  assign n37537 = n37229 & ~n37536 ;
  assign n37538 = ~n37229 & n37536 ;
  assign n37539 = n37537 | n37538 ;
  assign n37540 = n37423 & ~n37539 ;
  assign n37541 = ( n37426 & n37539 ) | ( n37426 & ~n37540 ) | ( n37539 & ~n37540 ) ;
  assign n37542 = ~n37539 & n37540 ;
  assign n37543 = ( n37418 & ~n37541 ) | ( n37418 & n37542 ) | ( ~n37541 & n37542 ) ;
  assign n37544 = n37529 & ~n37543 ;
  assign n37545 = x118 & n17146 ;
  assign n37546 = x117 & n17141 ;
  assign n37547 = x116 & ~n17140 ;
  assign n37548 = n17724 & n37547 ;
  assign n37549 = n37546 | n37548 ;
  assign n37550 = n37545 | n37549 ;
  assign n37551 = n17149 | n37545 ;
  assign n37552 = n37549 | n37551 ;
  assign n37553 = ( ~n14002 & n37550 ) | ( ~n14002 & n37552 ) | ( n37550 & n37552 ) ;
  assign n37554 = n37550 & n37552 ;
  assign n37555 = ( n13981 & n37553 ) | ( n13981 & n37554 ) | ( n37553 & n37554 ) ;
  assign n37556 = x62 & n37555 ;
  assign n37557 = x62 & ~n37555 ;
  assign n37558 = ( n37555 & ~n37556 ) | ( n37555 & n37557 ) | ( ~n37556 & n37557 ) ;
  assign n37559 = n37539 | n37540 ;
  assign n37560 = n37426 & ~n37539 ;
  assign n37561 = ~n37540 & n37560 ;
  assign n37562 = ( n37418 & n37559 ) | ( n37418 & ~n37561 ) | ( n37559 & ~n37561 ) ;
  assign n37563 = ~n37558 & n37562 ;
  assign n37564 = ~n37544 & n37563 ;
  assign n37565 = n37558 & ~n37562 ;
  assign n37566 = ( n37544 & n37558 ) | ( n37544 & n37565 ) | ( n37558 & n37565 ) ;
  assign n37567 = n37564 | n37566 ;
  assign n37568 = x121 & n15552 ;
  assign n37569 = x120 & n15547 ;
  assign n37570 = x119 & ~n15546 ;
  assign n37571 = n16123 & n37570 ;
  assign n37572 = n37569 | n37571 ;
  assign n37573 = n37568 | n37572 ;
  assign n37574 = n15555 | n37568 ;
  assign n37575 = n37572 | n37574 ;
  assign n37576 = ( n15501 & n37573 ) | ( n15501 & n37575 ) | ( n37573 & n37575 ) ;
  assign n37577 = x59 & n37575 ;
  assign n37578 = x59 & n37568 ;
  assign n37579 = ( x59 & n37572 ) | ( x59 & n37578 ) | ( n37572 & n37578 ) ;
  assign n37580 = ( n15501 & n37577 ) | ( n15501 & n37579 ) | ( n37577 & n37579 ) ;
  assign n37581 = x59 & ~n37579 ;
  assign n37582 = x59 & ~n37575 ;
  assign n37583 = ( ~n15501 & n37581 ) | ( ~n15501 & n37582 ) | ( n37581 & n37582 ) ;
  assign n37584 = ( n37576 & ~n37580 ) | ( n37576 & n37583 ) | ( ~n37580 & n37583 ) ;
  assign n37585 = ~n37567 & n37584 ;
  assign n37586 = n37567 | n37585 ;
  assign n37588 = n37431 | n37451 ;
  assign n37589 = ( ~n37429 & n37451 ) | ( ~n37429 & n37588 ) | ( n37451 & n37588 ) ;
  assign n37590 = ( n37433 & ~n37434 ) | ( n37433 & n37589 ) | ( ~n37434 & n37589 ) ;
  assign n37587 = n37567 & n37584 ;
  assign n37591 = n37587 & n37590 ;
  assign n37592 = ( ~n37586 & n37590 ) | ( ~n37586 & n37591 ) | ( n37590 & n37591 ) ;
  assign n37593 = n37587 | n37590 ;
  assign n37594 = n37586 & ~n37593 ;
  assign n37595 = n37592 | n37594 ;
  assign n37596 = x124 & n14045 ;
  assign n37597 = x123 & n14040 ;
  assign n37598 = x122 & ~n14039 ;
  assign n37599 = n14552 & n37598 ;
  assign n37600 = n37597 | n37599 ;
  assign n37601 = n37596 | n37600 ;
  assign n37602 = n14048 | n37596 ;
  assign n37603 = n37600 | n37602 ;
  assign n37604 = ( n17084 & n37601 ) | ( n17084 & n37603 ) | ( n37601 & n37603 ) ;
  assign n37605 = x56 & n37603 ;
  assign n37606 = x56 & n37596 ;
  assign n37607 = ( x56 & n37600 ) | ( x56 & n37606 ) | ( n37600 & n37606 ) ;
  assign n37608 = ( n17084 & n37605 ) | ( n17084 & n37607 ) | ( n37605 & n37607 ) ;
  assign n37609 = x56 & ~n37607 ;
  assign n37610 = x56 & ~n37603 ;
  assign n37611 = ( ~n17084 & n37609 ) | ( ~n17084 & n37610 ) | ( n37609 & n37610 ) ;
  assign n37612 = ( n37604 & ~n37608 ) | ( n37604 & n37611 ) | ( ~n37608 & n37611 ) ;
  assign n37613 = ~n37595 & n37612 ;
  assign n37614 = n37595 & ~n37612 ;
  assign n37615 = n37613 | n37614 ;
  assign n37616 = n37458 | n37477 ;
  assign n37617 = ( n37458 & ~n37460 ) | ( n37458 & n37616 ) | ( ~n37460 & n37616 ) ;
  assign n37618 = ~n37615 & n37617 ;
  assign n37619 = n37615 & ~n37617 ;
  assign n37620 = n37618 | n37619 ;
  assign n37621 = x127 & n12574 ;
  assign n37622 = x126 & n12569 ;
  assign n37623 = x125 & ~n12568 ;
  assign n37624 = n13076 & n37623 ;
  assign n37625 = n37622 | n37624 ;
  assign n37626 = n37621 | n37625 ;
  assign n37627 = n12577 | n37621 ;
  assign n37628 = n37625 | n37627 ;
  assign n37629 = ( n18763 & n37626 ) | ( n18763 & n37628 ) | ( n37626 & n37628 ) ;
  assign n37630 = x53 & n37628 ;
  assign n37631 = x53 & n37621 ;
  assign n37632 = ( x53 & n37625 ) | ( x53 & n37631 ) | ( n37625 & n37631 ) ;
  assign n37633 = ( n18763 & n37630 ) | ( n18763 & n37632 ) | ( n37630 & n37632 ) ;
  assign n37634 = x53 & ~n37632 ;
  assign n37635 = x53 & ~n37628 ;
  assign n37636 = ( ~n18763 & n37634 ) | ( ~n18763 & n37635 ) | ( n37634 & n37635 ) ;
  assign n37637 = ( n37629 & ~n37633 ) | ( n37629 & n37636 ) | ( ~n37633 & n37636 ) ;
  assign n37638 = ~n37620 & n37637 ;
  assign n37639 = n37620 | n37638 ;
  assign n37640 = n37620 & n37637 ;
  assign n37641 = n37639 & ~n37640 ;
  assign n37642 = n37483 | n37505 ;
  assign n37643 = n37479 & ~n37505 ;
  assign n37644 = ( n37484 & n37642 ) | ( n37484 & ~n37643 ) | ( n37642 & ~n37643 ) ;
  assign n37645 = ( n37485 & ~n37488 ) | ( n37485 & n37644 ) | ( ~n37488 & n37644 ) ;
  assign n37646 = n37641 & ~n37645 ;
  assign n37647 = ~n37641 & n37645 ;
  assign n37648 = n37646 | n37647 ;
  assign n37649 = n37394 | n37509 ;
  assign n37650 = n37648 & ~n37649 ;
  assign n37651 = ~n37648 & n37649 ;
  assign n37652 = n37650 | n37651 ;
  assign n37653 = ~n37515 & n37523 ;
  assign n37654 = ~n37515 & n37516 ;
  assign n37655 = ( n37358 & n37515 ) | ( n37358 & ~n37654 ) | ( n37515 & ~n37654 ) ;
  assign n37656 = ( n37362 & ~n37653 ) | ( n37362 & n37655 ) | ( ~n37653 & n37655 ) ;
  assign n37657 = ( n37371 & n37654 ) | ( n37371 & ~n37655 ) | ( n37654 & ~n37655 ) ;
  assign n37658 = ( n36715 & ~n37656 ) | ( n36715 & n37657 ) | ( ~n37656 & n37657 ) ;
  assign n37659 = n37652 & n37658 ;
  assign n37660 = ~n37652 & n37655 ;
  assign n37661 = n37515 & ~n37652 ;
  assign n37662 = ( n37523 & n37652 ) | ( n37523 & ~n37661 ) | ( n37652 & ~n37661 ) ;
  assign n37663 = ( n37362 & n37660 ) | ( n37362 & ~n37662 ) | ( n37660 & ~n37662 ) ;
  assign n37664 = ( n37516 & n37652 ) | ( n37516 & ~n37661 ) | ( n37652 & ~n37661 ) ;
  assign n37665 = ( n37371 & ~n37660 ) | ( n37371 & n37664 ) | ( ~n37660 & n37664 ) ;
  assign n37666 = ( n36715 & ~n37663 ) | ( n36715 & n37665 ) | ( ~n37663 & n37665 ) ;
  assign n37667 = ~n37659 & n37666 ;
  assign n37668 = n37585 | n37592 ;
  assign n37669 = x116 & n18290 ;
  assign n37670 = x63 & x115 ;
  assign n37671 = ~n18290 & n37670 ;
  assign n37672 = n37669 | n37671 ;
  assign n37673 = n37229 | n37534 ;
  assign n37674 = ( n37534 & ~n37536 ) | ( n37534 & n37673 ) | ( ~n37536 & n37673 ) ;
  assign n37675 = n37672 & ~n37674 ;
  assign n37676 = ~n37672 & n37674 ;
  assign n37677 = n37675 | n37676 ;
  assign n37678 = x118 & n17141 ;
  assign n37679 = x117 & ~n17140 ;
  assign n37680 = n17724 & n37679 ;
  assign n37681 = n37678 | n37680 ;
  assign n37682 = x119 & n17146 ;
  assign n37683 = n17149 | n37682 ;
  assign n37684 = n37681 | n37683 ;
  assign n37685 = x62 & ~n37684 ;
  assign n37686 = ~n37677 & n37685 ;
  assign n37687 = x62 & x119 ;
  assign n37688 = n17146 & n37687 ;
  assign n37689 = x62 & ~n37688 ;
  assign n37690 = ~n37681 & n37689 ;
  assign n37691 = ~n37677 & n37690 ;
  assign n37692 = ( ~n14496 & n37686 ) | ( ~n14496 & n37691 ) | ( n37686 & n37691 ) ;
  assign n37693 = ~x62 & n37684 ;
  assign n37694 = ~x62 & n37682 ;
  assign n37695 = ( ~x62 & n37681 ) | ( ~x62 & n37694 ) | ( n37681 & n37694 ) ;
  assign n37696 = ( n14496 & n37693 ) | ( n14496 & n37695 ) | ( n37693 & n37695 ) ;
  assign n37697 = ( ~n37677 & n37692 ) | ( ~n37677 & n37696 ) | ( n37692 & n37696 ) ;
  assign n37698 = n37677 & ~n37685 ;
  assign n37699 = n37677 & ~n37690 ;
  assign n37700 = ( n14496 & n37698 ) | ( n14496 & n37699 ) | ( n37698 & n37699 ) ;
  assign n37701 = ~n37696 & n37700 ;
  assign n37702 = n37697 | n37701 ;
  assign n37703 = n37543 & ~n37702 ;
  assign n37704 = ( n37566 & ~n37702 ) | ( n37566 & n37703 ) | ( ~n37702 & n37703 ) ;
  assign n37705 = ~n37543 & n37702 ;
  assign n37706 = ~n37566 & n37705 ;
  assign n37707 = n37704 | n37706 ;
  assign n37708 = x122 & n15552 ;
  assign n37709 = x121 & n15547 ;
  assign n37710 = x120 & ~n15546 ;
  assign n37711 = n16123 & n37710 ;
  assign n37712 = n37709 | n37711 ;
  assign n37713 = n37708 | n37712 ;
  assign n37714 = n15555 | n37708 ;
  assign n37715 = n37712 | n37714 ;
  assign n37716 = ( n16043 & n37713 ) | ( n16043 & n37715 ) | ( n37713 & n37715 ) ;
  assign n37717 = x59 & n37715 ;
  assign n37718 = x59 & n37708 ;
  assign n37719 = ( x59 & n37712 ) | ( x59 & n37718 ) | ( n37712 & n37718 ) ;
  assign n37720 = ( n16043 & n37717 ) | ( n16043 & n37719 ) | ( n37717 & n37719 ) ;
  assign n37721 = x59 & ~n37719 ;
  assign n37722 = x59 & ~n37715 ;
  assign n37723 = ( ~n16043 & n37721 ) | ( ~n16043 & n37722 ) | ( n37721 & n37722 ) ;
  assign n37724 = ( n37716 & ~n37720 ) | ( n37716 & n37723 ) | ( ~n37720 & n37723 ) ;
  assign n37725 = ~n37707 & n37724 ;
  assign n37726 = n37707 & ~n37724 ;
  assign n37727 = n37725 | n37726 ;
  assign n37728 = n37668 & ~n37727 ;
  assign n37729 = n37668 & ~n37728 ;
  assign n37730 = x125 & n14045 ;
  assign n37731 = x124 & n14040 ;
  assign n37732 = x123 & ~n14039 ;
  assign n37733 = n14552 & n37732 ;
  assign n37734 = n37731 | n37733 ;
  assign n37735 = n37730 | n37734 ;
  assign n37736 = n14048 | n37730 ;
  assign n37737 = n37734 | n37736 ;
  assign n37738 = ( n17670 & n37735 ) | ( n17670 & n37737 ) | ( n37735 & n37737 ) ;
  assign n37739 = x56 & n37737 ;
  assign n37740 = x56 & n37730 ;
  assign n37741 = ( x56 & n37734 ) | ( x56 & n37740 ) | ( n37734 & n37740 ) ;
  assign n37742 = ( n17670 & n37739 ) | ( n17670 & n37741 ) | ( n37739 & n37741 ) ;
  assign n37743 = x56 & ~n37741 ;
  assign n37744 = x56 & ~n37737 ;
  assign n37745 = ( ~n17670 & n37743 ) | ( ~n17670 & n37744 ) | ( n37743 & n37744 ) ;
  assign n37746 = ( n37738 & ~n37742 ) | ( n37738 & n37745 ) | ( ~n37742 & n37745 ) ;
  assign n37747 = n37727 & ~n37746 ;
  assign n37748 = ( n37668 & ~n37746 ) | ( n37668 & n37747 ) | ( ~n37746 & n37747 ) ;
  assign n37749 = ~n37729 & n37748 ;
  assign n37750 = ( n37668 & ~n37727 ) | ( n37668 & n37746 ) | ( ~n37727 & n37746 ) ;
  assign n37751 = ~n37728 & n37750 ;
  assign n37752 = n37749 | n37751 ;
  assign n37753 = n37613 | n37617 ;
  assign n37754 = ( n37613 & ~n37615 ) | ( n37613 & n37753 ) | ( ~n37615 & n37753 ) ;
  assign n37755 = ~n37752 & n37754 ;
  assign n37756 = n37752 & ~n37754 ;
  assign n37757 = n37755 | n37756 ;
  assign n37758 = x127 & n12569 ;
  assign n37759 = x126 & ~n12568 ;
  assign n37760 = n13076 & n37759 ;
  assign n37761 = n37758 | n37760 ;
  assign n37762 = n12577 | n37761 ;
  assign n37763 = ( n19328 & n37761 ) | ( n19328 & n37762 ) | ( n37761 & n37762 ) ;
  assign n37764 = x53 & n37761 ;
  assign n37765 = ( x53 & n16112 ) | ( x53 & n37761 ) | ( n16112 & n37761 ) ;
  assign n37766 = ( n19328 & n37764 ) | ( n19328 & n37765 ) | ( n37764 & n37765 ) ;
  assign n37767 = x53 & ~n16112 ;
  assign n37768 = ~n37761 & n37767 ;
  assign n37769 = x53 & ~n37761 ;
  assign n37770 = ( ~n19328 & n37768 ) | ( ~n19328 & n37769 ) | ( n37768 & n37769 ) ;
  assign n37771 = ( n37763 & ~n37766 ) | ( n37763 & n37770 ) | ( ~n37766 & n37770 ) ;
  assign n37772 = n37757 | n37771 ;
  assign n37773 = n37757 & ~n37771 ;
  assign n37774 = ( ~n37757 & n37772 ) | ( ~n37757 & n37773 ) | ( n37772 & n37773 ) ;
  assign n37775 = n37638 | n37645 ;
  assign n37776 = ( n37638 & ~n37641 ) | ( n37638 & n37775 ) | ( ~n37641 & n37775 ) ;
  assign n37777 = n37774 & ~n37776 ;
  assign n37778 = ~n37774 & n37776 ;
  assign n37779 = n37777 | n37778 ;
  assign n37780 = n37651 | n37661 ;
  assign n37781 = ~n37651 & n37652 ;
  assign n37782 = ( n37523 & ~n37780 ) | ( n37523 & n37781 ) | ( ~n37780 & n37781 ) ;
  assign n37783 = ( n37651 & n37655 ) | ( n37651 & ~n37781 ) | ( n37655 & ~n37781 ) ;
  assign n37784 = ( n37362 & ~n37782 ) | ( n37362 & n37783 ) | ( ~n37782 & n37783 ) ;
  assign n37785 = ~n37651 & n37664 ;
  assign n37786 = ( n37371 & ~n37783 ) | ( n37371 & n37785 ) | ( ~n37783 & n37785 ) ;
  assign n37787 = ( n36715 & ~n37784 ) | ( n36715 & n37786 ) | ( ~n37784 & n37786 ) ;
  assign n37788 = n37779 & n37787 ;
  assign n37789 = n37779 | n37781 ;
  assign n37790 = n37651 & ~n37779 ;
  assign n37791 = ( n37655 & ~n37789 ) | ( n37655 & n37790 ) | ( ~n37789 & n37790 ) ;
  assign n37792 = ( n37664 & n37779 ) | ( n37664 & ~n37790 ) | ( n37779 & ~n37790 ) ;
  assign n37793 = ( n37371 & ~n37791 ) | ( n37371 & n37792 ) | ( ~n37791 & n37792 ) ;
  assign n37794 = ~n37779 & n37780 ;
  assign n37795 = ( n37523 & n37789 ) | ( n37523 & ~n37794 ) | ( n37789 & ~n37794 ) ;
  assign n37796 = ( n37360 & ~n37791 ) | ( n37360 & n37795 ) | ( ~n37791 & n37795 ) ;
  assign n37797 = ( n37361 & n37791 ) | ( n37361 & ~n37795 ) | ( n37791 & ~n37795 ) ;
  assign n37798 = ( n37059 & ~n37796 ) | ( n37059 & n37797 ) | ( ~n37796 & n37797 ) ;
  assign n37799 = ( n36715 & n37793 ) | ( n36715 & ~n37798 ) | ( n37793 & ~n37798 ) ;
  assign n37800 = ~n37788 & n37799 ;
  assign n37801 = x127 & ~n12568 ;
  assign n37802 = n13076 & n37801 ;
  assign n37803 = n12577 | n37802 ;
  assign n37804 = n19877 | n37802 ;
  assign n37805 = n37803 & n37804 ;
  assign n37806 = n19880 | n37802 ;
  assign n37807 = n37803 & n37806 ;
  assign n37808 = ( n18202 & n37805 ) | ( n18202 & n37807 ) | ( n37805 & n37807 ) ;
  assign n37809 = n37805 & n37807 ;
  assign n37810 = ( n18212 & n37808 ) | ( n18212 & n37809 ) | ( n37808 & n37809 ) ;
  assign n37811 = ( n18214 & n37808 ) | ( n18214 & n37809 ) | ( n37808 & n37809 ) ;
  assign n37812 = ( n14002 & n37810 ) | ( n14002 & n37811 ) | ( n37810 & n37811 ) ;
  assign n37813 = x53 & n37810 ;
  assign n37814 = x53 & n37811 ;
  assign n37815 = ( n14002 & n37813 ) | ( n14002 & n37814 ) | ( n37813 & n37814 ) ;
  assign n37816 = x53 & ~n37814 ;
  assign n37817 = x53 & ~n37813 ;
  assign n37818 = ( ~n14002 & n37816 ) | ( ~n14002 & n37817 ) | ( n37816 & n37817 ) ;
  assign n37819 = ( n37812 & ~n37815 ) | ( n37812 & n37818 ) | ( ~n37815 & n37818 ) ;
  assign n37820 = ~n37727 & n37819 ;
  assign n37821 = n37668 & n37820 ;
  assign n37822 = ( n37751 & n37819 ) | ( n37751 & n37821 ) | ( n37819 & n37821 ) ;
  assign n37823 = n37727 & ~n37819 ;
  assign n37824 = ( n37668 & n37819 ) | ( n37668 & ~n37823 ) | ( n37819 & ~n37823 ) ;
  assign n37825 = n37751 | n37824 ;
  assign n37826 = ~n37822 & n37825 ;
  assign n37827 = n37676 | n37697 ;
  assign n37828 = x117 & n18290 ;
  assign n37829 = x63 & x116 ;
  assign n37830 = ~n18290 & n37829 ;
  assign n37831 = n37828 | n37830 ;
  assign n37832 = ~n37672 & n37831 ;
  assign n37833 = n37672 & ~n37831 ;
  assign n37834 = n37832 | n37833 ;
  assign n37835 = n37672 | n37834 ;
  assign n37836 = n37674 & ~n37835 ;
  assign n37837 = ( n37697 & ~n37834 ) | ( n37697 & n37836 ) | ( ~n37834 & n37836 ) ;
  assign n37838 = n37827 & ~n37837 ;
  assign n37839 = x120 & n17146 ;
  assign n37840 = x119 & n17141 ;
  assign n37841 = x118 & ~n17140 ;
  assign n37842 = n17724 & n37841 ;
  assign n37843 = n37840 | n37842 ;
  assign n37844 = n37839 | n37843 ;
  assign n37845 = n17149 | n37839 ;
  assign n37846 = n37843 | n37845 ;
  assign n37847 = ( n14991 & n37844 ) | ( n14991 & n37846 ) | ( n37844 & n37846 ) ;
  assign n37848 = x62 & n37846 ;
  assign n37849 = x62 & n37839 ;
  assign n37850 = ( x62 & n37843 ) | ( x62 & n37849 ) | ( n37843 & n37849 ) ;
  assign n37851 = ( n14991 & n37848 ) | ( n14991 & n37850 ) | ( n37848 & n37850 ) ;
  assign n37852 = x62 & ~n37850 ;
  assign n37853 = x62 & ~n37846 ;
  assign n37854 = ( ~n14991 & n37852 ) | ( ~n14991 & n37853 ) | ( n37852 & n37853 ) ;
  assign n37855 = ( n37847 & ~n37851 ) | ( n37847 & n37854 ) | ( ~n37851 & n37854 ) ;
  assign n37856 = n37834 | n37836 ;
  assign n37857 = n37697 | n37856 ;
  assign n37858 = n37855 | n37857 ;
  assign n37859 = ( ~n37838 & n37855 ) | ( ~n37838 & n37858 ) | ( n37855 & n37858 ) ;
  assign n37860 = n37855 & n37857 ;
  assign n37861 = ~n37838 & n37860 ;
  assign n37862 = n37859 & ~n37861 ;
  assign n37863 = x123 & n15552 ;
  assign n37864 = x122 & n15547 ;
  assign n37865 = x121 & ~n15546 ;
  assign n37866 = n16123 & n37865 ;
  assign n37867 = n37864 | n37866 ;
  assign n37868 = n37863 | n37867 ;
  assign n37869 = n15555 | n37863 ;
  assign n37870 = n37867 | n37869 ;
  assign n37871 = ( n16086 & n37868 ) | ( n16086 & n37870 ) | ( n37868 & n37870 ) ;
  assign n37872 = x59 & n37870 ;
  assign n37873 = x59 & n37863 ;
  assign n37874 = ( x59 & n37867 ) | ( x59 & n37873 ) | ( n37867 & n37873 ) ;
  assign n37875 = ( n16086 & n37872 ) | ( n16086 & n37874 ) | ( n37872 & n37874 ) ;
  assign n37876 = x59 & ~n37874 ;
  assign n37877 = x59 & ~n37870 ;
  assign n37878 = ( ~n16086 & n37876 ) | ( ~n16086 & n37877 ) | ( n37876 & n37877 ) ;
  assign n37879 = ( n37871 & ~n37875 ) | ( n37871 & n37878 ) | ( ~n37875 & n37878 ) ;
  assign n37880 = ~n37862 & n37879 ;
  assign n37881 = n37862 & ~n37879 ;
  assign n37882 = n37880 | n37881 ;
  assign n37883 = n37703 | n37724 ;
  assign n37884 = n37702 & ~n37724 ;
  assign n37885 = ( n37566 & n37883 ) | ( n37566 & ~n37884 ) | ( n37883 & ~n37884 ) ;
  assign n37886 = ( n37704 & ~n37707 ) | ( n37704 & n37885 ) | ( ~n37707 & n37885 ) ;
  assign n37887 = n37882 & ~n37886 ;
  assign n37888 = ~n37882 & n37886 ;
  assign n37889 = n37887 | n37888 ;
  assign n37890 = x126 & n14045 ;
  assign n37891 = x125 & n14040 ;
  assign n37892 = x124 & ~n14039 ;
  assign n37893 = n14552 & n37892 ;
  assign n37894 = n37891 | n37893 ;
  assign n37895 = n37890 | n37894 ;
  assign n37896 = n14048 | n37890 ;
  assign n37897 = n37894 | n37896 ;
  assign n37898 = ( n18220 & n37895 ) | ( n18220 & n37897 ) | ( n37895 & n37897 ) ;
  assign n37899 = x56 & n37897 ;
  assign n37900 = x56 & n37890 ;
  assign n37901 = ( x56 & n37894 ) | ( x56 & n37900 ) | ( n37894 & n37900 ) ;
  assign n37902 = ( n18220 & n37899 ) | ( n18220 & n37901 ) | ( n37899 & n37901 ) ;
  assign n37903 = x56 & ~n37901 ;
  assign n37904 = x56 & ~n37897 ;
  assign n37905 = ( ~n18220 & n37903 ) | ( ~n18220 & n37904 ) | ( n37903 & n37904 ) ;
  assign n37906 = ( n37898 & ~n37902 ) | ( n37898 & n37905 ) | ( ~n37902 & n37905 ) ;
  assign n37907 = n37889 & n37906 ;
  assign n37908 = n37888 | n37906 ;
  assign n37909 = n37887 | n37908 ;
  assign n37910 = ~n37907 & n37909 ;
  assign n37911 = n37826 & ~n37910 ;
  assign n37912 = n37826 | n37910 ;
  assign n37913 = ( ~n37826 & n37911 ) | ( ~n37826 & n37912 ) | ( n37911 & n37912 ) ;
  assign n37914 = n37754 | n37771 ;
  assign n37915 = ( ~n37752 & n37771 ) | ( ~n37752 & n37914 ) | ( n37771 & n37914 ) ;
  assign n37916 = ( n37755 & ~n37757 ) | ( n37755 & n37915 ) | ( ~n37757 & n37915 ) ;
  assign n37917 = n37913 & ~n37916 ;
  assign n37918 = ~n37913 & n37916 ;
  assign n37919 = n37917 | n37918 ;
  assign n37920 = n37778 | n37798 ;
  assign n37921 = ~n37778 & n37789 ;
  assign n37922 = n37778 | n37790 ;
  assign n37923 = ( n37655 & ~n37921 ) | ( n37655 & n37922 ) | ( ~n37921 & n37922 ) ;
  assign n37924 = ~n37778 & n37779 ;
  assign n37925 = ( n37664 & ~n37922 ) | ( n37664 & n37924 ) | ( ~n37922 & n37924 ) ;
  assign n37926 = ( n37369 & n37923 ) | ( n37369 & ~n37925 ) | ( n37923 & ~n37925 ) ;
  assign n37927 = ( n37370 & ~n37923 ) | ( n37370 & n37925 ) | ( ~n37923 & n37925 ) ;
  assign n37928 = ( n37064 & ~n37926 ) | ( n37064 & n37927 ) | ( ~n37926 & n37927 ) ;
  assign n37929 = ( n36715 & ~n37920 ) | ( n36715 & n37928 ) | ( ~n37920 & n37928 ) ;
  assign n37930 = n37919 & n37929 ;
  assign n37931 = n37919 | n37928 ;
  assign n37932 = n37778 & ~n37919 ;
  assign n37933 = ( n37798 & ~n37919 ) | ( n37798 & n37932 ) | ( ~n37919 & n37932 ) ;
  assign n37934 = ( n36715 & n37931 ) | ( n36715 & ~n37933 ) | ( n37931 & ~n37933 ) ;
  assign n37935 = ~n37930 & n37934 ;
  assign n37936 = n37833 | n37836 ;
  assign n37937 = ~n37833 & n37834 ;
  assign n37938 = ( n37697 & n37936 ) | ( n37697 & ~n37937 ) | ( n37936 & ~n37937 ) ;
  assign n37939 = x53 & n37831 ;
  assign n37940 = x53 | n37831 ;
  assign n37941 = ~n37939 & n37940 ;
  assign n37942 = x118 & n18290 ;
  assign n37943 = x63 & x117 ;
  assign n37944 = ~n18290 & n37943 ;
  assign n37945 = n37942 | n37944 ;
  assign n37946 = n37941 & ~n37945 ;
  assign n37947 = ~n37941 & n37945 ;
  assign n37948 = n37946 | n37947 ;
  assign n37949 = x120 & n17141 ;
  assign n37950 = x119 & ~n17140 ;
  assign n37951 = n17724 & n37950 ;
  assign n37952 = n37949 | n37951 ;
  assign n37953 = x121 & n17146 ;
  assign n37954 = n17149 | n37953 ;
  assign n37955 = n37952 | n37954 ;
  assign n37956 = ~x62 & n37955 ;
  assign n37957 = ~x62 & n37953 ;
  assign n37958 = ( ~x62 & n37952 ) | ( ~x62 & n37957 ) | ( n37952 & n37957 ) ;
  assign n37959 = ( n15501 & n37956 ) | ( n15501 & n37958 ) | ( n37956 & n37958 ) ;
  assign n37960 = x62 & ~n37955 ;
  assign n37961 = x62 & x121 ;
  assign n37962 = n17146 & n37961 ;
  assign n37963 = x62 & ~n37962 ;
  assign n37964 = ~n37952 & n37963 ;
  assign n37965 = ( ~n15501 & n37960 ) | ( ~n15501 & n37964 ) | ( n37960 & n37964 ) ;
  assign n37966 = n37959 | n37965 ;
  assign n37967 = ~n37948 & n37966 ;
  assign n37968 = n37948 & ~n37966 ;
  assign n37969 = n37967 | n37968 ;
  assign n37970 = n37938 & ~n37969 ;
  assign n37971 = ~n37938 & n37969 ;
  assign n37972 = n37970 | n37971 ;
  assign n37973 = x124 & n15552 ;
  assign n37974 = x123 & n15547 ;
  assign n37975 = x122 & ~n15546 ;
  assign n37976 = n16123 & n37975 ;
  assign n37977 = n37974 | n37976 ;
  assign n37978 = n37973 | n37977 ;
  assign n37979 = n15555 | n37973 ;
  assign n37980 = n37977 | n37979 ;
  assign n37981 = ( n17084 & n37978 ) | ( n17084 & n37980 ) | ( n37978 & n37980 ) ;
  assign n37982 = x59 & n37980 ;
  assign n37983 = x59 & n37973 ;
  assign n37984 = ( x59 & n37977 ) | ( x59 & n37983 ) | ( n37977 & n37983 ) ;
  assign n37985 = ( n17084 & n37982 ) | ( n17084 & n37984 ) | ( n37982 & n37984 ) ;
  assign n37986 = x59 & ~n37984 ;
  assign n37987 = x59 & ~n37980 ;
  assign n37988 = ( ~n17084 & n37986 ) | ( ~n17084 & n37987 ) | ( n37986 & n37987 ) ;
  assign n37989 = ( n37981 & ~n37985 ) | ( n37981 & n37988 ) | ( ~n37985 & n37988 ) ;
  assign n37990 = ~n37972 & n37989 ;
  assign n37991 = n37972 | n37990 ;
  assign n37992 = ( n37855 & ~n37857 ) | ( n37855 & n37879 ) | ( ~n37857 & n37879 ) ;
  assign n37993 = n37855 | n37879 ;
  assign n37994 = ( n37838 & n37992 ) | ( n37838 & n37993 ) | ( n37992 & n37993 ) ;
  assign n37995 = n37989 & n37994 ;
  assign n37996 = n37972 & n37995 ;
  assign n37997 = ( ~n37991 & n37994 ) | ( ~n37991 & n37996 ) | ( n37994 & n37996 ) ;
  assign n37998 = n37989 | n37994 ;
  assign n37999 = ( n37972 & n37994 ) | ( n37972 & n37998 ) | ( n37994 & n37998 ) ;
  assign n38000 = n37991 & ~n37999 ;
  assign n38001 = n37997 | n38000 ;
  assign n38002 = x127 & n14045 ;
  assign n38003 = x126 & n14040 ;
  assign n38004 = x125 & ~n14039 ;
  assign n38005 = n14552 & n38004 ;
  assign n38006 = n38003 | n38005 ;
  assign n38007 = n38002 | n38006 ;
  assign n38008 = n14048 | n38002 ;
  assign n38009 = n38006 | n38008 ;
  assign n38010 = ( n18763 & n38007 ) | ( n18763 & n38009 ) | ( n38007 & n38009 ) ;
  assign n38011 = x56 & n38009 ;
  assign n38012 = x56 & n38002 ;
  assign n38013 = ( x56 & n38006 ) | ( x56 & n38012 ) | ( n38006 & n38012 ) ;
  assign n38014 = ( n18763 & n38011 ) | ( n18763 & n38013 ) | ( n38011 & n38013 ) ;
  assign n38015 = x56 & ~n38013 ;
  assign n38016 = x56 & ~n38009 ;
  assign n38017 = ( ~n18763 & n38015 ) | ( ~n18763 & n38016 ) | ( n38015 & n38016 ) ;
  assign n38018 = ( n38010 & ~n38014 ) | ( n38010 & n38017 ) | ( ~n38014 & n38017 ) ;
  assign n38019 = ( n37888 & ~n37889 ) | ( n37888 & n37908 ) | ( ~n37889 & n37908 ) ;
  assign n38020 = ( n38001 & n38018 ) | ( n38001 & ~n38019 ) | ( n38018 & ~n38019 ) ;
  assign n38021 = ( ~n38018 & n38019 ) | ( ~n38018 & n38020 ) | ( n38019 & n38020 ) ;
  assign n38022 = ( ~n38001 & n38020 ) | ( ~n38001 & n38021 ) | ( n38020 & n38021 ) ;
  assign n38023 = ~n37822 & n37910 ;
  assign n38024 = ( n37822 & n37826 ) | ( n37822 & ~n38023 ) | ( n37826 & ~n38023 ) ;
  assign n38025 = ~n38022 & n38024 ;
  assign n38026 = n38022 & ~n38024 ;
  assign n38027 = n38025 | n38026 ;
  assign n38028 = n37918 | n37932 ;
  assign n38029 = ~n37918 & n37919 ;
  assign n38030 = ( n37798 & n38028 ) | ( n37798 & ~n38029 ) | ( n38028 & ~n38029 ) ;
  assign n38031 = ( ~n37918 & n37928 ) | ( ~n37918 & n38029 ) | ( n37928 & n38029 ) ;
  assign n38032 = ( n36715 & ~n38030 ) | ( n36715 & n38031 ) | ( ~n38030 & n38031 ) ;
  assign n38033 = n38027 & n38032 ;
  assign n38034 = n37918 & ~n38027 ;
  assign n38035 = ( n37932 & ~n38027 ) | ( n37932 & n38034 ) | ( ~n38027 & n38034 ) ;
  assign n38036 = ( n37919 & n38027 ) | ( n37919 & ~n38034 ) | ( n38027 & ~n38034 ) ;
  assign n38037 = ( n37798 & n38035 ) | ( n37798 & ~n38036 ) | ( n38035 & ~n38036 ) ;
  assign n38038 = ( n37928 & ~n38034 ) | ( n37928 & n38036 ) | ( ~n38034 & n38036 ) ;
  assign n38039 = ( n36715 & ~n38037 ) | ( n36715 & n38038 ) | ( ~n38037 & n38038 ) ;
  assign n38040 = ~n38033 & n38039 ;
  assign n38120 = n38018 & n38019 ;
  assign n38121 = n38019 & ~n38120 ;
  assign n38122 = n38001 | n38018 ;
  assign n38123 = ( n38001 & ~n38019 ) | ( n38001 & n38122 ) | ( ~n38019 & n38122 ) ;
  assign n38124 = ( ~n38001 & n38120 ) | ( ~n38001 & n38123 ) | ( n38120 & n38123 ) ;
  assign n38125 = n38001 & ~n38018 ;
  assign n38126 = ( n38001 & ~n38019 ) | ( n38001 & n38125 ) | ( ~n38019 & n38125 ) ;
  assign n38127 = ( n38121 & n38124 ) | ( n38121 & ~n38126 ) | ( n38124 & ~n38126 ) ;
  assign n38069 = n37938 | n37967 ;
  assign n38070 = ( n37967 & ~n37969 ) | ( n37967 & n38069 ) | ( ~n37969 & n38069 ) ;
  assign n38041 = x119 & n18290 ;
  assign n38042 = x63 & x118 ;
  assign n38043 = ~n18290 & n38042 ;
  assign n38044 = n38041 | n38043 ;
  assign n38045 = ( ~x53 & n37831 ) | ( ~x53 & n37945 ) | ( n37831 & n37945 ) ;
  assign n38046 = ~n38044 & n38045 ;
  assign n38047 = n38044 & ~n38045 ;
  assign n38048 = n38046 | n38047 ;
  assign n38050 = x121 & n17141 ;
  assign n38051 = x120 & ~n17140 ;
  assign n38052 = n17724 & n38051 ;
  assign n38053 = n38050 | n38052 ;
  assign n38049 = x122 & n17146 ;
  assign n38055 = n17149 | n38049 ;
  assign n38056 = n38053 | n38055 ;
  assign n38054 = n38049 | n38053 ;
  assign n38057 = n38054 & n38056 ;
  assign n38058 = ( n16043 & n38056 ) | ( n16043 & n38057 ) | ( n38056 & n38057 ) ;
  assign n38059 = x62 & n38057 ;
  assign n38060 = x62 & n38056 ;
  assign n38061 = ( n16043 & n38059 ) | ( n16043 & n38060 ) | ( n38059 & n38060 ) ;
  assign n38062 = x62 & ~n38057 ;
  assign n38063 = x62 & ~n38056 ;
  assign n38064 = ( ~n16043 & n38062 ) | ( ~n16043 & n38063 ) | ( n38062 & n38063 ) ;
  assign n38065 = ( n38058 & ~n38061 ) | ( n38058 & n38064 ) | ( ~n38061 & n38064 ) ;
  assign n38066 = ~n38048 & n38065 ;
  assign n38067 = n38048 & ~n38065 ;
  assign n38068 = n38066 | n38067 ;
  assign n38071 = ~n38068 & n38070 ;
  assign n38072 = n38070 & ~n38071 ;
  assign n38073 = x125 & n15552 ;
  assign n38074 = x124 & n15547 ;
  assign n38075 = x123 & ~n15546 ;
  assign n38076 = n16123 & n38075 ;
  assign n38077 = n38074 | n38076 ;
  assign n38078 = n38073 | n38077 ;
  assign n38079 = n15555 | n38073 ;
  assign n38080 = n38077 | n38079 ;
  assign n38081 = ( n17670 & n38078 ) | ( n17670 & n38080 ) | ( n38078 & n38080 ) ;
  assign n38082 = x59 & n38080 ;
  assign n38083 = x59 & n38073 ;
  assign n38084 = ( x59 & n38077 ) | ( x59 & n38083 ) | ( n38077 & n38083 ) ;
  assign n38085 = ( n17670 & n38082 ) | ( n17670 & n38084 ) | ( n38082 & n38084 ) ;
  assign n38086 = x59 & ~n38084 ;
  assign n38087 = x59 & ~n38080 ;
  assign n38088 = ( ~n17670 & n38086 ) | ( ~n17670 & n38087 ) | ( n38086 & n38087 ) ;
  assign n38089 = ( n38081 & ~n38085 ) | ( n38081 & n38088 ) | ( ~n38085 & n38088 ) ;
  assign n38090 = n38068 & ~n38089 ;
  assign n38091 = ( n38070 & ~n38089 ) | ( n38070 & n38090 ) | ( ~n38089 & n38090 ) ;
  assign n38092 = ~n38072 & n38091 ;
  assign n38093 = ~n38068 & n38089 ;
  assign n38094 = ~n38070 & n38093 ;
  assign n38095 = ( n38072 & n38089 ) | ( n38072 & n38094 ) | ( n38089 & n38094 ) ;
  assign n38096 = n38092 | n38095 ;
  assign n38097 = n37990 | n37996 ;
  assign n38098 = n37990 | n37994 ;
  assign n38099 = ( ~n37991 & n38097 ) | ( ~n37991 & n38098 ) | ( n38097 & n38098 ) ;
  assign n38100 = ~n38096 & n38099 ;
  assign n38101 = n38096 & ~n38099 ;
  assign n38102 = n38100 | n38101 ;
  assign n38103 = x127 & n14040 ;
  assign n38104 = x126 & ~n14039 ;
  assign n38105 = n14552 & n38104 ;
  assign n38106 = n38103 | n38105 ;
  assign n38107 = n14048 | n38106 ;
  assign n38108 = ( n19328 & n38106 ) | ( n19328 & n38107 ) | ( n38106 & n38107 ) ;
  assign n38109 = x56 & n38106 ;
  assign n38110 = ( x56 & n17713 ) | ( x56 & n38106 ) | ( n17713 & n38106 ) ;
  assign n38111 = ( n19328 & n38109 ) | ( n19328 & n38110 ) | ( n38109 & n38110 ) ;
  assign n38112 = x56 & ~n17713 ;
  assign n38113 = ~n38106 & n38112 ;
  assign n38114 = x56 & ~n38106 ;
  assign n38115 = ( ~n19328 & n38113 ) | ( ~n19328 & n38114 ) | ( n38113 & n38114 ) ;
  assign n38116 = ( n38108 & ~n38111 ) | ( n38108 & n38115 ) | ( ~n38111 & n38115 ) ;
  assign n38117 = n38102 | n38116 ;
  assign n38118 = n38102 & ~n38116 ;
  assign n38119 = ( ~n38102 & n38117 ) | ( ~n38102 & n38118 ) | ( n38117 & n38118 ) ;
  assign n38128 = ~n38119 & n38127 ;
  assign n38129 = n38127 & ~n38128 ;
  assign n38130 = n38119 | n38127 ;
  assign n38131 = ~n38129 & n38130 ;
  assign n38132 = ~n38025 & n38036 ;
  assign n38133 = ~n38025 & n38027 ;
  assign n38134 = ( n37918 & n38025 ) | ( n37918 & ~n38133 ) | ( n38025 & ~n38133 ) ;
  assign n38135 = ( n37932 & ~n38133 ) | ( n37932 & n38134 ) | ( ~n38133 & n38134 ) ;
  assign n38136 = ( n37798 & ~n38132 ) | ( n37798 & n38135 ) | ( ~n38132 & n38135 ) ;
  assign n38137 = ( n37928 & n38132 ) | ( n37928 & ~n38134 ) | ( n38132 & ~n38134 ) ;
  assign n38138 = ( n36715 & ~n38136 ) | ( n36715 & n38137 ) | ( ~n38136 & n38137 ) ;
  assign n38139 = n38131 & n38138 ;
  assign n38140 = ~n38131 & n38135 ;
  assign n38141 = n38025 & ~n38131 ;
  assign n38142 = ( n38036 & n38131 ) | ( n38036 & ~n38141 ) | ( n38131 & ~n38141 ) ;
  assign n38143 = ( n37798 & n38140 ) | ( n37798 & ~n38142 ) | ( n38140 & ~n38142 ) ;
  assign n38144 = ~n38131 & n38134 ;
  assign n38145 = ( n37928 & n38142 ) | ( n37928 & ~n38144 ) | ( n38142 & ~n38144 ) ;
  assign n38146 = ( n36715 & ~n38143 ) | ( n36715 & n38145 ) | ( ~n38143 & n38145 ) ;
  assign n38147 = ~n38139 & n38146 ;
  assign n38148 = x127 & ~n14039 ;
  assign n38149 = n14552 & n38148 ;
  assign n38150 = n14048 | n38149 ;
  assign n38151 = n19877 | n38149 ;
  assign n38152 = n38150 & n38151 ;
  assign n38153 = n19880 | n38149 ;
  assign n38154 = n38150 & n38153 ;
  assign n38155 = ( n18202 & n38152 ) | ( n18202 & n38154 ) | ( n38152 & n38154 ) ;
  assign n38156 = n38152 & n38154 ;
  assign n38157 = ( n18212 & n38155 ) | ( n18212 & n38156 ) | ( n38155 & n38156 ) ;
  assign n38158 = ( n18214 & n38155 ) | ( n18214 & n38156 ) | ( n38155 & n38156 ) ;
  assign n38159 = ( n14002 & n38157 ) | ( n14002 & n38158 ) | ( n38157 & n38158 ) ;
  assign n38160 = x56 & n38157 ;
  assign n38161 = x56 & n38158 ;
  assign n38162 = ( n14002 & n38160 ) | ( n14002 & n38161 ) | ( n38160 & n38161 ) ;
  assign n38163 = x56 & ~n38161 ;
  assign n38164 = x56 & ~n38160 ;
  assign n38165 = ( ~n14002 & n38163 ) | ( ~n14002 & n38164 ) | ( n38163 & n38164 ) ;
  assign n38166 = ( n38159 & ~n38162 ) | ( n38159 & n38165 ) | ( ~n38162 & n38165 ) ;
  assign n38167 = ~n38068 & n38166 ;
  assign n38168 = n38070 & n38167 ;
  assign n38169 = ( n38094 & n38166 ) | ( n38094 & n38168 ) | ( n38166 & n38168 ) ;
  assign n38170 = ( n38089 & n38166 ) | ( n38089 & n38168 ) | ( n38166 & n38168 ) ;
  assign n38171 = ( n38072 & n38169 ) | ( n38072 & n38170 ) | ( n38169 & n38170 ) ;
  assign n38172 = n38068 & ~n38166 ;
  assign n38173 = ( n38070 & n38166 ) | ( n38070 & ~n38172 ) | ( n38166 & ~n38172 ) ;
  assign n38174 = n38094 | n38173 ;
  assign n38175 = n38089 | n38173 ;
  assign n38176 = ( n38072 & n38174 ) | ( n38072 & n38175 ) | ( n38174 & n38175 ) ;
  assign n38177 = ~n38171 & n38176 ;
  assign n38178 = x122 & n17141 ;
  assign n38179 = x121 & ~n17140 ;
  assign n38180 = n17724 & n38179 ;
  assign n38181 = n38178 | n38180 ;
  assign n38182 = x123 & n17146 ;
  assign n38183 = n17149 | n38182 ;
  assign n38184 = n38181 | n38183 ;
  assign n38185 = ~x62 & n38184 ;
  assign n38186 = ~x62 & n38182 ;
  assign n38187 = ( ~x62 & n38181 ) | ( ~x62 & n38186 ) | ( n38181 & n38186 ) ;
  assign n38188 = ( n16086 & n38185 ) | ( n16086 & n38187 ) | ( n38185 & n38187 ) ;
  assign n38189 = x62 & ~n38184 ;
  assign n38190 = x62 & x123 ;
  assign n38191 = n17146 & n38190 ;
  assign n38192 = x62 & ~n38191 ;
  assign n38193 = ~n38181 & n38192 ;
  assign n38194 = ( ~n16086 & n38189 ) | ( ~n16086 & n38193 ) | ( n38189 & n38193 ) ;
  assign n38195 = n38188 | n38194 ;
  assign n38196 = x120 & n18290 ;
  assign n38197 = x63 & x119 ;
  assign n38198 = ~n18290 & n38197 ;
  assign n38199 = n38196 | n38198 ;
  assign n38200 = ~n38044 & n38199 ;
  assign n38201 = n38044 | n38200 ;
  assign n38202 = n38199 & ~n38200 ;
  assign n38203 = n38201 & ~n38202 ;
  assign n38204 = n38195 & ~n38203 ;
  assign n38205 = ~n38195 & n38203 ;
  assign n38206 = n38204 | n38205 ;
  assign n38207 = ~n38046 & n38048 ;
  assign n38208 = ( n38046 & n38065 ) | ( n38046 & ~n38207 ) | ( n38065 & ~n38207 ) ;
  assign n38209 = n38206 & ~n38208 ;
  assign n38210 = ~n38206 & n38208 ;
  assign n38211 = n38209 | n38210 ;
  assign n38212 = x126 & n15552 ;
  assign n38213 = x125 & n15547 ;
  assign n38214 = x124 & ~n15546 ;
  assign n38215 = n16123 & n38214 ;
  assign n38216 = n38213 | n38215 ;
  assign n38217 = n38212 | n38216 ;
  assign n38218 = n15555 | n38212 ;
  assign n38219 = n38216 | n38218 ;
  assign n38220 = ( n18220 & n38217 ) | ( n18220 & n38219 ) | ( n38217 & n38219 ) ;
  assign n38221 = x59 & n38219 ;
  assign n38222 = x59 & n38212 ;
  assign n38223 = ( x59 & n38216 ) | ( x59 & n38222 ) | ( n38216 & n38222 ) ;
  assign n38224 = ( n18220 & n38221 ) | ( n18220 & n38223 ) | ( n38221 & n38223 ) ;
  assign n38225 = x59 & ~n38223 ;
  assign n38226 = x59 & ~n38219 ;
  assign n38227 = ( ~n18220 & n38225 ) | ( ~n18220 & n38226 ) | ( n38225 & n38226 ) ;
  assign n38228 = ( n38220 & ~n38224 ) | ( n38220 & n38227 ) | ( ~n38224 & n38227 ) ;
  assign n38229 = n38211 & n38228 ;
  assign n38230 = n38208 | n38228 ;
  assign n38231 = ( ~n38206 & n38228 ) | ( ~n38206 & n38230 ) | ( n38228 & n38230 ) ;
  assign n38232 = n38209 | n38231 ;
  assign n38233 = ~n38229 & n38232 ;
  assign n38234 = n38177 & ~n38233 ;
  assign n38235 = n38177 | n38233 ;
  assign n38236 = ( ~n38177 & n38234 ) | ( ~n38177 & n38235 ) | ( n38234 & n38235 ) ;
  assign n38237 = n38100 | n38116 ;
  assign n38238 = ( n38100 & ~n38102 ) | ( n38100 & n38237 ) | ( ~n38102 & n38237 ) ;
  assign n38239 = n38236 & ~n38238 ;
  assign n38240 = ~n38236 & n38238 ;
  assign n38241 = n38239 | n38240 ;
  assign n38242 = ~n38128 & n38131 ;
  assign n38243 = ( n38128 & n38135 ) | ( n38128 & ~n38242 ) | ( n38135 & ~n38242 ) ;
  assign n38244 = n38128 | n38141 ;
  assign n38245 = ( n38036 & n38242 ) | ( n38036 & ~n38244 ) | ( n38242 & ~n38244 ) ;
  assign n38246 = ( n37798 & n38243 ) | ( n37798 & ~n38245 ) | ( n38243 & ~n38245 ) ;
  assign n38247 = ( n38128 & n38134 ) | ( n38128 & ~n38242 ) | ( n38134 & ~n38242 ) ;
  assign n38248 = ( n37928 & n38245 ) | ( n37928 & ~n38247 ) | ( n38245 & ~n38247 ) ;
  assign n38249 = ( n36715 & ~n38246 ) | ( n36715 & n38248 ) | ( ~n38246 & n38248 ) ;
  assign n38250 = n38241 & n38249 ;
  assign n38251 = n38241 | n38242 ;
  assign n38252 = n38128 & ~n38241 ;
  assign n38253 = ( n38135 & ~n38251 ) | ( n38135 & n38252 ) | ( ~n38251 & n38252 ) ;
  assign n38254 = ~n38241 & n38244 ;
  assign n38255 = ( n38036 & n38251 ) | ( n38036 & ~n38254 ) | ( n38251 & ~n38254 ) ;
  assign n38256 = ( n37798 & n38253 ) | ( n37798 & ~n38255 ) | ( n38253 & ~n38255 ) ;
  assign n38257 = ( n38134 & ~n38251 ) | ( n38134 & n38252 ) | ( ~n38251 & n38252 ) ;
  assign n38258 = ( n37928 & n38255 ) | ( n37928 & ~n38257 ) | ( n38255 & ~n38257 ) ;
  assign n38259 = ( n36715 & ~n38256 ) | ( n36715 & n38258 ) | ( ~n38256 & n38258 ) ;
  assign n38260 = ~n38250 & n38259 ;
  assign n38261 = ( n38210 & ~n38211 ) | ( n38210 & n38231 ) | ( ~n38211 & n38231 ) ;
  assign n38262 = x127 & n15552 ;
  assign n38263 = x126 & n15547 ;
  assign n38264 = x125 & ~n15546 ;
  assign n38265 = n16123 & n38264 ;
  assign n38266 = n38263 | n38265 ;
  assign n38267 = n38262 | n38266 ;
  assign n38268 = n15555 | n38262 ;
  assign n38269 = n38266 | n38268 ;
  assign n38270 = ( n18763 & n38267 ) | ( n18763 & n38269 ) | ( n38267 & n38269 ) ;
  assign n38271 = x59 & n38269 ;
  assign n38272 = x59 & n38262 ;
  assign n38273 = ( x59 & n38266 ) | ( x59 & n38272 ) | ( n38266 & n38272 ) ;
  assign n38274 = ( n18763 & n38271 ) | ( n18763 & n38273 ) | ( n38271 & n38273 ) ;
  assign n38275 = x59 & ~n38273 ;
  assign n38276 = x59 & ~n38269 ;
  assign n38277 = ( ~n18763 & n38275 ) | ( ~n18763 & n38276 ) | ( n38275 & n38276 ) ;
  assign n38278 = ( n38270 & ~n38274 ) | ( n38270 & n38277 ) | ( ~n38274 & n38277 ) ;
  assign n38279 = n38231 & n38278 ;
  assign n38280 = n38210 & n38278 ;
  assign n38281 = ( ~n38211 & n38279 ) | ( ~n38211 & n38280 ) | ( n38279 & n38280 ) ;
  assign n38282 = n38261 & ~n38281 ;
  assign n38283 = ~n38231 & n38278 ;
  assign n38284 = ~n38210 & n38278 ;
  assign n38285 = ( n38211 & n38283 ) | ( n38211 & n38284 ) | ( n38283 & n38284 ) ;
  assign n38286 = n38282 | n38285 ;
  assign n38287 = x121 & n18290 ;
  assign n38288 = x63 & x120 ;
  assign n38289 = ~n18290 & n38288 ;
  assign n38290 = n38287 | n38289 ;
  assign n38291 = ~x56 & n38290 ;
  assign n38292 = n38290 & ~n38291 ;
  assign n38293 = x56 | n38290 ;
  assign n38294 = n38044 & ~n38293 ;
  assign n38295 = ( n38044 & n38292 ) | ( n38044 & n38294 ) | ( n38292 & n38294 ) ;
  assign n38296 = ~n38044 & n38293 ;
  assign n38297 = ~n38292 & n38296 ;
  assign n38298 = n38295 | n38297 ;
  assign n38299 = n38200 & ~n38298 ;
  assign n38300 = ( n38203 & n38298 ) | ( n38203 & ~n38299 ) | ( n38298 & ~n38299 ) ;
  assign n38301 = ~n38298 & n38299 ;
  assign n38302 = ( n38195 & ~n38300 ) | ( n38195 & n38301 ) | ( ~n38300 & n38301 ) ;
  assign n38303 = ~n38200 & n38298 ;
  assign n38304 = ~n38200 & n38203 ;
  assign n38305 = n38298 & n38304 ;
  assign n38306 = ( ~n38195 & n38303 ) | ( ~n38195 & n38305 ) | ( n38303 & n38305 ) ;
  assign n38307 = n38302 | n38306 ;
  assign n38308 = x124 & n17146 ;
  assign n38309 = x123 & n17141 ;
  assign n38310 = x122 & ~n17140 ;
  assign n38311 = n17724 & n38310 ;
  assign n38312 = n38309 | n38311 ;
  assign n38313 = n38308 | n38312 ;
  assign n38314 = n17149 | n38308 ;
  assign n38315 = n38312 | n38314 ;
  assign n38316 = ( n17084 & n38313 ) | ( n17084 & n38315 ) | ( n38313 & n38315 ) ;
  assign n38317 = x62 & n38315 ;
  assign n38318 = x62 & n38308 ;
  assign n38319 = ( x62 & n38312 ) | ( x62 & n38318 ) | ( n38312 & n38318 ) ;
  assign n38320 = ( n17084 & n38317 ) | ( n17084 & n38319 ) | ( n38317 & n38319 ) ;
  assign n38321 = x62 & ~n38319 ;
  assign n38322 = x62 & ~n38315 ;
  assign n38323 = ( ~n17084 & n38321 ) | ( ~n17084 & n38322 ) | ( n38321 & n38322 ) ;
  assign n38324 = ( n38316 & ~n38320 ) | ( n38316 & n38323 ) | ( ~n38320 & n38323 ) ;
  assign n38325 = ~n38307 & n38324 ;
  assign n38326 = n38307 & ~n38324 ;
  assign n38327 = n38285 & ~n38326 ;
  assign n38328 = ( n38282 & ~n38326 ) | ( n38282 & n38327 ) | ( ~n38326 & n38327 ) ;
  assign n38329 = ~n38325 & n38328 ;
  assign n38330 = n38286 & ~n38329 ;
  assign n38331 = ~n38171 & n38233 ;
  assign n38332 = ( n38171 & n38177 ) | ( n38171 & ~n38331 ) | ( n38177 & ~n38331 ) ;
  assign n38333 = n38325 | n38326 ;
  assign n38334 = n38328 | n38333 ;
  assign n38335 = n38332 & ~n38334 ;
  assign n38336 = ( n38330 & n38332 ) | ( n38330 & n38335 ) | ( n38332 & n38335 ) ;
  assign n38337 = ~n38332 & n38334 ;
  assign n38338 = ~n38330 & n38337 ;
  assign n38339 = n38336 | n38338 ;
  assign n38340 = ~n38240 & n38255 ;
  assign n38341 = ~n38240 & n38251 ;
  assign n38342 = n38240 | n38252 ;
  assign n38343 = ( n38135 & ~n38341 ) | ( n38135 & n38342 ) | ( ~n38341 & n38342 ) ;
  assign n38344 = ( n37798 & ~n38340 ) | ( n37798 & n38343 ) | ( ~n38340 & n38343 ) ;
  assign n38345 = n38240 | n38257 ;
  assign n38346 = ( n37928 & n38340 ) | ( n37928 & ~n38345 ) | ( n38340 & ~n38345 ) ;
  assign n38347 = ( n36715 & ~n38344 ) | ( n36715 & n38346 ) | ( ~n38344 & n38346 ) ;
  assign n38348 = n38339 & n38347 ;
  assign n38349 = n38339 | n38341 ;
  assign n38350 = ~n38339 & n38342 ;
  assign n38351 = ( n38135 & ~n38349 ) | ( n38135 & n38350 ) | ( ~n38349 & n38350 ) ;
  assign n38352 = n38240 & ~n38339 ;
  assign n38353 = ( n38255 & n38339 ) | ( n38255 & ~n38352 ) | ( n38339 & ~n38352 ) ;
  assign n38354 = ( n37798 & n38351 ) | ( n37798 & ~n38353 ) | ( n38351 & ~n38353 ) ;
  assign n38355 = ( n38257 & ~n38339 ) | ( n38257 & n38352 ) | ( ~n38339 & n38352 ) ;
  assign n38356 = ( n37928 & n38353 ) | ( n37928 & ~n38355 ) | ( n38353 & ~n38355 ) ;
  assign n38357 = ( n36715 & ~n38354 ) | ( n36715 & n38356 ) | ( ~n38354 & n38356 ) ;
  assign n38358 = ~n38348 & n38357 ;
  assign n38359 = x122 & n18290 ;
  assign n38360 = x63 & x121 ;
  assign n38361 = ~n18290 & n38360 ;
  assign n38362 = n38359 | n38361 ;
  assign n38363 = n38291 & ~n38362 ;
  assign n38364 = ( n38295 & ~n38362 ) | ( n38295 & n38363 ) | ( ~n38362 & n38363 ) ;
  assign n38365 = ~n38291 & n38362 ;
  assign n38366 = ~n38295 & n38365 ;
  assign n38367 = n38364 | n38366 ;
  assign n38369 = x124 & n17141 ;
  assign n38370 = x123 & ~n17140 ;
  assign n38371 = n17724 & n38370 ;
  assign n38372 = n38369 | n38371 ;
  assign n38368 = x125 & n17146 ;
  assign n38374 = n17149 | n38368 ;
  assign n38375 = n38372 | n38374 ;
  assign n38373 = n38368 | n38372 ;
  assign n38376 = n38373 & n38375 ;
  assign n38377 = ( n17670 & n38375 ) | ( n17670 & n38376 ) | ( n38375 & n38376 ) ;
  assign n38378 = x62 & n38376 ;
  assign n38379 = x62 & n38375 ;
  assign n38380 = ( n17670 & n38378 ) | ( n17670 & n38379 ) | ( n38378 & n38379 ) ;
  assign n38381 = x62 & ~n38376 ;
  assign n38382 = x62 & ~n38375 ;
  assign n38383 = ( ~n17670 & n38381 ) | ( ~n17670 & n38382 ) | ( n38381 & n38382 ) ;
  assign n38384 = ( n38377 & ~n38380 ) | ( n38377 & n38383 ) | ( ~n38380 & n38383 ) ;
  assign n38385 = ~n38367 & n38384 ;
  assign n38386 = n38367 & ~n38384 ;
  assign n38387 = n38385 | n38386 ;
  assign n38388 = n38302 | n38324 ;
  assign n38389 = ( n38302 & ~n38307 ) | ( n38302 & n38388 ) | ( ~n38307 & n38388 ) ;
  assign n38390 = ~n38387 & n38389 ;
  assign n38391 = n38387 & ~n38389 ;
  assign n38392 = n38390 | n38391 ;
  assign n38393 = x127 & n15547 ;
  assign n38394 = x126 & ~n15546 ;
  assign n38395 = n16123 & n38394 ;
  assign n38396 = n38393 | n38395 ;
  assign n38397 = n15555 | n38396 ;
  assign n38398 = ( n19328 & n38396 ) | ( n19328 & n38397 ) | ( n38396 & n38397 ) ;
  assign n38399 = x59 & n38396 ;
  assign n38400 = ( x59 & n19404 ) | ( x59 & n38396 ) | ( n19404 & n38396 ) ;
  assign n38401 = ( n19328 & n38399 ) | ( n19328 & n38400 ) | ( n38399 & n38400 ) ;
  assign n38402 = x59 & ~n19404 ;
  assign n38403 = ~n38396 & n38402 ;
  assign n38404 = x59 & ~n38396 ;
  assign n38405 = ( ~n19328 & n38403 ) | ( ~n19328 & n38404 ) | ( n38403 & n38404 ) ;
  assign n38406 = ( n38398 & ~n38401 ) | ( n38398 & n38405 ) | ( ~n38401 & n38405 ) ;
  assign n38407 = n38392 | n38406 ;
  assign n38408 = n38392 & ~n38406 ;
  assign n38409 = ( ~n38392 & n38407 ) | ( ~n38392 & n38408 ) | ( n38407 & n38408 ) ;
  assign n38410 = ~n38281 & n38325 ;
  assign n38411 = n38409 | n38410 ;
  assign n38412 = n38281 & ~n38409 ;
  assign n38413 = ( n38328 & ~n38411 ) | ( n38328 & n38412 ) | ( ~n38411 & n38412 ) ;
  assign n38414 = n38409 & n38410 ;
  assign n38415 = ~n38281 & n38409 ;
  assign n38416 = ( ~n38328 & n38414 ) | ( ~n38328 & n38415 ) | ( n38414 & n38415 ) ;
  assign n38417 = n38413 | n38416 ;
  assign n38418 = n38336 | n38351 ;
  assign n38419 = n38336 | n38352 ;
  assign n38420 = ~n38336 & n38339 ;
  assign n38421 = ( n38255 & ~n38419 ) | ( n38255 & n38420 ) | ( ~n38419 & n38420 ) ;
  assign n38422 = ( n37798 & n38418 ) | ( n37798 & ~n38421 ) | ( n38418 & ~n38421 ) ;
  assign n38423 = ( n38257 & n38419 ) | ( n38257 & ~n38420 ) | ( n38419 & ~n38420 ) ;
  assign n38424 = ( n37928 & n38421 ) | ( n37928 & ~n38423 ) | ( n38421 & ~n38423 ) ;
  assign n38425 = ( n36715 & ~n38422 ) | ( n36715 & n38424 ) | ( ~n38422 & n38424 ) ;
  assign n38426 = n38417 & n38425 ;
  assign n38427 = n38336 & ~n38417 ;
  assign n38428 = ( n38351 & ~n38417 ) | ( n38351 & n38427 ) | ( ~n38417 & n38427 ) ;
  assign n38429 = ~n38417 & n38419 ;
  assign n38430 = n38417 | n38420 ;
  assign n38431 = ( n38255 & ~n38429 ) | ( n38255 & n38430 ) | ( ~n38429 & n38430 ) ;
  assign n38432 = ( n37798 & n38428 ) | ( n37798 & ~n38431 ) | ( n38428 & ~n38431 ) ;
  assign n38433 = ( n38257 & n38429 ) | ( n38257 & ~n38430 ) | ( n38429 & ~n38430 ) ;
  assign n38434 = ( n37928 & n38431 ) | ( n37928 & ~n38433 ) | ( n38431 & ~n38433 ) ;
  assign n38435 = ( n36715 & ~n38432 ) | ( n36715 & n38434 ) | ( ~n38432 & n38434 ) ;
  assign n38436 = ~n38426 & n38435 ;
  assign n38501 = n38387 & ~n38406 ;
  assign n38502 = ( n38389 & n38406 ) | ( n38389 & ~n38501 ) | ( n38406 & ~n38501 ) ;
  assign n38503 = ( n38390 & ~n38392 ) | ( n38390 & n38502 ) | ( ~n38392 & n38502 ) ;
  assign n38437 = x123 & n18290 ;
  assign n38438 = x63 & x122 ;
  assign n38439 = ~n18290 & n38438 ;
  assign n38440 = n38437 | n38439 ;
  assign n38441 = ~n38362 & n38440 ;
  assign n38442 = n38362 & ~n38440 ;
  assign n38443 = n38363 & ~n38442 ;
  assign n38444 = n38362 | n38442 ;
  assign n38445 = ( n38295 & n38443 ) | ( n38295 & ~n38444 ) | ( n38443 & ~n38444 ) ;
  assign n38446 = ~n38441 & n38445 ;
  assign n38447 = n38441 | n38442 ;
  assign n38448 = ( n38367 & ~n38446 ) | ( n38367 & n38447 ) | ( ~n38446 & n38447 ) ;
  assign n38449 = ( n38384 & n38446 ) | ( n38384 & ~n38448 ) | ( n38446 & ~n38448 ) ;
  assign n38450 = ( n38364 & n38385 ) | ( n38364 & ~n38449 ) | ( n38385 & ~n38449 ) ;
  assign n38451 = n38441 & ~n38442 ;
  assign n38452 = ( n38442 & n38445 ) | ( n38442 & ~n38451 ) | ( n38445 & ~n38451 ) ;
  assign n38453 = ( n38367 & n38451 ) | ( n38367 & ~n38452 ) | ( n38451 & ~n38452 ) ;
  assign n38454 = ~n38441 & n38453 ;
  assign n38455 = ~n38441 & n38451 ;
  assign n38456 = ( n38445 & n38447 ) | ( n38445 & ~n38455 ) | ( n38447 & ~n38455 ) ;
  assign n38457 = ( n38384 & ~n38454 ) | ( n38384 & n38456 ) | ( ~n38454 & n38456 ) ;
  assign n38458 = ~n38450 & n38457 ;
  assign n38459 = x126 & n17146 ;
  assign n38460 = x125 & n17141 ;
  assign n38461 = x124 & ~n17140 ;
  assign n38462 = n17724 & n38461 ;
  assign n38463 = n38460 | n38462 ;
  assign n38464 = n38459 | n38463 ;
  assign n38465 = n17149 | n38459 ;
  assign n38466 = n38463 | n38465 ;
  assign n38467 = ( n18220 & n38464 ) | ( n18220 & n38466 ) | ( n38464 & n38466 ) ;
  assign n38468 = x62 & n38466 ;
  assign n38469 = x62 & n38459 ;
  assign n38470 = ( x62 & n38463 ) | ( x62 & n38469 ) | ( n38463 & n38469 ) ;
  assign n38471 = ( n18220 & n38468 ) | ( n18220 & n38470 ) | ( n38468 & n38470 ) ;
  assign n38472 = x62 & ~n38470 ;
  assign n38473 = x62 & ~n38466 ;
  assign n38474 = ( ~n18220 & n38472 ) | ( ~n18220 & n38473 ) | ( n38472 & n38473 ) ;
  assign n38475 = ( n38467 & ~n38471 ) | ( n38467 & n38474 ) | ( ~n38471 & n38474 ) ;
  assign n38476 = x127 & ~n15546 ;
  assign n38477 = n16123 & n38476 ;
  assign n38478 = n15555 & n19877 ;
  assign n38479 = n38477 | n38478 ;
  assign n38480 = n15555 & n19880 ;
  assign n38481 = n38477 | n38480 ;
  assign n38482 = ( n18202 & n38479 ) | ( n18202 & n38481 ) | ( n38479 & n38481 ) ;
  assign n38483 = n38479 & n38481 ;
  assign n38484 = ( n18212 & n38482 ) | ( n18212 & n38483 ) | ( n38482 & n38483 ) ;
  assign n38485 = ( n18214 & n38482 ) | ( n18214 & n38483 ) | ( n38482 & n38483 ) ;
  assign n38486 = ( n14002 & n38484 ) | ( n14002 & n38485 ) | ( n38484 & n38485 ) ;
  assign n38487 = x59 & n38484 ;
  assign n38488 = x59 & n38485 ;
  assign n38489 = ( n14002 & n38487 ) | ( n14002 & n38488 ) | ( n38487 & n38488 ) ;
  assign n38490 = x59 & ~n38488 ;
  assign n38491 = x59 & ~n38487 ;
  assign n38492 = ( ~n14002 & n38490 ) | ( ~n14002 & n38491 ) | ( n38490 & n38491 ) ;
  assign n38493 = ( n38486 & ~n38489 ) | ( n38486 & n38492 ) | ( ~n38489 & n38492 ) ;
  assign n38494 = n38475 & n38493 ;
  assign n38495 = n38475 & ~n38494 ;
  assign n38496 = ~n38475 & n38493 ;
  assign n38497 = n38495 | n38496 ;
  assign n38498 = n38458 | n38497 ;
  assign n38499 = n38458 & n38497 ;
  assign n38500 = n38498 & ~n38499 ;
  assign n38504 = ~n38500 & n38503 ;
  assign n38505 = n38503 & ~n38504 ;
  assign n38506 = n38500 | n38503 ;
  assign n38507 = ~n38505 & n38506 ;
  assign n38508 = n38413 | n38427 ;
  assign n38509 = ~n38413 & n38417 ;
  assign n38510 = ( n38351 & n38508 ) | ( n38351 & ~n38509 ) | ( n38508 & ~n38509 ) ;
  assign n38511 = ~n38507 & n38510 ;
  assign n38512 = n38413 | n38429 ;
  assign n38513 = ~n38413 & n38430 ;
  assign n38514 = ( n38255 & ~n38512 ) | ( n38255 & n38513 ) | ( ~n38512 & n38513 ) ;
  assign n38515 = n38507 | n38514 ;
  assign n38516 = ( n37798 & n38511 ) | ( n37798 & ~n38515 ) | ( n38511 & ~n38515 ) ;
  assign n38517 = ( n38257 & n38512 ) | ( n38257 & ~n38513 ) | ( n38512 & ~n38513 ) ;
  assign n38518 = ~n38507 & n38517 ;
  assign n38519 = ( n37928 & n38515 ) | ( n37928 & ~n38518 ) | ( n38515 & ~n38518 ) ;
  assign n38520 = ( n36715 & ~n38516 ) | ( n36715 & n38519 ) | ( ~n38516 & n38519 ) ;
  assign n38521 = ( n37798 & n38510 ) | ( n37798 & ~n38514 ) | ( n38510 & ~n38514 ) ;
  assign n38522 = n38506 & ~n38521 ;
  assign n38523 = ~n38505 & n38522 ;
  assign n38524 = ( n37928 & n38514 ) | ( n37928 & ~n38517 ) | ( n38514 & ~n38517 ) ;
  assign n38525 = n38506 & n38524 ;
  assign n38526 = ~n38505 & n38525 ;
  assign n38527 = ( n36715 & n38523 ) | ( n36715 & n38526 ) | ( n38523 & n38526 ) ;
  assign n38528 = n38520 & ~n38527 ;
  assign n38529 = ( n38384 & n38452 ) | ( n38384 & ~n38453 ) | ( n38452 & ~n38453 ) ;
  assign n38530 = x59 & n38440 ;
  assign n38531 = x59 | n38440 ;
  assign n38532 = ~n38530 & n38531 ;
  assign n38533 = x124 & n18290 ;
  assign n38534 = x63 & x123 ;
  assign n38535 = ~n18290 & n38534 ;
  assign n38536 = n38533 | n38535 ;
  assign n38537 = n38532 & ~n38536 ;
  assign n38538 = ~n38532 & n38536 ;
  assign n38539 = n38537 | n38538 ;
  assign n38540 = x126 & n17141 ;
  assign n38541 = x125 & ~n17140 ;
  assign n38542 = n17724 & n38541 ;
  assign n38543 = n38540 | n38542 ;
  assign n38544 = x127 & n17146 ;
  assign n38545 = n17149 | n38544 ;
  assign n38546 = n38543 | n38545 ;
  assign n38547 = ~x62 & n38546 ;
  assign n38548 = n38543 | n38544 ;
  assign n38549 = ~x62 & n38548 ;
  assign n38550 = ( n18763 & n38547 ) | ( n18763 & n38549 ) | ( n38547 & n38549 ) ;
  assign n38551 = x62 & n38546 ;
  assign n38552 = x62 & ~n38551 ;
  assign n38553 = x62 & n38544 ;
  assign n38554 = ( x62 & n38543 ) | ( x62 & n38553 ) | ( n38543 & n38553 ) ;
  assign n38555 = x62 & ~n38554 ;
  assign n38556 = ( ~n18763 & n38552 ) | ( ~n18763 & n38555 ) | ( n38552 & n38555 ) ;
  assign n38557 = n38550 | n38556 ;
  assign n38558 = ~n38539 & n38557 ;
  assign n38559 = n38539 & ~n38557 ;
  assign n38560 = n38558 | n38559 ;
  assign n38561 = n38529 & ~n38560 ;
  assign n38562 = ~n38529 & n38560 ;
  assign n38563 = n38561 | n38562 ;
  assign n38564 = ( ~n38457 & n38475 ) | ( ~n38457 & n38493 ) | ( n38475 & n38493 ) ;
  assign n38565 = n38475 | n38493 ;
  assign n38566 = ( n38450 & n38564 ) | ( n38450 & n38565 ) | ( n38564 & n38565 ) ;
  assign n38567 = n38563 & n38566 ;
  assign n38568 = ~n38563 & n38566 ;
  assign n38569 = n38563 | n38568 ;
  assign n38570 = ~n38567 & n38569 ;
  assign n38571 = n38504 | n38511 ;
  assign n38572 = ~n38570 & n38571 ;
  assign n38573 = ~n38504 & n38515 ;
  assign n38574 = n38570 | n38573 ;
  assign n38575 = ( n37798 & n38572 ) | ( n37798 & ~n38574 ) | ( n38572 & ~n38574 ) ;
  assign n38576 = n38504 | n38518 ;
  assign n38577 = ~n38570 & n38576 ;
  assign n38578 = ( n37928 & n38574 ) | ( n37928 & ~n38577 ) | ( n38574 & ~n38577 ) ;
  assign n38579 = ( n36715 & ~n38575 ) | ( n36715 & n38578 ) | ( ~n38575 & n38578 ) ;
  assign n38580 = ( n37798 & n38571 ) | ( n37798 & ~n38573 ) | ( n38571 & ~n38573 ) ;
  assign n38581 = ( n37928 & n38573 ) | ( n37928 & ~n38576 ) | ( n38573 & ~n38576 ) ;
  assign n38582 = ( n36715 & ~n38580 ) | ( n36715 & n38581 ) | ( ~n38580 & n38581 ) ;
  assign n38583 = ( n38563 & n38566 ) | ( n38563 & n38582 ) | ( n38566 & n38582 ) ;
  assign n38584 = ( n38567 & n38579 ) | ( n38567 & ~n38583 ) | ( n38579 & ~n38583 ) ;
  assign n38585 = n38529 | n38558 ;
  assign n38586 = ( n38558 & ~n38560 ) | ( n38558 & n38585 ) | ( ~n38560 & n38585 ) ;
  assign n38587 = x125 & n18290 ;
  assign n38588 = x63 & x124 ;
  assign n38589 = ~n18290 & n38588 ;
  assign n38590 = n38587 | n38589 ;
  assign n38591 = ( ~x59 & n38440 ) | ( ~x59 & n38536 ) | ( n38440 & n38536 ) ;
  assign n38592 = ~n38590 & n38591 ;
  assign n38593 = n38590 & ~n38591 ;
  assign n38594 = n38592 | n38593 ;
  assign n38595 = x127 & n17141 ;
  assign n38596 = x126 & ~n17140 ;
  assign n38597 = n17724 & n38596 ;
  assign n38598 = n38595 | n38597 ;
  assign n38599 = n17149 | n38598 ;
  assign n38600 = ( n19328 & n38598 ) | ( n19328 & n38599 ) | ( n38598 & n38599 ) ;
  assign n38601 = x62 & n38599 ;
  assign n38602 = x62 & n38598 ;
  assign n38603 = ( n19328 & n38601 ) | ( n19328 & n38602 ) | ( n38601 & n38602 ) ;
  assign n38604 = x62 & ~n38601 ;
  assign n38605 = x62 & ~n38602 ;
  assign n38606 = ( ~n19328 & n38604 ) | ( ~n19328 & n38605 ) | ( n38604 & n38605 ) ;
  assign n38607 = ( n38600 & ~n38603 ) | ( n38600 & n38606 ) | ( ~n38603 & n38606 ) ;
  assign n38608 = ~n38594 & n38607 ;
  assign n38609 = n38594 & ~n38607 ;
  assign n38610 = n38608 | n38609 ;
  assign n38611 = n38586 & ~n38610 ;
  assign n38612 = n38586 & ~n38611 ;
  assign n38613 = n38586 | n38610 ;
  assign n38614 = ~n38612 & n38613 ;
  assign n38615 = n38568 | n38572 ;
  assign n38616 = ~n38614 & n38615 ;
  assign n38617 = ~n38568 & n38574 ;
  assign n38618 = n38614 | n38617 ;
  assign n38619 = ( n37798 & n38616 ) | ( n37798 & ~n38618 ) | ( n38616 & ~n38618 ) ;
  assign n38620 = n38568 | n38577 ;
  assign n38621 = ~n38614 & n38620 ;
  assign n38622 = ( n37928 & n38618 ) | ( n37928 & ~n38621 ) | ( n38618 & ~n38621 ) ;
  assign n38623 = ( n36715 & ~n38619 ) | ( n36715 & n38622 ) | ( ~n38619 & n38622 ) ;
  assign n38624 = ( n37798 & n38615 ) | ( n37798 & ~n38617 ) | ( n38615 & ~n38617 ) ;
  assign n38625 = ( n37928 & n38617 ) | ( n37928 & ~n38620 ) | ( n38617 & ~n38620 ) ;
  assign n38626 = ( n36715 & ~n38624 ) | ( n36715 & n38625 ) | ( ~n38624 & n38625 ) ;
  assign n38627 = n38623 & ~n38626 ;
  assign n38628 = ( ~n38614 & n38623 ) | ( ~n38614 & n38627 ) | ( n38623 & n38627 ) ;
  assign n38657 = ~n38592 & n38594 ;
  assign n38658 = ( n38592 & n38607 ) | ( n38592 & ~n38657 ) | ( n38607 & ~n38657 ) ;
  assign n38629 = x127 & ~n17140 ;
  assign n38630 = n17724 & n38629 ;
  assign n38631 = n17149 | n38630 ;
  assign n38632 = n19877 | n38630 ;
  assign n38633 = n38631 & n38632 ;
  assign n38634 = n19880 | n38630 ;
  assign n38635 = n38631 & n38634 ;
  assign n38636 = ( n18213 & n38633 ) | ( n18213 & n38635 ) | ( n38633 & n38635 ) ;
  assign n38637 = x62 & n38636 ;
  assign n38638 = ( n18215 & n38633 ) | ( n18215 & n38635 ) | ( n38633 & n38635 ) ;
  assign n38639 = x62 & n38638 ;
  assign n38640 = ( n14002 & n38637 ) | ( n14002 & n38639 ) | ( n38637 & n38639 ) ;
  assign n38641 = x62 & ~n38640 ;
  assign n38642 = x126 & n18290 ;
  assign n38643 = x63 & x125 ;
  assign n38644 = ~n18290 & n38643 ;
  assign n38645 = n38642 | n38644 ;
  assign n38646 = ~n38590 & n38645 ;
  assign n38647 = n38590 & ~n38645 ;
  assign n38648 = n38646 | n38647 ;
  assign n38649 = n38640 | n38648 ;
  assign n38650 = ( n14002 & n38636 ) | ( n14002 & n38638 ) | ( n38636 & n38638 ) ;
  assign n38651 = ~n38648 & n38650 ;
  assign n38652 = ( n38641 & ~n38649 ) | ( n38641 & n38651 ) | ( ~n38649 & n38651 ) ;
  assign n38653 = n38640 & n38648 ;
  assign n38654 = n38648 & ~n38650 ;
  assign n38655 = ( ~n38641 & n38653 ) | ( ~n38641 & n38654 ) | ( n38653 & n38654 ) ;
  assign n38656 = n38652 | n38655 ;
  assign n38659 = ~n38656 & n38658 ;
  assign n38660 = n38658 & ~n38659 ;
  assign n38661 = n38656 | n38658 ;
  assign n38662 = ~n38660 & n38661 ;
  assign n38663 = n38611 | n38616 ;
  assign n38664 = ~n38611 & n38618 ;
  assign n38665 = ( n37798 & n38663 ) | ( n37798 & ~n38664 ) | ( n38663 & ~n38664 ) ;
  assign n38666 = n38611 | n38621 ;
  assign n38667 = ( n37928 & n38664 ) | ( n37928 & ~n38666 ) | ( n38664 & ~n38666 ) ;
  assign n38668 = ( n36713 & ~n38665 ) | ( n36713 & n38667 ) | ( ~n38665 & n38667 ) ;
  assign n38669 = ( n36714 & ~n38665 ) | ( n36714 & n38667 ) | ( ~n38665 & n38667 ) ;
  assign n38670 = ( ~n21078 & n38668 ) | ( ~n21078 & n38669 ) | ( n38668 & n38669 ) ;
  assign n38671 = n38662 & n38670 ;
  assign n38672 = ~n38662 & n38663 ;
  assign n38673 = n38662 | n38664 ;
  assign n38674 = ( n37798 & n38672 ) | ( n37798 & ~n38673 ) | ( n38672 & ~n38673 ) ;
  assign n38675 = ~n38662 & n38666 ;
  assign n38676 = ( n37928 & n38673 ) | ( n37928 & ~n38675 ) | ( n38673 & ~n38675 ) ;
  assign n38677 = ( n36713 & ~n38674 ) | ( n36713 & n38676 ) | ( ~n38674 & n38676 ) ;
  assign n38678 = ( n36714 & ~n38674 ) | ( n36714 & n38676 ) | ( ~n38674 & n38676 ) ;
  assign n38679 = ( ~n21078 & n38677 ) | ( ~n21078 & n38678 ) | ( n38677 & n38678 ) ;
  assign n38680 = ~n38671 & n38679 ;
  assign n38681 = x127 & n18290 ;
  assign n38682 = x63 & x126 ;
  assign n38683 = ~n18290 & n38682 ;
  assign n38684 = n38681 | n38683 ;
  assign n38685 = ~x62 & n38684 ;
  assign n38686 = x62 & ~n38684 ;
  assign n38687 = n38685 | n38686 ;
  assign n38688 = n38590 & ~n38687 ;
  assign n38689 = ~n38590 & n38687 ;
  assign n38690 = n38688 | n38689 ;
  assign n38691 = ( n38646 & n38652 ) | ( n38646 & ~n38690 ) | ( n38652 & ~n38690 ) ;
  assign n38692 = ( ~n38640 & n38641 ) | ( ~n38640 & n38650 ) | ( n38641 & n38650 ) ;
  assign n38693 = ~n38646 & n38648 ;
  assign n38694 = ( n38646 & n38692 ) | ( n38646 & ~n38693 ) | ( n38692 & ~n38693 ) ;
  assign n38695 = n38690 & ~n38694 ;
  assign n38696 = n38691 | n38695 ;
  assign n38697 = n38659 | n38674 ;
  assign n38698 = ~n38659 & n38676 ;
  assign n38699 = ( n36715 & ~n38697 ) | ( n36715 & n38698 ) | ( ~n38697 & n38698 ) ;
  assign n38700 = n38696 & n38699 ;
  assign n38701 = ~n38696 & n38697 ;
  assign n38702 = n38696 | n38698 ;
  assign n38703 = ( n36715 & ~n38701 ) | ( n36715 & n38702 ) | ( ~n38701 & n38702 ) ;
  assign n38704 = ~n38700 & n38703 ;
  assign n38705 = n38691 | n38701 ;
  assign n38706 = ~n38691 & n38702 ;
  assign n38707 = ( n36715 & ~n38705 ) | ( n36715 & n38706 ) | ( ~n38705 & n38706 ) ;
  assign n38708 = x63 & x127 ;
  assign n38709 = ~n18290 & n38708 ;
  assign n38710 = n38685 | n38688 ;
  assign n38711 = n38709 & n38710 ;
  assign n38712 = n38709 | n38710 ;
  assign n38713 = ~n38711 & n38712 ;
  assign n38714 = n38707 & ~n38713 ;
  assign n38715 = n38713 | n38714 ;
  assign n38716 = ( ~n38707 & n38714 ) | ( ~n38707 & n38715 ) | ( n38714 & n38715 ) ;
  assign y0 = n132 ;
  assign y1 = n152 ;
  assign y2 = n175 ;
  assign y3 = n203 ;
  assign y4 = n265 ;
  assign y5 = n315 ;
  assign y6 = n366 ;
  assign y7 = n460 ;
  assign y8 = n539 ;
  assign y9 = n626 ;
  assign y10 = n731 ;
  assign y11 = n833 ;
  assign y12 = n951 ;
  assign y13 = n1086 ;
  assign y14 = n1215 ;
  assign y15 = n1357 ;
  assign y16 = n1523 ;
  assign y17 = n1674 ;
  assign y18 = n1834 ;
  assign y19 = n2034 ;
  assign y20 = n2218 ;
  assign y21 = n2404 ;
  assign y22 = n2628 ;
  assign y23 = n2840 ;
  assign y24 = n3060 ;
  assign y25 = n3305 ;
  assign y26 = n3541 ;
  assign y27 = n3791 ;
  assign y28 = n4063 ;
  assign y29 = n4326 ;
  assign y30 = n4606 ;
  assign y31 = n4921 ;
  assign y32 = n5225 ;
  assign y33 = n5527 ;
  assign y34 = n5872 ;
  assign y35 = n6188 ;
  assign y36 = n6510 ;
  assign y37 = n6867 ;
  assign y38 = n7202 ;
  assign y39 = n7552 ;
  assign y40 = n7932 ;
  assign y41 = n8296 ;
  assign y42 = n8679 ;
  assign y43 = n9107 ;
  assign y44 = n9500 ;
  assign y45 = n9902 ;
  assign y46 = n10354 ;
  assign y47 = n10773 ;
  assign y48 = n11193 ;
  assign y49 = n11656 ;
  assign y50 = n12110 ;
  assign y51 = n12563 ;
  assign y52 = n13054 ;
  assign y53 = n13534 ;
  assign y54 = n14017 ;
  assign y55 = n14519 ;
  assign y56 = n15015 ;
  assign y57 = n15526 ;
  assign y58 = n16066 ;
  assign y59 = n16582 ;
  assign y60 = n17119 ;
  assign y61 = n17702 ;
  assign y62 = n18253 ;
  assign y63 = n18794 ;
  assign y64 = n19352 ;
  assign y65 = n19933 ;
  assign y66 = n20503 ;
  assign y67 = n21079 ;
  assign y68 = n21666 ;
  assign y69 = n22230 ;
  assign y70 = n22797 ;
  assign y71 = n23365 ;
  assign y72 = n23894 ;
  assign y73 = n24475 ;
  assign y74 = n25008 ;
  assign y75 = n25524 ;
  assign y76 = n26033 ;
  assign y77 = n26501 ;
  assign y78 = n26959 ;
  assign y79 = n27392 ;
  assign y80 = n27858 ;
  assign y81 = n28323 ;
  assign y82 = n28761 ;
  assign y83 = n29176 ;
  assign y84 = n29591 ;
  assign y85 = n29975 ;
  assign y86 = n30371 ;
  assign y87 = n30755 ;
  assign y88 = n31120 ;
  assign y89 = n31479 ;
  assign y90 = n31829 ;
  assign y91 = n32159 ;
  assign y92 = n32514 ;
  assign y93 = n32853 ;
  assign y94 = n33163 ;
  assign y95 = n33479 ;
  assign y96 = n33798 ;
  assign y97 = n34077 ;
  assign y98 = n34362 ;
  assign y99 = n34641 ;
  assign y100 = n34901 ;
  assign y101 = n35161 ;
  assign y102 = n35417 ;
  assign y103 = n35636 ;
  assign y104 = n35867 ;
  assign y105 = n36088 ;
  assign y106 = n36290 ;
  assign y107 = n36506 ;
  assign y108 = n36716 ;
  assign y109 = n36889 ;
  assign y110 = n37066 ;
  assign y111 = n37225 ;
  assign y112 = n37373 ;
  assign y113 = n37527 ;
  assign y114 = n37667 ;
  assign y115 = n37800 ;
  assign y116 = n37935 ;
  assign y117 = n38040 ;
  assign y118 = n38147 ;
  assign y119 = n38260 ;
  assign y120 = n38358 ;
  assign y121 = n38436 ;
  assign y122 = n38528 ;
  assign y123 = n38584 ;
  assign y124 = n38628 ;
  assign y125 = n38680 ;
  assign y126 = n38704 ;
  assign y127 = n38716 ;
endmodule
