module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 ;
  assign n12 = ~x5 & x6 ;
  assign n13 = x5 & ~x6 ;
  assign n14 = ~x1 & x2 ;
  assign n15 = x7 | x8 ;
  assign n16 = n14 & ~n15 ;
  assign n17 = x9 | n16 ;
  assign n18 = x1 & ~x2 ;
  assign n19 = x4 & ~x8 ;
  assign n20 = ~x3 & n19 ;
  assign n21 = x4 | x7 ;
  assign n22 = ( n18 & n20 ) | ( n18 & ~n21 ) | ( n20 & ~n21 ) ;
  assign n23 = n18 & n22 ;
  assign n24 = ( n13 & n17 ) | ( n13 & n23 ) | ( n17 & n23 ) ;
  assign n25 = n13 & n24 ;
  assign n26 = ( x9 & n12 ) | ( x9 & n25 ) | ( n12 & n25 ) ;
  assign n27 = x4 & x8 ;
  assign n28 = x6 | x7 ;
  assign n29 = ( x0 & x1 ) | ( x0 & x4 ) | ( x1 & x4 ) ;
  assign n30 = x0 & x1 ;
  assign n31 = x4 | x8 ;
  assign n32 = x0 & ~n31 ;
  assign n33 = ( n29 & ~n30 ) | ( n29 & n32 ) | ( ~n30 & n32 ) ;
  assign n34 = n27 | n33 ;
  assign n35 = ( n27 & ~n28 ) | ( n27 & n34 ) | ( ~n28 & n34 ) ;
  assign n36 = ~x5 & n35 ;
  assign n37 = ~x4 & x5 ;
  assign n38 = ( x8 & n36 ) | ( x8 & n37 ) | ( n36 & n37 ) ;
  assign n39 = x3 & ~x4 ;
  assign n40 = ( x3 & x4 ) | ( x3 & x7 ) | ( x4 & x7 ) ;
  assign n41 = x5 & ~x7 ;
  assign n42 = n18 & n41 ;
  assign n43 = x3 & ~n42 ;
  assign n44 = ( n39 & n40 ) | ( n39 & ~n43 ) | ( n40 & ~n43 ) ;
  assign n45 = ( ~x8 & n36 ) | ( ~x8 & n44 ) | ( n36 & n44 ) ;
  assign n46 = n38 | n45 ;
  assign n47 = ( ~x9 & n25 ) | ( ~x9 & n46 ) | ( n25 & n46 ) ;
  assign n48 = n26 | n47 ;
  assign n49 = ~x10 & n48 ;
  assign n50 = x2 & x3 ;
  assign n51 = x8 | x9 ;
  assign n52 = ( x2 & x3 ) | ( x2 & ~n51 ) | ( x3 & ~n51 ) ;
  assign n53 = ( x10 & ~n50 ) | ( x10 & n52 ) | ( ~n50 & n52 ) ;
  assign n54 = ~x7 & n53 ;
  assign n55 = x9 & x10 ;
  assign n56 = x8 & n55 ;
  assign n57 = n54 | n56 ;
  assign n58 = x6 & n57 ;
  assign n59 = ~x6 & x10 ;
  assign n60 = x7 & n59 ;
  assign n61 = n58 | n60 ;
  assign n62 = n49 | n61 ;
  assign n63 = x4 | x9 ;
  assign n64 = x2 | x7 ;
  assign n65 = n63 & n64 ;
  assign n66 = x1 | n65 ;
  assign n67 = ( ~x0 & x2 ) | ( ~x0 & x7 ) | ( x2 & x7 ) ;
  assign n68 = x1 & x2 ;
  assign n69 = ( x0 & x7 ) | ( x0 & ~n68 ) | ( x7 & ~n68 ) ;
  assign n70 = n67 | n69 ;
  assign n71 = x4 & ~n70 ;
  assign n72 = x8 & ~x9 ;
  assign n73 = n71 | n72 ;
  assign n74 = n66 & ~n73 ;
  assign n75 = x6 | n74 ;
  assign n76 = ~x7 & x9 ;
  assign n77 = x3 & x4 ;
  assign n78 = x7 & ~n77 ;
  assign n79 = n76 | n78 ;
  assign n80 = ( ~n51 & n76 ) | ( ~n51 & n79 ) | ( n76 & n79 ) ;
  assign n81 = n75 & ~n80 ;
  assign n82 = ~x4 & n72 ;
  assign n83 = n76 | n82 ;
  assign n84 = ~x6 & n83 ;
  assign n85 = ( x5 & n81 ) | ( x5 & ~n84 ) | ( n81 & ~n84 ) ;
  assign n86 = x7 & ~x9 ;
  assign n87 = n19 & n86 ;
  assign n88 = x4 | n28 ;
  assign n89 = x9 & n88 ;
  assign n90 = ( ~n19 & n88 ) | ( ~n19 & n89 ) | ( n88 & n89 ) ;
  assign n91 = ( n68 & n87 ) | ( n68 & ~n90 ) | ( n87 & ~n90 ) ;
  assign n92 = x3 & n91 ;
  assign n93 = x4 & n72 ;
  assign n94 = x7 & x9 ;
  assign n95 = n93 | n94 ;
  assign n96 = x6 & n95 ;
  assign n97 = n92 | n96 ;
  assign n98 = ( x5 & n84 ) | ( x5 & n97 ) | ( n84 & n97 ) ;
  assign n99 = n85 & ~n98 ;
  assign n100 = x10 | n99 ;
  assign n101 = x6 & ~x9 ;
  assign n102 = x4 & ~x6 ;
  assign n103 = x4 & x6 ;
  assign n104 = n50 & n103 ;
  assign n105 = ( n101 & n102 ) | ( n101 & n104 ) | ( n102 & n104 ) ;
  assign n106 = x10 | n105 ;
  assign n107 = ~x4 & n101 ;
  assign n108 = ~x1 & n13 ;
  assign n109 = ( ~x3 & n107 ) | ( ~x3 & n108 ) | ( n107 & n108 ) ;
  assign n110 = n106 | n109 ;
  assign n111 = ~x3 & n13 ;
  assign n112 = ( ~x2 & n107 ) | ( ~x2 & n111 ) | ( n107 & n111 ) ;
  assign n113 = n110 | n112 ;
  assign n114 = ~x7 & n113 ;
  assign n115 = n59 | n114 ;
  assign n116 = ~x8 & n115 ;
  assign n117 = x6 & x7 ;
  assign n118 = ( x10 & n72 ) | ( x10 & ~n117 ) | ( n72 & ~n117 ) ;
  assign n119 = n117 & n118 ;
  assign n120 = n116 | n119 ;
  assign n121 = n100 & ~n120 ;
  assign n122 = ~x6 & x7 ;
  assign n123 = x3 & n122 ;
  assign n124 = x6 & ~x7 ;
  assign n125 = ~x2 & n124 ;
  assign n126 = n123 | n125 ;
  assign n127 = ( x5 & n37 ) | ( x5 & ~n126 ) | ( n37 & ~n126 ) ;
  assign n128 = ( ~x5 & n37 ) | ( ~x5 & n117 ) | ( n37 & n117 ) ;
  assign n129 = ( x5 & ~n127 ) | ( x5 & n128 ) | ( ~n127 & n128 ) ;
  assign n130 = x2 & n12 ;
  assign n131 = n108 | n130 ;
  assign n132 = x0 & ~x3 ;
  assign n133 = n102 & n132 ;
  assign n134 = x3 & n37 ;
  assign n135 = n133 | n134 ;
  assign n136 = x1 & n135 ;
  assign n137 = ~n30 & n77 ;
  assign n138 = x5 | x6 ;
  assign n139 = x4 | n138 ;
  assign n140 = ( x5 & ~n137 ) | ( x5 & n139 ) | ( ~n137 & n139 ) ;
  assign n141 = x2 & ~n140 ;
  assign n142 = ( x2 & n136 ) | ( x2 & n141 ) | ( n136 & n141 ) ;
  assign n143 = x3 & ~x6 ;
  assign n144 = ~x2 & n143 ;
  assign n145 = x4 & x5 ;
  assign n146 = ~x3 & n145 ;
  assign n147 = ( x4 & n144 ) | ( x4 & n146 ) | ( n144 & n146 ) ;
  assign n148 = ~x7 & n147 ;
  assign n149 = ( ~x7 & n142 ) | ( ~x7 & n148 ) | ( n142 & n148 ) ;
  assign n150 = ( n77 & n131 ) | ( n77 & n149 ) | ( n131 & n149 ) ;
  assign n151 = x5 & x6 ;
  assign n152 = ( ~n77 & n149 ) | ( ~n77 & n151 ) | ( n149 & n151 ) ;
  assign n153 = n150 | n152 ;
  assign n154 = ~n129 & n153 ;
  assign n155 = ~x8 & n154 ;
  assign n156 = ( ~x9 & n129 ) | ( ~x9 & n155 ) | ( n129 & n155 ) ;
  assign n157 = x10 | n156 ;
  assign n158 = ( n41 & n103 ) | ( n41 & n122 ) | ( n103 & n122 ) ;
  assign n159 = ( x8 & n122 ) | ( x8 & n158 ) | ( n122 & n158 ) ;
  assign n160 = n157 | n159 ;
  assign n161 = x5 & x7 ;
  assign n162 = x8 | x10 ;
  assign n163 = ( x10 & ~n161 ) | ( x10 & n162 ) | ( ~n161 & n162 ) ;
  assign n164 = x9 & n163 ;
  assign n165 = ~x8 & x9 ;
  assign n166 = x5 & n165 ;
  assign n167 = x8 & x10 ;
  assign n168 = ( n117 & n166 ) | ( n117 & n167 ) | ( n166 & n167 ) ;
  assign n169 = n164 | n168 ;
  assign n170 = ( ~x10 & n160 ) | ( ~x10 & n169 ) | ( n160 & n169 ) ;
  assign n171 = x9 | x10 ;
  assign n172 = ~x2 & n117 ;
  assign n173 = x5 & n27 ;
  assign n174 = n172 & n173 ;
  assign n175 = x5 | n15 ;
  assign n176 = ( ~x5 & n139 ) | ( ~x5 & n175 ) | ( n139 & n175 ) ;
  assign n177 = ( n171 & ~n174 ) | ( n171 & n176 ) | ( ~n174 & n176 ) ;
  assign n178 = n171 | n177 ;
  assign n179 = x3 | n178 ;
  assign n180 = x4 | n124 ;
  assign n181 = x7 & ~n151 ;
  assign n182 = ~x9 & n68 ;
  assign n183 = ( x9 & n13 ) | ( x9 & ~n182 ) | ( n13 & ~n182 ) ;
  assign n184 = n181 | n183 ;
  assign n185 = ( ~x3 & x7 ) | ( ~x3 & n111 ) | ( x7 & n111 ) ;
  assign n186 = n184 | n185 ;
  assign n187 = n180 & ~n186 ;
  assign n188 = n30 & ~n138 ;
  assign n189 = ( n50 & n158 ) | ( n50 & n188 ) | ( n158 & n188 ) ;
  assign n190 = n50 & n189 ;
  assign n191 = n187 & ~n190 ;
  assign n192 = x8 | n191 ;
  assign n193 = x4 & x7 ;
  assign n194 = x2 & ~x3 ;
  assign n195 = x3 & x8 ;
  assign n196 = ( n151 & n194 ) | ( n151 & n195 ) | ( n194 & n195 ) ;
  assign n197 = n151 & n196 ;
  assign n198 = ( x9 & n193 ) | ( x9 & ~n197 ) | ( n193 & ~n197 ) ;
  assign n199 = n193 & ~n198 ;
  assign n200 = ( x9 & n76 ) | ( x9 & ~n151 ) | ( n76 & ~n151 ) ;
  assign n201 = n199 | n200 ;
  assign n202 = n192 & ~n201 ;
  assign n203 = x10 | n202 ;
  assign n204 = x8 & n161 ;
  assign n205 = x6 & n204 ;
  assign n206 = ( ~x3 & n30 ) | ( ~x3 & n175 ) | ( n30 & n175 ) ;
  assign n207 = n30 & ~n206 ;
  assign n208 = n205 | n207 ;
  assign n209 = x2 & n208 ;
  assign n210 = ( x3 & n111 ) | ( x3 & n205 ) | ( n111 & n205 ) ;
  assign n211 = n209 | n210 ;
  assign n212 = x4 & n211 ;
  assign n213 = x5 & ~n104 ;
  assign n214 = ( n12 & ~n15 ) | ( n12 & n213 ) | ( ~n15 & n213 ) ;
  assign n215 = n171 | n214 ;
  assign n216 = n212 | n215 ;
  assign n217 = ( n106 & ~n130 ) | ( n106 & n171 ) | ( ~n130 & n171 ) ;
  assign n218 = ( x2 & n171 ) | ( x2 & n217 ) | ( n171 & n217 ) ;
  assign n219 = n15 | n218 ;
  assign y0 = n62 ;
  assign y1 = n121 ;
  assign y2 = n170 ;
  assign y3 = n179 ;
  assign y4 = n203 ;
  assign y5 = n216 ;
  assign y6 = n219 ;
endmodule
