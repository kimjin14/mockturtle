//Written by the Majority Logic Package Fri Nov 14 22:14:15 2014
module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, 
            po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60, po61, po62, po63, po64, po65);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255;
output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60, po61, po62, po63, po64, po65;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211;
assign w0 = ~w974 & ~w1547;
assign w1 = ~w1122 & ~w906;
assign w2 = ~pi231 & w1923;
assign w3 = ~w496 & ~w1051;
assign w4 = ~w69 & ~w1120;
assign w5 = (w1943 & w84) | (w1943 & w2083) | (w84 & w2083);
assign w6 = (~w678 & w1609) | (~w678 & w922) | (w1609 & w922);
assign w7 = ~w1649 & ~w149;
assign w8 = ~w731 & ~w660;
assign w9 = ~w606 & ~w563;
assign w10 = ~w599 & ~w2114;
assign w11 = ~pi180 & ~w233;
assign w12 = ~pi185 & ~w345;
assign w13 = ~w2037 & w450;
assign w14 = ~w1866 & ~w951;
assign w15 = ~w1705 & ~w1141;
assign w16 = ~pi184 & ~w257;
assign w17 = w1459 & ~w1431;
assign w18 = (w1870 & w1941) | (w1870 & w171) | (w1941 & w171);
assign w19 = ~pi147 & ~w1479;
assign w20 = ~w829 & ~w1843;
assign w21 = (~w416 & w1443) | (~w416 & w1836) | (w1443 & w1836);
assign w22 = (w863 & w1975) | (w863 & w447) | (w1975 & w447);
assign w23 = (w1164 & w1344) | (w1164 & w128) | (w1344 & w128);
assign w24 = ~w367 & ~w1955;
assign w25 = (w1237 & w1100) | (w1237 & w231) | (w1100 & w231);
assign w26 = (~w1680 & w783) | (~w1680 & w2210) | (w783 & w2210);
assign w27 = pi171 & w1461;
assign w28 = ~w149 & ~w1147;
assign w29 = ~w1536 & ~w1101;
assign w30 = ~w235 & ~w1257;
assign w31 = ~pi177 & ~w1463;
assign w32 = ~w688 & ~w583;
assign w33 = ~w1081 & ~w1337;
assign w34 = ~pi033 & ~pi097;
assign w35 = pi034 & pi098;
assign w36 = ~w161 & ~w165;
assign w37 = (w2028 & w631) | (w2028 & w806) | (w631 & w806);
assign w38 = pi208 & ~w2192;
assign w39 = (~w56 & w455) | (~w56 & w1573) | (w455 & w1573);
assign w40 = w104 & ~w1111;
assign w41 = ~w376 & w263;
assign w42 = (w489 & w1412) | (w489 & w1254) | (w1412 & w1254);
assign w43 = (~w1968 & w245) | (~w1968 & w920) | (w245 & w920);
assign w44 = ~w1136 & ~w330;
assign w45 = ~w1006 & ~w1599;
assign w46 = ~pi143 & ~w32;
assign w47 = ~w665 & w1584;
assign w48 = ~w838 & ~w628;
assign w49 = (~w301 & ~w1389) | (~w301 & w1902) | (~w1389 & w1902);
assign w50 = (~w980 & w1348) | (~w980 & w376) | (w1348 & w376);
assign w51 = pi139 & w1166;
assign w52 = ~pi176 & ~w1006;
assign w53 = w1134 & ~w1748;
assign w54 = ~w1720 & w1638;
assign w55 = w500 & ~w751;
assign w56 = (~w628 & w1726) | (~w628 & w48) | (w1726 & w48);
assign w57 = (w980 & w774) | (w980 & w404) | (w774 & w404);
assign w58 = w49 & ~w374;
assign w59 = ~w194 & ~w1462;
assign w60 = ~w674 & ~w2077;
assign w61 = ~w187 & w1819;
assign w62 = ~w351 & ~w89;
assign w63 = ~w1716 & ~w532;
assign w64 = pi196 & ~w668;
assign w65 = (~w1147 & ~w1649) | (~w1147 & w28) | (~w1649 & w28);
assign w66 = w1503 & w1906;
assign w67 = w833 & ~w1167;
assign w68 = pi239 & ~w1188;
assign w69 = ~w1120 & ~w1703;
assign w70 = (~w489 & w212) | (~w489 & w2171) | (w212 & w2171);
assign w71 = pi198 & ~w2194;
assign w72 = w1425 & ~w1677;
assign w73 = pi185 & w345;
assign w74 = ~w1261 & ~w260;
assign w75 = (~w2126 & ~w2183) | (~w2126 & w1102) | (~w2183 & w1102);
assign w76 = ~w2059 & ~w2034;
assign w77 = (~w813 & ~w1342) | (~w813 & w2127) | (~w1342 & w2127);
assign w78 = w1893 & w1607;
assign w79 = ~w1920 & ~w1165;
assign w80 = (~w65 & ~w1596) | (~w65 & ~w2088) | (~w1596 & ~w2088);
assign w81 = ~w169 & ~w370;
assign w82 = w1861 & ~w872;
assign w83 = ~w1269 & w318;
assign w84 = ~w275 & ~w1295;
assign w85 = pi203 & ~w1625;
assign w86 = ~w1962 & ~w296;
assign w87 = ~w2088 & ~w1819;
assign w88 = ~w648 & w1405;
assign w89 = w984 & ~w1103;
assign w90 = ~pi226 & w1564;
assign w91 = ~w141 & ~w1721;
assign w92 = (w2067 & w1578) | (w2067 & w916) | (w1578 & w916);
assign w93 = ~w1806 & w756;
assign w94 = (w1196 & w1785) | (w1196 & w1272) | (w1785 & w1272);
assign w95 = ~w1209 & ~w788;
assign w96 = w629 & ~w745;
assign w97 = ~w2143 & ~w312;
assign w98 = ~w2151 & ~w1238;
assign w99 = w440 & w1039;
assign w100 = (~w957 & ~w693) | (~w957 & w837) | (~w693 & w837);
assign w101 = w1680 & ~w217;
assign w102 = w1562 & w1342;
assign w103 = pi158 & w737;
assign w104 = (~w752 & ~w177) | (~w752 & w940) | (~w177 & w940);
assign w105 = (~w35 & ~w602) | (~w35 & w482) | (~w602 & w482);
assign w106 = w1072 & w2092;
assign w107 = ~w1562 & ~w288;
assign w108 = ~pi163 & ~w1315;
assign w109 = w1012 & ~w1556;
assign w110 = pi226 & ~w1564;
assign w111 = ~w424 & ~w29;
assign w112 = (w818 & w859) | (w818 & w416) | (w859 & w416);
assign w113 = ~pi174 & ~w1156;
assign w114 = ~w519 & ~w163;
assign w115 = ~w311 & ~w925;
assign w116 = pi238 & ~w170;
assign w117 = w780 & w36;
assign w118 = (~w584 & ~w1037) | (~w584 & w2196) | (~w1037 & w2196);
assign w119 = ~w1136 & w1991;
assign w120 = (w740 & w1312) | (w740 & ~w1602) | (w1312 & ~w1602);
assign w121 = ~w1756 & ~w1667;
assign w122 = ~w1055 & ~w818;
assign w123 = w391 & ~w822;
assign w124 = ~w1831 & ~w2;
assign w125 = pi219 & ~w875;
assign w126 = ~w1906 & ~w143;
assign w127 = (~w233 & ~w592) | (~w233 & w11) | (~w592 & w11);
assign w128 = ~w1269 & w410;
assign w129 = ~w1711 & ~w1804;
assign w130 = ~w866 & ~w1369;
assign w131 = (~w808 & ~w1650) | (~w808 & w2044) | (~w1650 & w2044);
assign w132 = w1002 & ~w223;
assign w133 = (~w561 & ~w634) | (~w561 & w1004) | (~w634 & w1004);
assign w134 = w2174 & w803;
assign w135 = w208 & ~w122;
assign w136 = (w1041 & w638) | (w1041 & w2064) | (w638 & w2064);
assign w137 = (w585 & ~w1785) | (w585 & ~w43) | (~w1785 & ~w43);
assign w138 = ~w398 & ~w545;
assign w139 = ~w297 & ~w232;
assign w140 = (~w2126 & ~w2183) | (~w2126 & w1677) | (~w2183 & w1677);
assign w141 = (w948 & w2021) | (w948 & w904) | (w2021 & w904);
assign w142 = (w1953 & w1882) | (w1953 & w1139) | (w1882 & w1139);
assign w143 = pi243 & ~w1158;
assign w144 = w985 & w695;
assign w145 = (w1682 & w586) | (w1682 & w500) | (w586 & w500);
assign w146 = ~w1131 & ~w870;
assign w147 = ~w1294 & ~w621;
assign w148 = ~pi139 & ~w1166;
assign w149 = ~w104 & w1111;
assign w150 = pi200 & ~w1290;
assign w151 = (~w1927 & w2026) | (~w1927 & w1591) | (w2026 & w1591);
assign w152 = (w801 & ~w258) | (w801 & ~w2028) | (~w258 & ~w2028);
assign w153 = ~w1295 & ~w88;
assign w154 = ~pi216 & w1173;
assign w155 = (w1098 & w1229) | (w1098 & w915) | (w1229 & w915);
assign w156 = ~w2043 & w1456;
assign w157 = (w553 & w216) | (w553 & ~w416) | (w216 & ~w416);
assign w158 = (w1528 & w1801) | (w1528 & w62) | (w1801 & w62);
assign w159 = ~w408 & ~w578;
assign w160 = ~w1281 & ~w1640;
assign w161 = pi155 & w185;
assign w162 = ~w351 & ~w1528;
assign w163 = ~pi059 & ~pi123;
assign w164 = pi060 & pi124;
assign w165 = ~pi155 & ~w185;
assign w166 = ~pi228 & w382;
assign w167 = (w2028 & w1887) | (w2028 & w598) | (w1887 & w598);
assign w168 = ~pi043 & ~pi107;
assign w169 = pi044 & pi108;
assign w170 = (~w371 & ~w426) | (~w371 & w386) | (~w426 & w386);
assign w171 = (~w1237 & w451) | (~w1237 & w572) | (w451 & w572);
assign w172 = (~w882 & w1532) | (~w882 & w294) | (w1532 & w294);
assign w173 = ~w1747 & w1187;
assign w174 = (w1655 & w2043) | (w1655 & w1808) | (w2043 & w1808);
assign w175 = ~w1453 & ~w650;
assign w176 = ~w2180 & ~w686;
assign w177 = ~w752 & ~w2008;
assign w178 = ~w1760 & ~w2157;
assign w179 = (w1680 & w308) | (w1680 & w1059) | (w308 & w1059);
assign w180 = w1425 & ~w1102;
assign w181 = ~pi187 & ~w519;
assign w182 = (w2047 & w2007) | (w2047 & w610) | (w2007 & w610);
assign w183 = ~w198 & ~w1176;
assign w184 = w1151 & w466;
assign w185 = ~w517 & ~w2032;
assign w186 = ~w995 & ~w1576;
assign w187 = ~w149 & ~w40;
assign w188 = ~w1249 & ~w1905;
assign w189 = ~w440 & ~w1039;
assign w190 = pi236 & ~w1749;
assign w191 = (~w1102 & w1212) | (~w1102 & w884) | (w1212 & w884);
assign w192 = w2094 & w1652;
assign w193 = (w1180 & w355) | (w1180 & w963) | (w355 & w963);
assign w194 = (~w1680 & w112) | (~w1680 & w1341) | (w112 & w1341);
assign w195 = ~w129 & w1870;
assign w196 = (~w190 & ~w2197) | (~w190 & w1288) | (~w2197 & w1288);
assign w197 = w1348 & ~w980;
assign w198 = pi230 & ~w564;
assign w199 = w609 & w1360;
assign w200 = ~pi163 & ~w2141;
assign w201 = w1050 & ~w2076;
assign w202 = w2168 & ~w1047;
assign w203 = (w1150 & w807) | (w1150 & w675) | (w807 & w675);
assign w204 = (~w953 & w947) | (~w953 & w1541) | (w947 & w1541);
assign w205 = ~w885 & ~w1986;
assign w206 = ~w900 & ~w459;
assign w207 = ~w878 & ~w1981;
assign w208 = ~w811 & ~w575;
assign w209 = w431 & w588;
assign w210 = ~pi025 & ~pi089;
assign w211 = pi026 & pi090;
assign w212 = (~w137 & w2158) | (~w137 & w735) | (w2158 & w735);
assign w213 = ~w2136 & ~w2081;
assign w214 = (~w667 & ~w1091) | (~w667 & w1154) | (~w1091 & w1154);
assign w215 = ~pi136 & ~w974;
assign w216 = (~w405 & w1350) | (~w405 & w399) | (w1350 & w399);
assign w217 = ~w1458 & ~w2030;
assign w218 = ~w1057 & ~w674;
assign w219 = w398 & w545;
assign w220 = w1535 & w1702;
assign w221 = ~w376 & w270;
assign w222 = (~w974 & ~w0) | (~w974 & w215) | (~w0 & w215);
assign w223 = ~w147 & ~w246;
assign w224 = w275 & ~w256;
assign w225 = (w2047 & w2007) | (w2047 & w2198) | (w2007 & w2198);
assign w226 = pi188 & w1745;
assign w227 = ~w1021 & ~w1439;
assign w228 = ~w1327 & ~w46;
assign w229 = ~pi011 & ~pi075;
assign w230 = pi012 & pi076;
assign w231 = w849 & ~w1635;
assign w232 = ~pi051 & ~pi115;
assign w233 = pi052 & pi116;
assign w234 = ~pi061 & ~pi125;
assign w235 = pi062 & pi126;
assign w236 = (~w2163 & w109) | (~w2163 & w2203) | (w109 & w2203);
assign w237 = ~pi149 & ~w1128;
assign w238 = (~w1825 & ~w1713) | (~w1825 & w1997) | (~w1713 & w1997);
assign w239 = pi241 & ~w1542;
assign w240 = ~pi220 & w754;
assign w241 = w1091 & w2123;
assign w242 = ~pi197 & w1665;
assign w243 = ~pi195 & w1464;
assign w244 = pi235 & ~w1877;
assign w245 = (~w265 & ~w1555) | (~w265 & w916) | (~w1555 & w916);
assign w246 = w1294 & w621;
assign w247 = ~w1437 & ~w529;
assign w248 = (w2120 & w1237) | (w2120 & ~w915) | (w1237 & ~w915);
assign w249 = (w1115 & w894) | (w1115 & ~w748) | (w894 & ~w748);
assign w250 = ~w1415 & ~w85;
assign w251 = w1759 & ~w1586;
assign w252 = w2143 & w1402;
assign w253 = ~w1295 & ~w1230;
assign w254 = ~w1499 & ~w1717;
assign w255 = (~w326 & w306) | (~w326 & w790) | (w306 & w790);
assign w256 = (~w1295 & w1762) | (~w1295 & w480) | (w1762 & w480);
assign w257 = ~w443 & ~w816;
assign w258 = (w1638 & w56) | (w1638 & w675) | (w56 & w675);
assign w259 = ~w651 & w1971;
assign w260 = ~w1261 & ~w510;
assign w261 = ~w285 & ~w625;
assign w262 = ~w1397 & ~w850;
assign w263 = (~w1711 & w947) | (~w1711 & w1800) | (w947 & w1800);
assign w264 = (~w1543 & w1638) | (~w1543 & w939) | (w1638 & w939);
assign w265 = ~w1837 & w1839;
assign w266 = ~w1548 & ~w1740;
assign w267 = (~w150 & ~w424) | (~w150 & w2086) | (~w424 & w2086);
assign w268 = (~w2028 & w712) | (~w2028 & w565) | (w712 & w565);
assign w269 = ~w2126 & ~w1256;
assign w270 = ~w840 & ~w1417;
assign w271 = ~pi006 & ~pi070;
assign w272 = pi007 & pi071;
assign w273 = ~w208 & ~w811;
assign w274 = ~w376 & w581;
assign w275 = ~w2151 & ~w689;
assign w276 = (~w1402 & ~w1875) | (~w1402 & ~w137) | (~w1875 & ~w137);
assign w277 = ~w2063 & ~w1261;
assign w278 = w908 & w539;
assign w279 = w832 & w782;
assign w280 = (~w2180 & ~w176) | (~w2180 & w1687) | (~w176 & w1687);
assign w281 = ~w1050 & w1313;
assign w282 = ~w970 & ~w1999;
assign w283 = ~w385 & ~w1688;
assign w284 = ~pi022 & ~pi086;
assign w285 = pi023 & pi087;
assign w286 = (~w477 & ~w987) | (~w477 & w732) | (~w987 & w732);
assign w287 = (w1345 & w1603) | (w1345 & w83) | (w1603 & w83);
assign w288 = w196 & ~w1645;
assign w289 = (w394 & w97) | (w394 & w1447) | (w97 & w1447);
assign w290 = (w489 & w1926) | (w489 & w714) | (w1926 & w714);
assign w291 = ~w62 & ~w1610;
assign w292 = ~w376 & ~w1711;
assign w293 = (w1680 & w21) | (w1680 & w1915) | (w21 & w1915);
assign w294 = w680 & ~w1177;
assign w295 = w107 & ~w1404;
assign w296 = ~pi050 & ~pi114;
assign w297 = pi051 & pi115;
assign w298 = ~pi142 & ~w176;
assign w299 = ~w1304 & w530;
assign w300 = ~w1069 & ~w991;
assign w301 = pi244 & ~w478;
assign w302 = ~w786 & ~w1357;
assign w303 = (~w1680 & w1558) | (~w1680 & w998) | (w1558 & w998);
assign w304 = (w1296 & w1919) | (w1296 & w873) | (w1919 & w873);
assign w305 = ~w389 & ~w1340;
assign w306 = ~w2134 & w1268;
assign w307 = ~w2134 & ~w1652;
assign w308 = (~w416 & w1672) | (~w416 & w1112) | (w1672 & w1112);
assign w309 = pi227 & ~w105;
assign w310 = (w792 & w2209) | (w792 & w1485) | (w2209 & w1485);
assign w311 = ~w1309 & ~w1000;
assign w312 = ~w1299 & w2105;
assign w313 = pi245 & ~w127;
assign w314 = ~pi184 & ~w443;
assign w315 = ~w1382 & ~w282;
assign w316 = (~w1688 & w741) | (~w1688 & w283) | (w741 & w283);
assign w317 = w1471 & ~w361;
assign w318 = ~w1181 & ~w507;
assign w319 = ~w1057 & ~w60;
assign w320 = (~w878 & ~w207) | (~w878 & w1840) | (~w207 & w1840);
assign w321 = (w1502 & w1691) | (w1502 & w1307) | (w1691 & w1307);
assign w322 = (~w953 & ~w376) | (~w953 & w2193) | (~w376 & w2193);
assign w323 = ~pi032 & ~pi096;
assign w324 = pi033 & pi097;
assign w325 = (w1680 & w1656) | (w1680 & w770) | (w1656 & w770);
assign w326 = (w881 & w819) | (w881 & ~w644) | (w819 & ~w644);
assign w327 = w62 & w1610;
assign w328 = (~w1870 & w903) | (~w1870 & w2024) | (w903 & w2024);
assign w329 = w2148 & w1088;
assign w330 = ~w391 & w822;
assign w331 = ~pi232 & w1467;
assign w332 = ~pi222 & w1978;
assign w333 = ~w1325 & ~w368;
assign w334 = (~w1185 & w1354) | (~w1185 & w1851) | (w1354 & w1851);
assign w335 = ~w1434 & w1918;
assign w336 = (w1680 & w1428) | (w1680 & w255) | (w1428 & w255);
assign w337 = ~w409 & ~w828;
assign w338 = ~pi204 & w1987;
assign w339 = ~w1458 & ~w360;
assign w340 = ~pi039 & ~pi103;
assign w341 = pi040 & pi104;
assign w342 = ~w1231 & ~w1029;
assign w343 = ~w2078 & ~w228;
assign w344 = ~w1996 & ~w2085;
assign w345 = ~w817 & ~w1034;
assign w346 = w2137 & ~w1161;
assign w347 = w481 & w1417;
assign w348 = ~pi134 & ~w437;
assign w349 = (~w406 & ~w733) | (~w406 & w1719) | (~w733 & w1719);
assign w350 = (w276 & w1590) | (w276 & w1563) | (w1590 & w1563);
assign w351 = ~w984 & w1103;
assign w352 = (~w1927 & w2046) | (~w1927 & w2113) | (w2046 & w2113);
assign w353 = pi202 & ~w1619;
assign w354 = ~w26 & ~w428;
assign w355 = ~w1438 & ~w1120;
assign w356 = ~w838 & ~w1655;
assign w357 = ~w341 & ~w1796;
assign w358 = ~w454 & ~w560;
assign w359 = ~w1852 & ~w2019;
assign w360 = ~w1048 & w1074;
assign w361 = ~w772 & ~w669;
assign w362 = (w489 & w1928) | (w489 & w142) | (w1928 & w142);
assign w363 = ~w1487 & ~w338;
assign w364 = pi161 & w1491;
assign w365 = ~w1893 & ~w1607;
assign w366 = ~pi137 & ~w266;
assign w367 = ~w2012 & ~w1938;
assign w368 = ~w267 & w1818;
assign w369 = (w1583 & w2185) | (w1583 & w6) | (w2185 & w6);
assign w370 = ~pi044 & ~pi108;
assign w371 = pi045 & pi109;
assign w372 = (~w489 & w1811) | (~w489 & w1481) | (w1811 & w1481);
assign w373 = ~w898 & ~w1879;
assign w374 = ~w550 & ~w1323;
assign w375 = pi177 & w1463;
assign w376 = ~w953 & ~w1992;
assign w377 = (~w1870 & w1778) | (~w1870 & w25) | (w1778 & w25);
assign w378 = w1010 & ~w706;
assign w379 = (~w309 & ~w544) | (~w309 & w1414) | (~w544 & w1414);
assign w380 = w2189 | w1635;
assign w381 = ~w2092 & ~w1514;
assign w382 = (~w2141 & ~w1315) | (~w2141 & w200) | (~w1315 & w200);
assign w383 = ~w505 & ~w997;
assign w384 = ~w813 & ~w1342;
assign w385 = ~w1688 & ~w1298;
assign w386 = ~pi173 & ~w371;
assign w387 = ~w743 & ~w1916;
assign w388 = ~w715 & ~w117;
assign w389 = ~w1823 & ~w2098;
assign w390 = pi195 & ~w1464;
assign w391 = (~w659 & ~w1866) | (~w659 & w1220) | (~w1866 & w1220);
assign w392 = ~pi000 & ~pi064;
assign w393 = pi001 & pi065;
assign w394 = ~w262 & w2109;
assign w395 = (~w2082 & ~w1493) | (~w2082 & w639) | (~w1493 & w639);
assign w396 = w1118 & ~w1960;
assign w397 = (~w2066 & ~w1984) | (~w2066 & w511) | (~w1984 & w511);
assign w398 = ~w244 & ~w1500;
assign w399 = ~w833 & w608;
assign w400 = (w1528 & w1801) | (w1528 & w1433) | (w1801 & w1433);
assign w401 = (w948 & w748) | (w948 & w1748) | (w748 & w1748);
assign w402 = ~w205 & ~w1487;
assign w403 = ~w2098 & ~w1699;
assign w404 = (w2074 & w910) | (w2074 & w915) | (w910 & w915);
assign w405 = (~w2064 & w192) | (~w2064 & w434) | (w192 & w434);
assign w406 = pi199 & ~w895;
assign w407 = ~pi019 & ~pi083;
assign w408 = pi020 & pi084;
assign w409 = (w1502 & w549) | (w1502 & w972) | (w549 & w972);
assign w410 = ~w1560 & ~w1045;
assign w411 = ~w1601 & ~w425;
assign w412 = (w135 & w645) | (w135 & w326) | (w645 & w326);
assign w413 = ~pi024 & ~pi088;
assign w414 = pi025 & pi089;
assign w415 = ~w262 & ~w585;
assign w416 = (w881 & w819) | (w881 & ~w1939) | (w819 & ~w1939);
assign w417 = ~w1459 & w1431;
assign w418 = ~pi189 & ~w1725;
assign w419 = ~w217 & ~w1458;
assign w420 = w238 & ~w508;
assign w421 = ~pi159 & ~w213;
assign w422 = ~w1371 & ~w2201;
assign w423 = ~w2052 & ~w555;
assign w424 = ~w150 & ~w515;
assign w425 = pi223 & ~w911;
assign w426 = ~w371 & ~w1155;
assign w427 = ~w2018 & ~w1543;
assign w428 = (w1680 & w1681) | (w1680 & w1683) | (w1681 & w1683);
assign w429 = (~w1197 & ~w642) | (~w1197 & w1608) | (~w642 & w1608);
assign w430 = ~pi169 & ~w1654;
assign w431 = ~w1744 & ~w2121;
assign w432 = w1837 & ~w1839;
assign w433 = (w1778 & w25) | (w1778 & ~w1250) | (w25 & ~w1250);
assign w434 = w2094 & ~w307;
assign w435 = ~w397 & w590;
assign w436 = (~w1748 & w1898) | (~w1748 & w571) | (w1898 & w571);
assign w437 = ~w2035 & ~w271;
assign w438 = ~w1269 & w1152;
assign w439 = (~w312 & ~w1942) | (~w312 & w2109) | (~w1942 & w2109);
assign w440 = ~w239 & ~w1140;
assign w441 = w1325 & ~w571;
assign w442 = ~pi055 & ~pi119;
assign w443 = pi056 & pi120;
assign w444 = ~w1466 & ~w1756;
assign w445 = (~w1502 & w119) | (~w1502 & w1119) | (w119 & w1119);
assign w446 = (w1602 & w2198) | (w1602 & ~w1715) | (w2198 & ~w1715);
assign w447 = (w1775 & w67) | (w1775 & w2094) | (w67 & w2094);
assign w448 = ~w1007 & ~w1617;
assign w449 = ~w838 & w1726;
assign w450 = ~w808 & ~w1650;
assign w451 = w1178 & ~w231;
assign w452 = w1134 & ~w748;
assign w453 = ~pi053 & ~pi117;
assign w454 = pi054 & pi118;
assign w455 = w2018 & w1543;
assign w456 = ~w651 & w1718;
assign w457 = w1511 & ~w1177;
assign w458 = (w1425 & w983) | (w1425 & w1876) | (w983 & w1876);
assign w459 = ~pi224 & w927;
assign w460 = ~w95 & ~w198;
assign w461 = w833 & w1585;
assign w462 = (~w1502 & w1019) | (~w1502 & w1544) | (w1019 & w1544);
assign w463 = w1912 & ~w1927;
assign w464 = (w975 & w1403) | (w975 & w644) | (w1403 & w644);
assign w465 = w642 & w1709;
assign w466 = ~w335 & ~w1339;
assign w467 = (~w1502 & w1929) | (~w1502 & w996) | (w1929 & w996);
assign w468 = ~w1008 & w1495;
assign w469 = ~w73 & ~w12;
assign w470 = ~w1716 & ~w1090;
assign w471 = ~w1397 & ~w1942;
assign w472 = w187 & ~w2088;
assign w473 = ~pi017 & ~pi081;
assign w474 = pi018 & pi082;
assign w475 = (~w489 & w1478) | (~w489 & w2010) | (w1478 & w2010);
assign w476 = pi141 & w600;
assign w477 = pi215 & ~w1246;
assign w478 = (~w297 & ~w139) | (~w297 & w1075) | (~w139 & w1075);
assign w479 = ~w567 & ~w1595;
assign w480 = ~w2143 & ~w88;
assign w481 = ~w49 & w374;
assign w482 = ~pi162 & ~w35;
assign w483 = (~w519 & ~w114) | (~w519 & w181) | (~w114 & w181);
assign w484 = (w6 & w80) | (w6 & w1204) | (w80 & w1204);
assign w485 = (w1911 & w2003) | (w1911 & w622) | (w2003 & w622);
assign w486 = pi207 & ~w280;
assign w487 = (w173 & w730) | (w173 & ~w1100) | (w730 & ~w1100);
assign w488 = (w1502 & w1631) | (w1502 & w610) | (w1631 & w610);
assign w489 = (~w2028 & w1913) | (~w2028 & w2025) | (w1913 & w2025);
assign w490 = (~w276 & w224) | (~w276 & w1200) | (w224 & w1200);
assign w491 = (w2044 & w595) | (w2044 & w551) | (w595 & w551);
assign w492 = w1720 & w152;
assign w493 = ~w2167 & ~w110;
assign w494 = ~w763 & ~w1731;
assign w495 = ~pi181 & ~w1452;
assign w496 = pi252 & ~w483;
assign w497 = pi163 & w1315;
assign w498 = (w980 & w708) | (w980 & w1627) | (w708 & w1627);
assign w499 = (~w980 & w1227) | (~w980 & w1545) | (w1227 & w1545);
assign w500 = ~w1386 & ~w1789;
assign w501 = (~w408 & ~w159) | (~w408 & w1886) | (~w159 & w1886);
assign w502 = ~w1218 & ~w331;
assign w503 = (~w390 & ~w1382) | (~w390 & w1056) | (~w1382 & w1056);
assign w504 = w206 & w1930;
assign w505 = (w1502 & w798) | (w1502 & w2084) | (w798 & w2084);
assign w506 = ~w849 & w1635;
assign w507 = ~w759 & w522;
assign w508 = ~w2147 & ~w1076;
assign w509 = w887 & w1283;
assign w510 = w968 & ~w853;
assign w511 = ~w1149 & ~w2066;
assign w512 = w2078 & w228;
assign w513 = ~w2094 & w1792;
assign w514 = ~w1984 & ~w1149;
assign w515 = ~pi200 & w1290;
assign w516 = ~pi026 & ~pi090;
assign w517 = pi027 & pi091;
assign w518 = ~pi058 & ~pi122;
assign w519 = pi059 & pi123;
assign w520 = ~pi012 & ~pi076;
assign w521 = pi013 & pi077;
assign w522 = ~w1117 & ~w106;
assign w523 = w187 & w826;
assign w524 = (w1179 & w1345) | (w1179 & w1102) | (w1345 & w1102);
assign w525 = w335 & w1950;
assign w526 = ~w1469 & ~w1429;
assign w527 = (w1735 & w723) | (w1735 & ~w644) | (w723 & ~w644);
assign w528 = ~w124 & ~w1399;
assign w529 = w987 & w2133;
assign w530 = ~w1712 & ~w241;
assign w531 = w2063 & w260;
assign w532 = ~pi255 & ~w949;
assign w533 = pi213 & ~w501;
assign w534 = ~pi001 & ~pi065;
assign w535 = pi002 & pi066;
assign w536 = ~w695 & ~w1890;
assign w537 = ~w1225 & ~w279;
assign w538 = ~w1286 & ~w599;
assign w539 = ~w1501 & ~w2181;
assign w540 = w262 & w585;
assign w541 = ~pi173 & ~w426;
assign w542 = pi173 & w426;
assign w543 = (w980 & w1489) | (w980 & w404) | (w1489 & w404);
assign w544 = ~w309 & ~w2172;
assign w545 = ~w27 & ~w842;
assign w546 = (w98 & w2162) | (w98 & ~w1329) | (w2162 & ~w1329);
assign w547 = ~pi239 & w1188;
assign w548 = (~w1410 & ~w1893) | (~w1410 & w1401) | (~w1893 & w1401);
assign w549 = (w882 & w1177) | (w882 & w1876) | (w1177 & w1876);
assign w550 = ~w697 & ~w1692;
assign w551 = ~w651 & w2044;
assign w552 = ~w2073 & ~w2177;
assign w553 = (~w1108 & w399) | (~w1108 & w1284) | (w399 & w1284);
assign w554 = ~w376 & w947;
assign w555 = (w1680 & w1003) | (w1680 & w1248) | (w1003 & w1248);
assign w556 = ~w485 & ~w179;
assign w557 = ~w62 & w162;
assign w558 = w838 & w1655;
assign w559 = (w1502 & w717) | (w1502 & w800) | (w717 & w800);
assign w560 = ~pi054 & ~pi118;
assign w561 = pi055 & pi119;
assign w562 = w424 & w29;
assign w563 = ~pi210 & w883;
assign w564 = (~w1566 & ~w1727) | (~w1566 & w958) | (~w1727 & w958);
assign w565 = (~w1320 & w670) | (~w1320 & w1704) | (w670 & w1704);
assign w566 = ~w1088 & ~w68;
assign w567 = pi183 & w634;
assign w568 = (~w1494 & ~w1965) | (~w1494 & w1297) | (~w1965 & w1297);
assign w569 = ~pi158 & ~w1880;
assign w570 = ~w630 & w1734;
assign w571 = (~w599 & ~w10) | (~w599 & w538) | (~w10 & w538);
assign w572 = w1178 & ~w1100;
assign w573 = (w1655 & ~w1726) | (w1655 & ~w1456) | (~w1726 & ~w1456);
assign w574 = w1269 & w1705;
assign w575 = w1205 & ~w704;
assign w576 = ~w129 & w915;
assign w577 = ~w1496 & ~w656;
assign w578 = ~pi020 & ~pi084;
assign w579 = pi021 & pi085;
assign w580 = ~w1259 & ~w1601;
assign w581 = (~w840 & ~w1417) | (~w840 & w2093) | (~w1417 & w2093);
assign w582 = ~w762 & ~w2058;
assign w583 = ~pi015 & ~pi079;
assign w584 = pi016 & pi080;
assign w585 = ~w1002 & w223;
assign w586 = ~w187 & ~w1789;
assign w587 = w3 & w1333;
assign w588 = ~w542 & ~w541;
assign w589 = ~pi190 & ~w235;
assign w590 = ~w315 & ~w1579;
assign w591 = (w1311 & w1380) | (w1311 & w1033) | (w1380 & w1033);
assign w592 = ~w233 & ~w1317;
assign w593 = ~pi190 & ~w30;
assign w594 = w1521 & ~w2182;
assign w595 = (~w1606 & w65) | (~w1606 & w1718) | (w65 & w1718);
assign w596 = ~w1022 & ~w1270;
assign w597 = (w1502 & w400) | (w1502 & w1400) | (w400 & w1400);
assign w598 = (w1320 & w1957) | (w1320 & w156) | (w1957 & w156);
assign w599 = ~w349 & w805;
assign w600 = ~w521 & ~w2179;
assign w601 = w1894 & w2101;
assign w602 = ~w35 & ~w2140;
assign w603 = (w1041 & w638) | (w1041 & w1268) | (w638 & w1268);
assign w604 = ~w1095 & ~w1998;
assign w605 = ~w2042 & ~w943;
assign w606 = pi210 & ~w883;
assign w607 = ~w211 & ~w516;
assign w608 = (~w47 & ~w2208) | (~w47 & w1792) | (~w2208 & w1792);
assign w609 = ~w1700 & ~w1023;
assign w610 = (~w980 & w446) | (~w980 & w1262) | (w446 & w1262);
assign w611 = ~w1803 & ~w1228;
assign w612 = ~pi188 & ~w164;
assign w613 = w1325 & ~w1898;
assign w614 = (w1342 & w1927) | (w1342 & w102) | (w1927 & w102);
assign w615 = ~w290 & ~w1799;
assign w616 = ~w804 & ~w311;
assign w617 = ~pi164 & ~w693;
assign w618 = (~w1502 & w18) | (~w1502 & w2206) | (w18 & w2206);
assign w619 = (~w1680 & w1976) | (~w1680 & w6) | (w1976 & w6);
assign w620 = (w1650 & w1815) | (w1650 & w651) | (w1815 & w651);
assign w621 = ~w1626 & ~w19;
assign w622 = (w326 & w1114) | (w326 & w967) | (w1114 & w967);
assign w623 = ~w1937 & ~w1763;
assign w624 = ~w93 & ~w1087;
assign w625 = ~pi023 & ~pi087;
assign w626 = pi024 & pi088;
assign w627 = w1832 & w2208;
assign w628 = ~w238 & w508;
assign w629 = (~w353 & ~w908) | (~w353 & w858) | (~w908 & w858);
assign w630 = ~w1286 & ~w1706;
assign w631 = ~w809 & w1871;
assign w632 = ~pi180 & ~w592;
assign w633 = (w1502 & w692) | (w1502 & w2154) | (w692 & w2154);
assign w634 = ~w561 & ~w442;
assign w635 = ~w15 & ~w813;
assign w636 = (~w1502 & w1914) | (~w1502 & w1217) | (w1914 & w1217);
assign w637 = ~w1362 & ~w360;
assign w638 = ~w2094 & w307;
assign w639 = ~pi160 & ~w2082;
assign w640 = (~w1514 & ~w1072) | (~w1514 & w381) | (~w1072 & w381);
assign w641 = w62 & ~w1071;
assign w642 = ~w1197 & ~w1506;
assign w643 = (w678 & w1621) | (w678 & w847) | (w1621 & w847);
assign w644 = (~w6 & w1819) | (~w6 & w2088) | (w1819 & w2088);
assign w645 = w208 & ~w1597;
assign w646 = w1181 & w1705;
assign w647 = (w1164 & w1344) | (w1164 & w410) | (w1344 & w410);
assign w648 = (~w533 & ~w1894) | (~w533 & w1907) | (~w1894 & w1907);
assign w649 = ~w262 & w1785;
assign w650 = pi248 & ~w133;
assign w651 = ~w299 & ~w2017;
assign w652 = (w231 & w753) | (w231 & w1375) | (w753 & w1375);
assign w653 = ~w359 & ~w2089;
assign w654 = ~pi171 & ~w1216;
assign w655 = (~w650 & ~w1570) | (~w650 & w175) | (~w1570 & w175);
assign w656 = ~w1512 & ~w348;
assign w657 = ~w1968 & ~w265;
assign w658 = ~w982 & ~w475;
assign w659 = pi234 & ~w1169;
assign w660 = w1036 & w302;
assign w661 = w1390 & ~w868;
assign w662 = ~pi135 & ~w1419;
assign w663 = ~w950 & ~w1865;
assign w664 = (w1303 & w913) | (w1303 & ~w1875) | (w913 & ~w1875);
assign w665 = (~w1831 & ~w124) | (~w1831 & w1540) | (~w124 & w1540);
assign w666 = (w1502 & w1433) | (w1502 & w1810) | (w1433 & w1810);
assign w667 = pi225 & ~w395;
assign w668 = (~w857 & ~w1842) | (~w857 & w775) | (~w1842 & w775);
assign w669 = w363 & w205;
assign w670 = w2043 & w1974;
assign w671 = ~w535 & ~w856;
assign w672 = ~w160 & ~w1319;
assign w673 = (~w817 & ~w345) | (~w817 & w929) | (~w345 & w929);
assign w674 = ~w1782 & w749;
assign w675 = (~w1974 & w1320) | (~w1974 & w1456) | (w1320 & w1456);
assign w676 = w648 & ~w1405;
assign w677 = ~pi206 & w1015;
assign w678 = (~w360 & w419) | (~w360 & w637) | (w419 & w637);
assign w679 = ~w1560 & ~w931;
assign w680 = ~w1181 & ~w1705;
assign w681 = (w260 & w531) | (w260 & w231) | (w531 & w231);
assign w682 = ~pi181 & ~w1318;
assign w683 = w1180 & ~w69;
assign w684 = w928 & ~w204;
assign w685 = w2126 | w1705;
assign w686 = ~pi014 & ~pi078;
assign w687 = (~w1320 & w174) | (~w1320 & w573) | (w174 & w573);
assign w688 = pi015 & pi079;
assign w689 = w286 & ~w1;
assign w690 = (w1696 & w1144) | (w1696 & w1939) | (w1144 & w1939);
assign w691 = (~w1742 & ~w1294) | (~w1742 & w1001) | (~w1294 & w1001);
assign w692 = (~w1715 & w1812) | (~w1715 & w1080) | (w1812 & w1080);
assign w693 = ~w957 & ~w1565;
assign w694 = ~w230 & ~w520;
assign w695 = ~w1366 & ~w2129;
assign w696 = ~pi143 & ~w688;
assign w697 = ~w313 & ~w1863;
assign w698 = (w1555 & w489) | (w1555 & w2202) | (w489 & w2202);
assign w699 = (w1179 & w1345) | (w1179 & w1677) | (w1345 & w1677);
assign w700 = ~w1042 & ~w392;
assign w701 = ~w1894 & ~w2101;
assign w702 = ~w864 & ~w632;
assign w703 = (~w1133 & w1061) | (~w1133 & w158) | (w1061 & w158);
assign w704 = ~w1301 & ~w465;
assign w705 = ~w1282 & ~w1820;
assign w706 = (~w1268 & w192) | (~w1268 & w434) | (w192 & w434);
assign w707 = w787 & w2170;
assign w708 = (w1518 & w41) | (w1518 & w971) | (w41 & w971);
assign w709 = ~pi188 & ~w1745;
assign w710 = ~pi179 & ~w139;
assign w711 = ~w867 & ~w329;
assign w712 = w2043 & ~w1980;
assign w713 = ~pi201 & w222;
assign w714 = w1901 & ~w245;
assign w715 = ~w780 & ~w36;
assign w716 = ~w1649 & ~w1967;
assign w717 = (w1927 & w180) | (w1927 & w72) | (w180 & w72);
assign w718 = (w204 & w1326) | (w204 & w1387) | (w1326 & w1387);
assign w719 = (~w1680 & w896) | (~w1680 & w1567) | (w896 & w1567);
assign w720 = ~pi212 & w1660;
assign w721 = ~pi133 & ~w76;
assign w722 = ~pi133 & ~w2059;
assign w723 = (w1650 & w1815) | (w1650 & w1538) | (w1815 & w1538);
assign w724 = (w1735 & w723) | (w1735 & ~w1939) | (w723 & ~w1939);
assign w725 = (w1528 & w1801) | (w1528 & w2120) | (w1801 & w2120);
assign w726 = w1397 & w1942;
assign w727 = (w915 & w1387) | (w915 & w1646) | (w1387 & w1646);
assign w728 = (~w2033 & ~w1813) | (~w2033 & w1376) | (~w1813 & w1376);
assign w729 = w1560 & w931;
assign w730 = ~w1747 & w74;
assign w731 = ~w1036 & ~w302;
assign w732 = ~w2133 & ~w477;
assign w733 = ~w406 & ~w2125;
assign w734 = w1211 & w1415;
assign w735 = ~w2143 & ~w1875;
assign w736 = ~pi165 & ~w1727;
assign w737 = ~w1880 & ~w2135;
assign w738 = (w1583 & w2185) | (w1583 & w751) | (w2185 & w751);
assign w739 = ~w1753 & ~w1969;
assign w740 = ~w466 & w1454;
assign w741 = (~w360 & ~w1362) | (~w360 & w339) | (~w1362 & w339);
assign w742 = ~w633 & ~w1391;
assign w743 = (w1502 & w776) | (w1502 & w614) | (w776 & w614);
assign w744 = (w236 & w760) | (w236 & w1715) | (w760 & w1715);
assign w745 = ~w1829 & ~w734;
assign w746 = ~pi202 & w1619;
assign w747 = (~w532 & ~w1090) | (~w532 & w63) | (~w1090 & w63);
assign w748 = w630 & ~w1734;
assign w749 = ~w577 & ~w1432;
assign w750 = (~w1261 & ~w260) | (~w1261 & w944) | (~w260 & w944);
assign w751 = ~w1386 & ~w988;
assign w752 = pi221 & ~w728;
assign w753 = w1747 & ~w1187;
assign w754 = (~w517 & ~w185) | (~w517 & w1046) | (~w185 & w1046);
assign w755 = ~w1104 & ~w2205;
assign w756 = ~w435 & ~w1896;
assign w757 = w207 & w1888;
assign w758 = w1866 & w951;
assign w759 = (~w239 & ~w440) | (~w239 & w1791) | (~w440 & w1791);
assign w760 = (~w792 & w1193) | (~w792 & w1824) | (w1193 & w1824);
assign w761 = ~pi003 & ~pi067;
assign w762 = pi004 & pi068;
assign w763 = pi233 & ~w1279;
assign w764 = ~w2000 & ~w763;
assign w765 = ~w1569 & w65;
assign w766 = (~w995 & ~w186) | (~w995 & w926) | (~w186 & w926);
assign w767 = (w1556 & w2107) | (w1556 & w1385) | (w2107 & w1385);
assign w768 = (~w169 & ~w81) | (~w169 & w1534) | (~w81 & w1534);
assign w769 = ~w1710 & ~w359;
assign w770 = ~w6 & w1857;
assign w771 = pi178 & w86;
assign w772 = ~w363 & ~w205;
assign w773 = ~w1194 & ~w2122;
assign w774 = (w2074 & w910) | (w2074 & w1715) | (w910 & w1715);
assign w775 = ~pi131 & ~w857;
assign w776 = (w1342 & w882) | (w1342 & w102) | (w882 & w102);
assign w777 = ~w803 & ~w1052;
assign w778 = (w1682 & w586) | (w1682 & w55) | (w586 & w55);
assign w779 = ~w42 & ~w1571;
assign w780 = ~w125 & ~w1934;
assign w781 = ~w663 & ~w1218;
assign w782 = ~w1292 & ~w617;
assign w783 = w1362 & w1458;
assign w784 = ~pi018 & ~pi082;
assign w785 = pi019 & pi083;
assign w786 = pi132 & w582;
assign w787 = w2143 & ~w439;
assign w788 = ~pi166 & ~w526;
assign w789 = ~pi196 & w668;
assign w790 = ~w2134 & w2064;
assign w791 = w635 & w2146;
assign w792 = (~w1345 & w1910) | (~w1345 & w1332) | (w1910 & w1332);
assign w793 = (w1870 & w1387) | (w1870 & w1646) | (w1387 & w1646);
assign w794 = ~w351 & ~w1795;
assign w795 = w1649 & w1967;
assign w796 = ~w1930 & ~w900;
assign w797 = (~w1275 & ~w2103) | (~w1275 & w1848) | (~w2103 & w1848);
assign w798 = (~w1870 & w1212) | (~w1870 & w884) | (w1212 & w884);
assign w799 = w1844 & ~w976;
assign w800 = (w882 & w458) | (w882 & w901) | (w458 & w901);
assign w801 = (~w1638 & ~w56) | (~w1638 & ~w1980) | (~w56 & ~w1980);
assign w802 = (~w1185 & w1130) | (~w1185 & w812) | (w1130 & w812);
assign w803 = ~w1135 & ~w366;
assign w804 = ~w925 & ~w720;
assign w805 = ~w562 & ~w111;
assign w806 = ~w809 & w1320;
assign w807 = ~w2018 & w264;
assign w808 = ~w214 & w1381;
assign w809 = ~w1974 & ~w317;
assign w810 = ~pi150 & ~w979;
assign w811 = ~w1205 & w704;
assign w812 = (w396 & w1556) | (w396 & w792) | (w1556 & w792);
assign w813 = ~w1761 & w254;
assign w814 = (~w882 & w1689) | (~w882 & w1728) | (w1689 & w1728);
assign w815 = (w1334 & w1919) | (w1334 & w873) | (w1919 & w873);
assign w816 = ~pi056 & ~pi120;
assign w817 = pi057 & pi121;
assign w818 = ~w1055 & ~w1276;
assign w819 = (w1040 & w1407) | (w1040 & w1510) | (w1407 & w1510);
assign w820 = (w2076 & w941) | (w2076 & w1959) | (w941 & w1959);
assign w821 = (~w1329 & w1247) | (~w1329 & w5) | (w1247 & w5);
assign w822 = ~w138 & ~w219;
assign w823 = (~w335 & ~w466) | (~w335 & w889) | (~w466 & w889);
assign w824 = w2018 & ~w264;
assign w825 = w1984 & w1149;
assign w826 = (~w316 & w87) | (~w316 & w1393) | (w87 & w1393);
assign w827 = w1449 & ~w942;
assign w828 = (~w1502 & w986) | (~w1502 & w845) | (w986 & w845);
assign w829 = ~w1794 & ~w367;
assign w830 = pi184 & w257;
assign w831 = (w204 & w1588) | (w204 & w1387) | (w1588 & w1387);
assign w832 = ~w2002 & ~w166;
assign w833 = ~w1249 & ~w1629;
assign w834 = ~pi243 & w1158;
assign w835 = ~w1118 & w1012;
assign w836 = ~w782 & ~w2002;
assign w837 = ~pi164 & ~w957;
assign w838 = ~w628 & ~w420;
assign w839 = ~pi178 & ~w1962;
assign w840 = ~w1390 & w868;
assign w841 = ~pi153 & ~w959;
assign w842 = ~pi171 & ~w1461;
assign w843 = pi160 & w1493;
assign w844 = ~w849 & w1736;
assign w845 = (~w1927 & w1841) | (~w1927 & w1527) | (w1841 & w1527);
assign w846 = (~w393 & ~w2117) | (~w393 & w1482) | (~w2117 & w1482);
assign w847 = ~w751 & w283;
assign w848 = (~w1518 & w1043) | (~w1518 & w1531) | (w1043 & w1531);
assign w849 = ~w2063 & ~w1550;
assign w850 = w691 & ~w2142;
assign w851 = ~w877 & ~w1486;
assign w852 = ~pi135 & ~w272;
assign w853 = ~w1771 & ~w1208;
assign w854 = (w1313 & w941) | (w1313 & w1959) | (w941 & w1959);
assign w855 = (~w1890 & ~w985) | (~w1890 & w536) | (~w985 & w536);
assign w856 = ~pi002 & ~pi066;
assign w857 = pi003 & pi067;
assign w858 = ~w539 & ~w353;
assign w859 = w1868 & w818;
assign w860 = ~w2037 & w131;
assign w861 = ~w1684 & ~w293;
assign w862 = ~w849 & w277;
assign w863 = (w1652 & ~w307) | (w1652 & ~w2064) | (~w307 & ~w2064);
assign w864 = pi180 & w592;
assign w865 = (~w88 & w439) | (~w88 & w480) | (w439 & w480);
assign w866 = (~w1680 & ~w2051) | (~w1680 & w1977) | (~w2051 & w1977);
assign w867 = ~w2148 & ~w1088;
assign w868 = ~w769 & ~w2176;
assign w869 = (w489 & w799) | (w489 & w965) | (w799 & w965);
assign w870 = (w1502 & w182) | (w1502 & w1552) | (w182 & w1552);
assign w871 = (w1368 & w795) | (w1368 & w6) | (w795 & w6);
assign w872 = ~w2099 & ~w1058;
assign w873 = (w1417 & w347) | (w1417 & w1118) | (w347 & w1118);
assign w874 = ~w1985 & ~w462;
assign w875 = (~w211 & ~w607) | (~w211 & w1854) | (~w607 & w1854);
assign w876 = ~w833 & ~w47;
assign w877 = ~w981 & ~w1374;
assign w878 = pi218 & ~w1990;
assign w879 = w809 & ~w1871;
assign w880 = (w1423 & w1196) | (w1423 & w916) | (w1196 & w916);
assign w881 = (w1538 & w1407) | (w1538 & w1510) | (w1407 & w1510);
assign w882 = (~w2076 & w2080) | (~w2076 & w295) | (w2080 & w295);
assign w883 = (~w1989 & ~w1054) | (~w1989 & w1241) | (~w1054 & w1241);
assign w884 = w376 & ~w947;
assign w885 = pi140 & w694;
assign w886 = (w1303 & w913) | (w1303 & ~w1402) | (w913 & ~w1402);
assign w887 = ~w1769 & ~w332;
assign w888 = (~w316 & w1809) | (~w316 & w738) | (w1809 & w738);
assign w889 = ~w1151 & ~w335;
assign w890 = ~w1702 & ~w1949;
assign w891 = ~w1722 & ~w1258;
assign w892 = (w1696 & w1144) | (w1696 & w644) | (w1144 & w644);
assign w893 = ~pi246 & w1083;
assign w894 = (~w368 & w1898) | (~w368 & w333) | (w1898 & w333);
assign w895 = (~w2035 & ~w437) | (~w2035 & w1770) | (~w437 & w1770);
assign w896 = w385 & ~w741;
assign w897 = ~pi028 & ~pi092;
assign w898 = pi029 & pi093;
assign w899 = pi217 & ~w2106;
assign w900 = pi224 & ~w927;
assign w901 = (w1425 & w983) | (w1425 & w1177) | (w983 & w1177);
assign w902 = (w1870 & w844) | (w1870 & w1676) | (w844 & w1676);
assign w903 = (w466 & w184) | (w466 & w1602) | (w184 & w1602);
assign w904 = (w748 & w441) | (w748 & w613) | (w441 & w613);
assign w905 = ~w1711 & ~w1705;
assign w906 = w2138 & w1786;
assign w907 = w2050 & ~w2198;
assign w908 = ~w353 & ~w746;
assign w909 = (w1518 & w831) | (w1518 & w718) | (w831 & w718);
assign w910 = ~w62 & w1133;
assign w911 = (~w1880 & ~w737) | (~w1880 & w569) | (~w737 & w569);
assign w912 = (w980 & w1436) | (w980 & w1698) | (w1436 & w1698);
assign w913 = ~w253 & w480;
assign w914 = ~w1118 & w1768;
assign w915 = (~w792 & w1530) | (~w792 & w2144) | (w1530 & w2144);
assign w916 = ~w468 & ~w265;
assign w917 = w855 & ~w1505;
assign w918 = ~w1249 & ~w1932;
assign w919 = ~pi151 & ~w261;
assign w920 = ~w1901 & ~w1968;
assign w921 = (~w1502 & w1126) | (~w1502 & w1421) | (w1126 & w1421);
assign w922 = w751 & ~w283;
assign w923 = (w675 & w356) | (w675 & w449) | (w356 & w449);
assign w924 = ~w1786 & ~w1517;
assign w925 = pi212 & ~w1660;
assign w926 = ~w479 & ~w995;
assign w927 = (~w2136 & ~w213) | (~w2136 & w1038) | (~w213 & w1038);
assign w928 = ~w1610 & ~w1236;
assign w929 = ~pi185 & ~w817;
assign w930 = w429 & ~w705;
assign w931 = ~w1045 & ~w1524;
assign w932 = ~w401 & ~w1264;
assign w933 = (~w1943 & w1198) | (~w1943 & w1420) | (w1198 & w1420);
assign w934 = ~w116 & ~w1921;
assign w935 = ~w1756 & ~w1884;
assign w936 = (w1953 & w707) | (w1953 & w1192) | (w707 & w1192);
assign w937 = (w1502 & w992) | (w1502 & w977) | (w992 & w977);
assign w938 = ~w1097 & ~w1838;
assign w939 = ~w1720 & ~w1543;
assign w940 = ~w1663 & ~w752;
assign w941 = ~w107 & ~w417;
assign w942 = ~w14 & ~w758;
assign w943 = w733 & w1701;
assign w944 = (w277 & w2189) | (w277 & w862) | (w2189 & w862);
assign w945 = (w1100 & w753) | (w1100 & w1375) | (w753 & w1375);
assign w946 = w838 & ~w1726;
assign w947 = ~w129 & ~w1711;
assign w948 = (~w1180 & w1189) | (~w1180 & w1822) | (w1189 & w1822);
assign w949 = (~w235 & ~w30) | (~w235 & w589) | (~w30 & w589);
assign w950 = pi168 & w357;
assign w951 = ~w1105 & ~w1448;
assign w952 = (~w980 & w848) | (~w980 & w2155) | (w848 & w2155);
assign w953 = ~w766 & w1028;
assign w954 = (w466 & w184) | (w466 & w610) | (w184 & w610);
assign w955 = ~w489 & ~w1513;
assign w956 = ~pi035 & ~pi099;
assign w957 = pi036 & pi100;
assign w958 = ~pi165 & ~w1566;
assign w959 = ~w414 & ~w210;
assign w960 = (w1416 & w1919) | (w1416 & w873) | (w1919 & w873);
assign w961 = pi157 & w373;
assign w962 = (~w1953 & w886) | (~w1953 & w664) | (w886 & w664);
assign w963 = ~w1438 & w4;
assign w964 = (~w1789 & ~w1583) | (~w1789 & w55) | (~w1583 & w55);
assign w965 = w1844 & ~w43;
assign w966 = ~w1156 & ~w1274;
assign w967 = (w2208 & w1832) | (w2208 & w706) | (w1832 & w706);
assign w968 = (~w496 & ~w3) | (~w496 & w1529) | (~w3 & w1529);
assign w969 = ~w908 & ~w539;
assign w970 = pi131 & w1842;
assign w971 = ~w376 & w2195;
assign w972 = (w1927 & w1177) | (w1927 & w1876) | (w1177 & w1876);
assign w973 = ~pi007 & ~pi071;
assign w974 = pi008 & pi072;
assign w975 = (w1971 & w595) | (w1971 & w259) | (w595 & w259);
assign w976 = (~w1968 & w1604) | (~w1968 & w920) | (w1604 & w920);
assign w977 = (~w980 & w1678) | (~w980 & w2016) | (w1678 & w2016);
assign w978 = pi142 & w176;
assign w979 = ~w1191 & ~w284;
assign w980 = (~w2163 & w1530) | (~w2163 & w2144) | (w1530 & w2144);
assign w981 = pi254 & ~w1222;
assign w982 = (w489 & w1329) | (w489 & w1253) | (w1329 & w1253);
assign w983 = w1705 & w1425;
assign w984 = (~w1007 & ~w448) | (~w1007 & w1160) | (~w448 & w1160);
assign w985 = ~w1890 & ~w2161;
assign w986 = (~w882 & w791) | (~w882 & w1730) | (w791 & w1730);
assign w987 = ~w477 & ~w2053;
assign w988 = w2156 & ~w305;
assign w989 = (w1108 & w461) | (w1108 & w1214) | (w461 & w1214);
assign w990 = ~w2204 & ~w199;
assign w991 = ~w1502 & w188;
assign w992 = (~w1870 & w1328) | (~w1870 & w1251) | (w1328 & w1251);
assign w993 = w838 & w687;
assign w994 = ~w1868 & ~w1055;
assign w995 = pi247 & ~w1816;
assign w996 = (w1070 & w1345) | (w1070 & w172) | (w1345 & w172);
assign w997 = (~w1502 & w1729) | (~w1502 & w498) | (w1729 & w498);
assign w998 = (w326 & w2020) | (w326 & w1966) | (w2020 & w1966);
assign w999 = ~w833 & ~w2208;
assign w1000 = ~pi148 & ~w159;
assign w1001 = ~w621 & ~w1742;
assign w1002 = (~w606 & ~w9) | (~w606 & w1378) | (~w9 & w1378);
assign w1003 = (~w416 & w136) | (~w416 & w603) | (w136 & w603);
assign w1004 = ~pi183 & ~w561;
assign w1005 = ~pi047 & ~pi111;
assign w1006 = pi048 & pi112;
assign w1007 = pi249 & ~w1671;
assign w1008 = (~w486 & ~w2078) | (~w486 & w2031) | (~w2078 & w2031);
assign w1009 = w651 & ~w1718;
assign w1010 = ~w1539 & ~w2208;
assign w1011 = ~w985 & ~w695;
assign w1012 = ~w481 & ~w1417;
assign w1013 = w651 & w1606;
assign w1014 = pi162 & w602;
assign w1015 = (~w521 & ~w600) | (~w521 & w1308) | (~w600 & w1308);
assign w1016 = ~w1814 & ~w325;
assign w1017 = w1714 & ~w990;
assign w1018 = (~w2120 & w2189) | (~w2120 & w1635) | (w2189 & w1635);
assign w1019 = (w1715 & w1426) | (w1715 & w1858) | (w1426 & w1858);
assign w1020 = ~pi217 & w2106;
assign w1021 = (w1502 & w882) | (w1502 & w1927) | (w882 & w1927);
assign w1022 = (w1502 & w1946) | (w1502 & w499) | (w1946 & w499);
assign w1023 = ~pi240 & w797;
assign w1024 = w2050 & ~w1602;
assign w1025 = w2028 & ~w1845;
assign w1026 = ~w887 & ~w1283;
assign w1027 = (~w1218 & ~w502) | (~w1218 & w781) | (~w502 & w781);
assign w1028 = ~w1336 & ~w2011;
assign w1029 = ~pi172 & ~w81;
assign w1030 = (~w1927 & w524) | (~w1927 & w699) | (w524 & w699);
assign w1031 = ~w629 & w745;
assign w1032 = pi176 & w45;
assign w1033 = ~w2037 & ~w1650;
assign w1034 = ~pi057 & ~pi121;
assign w1035 = pi058 & pi122;
assign w1036 = ~w64 & ~w789;
assign w1037 = ~w584 & ~w1988;
assign w1038 = ~pi159 & ~w2136;
assign w1039 = ~w375 & ~w31;
assign w1040 = w651 & ~w595;
assign w1041 = ~w2094 & ~w1652;
assign w1042 = pi000 & pi064;
assign w1043 = (~w204 & w1504) | (~w204 & w1472) | (w1504 & w1472);
assign w1044 = ~pi158 & ~w737;
assign w1045 = ~w1873 & w611;
assign w1046 = ~pi155 & ~w517;
assign w1047 = (~w1927 & w75) | (~w1927 & w140) | (w75 & w140);
assign w1048 = (~w899 & ~w1568) | (~w899 & w1306) | (~w1568 & w1306);
assign w1049 = w1010 & ~w405;
assign w1050 = ~w417 & ~w17;
assign w1051 = ~pi252 & w483;
assign w1052 = pi201 & ~w222;
assign w1053 = ~w476 & ~w1316;
assign w1054 = ~w1989 & ~w473;
assign w1055 = ~w379 & w537;
assign w1056 = ~w282 & ~w390;
assign w1057 = ~w2137 & w1161;
assign w1058 = w544 & w1632;
assign w1059 = (~w326 & w1049) | (~w326 & w378) | (w1049 & w378);
assign w1060 = ~w1473 & ~w79;
assign w1061 = w1801 & w1528;
assign w1062 = w1917 & w747;
assign w1063 = w471 & ~w1253;
assign w1064 = (w740 & w1312) | (w740 & ~w2198) | (w1312 & ~w2198);
assign w1065 = (~w6 & w1203) | (~w6 & w716) | (w1203 & w716);
assign w1066 = (~w1715 & w812) | (~w1715 & w1130) | (w812 & w1130);
assign w1067 = ~w849 & w1677;
assign w1068 = w1008 & ~w1495;
assign w1069 = (w1905 & w1502) | (w1905 & w1331) | (w1502 & w1331);
assign w1070 = ~w1181 & w1179;
assign w1071 = ~w928 & ~w1610;
assign w1072 = ~w1514 & ~w2072;
assign w1073 = ~pi198 & w2194;
assign w1074 = ~w1129 & ~w757;
assign w1075 = ~pi179 & ~w297;
assign w1076 = w1965 & w1947;
assign w1077 = ~w1720 & ~w801;
assign w1078 = ~w1557 & ~w38;
assign w1079 = ~pi132 & ~w762;
assign w1080 = (w960 & w304) | (w960 & w1533) | (w304 & w1533);
assign w1081 = (w948 & w1878) | (w948 & w2118) | (w1878 & w2118);
assign w1082 = ~w1845 & ~w1206;
assign w1083 = (~w1318 & ~w1452) | (~w1318 & w682) | (~w1452 & w682);
assign w1084 = w1561 & w1557;
assign w1085 = w2143 & w1875;
assign w1086 = w267 & ~w1818;
assign w1087 = w1806 & ~w756;
assign w1088 = ~w1523 & ~w1110;
assign w1089 = (w980 & w151) | (w980 & w576) | (w151 & w576);
assign w1090 = ~w532 & ~w1774;
assign w1091 = ~w667 & ~w1445;
assign w1092 = w1569 & ~w65;
assign w1093 = ~w1720 & w56;
assign w1094 = ~w1474 & ~w2091;
assign w1095 = (~w2028 & w2029) | (~w2028 & w1234) | (w2029 & w1234);
assign w1096 = pi190 & w30;
assign w1097 = (~w1680 & w416) | (~w1680 & w326) | (w416 & w326);
assign w1098 = (w162 & w1133) | (w162 & w557) | (w1133 & w557);
assign w1099 = ~w1569 & w1596;
assign w1100 = w849 & ~w2189;
assign w1101 = ~pi136 & ~w0;
assign w1102 = (~w1705 & w384) | (~w1705 & w1800) | (w384 & w1800);
assign w1103 = ~w365 & ~w78;
assign w1104 = ~w1568 & ~w1409;
assign w1105 = pi170 & w2150;
assign w1106 = ~w448 & ~w469;
assign w1107 = w187 & ~w1819;
assign w1108 = (w1652 & ~w307) | (w1652 & ~w1268) | (~w307 & ~w1268);
assign w1109 = (~w1295 & ~w253) | (~w1295 & w153) | (~w253 & w153);
assign w1110 = ~pi175 & ~w2103;
assign w1111 = ~w1026 & ~w509;
assign w1112 = (w1010 & w2211) | (w1010 & ~w1108) | (w2211 & ~w1108);
assign w1113 = ~w1450 & ~w70;
assign w1114 = (w863 & w627) | (w863 & w2069) | (w627 & w2069);
assign w1115 = (~w368 & w571) | (~w368 & w333) | (w571 & w333);
assign w1116 = ~pi203 & w1625;
assign w1117 = ~w1072 & ~w2092;
assign w1118 = ~w481 & ~w58;
assign w1119 = ~w1136 & w1673;
assign w1120 = ~w503 & w8;
assign w1121 = w1578 & w2067;
assign w1122 = ~w2138 & ~w1786;
assign w1123 = ~w385 & w678;
assign w1124 = pi192 & w1903;
assign w1125 = w129 & ~w1102;
assign w1126 = (w1924 & w2153) | (w1924 & w1715) | (w2153 & w1715);
assign w1127 = (~w674 & ~w60) | (~w674 & w218) | (~w60 & w218);
assign w1128 = ~w579 & ~w1190;
assign w1129 = ~w207 & ~w1888;
assign w1130 = (w396 & w1556) | (w396 & w2163) | (w1556 & w2163);
assign w1131 = ~w1917 & ~w747;
assign w1132 = ~pi236 & w1749;
assign w1133 = (~w1610 & w322) | (~w1610 & w1071) | (w322 & w1071);
assign w1134 = ~w1286 & ~w10;
assign w1135 = pi137 & w266;
assign w1136 = ~w330 & ~w123;
assign w1137 = ~w1864 & ~w1519;
assign w1138 = ~w666 & ~w1537;
assign w1139 = (w1942 & w726) | (w1942 & w262) | (w726 & w262);
assign w1140 = ~pi241 & w1542;
assign w1141 = w2175 & ~w711;
assign w1142 = ~w1352 & ~w121;
assign w1143 = w2116 & ~w1767;
assign w1144 = ~w651 & w595;
assign w1145 = w448 & w469;
assign w1146 = ~pi157 & ~w898;
assign w1147 = ~w1522 & w1659;
assign w1148 = ~w651 & ~w1606;
assign w1149 = ~w1302 & ~w1624;
assign w1150 = (w56 & w427) | (w56 & w1889) | (w427 & w1889);
assign w1151 = ~w1470 & w1388;
assign w1152 = (~w507 & w1179) | (~w507 & w318) | (w1179 & w318);
assign w1153 = ~w1725 & ~w234;
assign w1154 = ~w2123 & ~w667;
assign w1155 = ~pi045 & ~pi109;
assign w1156 = pi046 & pi110;
assign w1157 = ~w2174 & ~w803;
assign w1158 = (~w1962 & ~w86) | (~w1962 & w839) | (~w86 & w839);
assign w1159 = (~w882 & w1492) | (~w882 & w457) | (w1492 & w457);
assign w1160 = ~w469 & ~w1007;
assign w1161 = ~w1757 & ~w220;
assign w1162 = (w1115 & w894) | (w1115 & ~w1748) | (w894 & ~w1748);
assign w1163 = w253 & ~w480;
assign w1164 = ~w1118 & ~w931;
assign w1165 = ~w1411 & ~w1507;
assign w1166 = ~w1347 & ~w229;
assign w1167 = ~w47 & ~w2208;
assign w1168 = ~w62 & w1071;
assign w1169 = (~w1797 & ~w1654) | (~w1797 & w1422) | (~w1654 & w1422);
assign w1170 = ~w1319 & ~w1281;
assign w1171 = ~w1995 & ~w1935;
assign w1172 = ~w1050 & w2076;
assign w1173 = (~w285 & ~w261) | (~w285 & w1853) | (~w261 & w1853);
assign w1174 = (~w2120 & w1598) | (~w2120 & w506) | (w1598 & w506);
assign w1175 = (~w6 & w2111) | (~w6 & w61) | (w2111 & w61);
assign w1176 = ~pi230 & w564;
assign w1177 = w15 & ~w384;
assign w1178 = ~w2063 & ~w260;
assign w1179 = (~w1256 & ~w2168) | (~w1256 & w269) | (~w2168 & w269);
assign w1180 = (~w435 & w1806) | (~w435 & w1444) | (w1806 & w1444);
assign w1181 = ~w507 & ~w2119;
assign w1182 = (w135 & w645) | (w135 & w416) | (w645 & w416);
assign w1183 = w1569 & w484;
assign w1184 = (w2028 & w1195) | (w2028 & w923) | (w1195 & w923);
assign w1185 = (~w882 & w1677) | (~w882 & w1102) | (w1677 & w1102);
assign w1186 = (w1533 & w574) | (w1533 & w2163) | (w574 & w2163);
assign w1187 = (~w1261 & ~w260) | (~w1261 & w277) | (~w260 & w277);
assign w1188 = (~w1156 & ~w966) | (~w1156 & w113) | (~w966 & w113);
assign w1189 = w1438 & w1120;
assign w1190 = ~pi021 & ~pi085;
assign w1191 = pi022 & pi086;
assign w1192 = (w2170 & w787) | (w2170 & w262) | (w787 & w262);
assign w1193 = (w1012 & w835) | (w1012 & w1768) | (w835 & w1768);
assign w1194 = pi189 & w1153;
assign w1195 = (w1980 & w356) | (w1980 & w449) | (w356 & w449);
assign w1196 = (~w1968 & w920) | (~w1968 & ~w1555) | (w920 & ~w1555);
assign w1197 = pi229 & ~w100;
assign w1198 = w275 & w1295;
assign w1199 = ~pi153 & ~w414;
assign w1200 = w275 & ~w1109;
assign w1201 = (~w1502 & w1958) | (~w1502 & w1908) | (w1958 & w1908);
assign w1202 = w494 & w2000;
assign w1203 = ~w1649 & ~w2062;
assign w1204 = (~w65 & ~w1596) | (~w65 & ~w1819) | (~w1596 & ~w1819);
assign w1205 = (~w2002 & ~w832) | (~w2002 & w836) | (~w832 & w836);
assign w1206 = ~w1521 & w2182;
assign w1207 = (~w326 & w216) | (~w326 & w1779) | (w216 & w1779);
assign w1208 = w422 & w773;
assign w1209 = pi166 & w526;
assign w1210 = ~w2168 & ~w1256;
assign w1211 = ~w85 & ~w1116;
assign w1212 = w376 & w1711;
assign w1213 = (w681 & w1835) | (w681 & w1237) | (w1835 & w1237);
assign w1214 = w833 & w1885;
assign w1215 = ~pi042 & ~pi106;
assign w1216 = pi043 & pi107;
assign w1217 = (w287 & w438) | (w287 & w1185) | (w438 & w1185);
assign w1218 = pi232 & ~w1467;
assign w1219 = pi169 & w1654;
assign w1220 = ~w951 & ~w659;
assign w1221 = (w1711 & ~w947) | (w1711 & w792) | (~w947 & w792);
assign w1222 = (~w1725 & ~w1153) | (~w1725 & w418) | (~w1153 & w418);
assign w1223 = ~w1180 & w69;
assign w1224 = ~w597 & ~w1377;
assign w1225 = ~w832 & ~w782;
assign w1226 = ~pi160 & ~w1493;
assign w1227 = (w1927 & w1125) | (w1927 & w2013) | (w1125 & w2013);
assign w1228 = w1389 & w702;
assign w1229 = ~w2120 & w162;
assign w1230 = w2006 & ~w247;
assign w1231 = pi172 & w81;
assign w1232 = ~w1106 & ~w1145;
assign w1233 = ~pi191 & w891;
assign w1234 = w2115 & ~w1082;
assign w1235 = ~w489 & w2104;
assign w1236 = w655 & ~w1232;
assign w1237 = w62 & ~w1133;
assign w1238 = (~w865 & w1198) | (~w865 & w1420) | (w1198 & w1420);
assign w1239 = ~w937 & ~w618;
assign w1240 = (~w1187 & ~w74) | (~w1187 & w231) | (~w74 & w231);
assign w1241 = ~pi145 & ~w1989;
assign w1242 = (w1502 & w2164) | (w1502 & w2186) | (w2164 & w2186);
assign w1243 = w9 & w1171;
assign w1244 = ~w1844 & ~w1555;
assign w1245 = ~pi193 & w1685;
assign w1246 = (~w1191 & ~w979) | (~w1191 & w1353) | (~w979 & w1353);
assign w1247 = (w865 & w84) | (w865 & w2083) | (w84 & w2083);
assign w1248 = (~w326 & w603) | (~w326 & w136) | (w603 & w136);
assign w1249 = ~w1027 & w1613;
assign w1250 = (w1715 & w915) | (w1715 & w980) | (w915 & w980);
assign w1251 = (w1237 & w681) | (w1237 & w1835) | (w681 & w1835);
assign w1252 = (w137 & w252) | (w137 & w1085) | (w252 & w1085);
assign w1253 = (~w43 & w540) | (~w43 & w1834) | (w540 & w1834);
assign w1254 = (w1329 & w1394) | (w1329 & w1925) | (w1394 & w1925);
assign w1255 = pi128 & w700;
assign w1256 = ~w1862 & w1440;
assign w1257 = ~pi062 & ~pi126;
assign w1258 = pi063 & pi127;
assign w1259 = ~w425 & ~w1892;
assign w1260 = w665 & ~w1584;
assign w1261 = ~w968 & w853;
assign w1262 = (w1602 & w2198) | (w1602 & ~w915) | (w2198 & ~w915);
assign w1263 = ~pi166 & ~w1469;
assign w1264 = (~w948 & w2036) | (~w948 & w570) | (w2036 & w570);
assign w1265 = (~w571 & ~w1898) | (~w571 & w748) | (~w1898 & w748);
assign w1266 = pi165 & w1727;
assign w1267 = (w882 & w1615) | (w882 & w1849) | (w1615 & w1849);
assign w1268 = (~w811 & w122) | (~w811 & w273) | (w122 & w273);
assign w1269 = ~w1560 & ~w1790;
assign w1270 = (~w1502 & w195) | (~w1502 & w1089) | (w195 & w1089);
assign w1271 = (w1368 & w795) | (w1368 & w1976) | (w795 & w1976);
assign w1272 = (~w585 & w1785) | (~w585 & w1423) | (w1785 & w1423);
assign w1273 = ~w1118 & w1960;
assign w1274 = ~pi046 & ~pi110;
assign w1275 = pi047 & pi111;
assign w1276 = w379 & ~w537;
assign w1277 = ~w2197 & ~w342;
assign w1278 = w548 & ~w20;
assign w1279 = (~w341 & ~w357) | (~w341 & w1642) | (~w357 & w1642);
assign w1280 = ~w1242 & ~w636;
assign w1281 = pi214 & ~w1781;
assign w1282 = ~w183 & ~w95;
assign w1283 = ~w103 & ~w1044;
assign w1284 = (w513 & w876) | (w513 & w999) | (w876 & w999);
assign w1285 = ~w110 & ~w90;
assign w1286 = ~w1546 & w605;
assign w1287 = (w173 & w730) | (w173 & ~w231) | (w730 & ~w231);
assign w1288 = ~w342 & ~w190;
assign w1289 = ~w1713 & ~w1053;
assign w1290 = (~w272 & ~w1419) | (~w272 & w852) | (~w1419 & w852);
assign w1291 = (~w1980 & w558) | (~w1980 & w946) | (w558 & w946);
assign w1292 = pi164 & w693;
assign w1293 = (w436 & ~w1265) | (w436 & ~w948) | (~w1265 & ~w948);
assign w1294 = ~w1742 & ~w1708;
assign w1295 = ~w2006 & w247;
assign w1296 = ~w1768 & ~w1960;
assign w1297 = ~w1947 & ~w1494;
assign w1298 = w320 & ~w388;
assign w1299 = (~w925 & ~w804) | (~w925 & w115) | (~w804 & w115);
assign w1300 = pi181 & w1452;
assign w1301 = ~w642 & ~w1709;
assign w1302 = pi130 & w671;
assign w1303 = ~w253 & ~w88;
assign w1304 = (~w900 & ~w206) | (~w900 & w796) | (~w206 & w796);
assign w1305 = (w2051 & w860) | (w2051 & w13) | (w860 & w13);
assign w1306 = ~w1409 & ~w899;
assign w1307 = w1136 & ~w1673;
assign w1308 = ~pi141 & ~w521;
assign w1309 = pi148 & w159;
assign w1310 = ~w751 & w1857;
assign w1311 = (w644 & w1605) | (w644 & w491) | (w1605 & w491);
assign w1312 = ~w1950 & w823;
assign w1313 = (~w330 & w1673) | (~w330 & w44) | (w1673 & w44);
assign w1314 = (w975 & w1403) | (w975 & w1939) | (w1403 & w1939);
assign w1315 = ~w2141 & ~w956;
assign w1316 = ~pi141 & ~w600;
assign w1317 = ~pi052 & ~pi116;
assign w1318 = pi053 & pi117;
assign w1319 = ~w1455 & ~w810;
assign w1320 = (~w1031 & w1082) | (~w1031 & w2041) | (w1082 & w2041);
assign w1321 = (~w474 & ~w1589) | (~w474 & w1639) | (~w1589 & w1639);
assign w1322 = ~w870 & ~w1628;
assign w1323 = w697 & w1692;
assign w1324 = ~pi152 & ~w1633;
assign w1325 = ~w368 & ~w1086;
assign w1326 = ~w928 & ~w1705;
assign w1327 = pi143 & w32;
assign w1328 = (w2120 & w681) | (w2120 & w1835) | (w681 & w1835);
assign w1329 = (~w976 & w540) | (~w976 & w1834) | (w540 & w1834);
assign w1330 = (w1939 & w765) | (w1939 & w1099) | (w765 & w1099);
assign w1331 = w1249 & w1905;
assign w1332 = w1269 & ~w318;
assign w1333 = ~w226 & ~w709;
assign w1334 = (~w1152 & w1296) | (~w1152 & w1416) | (w1296 & w1416);
assign w1335 = ~pi154 & ~w607;
assign w1336 = ~w1570 & ~w1453;
assign w1337 = (~w948 & w53) | (~w948 & w452) | (w53 & w452);
assign w1338 = ~w502 & ~w663;
assign w1339 = w1434 & ~w1918;
assign w1340 = w1823 & w2098;
assign w1341 = (w818 & w859) | (w818 & w326) | (w859 & w326);
assign w1342 = ~w813 & ~w2045;
assign w1343 = (w1502 & w202) | (w1502 & w1267) | (w202 & w1267);
assign w1344 = ~w1118 & ~w1045;
assign w1345 = (~w1256 & ~w2183) | (~w1256 & w1210) | (~w2183 & w1210);
assign w1346 = ~pi010 & ~pi074;
assign w1347 = pi011 & pi075;
assign w1348 = (w1927 & w191) | (w1927 & w1525) | (w191 & w1525);
assign w1349 = w1856 & ~w326;
assign w1350 = ~w833 & w1167;
assign w1351 = ~w1430 & ~w340;
assign w1352 = w1756 & w1667;
assign w1353 = ~pi150 & ~w1191;
assign w1354 = (~w1152 & w1883) | (~w1152 & w1783) | (w1883 & w1783);
assign w1355 = (w1680 & w1574) | (w1680 & w643) | (w1574 & w643);
assign w1356 = ~w1285 & ~w2167;
assign w1357 = ~pi132 & ~w582;
assign w1358 = ~w1828 & ~w467;
assign w1359 = (w98 & w2162) | (w98 & ~w1253) | (w2162 & ~w1253);
assign w1360 = ~w1032 & ~w1367;
assign w1361 = ~w268 & ~w167;
assign w1362 = ~w360 & ~w1644;
assign w1363 = ~w1360 & ~w1700;
assign w1364 = (~w2089 & ~w1710) | (~w2089 & w653) | (~w1710 & w653);
assign w1365 = (~w425 & ~w1259) | (~w425 & w411) | (~w1259 & w411);
assign w1366 = pi145 & w1054;
assign w1367 = ~pi176 & ~w45;
assign w1368 = w1649 & w2062;
assign w1369 = (w1680 & w892) | (w1680 & w690) | (w892 & w690);
assign w1370 = ~pi234 & w1169;
assign w1371 = pi253 & ~w2097;
assign w1372 = w186 & w479;
assign w1373 = ~w376 & ~w767;
assign w1374 = ~pi254 & w1222;
assign w1375 = w1747 & ~w74;
assign w1376 = ~pi156 & ~w2033;
assign w1377 = (~w1502 & w1766) | (~w1502 & w1983) | (w1766 & w1983);
assign w1378 = ~w1171 & ~w606;
assign w1379 = (w236 & w760) | (w236 & w1185) | (w760 & w1185);
assign w1380 = ~w2037 & ~w808;
assign w1381 = ~w1356 & ~w1690;
assign w1382 = ~w390 & ~w243;
assign w1383 = ~w1780 & ~w1184;
assign w1384 = w2197 & w342;
assign w1385 = (w1711 & ~w947) | (w1711 & ~w270) | (~w947 & ~w270);
assign w1386 = ~w2156 & w305;
assign w1387 = ~w928 & w322;
assign w1388 = ~w851 & ~w1424;
assign w1389 = ~w301 & ~w1833;
assign w1390 = (~w313 & ~w697) | (~w313 & w1594) | (~w697 & w1594);
assign w1391 = (~w1502 & w744) | (~w1502 & w1379) | (w744 & w1379);
assign w1392 = pi159 & w213;
assign w1393 = (~w1819 & ~w2088) | (~w1819 & w751) | (~w2088 & w751);
assign w1394 = w253 & ~w1943;
assign w1395 = ~w1680 & w217;
assign w1396 = ~pi178 & ~w86;
assign w1397 = ~w691 & w2142;
assign w1398 = ~pi156 & ~w1813;
assign w1399 = ~w2023 & ~w1647;
assign w1400 = (~w1250 & w725) | (~w1250 & w703) | (w725 & w703);
assign w1401 = ~w1607 & ~w1410;
assign w1402 = (~w439 & ~w1636) | (~w439 & w262) | (~w1636 & w262);
assign w1403 = ~w1538 & w1971;
assign w1404 = ~w1050 & ~w417;
assign w1405 = ~w672 & ~w2079;
assign w1406 = ~w1124 & ~w1614;
assign w1407 = w2037 & ~w450;
assign w1408 = (w1502 & w201) | (w1502 & w1651) | (w201 & w1651);
assign w1409 = ~w1695 & ~w841;
assign w1410 = pi250 & ~w673;
assign w1411 = pi129 & w2117;
assign w1412 = (w137 & w1572) | (w137 & w1674) | (w1572 & w1674);
assign w1413 = (w2168 & w2183) | (w2168 & w2130) | (w2183 & w2130);
assign w1414 = ~w1632 & ~w309;
assign w1415 = ~w51 & ~w148;
assign w1416 = (~w1960 & ~w1768) | (~w1960 & w1269) | (~w1768 & w1269);
assign w1417 = ~w840 & ~w661;
assign w1418 = ~w1395 & ~w101;
assign w1419 = ~w272 & ~w973;
assign w1420 = w275 & ~w1762;
assign w1421 = (w1924 & w2153) | (w1924 & w1185) | (w2153 & w1185);
assign w1422 = ~pi169 & ~w1797;
assign w1423 = (~w1968 & ~w1901) | (~w1968 & w657) | (~w1901 & w657);
assign w1424 = w877 & w1486;
assign w1425 = ~w2126 & ~w1017;
assign w1426 = (~w792 & w914) | (~w792 & w1273) | (w914 & w1273);
assign w1427 = ~w948 & ~w193;
assign w1428 = (~w416 & w790) | (~w416 & w306) | (w790 & w306);
assign w1429 = ~pi038 & ~pi102;
assign w1430 = pi039 & pi103;
assign w1431 = ~w1277 & ~w1384;
assign w1432 = w1496 & w656;
assign w1433 = (~w980 & w1520) | (~w980 & w248) | (w1520 & w248);
assign w1434 = (~w981 & ~w877) | (~w981 & w1869) | (~w877 & w1869);
assign w1435 = w1912 & ~w882;
assign w1436 = (w1018 & w1954) | (w1018 & w844) | (w1954 & w844);
assign w1437 = ~w987 & ~w2133;
assign w1438 = ~w1057 & ~w346;
assign w1439 = (~w1502 & w820) | (~w1502 & w854) | (w820 & w854);
assign w1440 = ~w189 & ~w99;
assign w1441 = ~w619 & ~w1355;
assign w1442 = (w1098 & w1229) | (w1098 & w1715) | (w1229 & w1715);
assign w1443 = ~w208 & w1597;
assign w1444 = ~w756 & ~w435;
assign w1445 = ~pi225 & w395;
assign w1446 = pi133 & w76;
assign w1447 = ~w2143 & ~w1942;
assign w1448 = ~pi170 & ~w2150;
assign w1449 = (~w763 & ~w494) | (~w763 & w764) | (~w494 & w764);
assign w1450 = (w489 & w1252) | (w489 & w936) | (w1252 & w936);
assign w1451 = (~w2028 & w879) | (~w2028 & w1662) | (w879 & w1662);
assign w1452 = ~w1318 & ~w453;
assign w1453 = ~w830 & ~w16;
assign w1454 = ~w335 & ~w1950;
assign w1455 = pi150 & w979;
assign w1456 = ~w809 & ~w1974;
assign w1457 = ~w1844 & w1423;
assign w1458 = ~w1764 & w755;
assign w1459 = (~w244 & ~w398) | (~w244 & w1881) | (~w398 & w1881);
assign w1460 = ~w559 & ~w1994;
assign w1461 = ~w1216 & ~w168;
assign w1462 = (w1680 & w1475) | (w1680 & w1349) | (w1475 & w1349);
assign w1463 = ~w1600 & ~w1961;
assign w1464 = (~w535 & ~w671) | (~w535 & w2178) | (~w671 & w2178);
assign w1465 = ~w2071 & ~w1025;
assign w1466 = ~w1124 & ~w1060;
assign w1467 = (~w1430 & ~w1351) | (~w1430 & w2152) | (~w1351 & w2152);
assign w1468 = ~pi037 & ~pi101;
assign w1469 = pi038 & pi102;
assign w1470 = (~w1371 & ~w422) | (~w1371 & w2014) | (~w422 & w2014);
assign w1471 = (~w85 & ~w1211) | (~w85 & w250) | (~w1211 & w250);
assign w1472 = w928 & w1705;
assign w1473 = w1920 & w1165;
assign w1474 = ~w177 & ~w1663;
assign w1475 = w1856 & ~w416;
assign w1476 = w1569 & ~w1596;
assign w1477 = ~w1206 & ~w1031;
assign w1478 = (w880 & w415) | (w880 & w649) | (w415 & w649);
assign w1479 = ~w785 & ~w407;
assign w1480 = ~pi140 & ~w230;
assign w1481 = (w1457 & w1666) | (w1457 & w916) | (w1666 & w916);
assign w1482 = ~pi129 & ~w393;
assign w1483 = ~w488 & ~w1201;
assign w1484 = w2050 & ~w610;
assign w1485 = (w873 & w1919) | (w873 & ~w1960) | (w1919 & ~w1960);
assign w1486 = ~w1096 & ~w593;
assign w1487 = pi204 & ~w1987;
assign w1488 = ~w698 & ~w1235;
assign w1489 = (w2074 & w910) | (w2074 & w1185) | (w910 & w1185);
assign w1490 = (w1870 & w120) | (w1870 & w1064) | (w120 & w1064);
assign w1491 = ~w324 & ~w34;
assign w1492 = w1511 & ~w1876;
assign w1493 = ~w2082 & ~w323;
assign w1494 = pi206 & ~w1015;
assign w1495 = ~w2096 & ~w1084;
assign w1496 = ~w71 & ~w1073;
assign w1497 = (w1870 & w1024) | (w1870 & w907) | (w1024 & w907);
assign w1498 = w214 & ~w1381;
assign w1499 = ~w934 & ~w344;
assign w1500 = ~pi235 & w1877;
assign w1501 = pi138 & w1637;
assign w1502 = (~w1680 & w2173) | (~w1680 & w1821) | (w2173 & w1821);
assign w1503 = ~w143 & ~w834;
assign w1504 = w928 & ~w322;
assign w1505 = ~w1891 & ~w1243;
assign w1506 = ~pi229 & w100;
assign w1507 = ~pi129 & ~w2117;
assign w1508 = pi193 & ~w1685;
assign w1509 = w124 & w1399;
assign w1510 = w2037 & ~w131;
assign w1511 = ~w1705 & ~w1425;
assign w1512 = pi134 & w437;
assign w1513 = (w2028 & w1847) | (w2028 & w203) | (w1847 & w203);
assign w1514 = pi242 & ~w1670;
assign w1515 = ~w362 & ~w1773;
assign w1516 = ~w303 & ~w336;
assign w1517 = pi216 & ~w1173;
assign w1518 = (w77 & w384) | (w77 & ~w1927) | (w384 & ~w1927);
assign w1519 = (~w1502 & w793) | (~w1502 & w1737) | (w793 & w1737);
assign w1520 = (w2120 & w1237) | (w2120 & ~w1185) | (w1237 & ~w1185);
assign w1521 = (~w1052 & ~w2174) | (~w1052 & w777) | (~w2174 & w777);
assign w1522 = (~w1769 & ~w887) | (~w1769 & w1860) | (~w887 & w1860);
assign w1523 = pi175 & w2103;
assign w1524 = w1873 & ~w611;
assign w1525 = (~w1677 & w1212) | (~w1677 & w884) | (w1212 & w884);
assign w1526 = (w1329 & w1238) | (w1329 & w933) | (w1238 & w933);
assign w1527 = ~w15 & w384;
assign w1528 = ~w1795 & ~w1278;
assign w1529 = ~w1333 & ~w496;
assign w1530 = (~w396 & w270) | (~w396 & w581) | (w270 & w581);
assign w1531 = (~w204 & w1504) | (~w204 & w1948) | (w1504 & w1948);
assign w1532 = w680 & ~w1876;
assign w1533 = (w507 & ~w318) | (w507 & ~w1345) | (~w318 & ~w1345);
assign w1534 = ~pi172 & ~w169;
assign w1535 = ~w1949 & ~w242;
assign w1536 = pi136 & w0;
assign w1537 = (~w1502 & w543) | (~w1502 & w57) | (w543 & w57);
assign w1538 = (~w1596 & w1013) | (~w1596 & w1009) | (w1013 & w1009);
assign w1539 = ~w2116 & w1767;
assign w1540 = ~w1399 & ~w1831;
assign w1541 = ~w376 & ~w953;
assign w1542 = (~w1006 & ~w45) | (~w1006 & w52) | (~w45 & w52);
assign w1543 = ~w568 & w1653;
assign w1544 = (w1185 & w1858) | (w1185 & w1426) | (w1858 & w1426);
assign w1545 = w129 & ~w915;
assign w1546 = (~w71 & ~w1496) | (~w71 & w2009) | (~w1496 & w2009);
assign w1547 = ~pi008 & ~pi072;
assign w1548 = pi009 & pi073;
assign w1549 = (~w1345 & w646) | (~w1345 & w1739) | (w646 & w1739);
assign w1550 = w1754 & ~w2027;
assign w1551 = w253 & w88;
assign w1552 = (~w1870 & w2070) | (~w1870 & w225) | (w2070 & w225);
assign w1553 = ~pi149 & ~w579;
assign w1554 = ~pi128 & ~w700;
assign w1555 = ~w265 & ~w432;
assign w1556 = w1118 & ~w1768;
assign w1557 = ~w1777 & ~w2090;
assign w1558 = (w416 & w1966) | (w416 & w2020) | (w1966 & w2020);
assign w1559 = (~w1530 & w767) | (~w1530 & w1221) | (w767 & w1221);
assign w1560 = ~w640 & w2100;
assign w1561 = ~w38 & ~w1657;
assign w1562 = ~w196 & w1645;
assign w1563 = ~w275 & w1109;
assign w1564 = (~w324 & ~w1491) | (~w324 & w1765) | (~w1491 & w1765);
assign w1565 = ~pi036 & ~pi100;
assign w1566 = pi037 & pi101;
assign w1567 = w385 & ~w678;
assign w1568 = ~w899 & ~w1020;
assign w1569 = ~w1606 & ~w1611;
assign w1570 = ~w650 & ~w2038;
assign w1571 = (~w489 & w1830) | (~w489 & w962) | (w1830 & w962);
assign w1572 = (w1402 & w1551) | (w1402 & w1163) | (w1551 & w1163);
assign w1573 = w2018 & ~w939;
assign w1574 = ~w751 & w316;
assign w1575 = ~w1569 & ~w484;
assign w1576 = ~pi247 & w1816;
assign w1577 = pi186 & w1750;
assign w1578 = ~w1901 & ~w265;
assign w1579 = w1382 & w282;
assign w1580 = w804 & w311;
assign w1581 = ~w1451 & ~w37;
assign w1582 = ~pi147 & ~w785;
assign w1583 = ~w1789 & ~w1993;
assign w1584 = ~w1338 & ~w1634;
assign w1585 = ~w1167 & ~w608;
assign w1586 = ~w1289 & ~w1612;
assign w1587 = ~w1649 & w1899;
assign w1588 = ~w928 & w1800;
assign w1589 = ~w474 & ~w784;
assign w1590 = ~w275 & w256;
assign w1591 = ~w129 & w1677;
assign w1592 = pi179 & w139;
assign w1593 = w1299 & ~w2105;
assign w1594 = ~w1692 & ~w313;
assign w1595 = ~pi183 & ~w634;
assign w1596 = (~w1147 & w1899) | (~w1147 & w1732) | (w1899 & w1732);
assign w1597 = (~w1055 & ~w818) | (~w1055 & w994) | (~w818 & w994);
assign w1598 = ~w849 & w2189;
assign w1599 = ~pi048 & ~pi112;
assign w1600 = pi049 & pi113;
assign w1601 = ~w1392 & ~w421;
assign w1602 = (w2120 & w652) | (w2120 & w945) | (w652 & w945);
assign w1603 = ~w1269 & ~w507;
assign w1604 = ~w265 & ~w1555;
assign w1605 = w2044 & ~w1538;
assign w1606 = ~w1365 & w2207;
assign w1607 = ~w1577 & ~w1963;
assign w1608 = ~w1709 & ~w1197;
assign w1609 = w751 & w1688;
assign w1610 = ~w655 & w1232;
assign w1611 = w1365 & ~w2207;
assign w1612 = w1713 & w1053;
assign w1613 = ~w1895 & ~w1202;
assign w1614 = ~pi192 & ~w1903;
assign w1615 = (w2131 & w1413) | (w2131 & w1876) | (w1413 & w1876);
assign w1616 = ~pi250 & w673;
assign w1617 = ~pi249 & w1671;
assign w1618 = ~w3 & ~w1333;
assign w1619 = (~w1548 & ~w266) | (~w1548 & w2004) | (~w266 & w2004);
assign w1620 = pi156 & w1813;
assign w1621 = ~w751 & ~w1688;
assign w1622 = w1259 & w1601;
assign w1623 = w1522 & ~w1659;
assign w1624 = ~pi130 & ~w671;
assign w1625 = (~w1741 & ~w1637) | (~w1741 & w1952) | (~w1637 & w1952);
assign w1626 = pi147 & w1479;
assign w1627 = (~w1221 & w1755) | (~w1221 & w1373) | (w1755 & w1373);
assign w1628 = (~w1502 & w2199) | (~w1502 & w1490) | (w2199 & w1490);
assign w1629 = w1027 & ~w1613;
assign w1630 = pi191 & ~w1722;
assign w1631 = (~w1870 & w1602) | (~w1870 & w2198) | (w1602 & w2198);
assign w1632 = ~w497 & ~w108;
assign w1633 = ~w626 & ~w413;
assign w1634 = w502 & w663;
assign w1635 = (~w1795 & ~w1528) | (~w1795 & w794) | (~w1528 & w794);
assign w1636 = ~w312 & ~w1942;
assign w1637 = ~w1741 & ~w1346;
assign w1638 = (~w628 & ~w838) | (~w628 & w2169) | (~w838 & w2169);
assign w1639 = ~pi146 & ~w474;
assign w1640 = ~pi214 & w1781;
assign w1641 = (w1680 & w157) | (w1680 & w1207) | (w157 & w1207);
assign w1642 = ~pi168 & ~w341;
assign w1643 = ~w849 & w1102;
assign w1644 = w1048 & ~w1074;
assign w1645 = ~w1751 & ~w209;
assign w1646 = ~w928 & w204;
assign w1647 = ~pi167 & ~w1351;
assign w1648 = (w1181 & ~w1345) | (w1181 & w1739) | (~w1345 & w1739);
assign w1649 = ~w1147 & ~w1623;
assign w1650 = ~w808 & ~w1498;
assign w1651 = w1050 & ~w1313;
assign w1652 = ~w429 & w705;
assign w1653 = ~w343 & ~w512;
assign w1654 = ~w1797 & ~w2055;
assign w1655 = ~w1759 & w1586;
assign w1656 = (w1857 & w316) | (w1857 & w1310) | (w316 & w1310);
assign w1657 = ~pi208 & w2192;
assign w1658 = pi149 & w1128;
assign w1659 = ~w580 & ~w1622;
assign w1660 = (~w785 & ~w1479) | (~w785 & w1582) | (~w1479 & w1582);
assign w1661 = ~w1408 & ~w2110;
assign w1662 = w809 & ~w1320;
assign w1663 = ~w961 & ~w1973;
assign w1664 = w1470 & ~w1388;
assign w1665 = (~w762 & ~w582) | (~w762 & w1079) | (~w582 & w1079);
assign w1666 = (w1244 & w920) | (w1244 & w2022) | (w920 & w2022);
assign w1667 = ~w1884 & ~w2188;
assign w1668 = ~pi162 & ~w602;
assign w1669 = w1181 & ~w1030;
assign w1670 = (~w1600 & ~w1463) | (~w1600 & w1850) | (~w1463 & w1850);
assign w1671 = (~w443 & ~w257) | (~w443 & w314) | (~w257 & w314);
assign w1672 = (w1010 & w2211) | (w1010 & ~w863) | (w2211 & ~w863);
assign w1673 = (~w1932 & ~w1905) | (~w1932 & w918) | (~w1905 & w918);
assign w1674 = (w1875 & w1551) | (w1875 & w1163) | (w1551 & w1163);
assign w1675 = (w1635 & w2189) | (w1635 & ~w62) | (w2189 & ~w62);
assign w1676 = (~w2120 & w506) | (~w2120 & w1598) | (w506 & w1598);
assign w1677 = (~w1705 & w77) | (~w1705 & w1800) | (w77 & w1800);
assign w1678 = (~w1715 & w1936) | (~w1715 & w1213) | (w1936 & w1213);
assign w1679 = ~w302 & ~w64;
assign w1680 = (~w489 & w1359) | (~w489 & w546) | (w1359 & w546);
assign w1681 = ~w1362 & ~w1458;
assign w1682 = ~w187 & ~w1583;
assign w1683 = ~w1362 & w419;
assign w1684 = (~w1680 & w1182) | (~w1680 & w412) | (w1182 & w412);
assign w1685 = (~w1042 & ~w700) | (~w1042 & w1798) | (~w700 & w1798);
assign w1686 = w1862 & ~w1440;
assign w1687 = ~pi142 & ~w2180;
assign w1688 = ~w320 & w388;
assign w1689 = (~w2183 & ~w1951) | (~w2183 & ~w1876) | (~w1951 & ~w1876);
assign w1690 = w1285 & w2167;
assign w1691 = w1136 & ~w1991;
assign w1692 = ~w1300 & ~w495;
assign w1693 = ~w1982 & ~w2015;
assign w1694 = pi135 & w1419;
assign w1695 = pi153 & w959;
assign w1696 = (w1596 & w1148) | (w1596 & w456) | (w1148 & w456);
assign w1697 = ~w1970 & ~w1372;
assign w1698 = (w844 & w1174) | (w844 & w915) | (w1174 & w915);
assign w1699 = pi220 & ~w754;
assign w1700 = pi240 & ~w797;
assign w1701 = ~w1694 & ~w662;
assign w1702 = ~w1446 & ~w721;
assign w1703 = w503 & ~w8;
assign w1704 = w2043 & ~w1456;
assign w1705 = ~w2175 & w711;
assign w1706 = w1546 & ~w605;
assign w1707 = ~w344 & ~w116;
assign w1708 = ~pi211 & w1321;
assign w1709 = ~w1266 & ~w736;
assign w1710 = ~w2089 & ~w893;
assign w1711 = ~w1364 & w1697;
assign w1712 = ~w1091 & ~w2123;
assign w1713 = ~w1825 & ~w2001;
assign w1714 = (~w68 & ~w2148) | (~w68 & w566) | (~w2148 & w566);
assign w1715 = (~w1927 & w1677) | (~w1927 & w1102) | (w1677 & w1102);
assign w1716 = ~w2040 & ~w1233;
assign w1717 = w934 & w344;
assign w1718 = ~w1569 & ~w1606;
assign w1719 = ~w1701 & ~w406;
assign w1720 = ~w1543 & ~w1784;
assign w1721 = ~w1325 & w1293;
assign w1722 = ~pi063 & ~pi127;
assign w1723 = ~w1165 & ~w1508;
assign w1724 = ~pi060 & ~pi124;
assign w1725 = pi061 & pi125;
assign w1726 = ~w2043 & ~w1655;
assign w1727 = ~w1566 & ~w1468;
assign w1728 = (~w2183 & ~w1951) | (~w2183 & ~w1177) | (~w1951 & ~w1177);
assign w1729 = (w1870 & w292) | (w1870 & w554) | (w292 & w554);
assign w1730 = (w2146 & w635) | (w2146 & w2127) | (w635 & w2127);
assign w1731 = ~pi233 & w1279;
assign w1732 = ~w1649 & ~w1147;
assign w1733 = ~pi182 & ~w454;
assign w1734 = ~w674 & ~w60;
assign w1735 = (~w595 & w2165) | (~w595 & w620) | (w2165 & w620);
assign w1736 = (w1133 & w380) | (w1133 & w1675) | (w380 & w1675);
assign w1737 = (w980 & w909) | (w980 & w727) | (w909 & w727);
assign w1738 = w1716 & w1090;
assign w1739 = ~w1179 & w1181;
assign w1740 = ~pi009 & ~pi073;
assign w1741 = pi010 & pi074;
assign w1742 = pi211 & ~w1321;
assign w1743 = (~w489 & w821) | (~w489 & w350) | (w821 & w350);
assign w1744 = pi237 & ~w768;
assign w1745 = ~w164 & ~w1724;
assign w1746 = ~w492 & ~w2187;
assign w1747 = ~w1151 & ~w1664;
assign w1748 = w630 & ~w1127;
assign w1749 = (~w1216 & ~w1461) | (~w1216 & w654) | (~w1461 & w654);
assign w1750 = ~w1035 & ~w518;
assign w1751 = ~w431 & ~w588;
assign w1752 = ~w1503 & ~w1906;
assign w1753 = (~w1680 & w871) | (~w1680 & w1271) | (w871 & w1271);
assign w1754 = (~w1955 & ~w1794) | (~w1955 & w24) | (~w1794 & w24);
assign w1755 = (~w396 & w274) | (~w396 & w221) | (w274 & w221);
assign w1756 = w1124 & w1060;
assign w1757 = ~w1535 & ~w1702;
assign w1758 = ~w321 & ~w445;
assign w1759 = (~w1487 & ~w363) | (~w1487 & w402) | (~w363 & w402);
assign w1760 = (~w1680 & w1183) | (~w1680 & w1944) | (w1183 & w1944);
assign w1761 = (~w1744 & ~w431) | (~w1744 & w1931) | (~w431 & w1931);
assign w1762 = ~w253 & ~w1295;
assign w1763 = (~w1502 & w1484) | (~w1502 & w1497) | (w1484 & w1497);
assign w1764 = (~w1517 & ~w2138) | (~w1517 & w924) | (~w2138 & w924);
assign w1765 = ~pi161 & ~w324;
assign w1766 = (w1098 & w1229) | (w1098 & w1870) | (w1229 & w1870);
assign w1767 = ~w528 & ~w1509;
assign w1768 = ~w1045 & ~w931;
assign w1769 = pi222 & ~w1978;
assign w1770 = ~pi134 & ~w2035;
assign w1771 = ~w422 & ~w773;
assign w1772 = (~w1502 & w902) | (~w1502 & w912) | (w902 & w912);
assign w1773 = (~w489 & w1063) | (~w489 & w1793) | (w1063 & w1793);
assign w1774 = pi255 & w949;
assign w1775 = w833 & ~w608;
assign w1776 = ~w948 & w319;
assign w1777 = pi144 & w1037;
assign w1778 = (w2120 & w1100) | (w2120 & w231) | (w1100 & w231);
assign w1779 = (w1350 & w399) | (w1350 & ~w706) | (w399 & ~w706);
assign w1780 = (~w2028 & w993) | (~w2028 & w1291) | (w993 & w1291);
assign w1781 = (~w579 & ~w1128) | (~w579 & w1553) | (~w1128 & w1553);
assign w1782 = (~w1949 & ~w1535) | (~w1949 & w890) | (~w1535 & w890);
assign w1783 = (w931 & w729) | (w931 & w1269) | (w729 & w1269);
assign w1784 = w568 & ~w1653;
assign w1785 = ~w1844 & ~w585;
assign w1786 = ~w2145 & ~w1324;
assign w1787 = ~pi186 & ~w1035;
assign w1788 = ~w1343 & ~w2060;
assign w1789 = ~w2159 & w1094;
assign w1790 = w640 & ~w2100;
assign w1791 = ~w1039 & ~w239;
assign w1792 = ~w1539 & ~w47;
assign w1793 = w471 & ~w1329;
assign w1794 = ~w1955 & ~w2190;
assign w1795 = ~w548 & w20;
assign w1796 = ~pi040 & ~pi104;
assign w1797 = pi041 & pi105;
assign w1798 = ~pi128 & ~w1042;
assign w1799 = (~w489 & w1121) | (~w489 & w92) | (w1121 & w92);
assign w1800 = ~w15 & ~w1705;
assign w1801 = w351 & w1528;
assign w1802 = ~pi139 & ~w1347;
assign w1803 = ~w1389 & ~w702;
assign w1804 = w1364 & ~w1697;
assign w1805 = ~pi170 & ~w2056;
assign w1806 = (~w1884 & ~w1667) | (~w1884 & w935) | (~w1667 & w935);
assign w1807 = (~w230 & ~w694) | (~w230 & w1480) | (~w694 & w1480);
assign w1808 = w1655 | w1974;
assign w1809 = w2185 & w1583;
assign w1810 = (w2120 & w1237) | (w2120 & ~w1250) | (w1237 & ~w1250);
assign w1811 = w1666 & w1457;
assign w1812 = (w960 & w304) | (w960 & ~w1152) | (w304 & ~w1152);
assign w1813 = ~w2033 & ~w897;
assign w1814 = (~w1680 & w369) | (~w1680 & w888) | (w369 & w888);
assign w1815 = w299 & w1650;
assign w1816 = (~w454 & ~w358) | (~w454 & w1733) | (~w358 & w1733);
assign w1817 = (w1502 & w377) | (w1502 & w433) | (w377 & w433);
assign w1818 = ~w1157 & ~w134;
assign w1819 = ~w1789 & ~w1583;
assign w1820 = w183 & w95;
assign w1821 = (w22 & w989) | (w22 & w326) | (w989 & w326);
assign w1822 = w1438 & ~w4;
assign w1823 = ~w1699 & ~w240;
assign w1824 = (w1012 & w835) | (w1012 & w1960) | (w835 & w1960);
assign w1825 = pi205 & ~w1807;
assign w1826 = ~w385 & w741;
assign w1827 = ~w1502 & ~w1641;
assign w1828 = (w1502 & w1669) | (w1502 & w2048) | (w1669 & w2048);
assign w1829 = ~w1211 & ~w1415;
assign w1830 = (~w137 & w886) | (~w137 & w664) | (w886 & w664);
assign w1831 = pi231 & ~w1923;
assign w1832 = w1539 & w2208;
assign w1833 = ~pi244 & w478;
assign w1834 = w262 & ~w1785;
assign w1835 = (w260 & w531) | (w260 & w1100) | (w531 & w1100);
assign w1836 = ~w208 & w122;
assign w1837 = (~w38 & ~w1561) | (~w38 & w1078) | (~w1561 & w1078);
assign w1838 = (w1680 & w591) | (w1680 & w1305) | (w591 & w1305);
assign w1839 = ~w1011 & ~w144;
assign w1840 = ~w1888 & ~w878;
assign w1841 = ~w15 & w77;
assign w1842 = ~w857 & ~w761;
assign w1843 = w1794 & w367;
assign w1844 = ~w585 & ~w132;
assign w1845 = ~w1206 & ~w594;
assign w1846 = ~w2087 & ~w1743;
assign w1847 = (w1150 & w807) | (w1150 & w1980) | (w807 & w1980);
assign w1848 = ~pi175 & ~w1275;
assign w1849 = (w2131 & w1413) | (w2131 & w1177) | (w1413 & w1177);
assign w1850 = ~pi177 & ~w1600;
assign w1851 = (w931 & w729) | (w931 & w792) | (w729 & w792);
assign w1852 = pi182 & w358;
assign w1853 = ~pi151 & ~w285;
assign w1854 = ~pi154 & ~w211;
assign w1855 = (w1680 & w1826) | (w1680 & w1123) | (w1826 & w1123);
assign w1856 = ~w1868 & ~w818;
assign w1857 = ~w1386 & ~w1583;
assign w1858 = (w1152 & w647) | (w1152 & w23) | (w647 & w23);
assign w1859 = (~w1240 & w750) | (~w1240 & ~w1237) | (w750 & ~w1237);
assign w1860 = ~w1283 & ~w1769;
assign w1861 = (~w110 & ~w1285) | (~w110 & w493) | (~w1285 & w493);
assign w1862 = (~w1700 & ~w609) | (~w1700 & w1363) | (~w609 & w1363);
assign w1863 = ~pi245 & w127;
assign w1864 = (w1502 & w2112) | (w1502 & w952) | (w2112 & w952);
assign w1865 = ~pi168 & ~w357;
assign w1866 = ~w659 & ~w1370;
assign w1867 = pi151 & w261;
assign w1868 = ~w1861 & w872;
assign w1869 = ~w1486 & ~w981;
assign w1870 = (w915 & w980) | (w915 & w1185) | (w980 & w1185);
assign w1871 = (~w1031 & ~w2115) | (~w1031 & w1477) | (~w2115 & w1477);
assign w1872 = ~w1747 & w1859;
assign w1873 = (~w143 & ~w1503) | (~w143 & w126) | (~w1503 & w126);
assign w1874 = ~w719 & ~w1855;
assign w1875 = ~w1636 & ~w439;
assign w1876 = w15 & ~w77;
assign w1877 = (~w2056 & ~w2150) | (~w2056 & w1805) | (~w2150 & w1805);
assign w1878 = (w10 & w2049) | (w10 & w1748) | (w2049 & w1748);
assign w1879 = ~pi029 & ~pi093;
assign w1880 = pi030 & pi094;
assign w1881 = ~w545 & ~w244;
assign w1882 = w726 & w1942;
assign w1883 = w729 & w931;
assign w1884 = ~w2061 & w2132;
assign w1885 = (~w608 & ~w1167) | (~w608 & w2094) | (~w1167 & w2094);
assign w1886 = ~pi148 & ~w408;
assign w1887 = ~w2043 & w1980;
assign w1888 = ~w2149 & ~w1335;
assign w1889 = ~w2018 & w939;
assign w1890 = pi209 & ~w118;
assign w1891 = ~w9 & ~w1171;
assign w1892 = ~pi223 & w911;
assign w1893 = ~w1410 & ~w1616;
assign w1894 = ~w533 & ~w2065;
assign w1895 = ~w494 & ~w2000;
assign w1896 = w397 & ~w590;
assign w1897 = ~w206 & ~w1930;
assign w1898 = ~w599 & ~w10;
assign w1899 = ~w187 & ~w149;
assign w1900 = ~w1269 & w679;
assign w1901 = ~w1968 & ~w917;
assign w1902 = ~w702 & ~w301;
assign w1903 = ~w1255 & ~w1554;
assign w1904 = ~w2143 & w439;
assign w1905 = ~w1932 & ~w827;
assign w1906 = ~w1592 & ~w710;
assign w1907 = ~w2101 & ~w533;
assign w1908 = (w1872 & w2124) | (w1872 & w1250) | (w2124 & w1250);
assign w1909 = ~w1817 & ~w1772;
assign w1910 = w1269 & w507;
assign w1911 = (w416 & w405) | (w416 & w706) | (w405 & w706);
assign w1912 = ~w1562 & ~w1342;
assign w1913 = (w39 & w824) | (w39 & ~w1980) | (w824 & ~w1980);
assign w1914 = (w287 & w438) | (w287 & w1715) | (w438 & w1715);
assign w1915 = (~w326 & w1443) | (~w326 & w1836) | (w1443 & w1836);
assign w1916 = (~w1502 & w463) | (~w1502 & w1435) | (w463 & w1435);
assign w1917 = (~w1722 & ~w891) | (~w1722 & w1630) | (~w891 & w1630);
assign w1918 = ~w1738 & ~w470;
assign w1919 = w347 & w1417;
assign w1920 = ~w1508 & ~w1245;
assign w1921 = ~pi238 & w170;
assign w1922 = w1057 & w60;
assign w1923 = (~w1469 & ~w526) | (~w1469 & w1263) | (~w526 & w1263);
assign w1924 = (w679 & w1152) | (w679 & w1900) | (w1152 & w1900);
assign w1925 = w253 & ~w865;
assign w1926 = w1901 & ~w1604;
assign w1927 = (~w1313 & w2080) | (~w1313 & w295) | (w2080 & w295);
assign w1928 = (w137 & w1882) | (w137 & w1139) | (w1882 & w1139);
assign w1929 = ~w1181 & w1030;
assign w1930 = ~w843 & ~w1226;
assign w1931 = ~w588 & ~w1744;
assign w1932 = ~w1449 & w942;
assign w1933 = (w675 & w54) | (w675 & w1093) | (w54 & w1093);
assign w1934 = ~pi219 & w875;
assign w1935 = ~pi146 & ~w1589;
assign w1936 = (w681 & w1835) | (w681 & w2120) | (w1835 & w2120);
assign w1937 = (w1502 & w954) | (w1502 & w328) | (w954 & w328);
assign w1938 = ~pi187 & ~w114;
assign w1939 = (w316 & w2088) | (w316 & w964) | (w2088 & w964);
assign w1940 = (~w1035 & ~w1750) | (~w1035 & w1787) | (~w1750 & w1787);
assign w1941 = (~w2120 & w451) | (~w2120 & w572) | (w451 & w572);
assign w1942 = ~w312 & ~w1593;
assign w1943 = (~w88 & w1636) | (~w88 & w480) | (w1636 & w480);
assign w1944 = (~w1939 & w1092) | (~w1939 & w1476) | (w1092 & w1476);
assign w1945 = ~w2168 & w814;
assign w1946 = w129 & ~w1870;
assign w1947 = ~w978 & ~w298;
assign w1948 = w928 & ~w1800;
assign w1949 = pi197 & ~w1665;
assign w1950 = ~w1131 & ~w1062;
assign w1951 = (w2126 & w1425) | (w2126 & w685) | (w1425 & w685);
assign w1952 = ~pi138 & ~w1741;
assign w1953 = (w585 & ~w1785) | (w585 & ~w976) | (~w1785 & ~w976);
assign w1954 = (~w1927 & w1643) | (~w1927 & w1067) | (w1643 & w1067);
assign w1955 = pi251 & ~w1940;
assign w1956 = (w60 & w948) | (w60 & w1922) | (w948 & w1922);
assign w1957 = ~w2043 & ~w1974;
assign w1958 = (w1872 & w2124) | (w1872 & w1870) | (w2124 & w1870);
assign w1959 = ~w107 & w1404;
assign w1960 = (~w1045 & ~w931) | (~w1045 & w410) | (~w931 & w410);
assign w1961 = ~pi049 & ~pi113;
assign w1962 = pi050 & pi114;
assign w1963 = ~pi186 & ~w1750;
assign w1964 = ~w2160 & ~w921;
assign w1965 = ~w1494 & ~w677;
assign w1966 = w2134 & ~w2064;
assign w1967 = (w149 & ~w1899) | (w149 & ~w1819) | (~w1899 & ~w1819);
assign w1968 = ~w855 & w1505;
assign w1969 = (w1680 & w1065) | (w1680 & w2166) | (w1065 & w2166);
assign w1970 = ~w186 & ~w479;
assign w1971 = ~w299 & ~w1650;
assign w1972 = ~w1956 & ~w1776;
assign w1973 = ~pi157 & ~w373;
assign w1974 = ~w1471 & w361;
assign w1975 = w67 & w1775;
assign w1976 = w751 & ~w316;
assign w1977 = (w1538 & w1040) | (w1538 & ~w644) | (w1040 & ~w644);
assign w1978 = (~w898 & ~w373) | (~w898 & w1146) | (~w373 & w1146);
assign w1979 = ~pi194 & w846;
assign w1980 = (~w1974 & w1871) | (~w1974 & w1456) | (w1871 & w1456);
assign w1981 = ~pi218 & w1990;
assign w1982 = (~w1680 & w2068) | (~w1680 & w523) | (w2068 & w523);
assign w1983 = (w980 & w1442) | (w980 & w155) | (w1442 & w155);
assign w1984 = ~w2066 & ~w1979;
assign w1985 = (w1502 & w1066) | (w1502 & w802) | (w1066 & w802);
assign w1986 = ~pi140 & ~w694;
assign w1987 = (~w1347 & ~w1166) | (~w1347 & w1802) | (~w1166 & w1802);
assign w1988 = ~pi016 & ~pi080;
assign w1989 = pi017 & pi081;
assign w1990 = (~w414 & ~w959) | (~w414 & w1199) | (~w959 & w1199);
assign w1991 = ~w1932 & ~w1905;
assign w1992 = w766 & ~w1028;
assign w1993 = w2159 & ~w1094;
assign w1994 = (~w1502 & w352) | (~w1502 & w1159) | (w352 & w1159);
assign w1995 = pi146 & w1589;
assign w1996 = pi174 & w966;
assign w1997 = ~w1053 & ~w1825;
assign w1998 = (w2028 & w2108) | (w2028 & w2191) | (w2108 & w2191);
assign w1999 = ~pi131 & ~w1842;
assign w2000 = ~w1219 & ~w430;
assign w2001 = ~pi205 & w1807;
assign w2002 = pi228 & ~w382;
assign w2003 = (w2208 & w1832) | (w2208 & ~w1680) | (w1832 & ~w1680);
assign w2004 = ~pi137 & ~w1548;
assign w2005 = (~w1715 & w1851) | (~w1715 & w1354) | (w1851 & w1354);
assign w2006 = (~w1281 & ~w160) | (~w1281 & w1170) | (~w160 & w1170);
assign w2007 = w1950 & ~w823;
assign w2008 = ~pi221 & w728;
assign w2009 = ~w656 & ~w71;
assign w2010 = ~w262 & w94;
assign w2011 = w1570 & w1453;
assign w2012 = pi187 & w114;
assign w2013 = w129 & ~w1677;
assign w2014 = ~w773 & ~w1371;
assign w2015 = (w1680 & w1175) | (w1680 & w2139) | (w1175 & w2139);
assign w2016 = (~w915 & w1936) | (~w915 & w1213) | (w1936 & w1213);
assign w2017 = w1304 & ~w530;
assign w2018 = ~w468 & ~w1068;
assign w2019 = ~pi182 & ~w358;
assign w2020 = w2134 & ~w1268;
assign w2021 = (w1748 & w441) | (w1748 & w613) | (w441 & w613);
assign w2022 = ~w1968 & ~w1844;
assign w2023 = pi167 & w1351;
assign w2024 = (w466 & w184) | (w466 & w2198) | (w184 & w2198);
assign w2025 = (w39 & w824) | (w39 & ~w675) | (w824 & ~w675);
assign w2026 = ~w129 & w1102;
assign w2027 = ~w1618 & ~w587;
assign w2028 = (~w948 & w1162) | (~w948 & w249) | (w1162 & w249);
assign w2029 = w2115 & w1206;
assign w2030 = w1764 & ~w755;
assign w2031 = ~w228 & ~w486;
assign w2032 = ~pi027 & ~pi091;
assign w2033 = pi028 & pi092;
assign w2034 = ~pi005 & ~pi069;
assign w2035 = pi006 & pi070;
assign w2036 = ~w630 & w1127;
assign w2037 = ~w1868 & ~w82;
assign w2038 = ~pi248 & w133;
assign w2039 = (w1269 & w1533) | (w1269 & w2163) | (w1533 & w2163);
assign w2040 = pi191 & ~w891;
assign w2041 = ~w2115 & ~w1031;
assign w2042 = ~w733 & ~w1701;
assign w2043 = ~w1655 & ~w251;
assign w2044 = ~w299 & ~w808;
assign w2045 = w1761 & ~w254;
assign w2046 = ~w1425 & w1102;
assign w2047 = (w1950 & w466) | (w1950 & w525) | (w466 & w525);
assign w2048 = (w549 & w1648) | (w549 & w1549) | (w1648 & w1549);
assign w2049 = w1286 & w10;
assign w2050 = ~w1151 & ~w466;
assign w2051 = (~w1040 & ~w1538) | (~w1040 & w1939) | (~w1538 & w1939);
assign w2052 = (~w1680 & w1911) | (~w1680 & ~w2054) | (w1911 & ~w2054);
assign w2053 = ~pi215 & w1246;
assign w2054 = (~w405 & ~w706) | (~w405 & ~w326) | (~w706 & ~w326);
assign w2055 = ~pi041 & ~pi105;
assign w2056 = pi042 & pi106;
assign w2057 = ~pi161 & ~w1491;
assign w2058 = ~pi004 & ~pi068;
assign w2059 = pi005 & pi069;
assign w2060 = (~w1502 & w2095) | (~w1502 & w1945) | (w2095 & w1945);
assign w2061 = (~w1508 & ~w1920) | (~w1508 & w1723) | (~w1920 & w1723);
assign w2062 = (w149 & ~w1899) | (w149 & ~w2088) | (~w1899 & ~w2088);
assign w2063 = ~w1754 & w2027;
assign w2064 = (~w811 & w1597) | (~w811 & w273) | (w1597 & w273);
assign w2065 = ~pi213 & w501;
assign w2066 = pi194 & ~w846;
assign w2067 = ~w1901 & ~w1555;
assign w2068 = (w6 & w472) | (w6 & w1107) | (w472 & w1107);
assign w2069 = (w2208 & w1832) | (w2208 & w2094) | (w1832 & w2094);
assign w2070 = (w2047 & w2007) | (w2047 & w1602) | (w2007 & w1602);
assign w2071 = ~w2028 & w1845;
assign w2072 = ~pi242 & w1670;
assign w2073 = (~w1680 & w724) | (~w1680 & w527) | (w724 & w527);
assign w2074 = (w204 & w291) | (w204 & w1168) | (w291 & w1168);
assign w2075 = ~pi152 & ~w626;
assign w2076 = (~w330 & w1991) | (~w330 & w44) | (w1991 & w44);
assign w2077 = w1782 & ~w749;
assign w2078 = ~w486 & ~w2184;
assign w2079 = w160 & w1319;
assign w2080 = w107 & w417;
assign w2081 = ~pi031 & ~pi095;
assign w2082 = pi032 & pi096;
assign w2083 = ~w275 & w1762;
assign w2084 = (w1559 & w197) | (w1559 & w50) | (w197 & w50);
assign w2085 = ~pi174 & ~w966;
assign w2086 = ~w29 & ~w150;
assign w2087 = (w489 & w490) | (w489 & w1526) | (w490 & w1526);
assign w2088 = (~w1789 & ~w1583) | (~w1789 & w500) | (~w1583 & w500);
assign w2089 = pi246 & ~w1083;
assign w2090 = ~pi144 & ~w1037;
assign w2091 = w177 & w1663;
assign w2092 = ~w771 & ~w1396;
assign w2093 = ~w481 & ~w840;
assign w2094 = ~w1539 & ~w1143;
assign w2095 = ~w2168 & w1047;
assign w2096 = ~w1561 & ~w1557;
assign w2097 = (~w164 & ~w1745) | (~w164 & w612) | (~w1745 & w612);
assign w2098 = ~w1620 & ~w1398;
assign w2099 = ~w544 & ~w1632;
assign w2100 = ~w1752 & ~w66;
assign w2101 = ~w1658 & ~w237;
assign w2102 = ~w36 & ~w125;
assign w2103 = ~w1275 & ~w1005;
assign w2104 = ~w468 & ~w1555;
assign w2105 = ~w701 & ~w601;
assign w2106 = (~w626 & ~w1633) | (~w626 & w2075) | (~w1633 & w2075);
assign w2107 = (w1711 & ~w947) | (w1711 & ~w581) | (~w947 & ~w581);
assign w2108 = ~w2115 & ~w1206;
assign w2109 = ~w1397 & ~w312;
assign w2110 = (~w1502 & w1172) | (~w1502 & w281) | (w1172 & w281);
assign w2111 = ~w187 & w2088;
assign w2112 = (~w1870 & w1504) | (~w1870 & w684) | (w1504 & w684);
assign w2113 = ~w1425 & w1677;
assign w2114 = w349 & ~w805;
assign w2115 = ~w1031 & ~w96;
assign w2116 = (~w198 & ~w183) | (~w198 & w460) | (~w183 & w460);
assign w2117 = ~w393 & ~w534;
assign w2118 = (w10 & w2049) | (w10 & w748) | (w2049 & w748);
assign w2119 = w759 & ~w522;
assign w2120 = (~w204 & w327) | (~w204 & w641) | (w327 & w641);
assign w2121 = ~pi237 & w768;
assign w2122 = ~pi189 & ~w1153;
assign w2123 = ~w364 & ~w2057;
assign w2124 = (~w2120 & w1287) | (~w2120 & w487) | (w1287 & w487);
assign w2125 = ~pi199 & w895;
assign w2126 = ~w1714 & w990;
assign w2127 = ~w1562 & ~w813;
assign w2128 = ~w869 & ~w372;
assign w2129 = ~pi145 & ~w1054;
assign w2130 = w2168 & w2126;
assign w2131 = w2168 & w1951;
assign w2132 = ~w514 & ~w825;
assign w2133 = ~w1867 & ~w919;
assign w2134 = ~w1652 & ~w930;
assign w2135 = ~pi030 & ~pi094;
assign w2136 = pi031 & pi095;
assign w2137 = (~w64 & ~w1036) | (~w64 & w1679) | (~w1036 & w1679);
assign w2138 = ~w1517 & ~w154;
assign w2139 = (w316 & w145) | (w316 & w778) | (w145 & w778);
assign w2140 = ~pi034 & ~pi098;
assign w2141 = pi035 & pi099;
assign w2142 = ~w616 & ~w1580;
assign w2143 = ~w88 & ~w676;
assign w2144 = (~w1556 & w270) | (~w1556 & w581) | (w270 & w581);
assign w2145 = pi152 & w1633;
assign w2146 = ~w15 & ~w1342;
assign w2147 = ~w1965 & ~w1947;
assign w2148 = ~w68 & ~w547;
assign w2149 = pi154 & w607;
assign w2150 = ~w2056 & ~w1215;
assign w2151 = ~w286 & w1;
assign w2152 = ~pi167 & ~w1430;
assign w2153 = ~w792 & w679;
assign w2154 = (~w1185 & w815) | (~w1185 & w310) | (w815 & w310);
assign w2155 = (~w915 & w1504) | (~w915 & w684) | (w1504 & w684);
assign w2156 = (~w125 & ~w780) | (~w125 & w2102) | (~w780 & w2102);
assign w2157 = (w1680 & w1575) | (w1680 & w1330) | (w1575 & w1330);
assign w2158 = ~w2143 & ~w1402;
assign w2159 = (~w1699 & ~w1823) | (~w1699 & w403) | (~w1823 & w403);
assign w2160 = (w1502 & w2005) | (w1502 & w334) | (w2005 & w334);
assign w2161 = ~pi209 & w118;
assign w2162 = ~w2151 & ~w933;
assign w2163 = w1269 & ~w1152;
assign w2164 = (~w1715 & w2163) | (~w1715 & w792) | (w2163 & w792);
assign w2165 = w1815 & w1650;
assign w2166 = (w1939 & w7) | (w1939 & w1587) | (w7 & w1587);
assign w2167 = ~w1014 & ~w1668;
assign w2168 = ~w1256 & ~w1686;
assign w2169 = ~w1655 & ~w628;
assign w2170 = w2143 & ~w1636;
assign w2171 = (~w1953 & w1904) | (~w1953 & w289) | (w1904 & w289);
assign w2172 = ~pi227 & w105;
assign w2173 = (w22 & w989) | (w22 & w416) | (w989 & w416);
assign w2174 = ~w1052 & ~w713;
assign w2175 = (~w116 & ~w934) | (~w116 & w1707) | (~w934 & w1707);
assign w2176 = w1710 & w359;
assign w2177 = (w1680 & w464) | (w1680 & w1314) | (w464 & w1314);
assign w2178 = ~pi130 & ~w535;
assign w2179 = ~pi013 & ~pi077;
assign w2180 = pi014 & pi078;
assign w2181 = ~pi138 & ~w1637;
assign w2182 = ~w969 & ~w278;
assign w2183 = w1425 | w2126;
assign w2184 = ~pi207 & w280;
assign w2185 = w1386 & w1583;
assign w2186 = (w549 & w2039) | (w549 & w1186) | (w2039 & w1186);
assign w2187 = (w2028 & w1077) | (w2028 & w1933) | (w1077 & w1933);
assign w2188 = w2061 & ~w2132;
assign w2189 = ~w1795 & ~w1528;
assign w2190 = ~pi251 & w1940;
assign w2191 = ~w2115 & w1082;
assign w2192 = (~w688 & ~w32) | (~w688 & w696) | (~w32 & w696);
assign w2193 = ~w1711 & ~w953;
assign w2194 = (~w2059 & ~w76) | (~w2059 & w722) | (~w76 & w722);
assign w2195 = (~w1711 & ~w129) | (~w1711 & w905) | (~w129 & w905);
assign w2196 = ~pi144 & ~w584;
assign w2197 = ~w190 & ~w1132;
assign w2198 = (w1237 & w652) | (w1237 & w945) | (w652 & w945);
assign w2199 = (w740 & w1312) | (w740 & ~w610) | (w1312 & ~w610);
assign w2200 = ~w1223 & ~w683;
assign w2201 = ~pi253 & w2097;
assign w2202 = w468 & w1555;
assign w2203 = w1012 & ~w396;
assign w2204 = ~w609 & ~w1360;
assign w2205 = w1568 & w1409;
assign w2206 = (w1250 & w1941) | (w1250 & w171) | (w1941 & w171);
assign w2207 = ~w1897 & ~w504;
assign w2208 = ~w47 & ~w1260;
assign w2209 = (w873 & w1919) | (w873 & ~w1768) | (w1919 & ~w1768);
assign w2210 = w1362 & ~w419;
assign w2211 = ~w2094 & w1010;
assign one = 1;
assign po00 = w1406;// level 6
assign po01 = w444;// level 9
assign po02 = w1142;// level 11
assign po03 = w624;// level 12
assign po04 = w2200;// level 13
assign po05 = w1427;// level 13
assign po06 = w1972;// level 14
assign po07 = w932;// level 14
assign po08 = w33;// level 14
assign po09 = w91;// level 15
assign po10 = w1465;// level 15
assign po11 = w604;// level 15
assign po12 = w1581;// level 15
assign po13 = w1361;// level 15
assign po14 = w1383;// level 15
assign po15 = w1746;// level 16
assign po16 = w955;// level 15
assign po17 = w1488;// level 16
assign po18 = w615;// level 16
assign po19 = w2128;// level 16
assign po20 = w658;// level 16
assign po21 = w1515;// level 16
assign po22 = w1113;// level 16
assign po23 = w779;// level 16
assign po24 = w1846;// level 16
assign po25 = w1418;// level 17
assign po26 = w354;// level 17
assign po27 = w1874;// level 17
assign po28 = w1441;// level 17
assign po29 = w1016;// level 17
assign po30 = w1693;// level 17
assign po31 = w739;// level 17
assign po32 = w178;// level 17
assign po33 = w130;// level 17
assign po34 = w552;// level 17
assign po35 = w938;// level 17
assign po36 = w59;// level 17
assign po37 = w861;// level 17
assign po38 = w1516;// level 17
assign po39 = w423;// level 17
assign po40 = w556;// level 18
assign po41 = w1827;// level 17
assign po42 = w300;// level 18
assign po43 = w1758;// level 18
assign po44 = w1661;// level 18
assign po45 = w227;// level 18
assign po46 = w387;// level 18
assign po47 = w337;// level 18
assign po48 = w1460;// level 18
assign po49 = w1788;// level 18
assign po50 = w1358;// level 18
assign po51 = w1280;// level 18
assign po52 = w1964;// level 18
assign po53 = w874;// level 18
assign po54 = w742;// level 18
assign po55 = w596;// level 18
assign po56 = w383;// level 18
assign po57 = w1137;// level 18
assign po58 = w1138;// level 18
assign po59 = w1224;// level 18
assign po60 = w1909;// level 18
assign po61 = w1239;// level 18
assign po62 = w1483;// level 18
assign po63 = w623;// level 18
assign po64 = w1322;// level 18
assign po65 = w146;// level 18
endmodule
