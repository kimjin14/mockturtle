module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 ;
  assign n257 = x0 & ~x128 ;
  assign n258 = ~x0 & x128 ;
  assign n259 = n257 | n258 ;
  assign n260 = x0 & x128 ;
  assign n261 = ( x1 & ~x129 ) | ( x1 & n260 ) | ( ~x129 & n260 ) ;
  assign n262 = ( ~x1 & x129 ) | ( ~x1 & n261 ) | ( x129 & n261 ) ;
  assign n263 = ( ~n260 & n261 ) | ( ~n260 & n262 ) | ( n261 & n262 ) ;
  assign n264 = ( x1 & x129 ) | ( x1 & n260 ) | ( x129 & n260 ) ;
  assign n265 = ( x2 & ~x130 ) | ( x2 & n264 ) | ( ~x130 & n264 ) ;
  assign n266 = ( ~x2 & x130 ) | ( ~x2 & n265 ) | ( x130 & n265 ) ;
  assign n267 = ( ~n264 & n265 ) | ( ~n264 & n266 ) | ( n265 & n266 ) ;
  assign n268 = ( x2 & x130 ) | ( x2 & n264 ) | ( x130 & n264 ) ;
  assign n269 = ( x3 & ~x131 ) | ( x3 & n268 ) | ( ~x131 & n268 ) ;
  assign n270 = ( ~x3 & x131 ) | ( ~x3 & n269 ) | ( x131 & n269 ) ;
  assign n271 = ( ~n268 & n269 ) | ( ~n268 & n270 ) | ( n269 & n270 ) ;
  assign n272 = ( x3 & x131 ) | ( x3 & n268 ) | ( x131 & n268 ) ;
  assign n273 = ( x4 & ~x132 ) | ( x4 & n272 ) | ( ~x132 & n272 ) ;
  assign n274 = ( ~x4 & x132 ) | ( ~x4 & n273 ) | ( x132 & n273 ) ;
  assign n275 = ( ~n272 & n273 ) | ( ~n272 & n274 ) | ( n273 & n274 ) ;
  assign n276 = x4 & x132 ;
  assign n277 = x4 | x132 ;
  assign n278 = n276 | n277 ;
  assign n279 = ( n272 & n276 ) | ( n272 & n278 ) | ( n276 & n278 ) ;
  assign n280 = ( x5 & ~x133 ) | ( x5 & n279 ) | ( ~x133 & n279 ) ;
  assign n281 = ( ~x5 & x133 ) | ( ~x5 & n280 ) | ( x133 & n280 ) ;
  assign n282 = ( ~n279 & n280 ) | ( ~n279 & n281 ) | ( n280 & n281 ) ;
  assign n283 = ( x5 & x133 ) | ( x5 & n279 ) | ( x133 & n279 ) ;
  assign n284 = ( x6 & ~x134 ) | ( x6 & n283 ) | ( ~x134 & n283 ) ;
  assign n285 = ( ~x6 & x134 ) | ( ~x6 & n284 ) | ( x134 & n284 ) ;
  assign n286 = ( ~n283 & n284 ) | ( ~n283 & n285 ) | ( n284 & n285 ) ;
  assign n287 = x6 & x134 ;
  assign n288 = x6 | x134 ;
  assign n289 = n287 | n288 ;
  assign n290 = ( n283 & n287 ) | ( n283 & n289 ) | ( n287 & n289 ) ;
  assign n291 = ( x7 & ~x135 ) | ( x7 & n290 ) | ( ~x135 & n290 ) ;
  assign n292 = ( ~x7 & x135 ) | ( ~x7 & n291 ) | ( x135 & n291 ) ;
  assign n293 = ( ~n290 & n291 ) | ( ~n290 & n292 ) | ( n291 & n292 ) ;
  assign n294 = ( x7 & x135 ) | ( x7 & n287 ) | ( x135 & n287 ) ;
  assign n295 = ( x7 & x135 ) | ( x7 & n289 ) | ( x135 & n289 ) ;
  assign n296 = ( n283 & n294 ) | ( n283 & n295 ) | ( n294 & n295 ) ;
  assign n297 = ( x8 & ~x136 ) | ( x8 & n296 ) | ( ~x136 & n296 ) ;
  assign n298 = ( ~x8 & x136 ) | ( ~x8 & n297 ) | ( x136 & n297 ) ;
  assign n299 = ( ~n296 & n297 ) | ( ~n296 & n298 ) | ( n297 & n298 ) ;
  assign n300 = x9 | x137 ;
  assign n301 = x9 & x137 ;
  assign n302 = x8 & x136 ;
  assign n303 = x8 | x136 ;
  assign n304 = n295 & n303 ;
  assign n305 = n294 & n303 ;
  assign n306 = ( n283 & n304 ) | ( n283 & n305 ) | ( n304 & n305 ) ;
  assign n307 = n302 | n306 ;
  assign n308 = ( ~n300 & n301 ) | ( ~n300 & n307 ) | ( n301 & n307 ) ;
  assign n309 = ( n300 & n301 ) | ( n300 & n307 ) | ( n301 & n307 ) ;
  assign n310 = ( n300 & n308 ) | ( n300 & ~n309 ) | ( n308 & ~n309 ) ;
  assign n311 = ( x10 & ~x138 ) | ( x10 & n309 ) | ( ~x138 & n309 ) ;
  assign n312 = ( ~x10 & x138 ) | ( ~x10 & n311 ) | ( x138 & n311 ) ;
  assign n313 = ( ~n309 & n311 ) | ( ~n309 & n312 ) | ( n311 & n312 ) ;
  assign n314 = x10 & x138 ;
  assign n315 = x10 | x138 ;
  assign n316 = ( n300 & n314 ) | ( n300 & n315 ) | ( n314 & n315 ) ;
  assign n317 = ( n302 & n314 ) | ( n302 & n316 ) | ( n314 & n316 ) ;
  assign n318 = ( n301 & n315 ) | ( n301 & n317 ) | ( n315 & n317 ) ;
  assign n319 = ( n306 & n316 ) | ( n306 & n318 ) | ( n316 & n318 ) ;
  assign n320 = ( x11 & ~x139 ) | ( x11 & n319 ) | ( ~x139 & n319 ) ;
  assign n321 = ( ~x11 & x139 ) | ( ~x11 & n320 ) | ( x139 & n320 ) ;
  assign n322 = ( ~n319 & n320 ) | ( ~n319 & n321 ) | ( n320 & n321 ) ;
  assign n323 = x12 | x140 ;
  assign n324 = x12 & x140 ;
  assign n325 = x11 & x139 ;
  assign n326 = x11 | x139 ;
  assign n327 = n316 & n326 ;
  assign n328 = n318 & n326 ;
  assign n329 = ( n306 & n327 ) | ( n306 & n328 ) | ( n327 & n328 ) ;
  assign n330 = n325 | n329 ;
  assign n331 = ( ~n323 & n324 ) | ( ~n323 & n330 ) | ( n324 & n330 ) ;
  assign n332 = ( n323 & n324 ) | ( n323 & n330 ) | ( n324 & n330 ) ;
  assign n333 = ( n323 & n331 ) | ( n323 & ~n332 ) | ( n331 & ~n332 ) ;
  assign n334 = ( x13 & ~x141 ) | ( x13 & n332 ) | ( ~x141 & n332 ) ;
  assign n335 = ( ~x13 & x141 ) | ( ~x13 & n334 ) | ( x141 & n334 ) ;
  assign n336 = ( ~n332 & n334 ) | ( ~n332 & n335 ) | ( n334 & n335 ) ;
  assign n337 = x13 & x141 ;
  assign n338 = x13 | x141 ;
  assign n339 = ( n323 & n337 ) | ( n323 & n338 ) | ( n337 & n338 ) ;
  assign n340 = ( n325 & n337 ) | ( n325 & n339 ) | ( n337 & n339 ) ;
  assign n341 = ( n324 & n338 ) | ( n324 & n340 ) | ( n338 & n340 ) ;
  assign n342 = ( n329 & n339 ) | ( n329 & n341 ) | ( n339 & n341 ) ;
  assign n343 = ( x14 & ~x142 ) | ( x14 & n342 ) | ( ~x142 & n342 ) ;
  assign n344 = ( ~x14 & x142 ) | ( ~x14 & n343 ) | ( x142 & n343 ) ;
  assign n345 = ( ~n342 & n343 ) | ( ~n342 & n344 ) | ( n343 & n344 ) ;
  assign n346 = ( x14 & x142 ) | ( x14 & n341 ) | ( x142 & n341 ) ;
  assign n347 = ( x14 & x142 ) | ( x14 & n339 ) | ( x142 & n339 ) ;
  assign n348 = ( n329 & n346 ) | ( n329 & n347 ) | ( n346 & n347 ) ;
  assign n349 = ( x15 & ~x143 ) | ( x15 & n348 ) | ( ~x143 & n348 ) ;
  assign n350 = ( ~x15 & x143 ) | ( ~x15 & n349 ) | ( x143 & n349 ) ;
  assign n351 = ( ~n348 & n349 ) | ( ~n348 & n350 ) | ( n349 & n350 ) ;
  assign n352 = x15 & x143 ;
  assign n353 = x15 | x143 ;
  assign n354 = n352 | n353 ;
  assign n355 = ( n348 & n352 ) | ( n348 & n354 ) | ( n352 & n354 ) ;
  assign n356 = ( x16 & ~x144 ) | ( x16 & n355 ) | ( ~x144 & n355 ) ;
  assign n357 = ( ~x16 & x144 ) | ( ~x16 & n356 ) | ( x144 & n356 ) ;
  assign n358 = ( ~n355 & n356 ) | ( ~n355 & n357 ) | ( n356 & n357 ) ;
  assign n359 = ( x16 & x144 ) | ( x16 & n352 ) | ( x144 & n352 ) ;
  assign n360 = ( x16 & x144 ) | ( x16 & n354 ) | ( x144 & n354 ) ;
  assign n361 = ( n348 & n359 ) | ( n348 & n360 ) | ( n359 & n360 ) ;
  assign n362 = ( x17 & ~x145 ) | ( x17 & n361 ) | ( ~x145 & n361 ) ;
  assign n363 = ( ~x17 & x145 ) | ( ~x17 & n362 ) | ( x145 & n362 ) ;
  assign n364 = ( ~n361 & n362 ) | ( ~n361 & n363 ) | ( n362 & n363 ) ;
  assign n365 = ( x17 & x145 ) | ( x17 & n359 ) | ( x145 & n359 ) ;
  assign n366 = x17 | x145 ;
  assign n367 = ( n360 & n365 ) | ( n360 & n366 ) | ( n365 & n366 ) ;
  assign n368 = ( n348 & n365 ) | ( n348 & n367 ) | ( n365 & n367 ) ;
  assign n369 = ( x18 & ~x146 ) | ( x18 & n368 ) | ( ~x146 & n368 ) ;
  assign n370 = ( ~x18 & x146 ) | ( ~x18 & n369 ) | ( x146 & n369 ) ;
  assign n371 = ( ~n368 & n369 ) | ( ~n368 & n370 ) | ( n369 & n370 ) ;
  assign n372 = x18 & x146 ;
  assign n373 = x18 | x146 ;
  assign n374 = n367 & n373 ;
  assign n375 = n372 | n374 ;
  assign n376 = ( x18 & x146 ) | ( x18 & n365 ) | ( x146 & n365 ) ;
  assign n377 = ( n348 & n375 ) | ( n348 & n376 ) | ( n375 & n376 ) ;
  assign n378 = ( x19 & ~x147 ) | ( x19 & n377 ) | ( ~x147 & n377 ) ;
  assign n379 = ( ~x19 & x147 ) | ( ~x19 & n378 ) | ( x147 & n378 ) ;
  assign n380 = ( ~n377 & n378 ) | ( ~n377 & n379 ) | ( n378 & n379 ) ;
  assign n381 = x19 & x147 ;
  assign n382 = x19 | x147 ;
  assign n383 = n381 | n382 ;
  assign n384 = ( n377 & n381 ) | ( n377 & n383 ) | ( n381 & n383 ) ;
  assign n385 = ( x20 & ~x148 ) | ( x20 & n384 ) | ( ~x148 & n384 ) ;
  assign n386 = ( ~x20 & x148 ) | ( ~x20 & n385 ) | ( x148 & n385 ) ;
  assign n387 = ( ~n384 & n385 ) | ( ~n384 & n386 ) | ( n385 & n386 ) ;
  assign n388 = ( x20 & x148 ) | ( x20 & n381 ) | ( x148 & n381 ) ;
  assign n389 = ( x20 & x148 ) | ( x20 & n383 ) | ( x148 & n383 ) ;
  assign n390 = ( n377 & n388 ) | ( n377 & n389 ) | ( n388 & n389 ) ;
  assign n391 = ( x21 & ~x149 ) | ( x21 & n390 ) | ( ~x149 & n390 ) ;
  assign n392 = ( ~x21 & x149 ) | ( ~x21 & n391 ) | ( x149 & n391 ) ;
  assign n393 = ( ~n390 & n391 ) | ( ~n390 & n392 ) | ( n391 & n392 ) ;
  assign n394 = ( x21 & x149 ) | ( x21 & n388 ) | ( x149 & n388 ) ;
  assign n395 = x21 | x149 ;
  assign n396 = ( n389 & n394 ) | ( n389 & n395 ) | ( n394 & n395 ) ;
  assign n397 = ( n377 & n394 ) | ( n377 & n396 ) | ( n394 & n396 ) ;
  assign n398 = ( x22 & ~x150 ) | ( x22 & n397 ) | ( ~x150 & n397 ) ;
  assign n399 = ( ~x22 & x150 ) | ( ~x22 & n398 ) | ( x150 & n398 ) ;
  assign n400 = ( ~n397 & n398 ) | ( ~n397 & n399 ) | ( n398 & n399 ) ;
  assign n401 = x22 & x150 ;
  assign n402 = x22 | x150 ;
  assign n403 = n396 & n402 ;
  assign n404 = n401 | n403 ;
  assign n405 = ( x22 & x150 ) | ( x22 & n394 ) | ( x150 & n394 ) ;
  assign n406 = ( n377 & n404 ) | ( n377 & n405 ) | ( n404 & n405 ) ;
  assign n407 = ( x23 & ~x151 ) | ( x23 & n406 ) | ( ~x151 & n406 ) ;
  assign n408 = ( ~x23 & x151 ) | ( ~x23 & n407 ) | ( x151 & n407 ) ;
  assign n409 = ( ~n406 & n407 ) | ( ~n406 & n408 ) | ( n407 & n408 ) ;
  assign n410 = x24 | x152 ;
  assign n411 = x24 & x152 ;
  assign n412 = x23 & x151 ;
  assign n413 = x23 | x151 ;
  assign n414 = n405 & n413 ;
  assign n415 = n404 & n413 ;
  assign n416 = ( n377 & n414 ) | ( n377 & n415 ) | ( n414 & n415 ) ;
  assign n417 = n412 | n416 ;
  assign n418 = ( ~n410 & n411 ) | ( ~n410 & n417 ) | ( n411 & n417 ) ;
  assign n419 = ( n410 & n411 ) | ( n410 & n417 ) | ( n411 & n417 ) ;
  assign n420 = ( n410 & n418 ) | ( n410 & ~n419 ) | ( n418 & ~n419 ) ;
  assign n421 = ( x25 & ~x153 ) | ( x25 & n419 ) | ( ~x153 & n419 ) ;
  assign n422 = ( ~x25 & x153 ) | ( ~x25 & n421 ) | ( x153 & n421 ) ;
  assign n423 = ( ~n419 & n421 ) | ( ~n419 & n422 ) | ( n421 & n422 ) ;
  assign n424 = x25 & x153 ;
  assign n425 = x25 | x153 ;
  assign n426 = ( n410 & n424 ) | ( n410 & n425 ) | ( n424 & n425 ) ;
  assign n427 = ( n412 & n424 ) | ( n412 & n426 ) | ( n424 & n426 ) ;
  assign n428 = ( n411 & n425 ) | ( n411 & n427 ) | ( n425 & n427 ) ;
  assign n429 = ( n416 & n426 ) | ( n416 & n428 ) | ( n426 & n428 ) ;
  assign n430 = ( x26 & ~x154 ) | ( x26 & n429 ) | ( ~x154 & n429 ) ;
  assign n431 = ( ~x26 & x154 ) | ( ~x26 & n430 ) | ( x154 & n430 ) ;
  assign n432 = ( ~n429 & n430 ) | ( ~n429 & n431 ) | ( n430 & n431 ) ;
  assign n433 = ( x26 & x154 ) | ( x26 & n428 ) | ( x154 & n428 ) ;
  assign n434 = ( x26 & x154 ) | ( x26 & n426 ) | ( x154 & n426 ) ;
  assign n435 = ( n416 & n433 ) | ( n416 & n434 ) | ( n433 & n434 ) ;
  assign n436 = ( x27 & ~x155 ) | ( x27 & n435 ) | ( ~x155 & n435 ) ;
  assign n437 = ( ~x27 & x155 ) | ( ~x27 & n436 ) | ( x155 & n436 ) ;
  assign n438 = ( ~n435 & n436 ) | ( ~n435 & n437 ) | ( n436 & n437 ) ;
  assign n439 = x27 & x155 ;
  assign n440 = x27 | x155 ;
  assign n441 = n434 & n440 ;
  assign n442 = n439 | n441 ;
  assign n443 = ( n433 & n439 ) | ( n433 & n440 ) | ( n439 & n440 ) ;
  assign n444 = ( n416 & n442 ) | ( n416 & n443 ) | ( n442 & n443 ) ;
  assign n445 = ( x28 & ~x156 ) | ( x28 & n444 ) | ( ~x156 & n444 ) ;
  assign n446 = ( ~x28 & x156 ) | ( ~x28 & n445 ) | ( x156 & n445 ) ;
  assign n447 = ( ~n444 & n445 ) | ( ~n444 & n446 ) | ( n445 & n446 ) ;
  assign n448 = x29 | x157 ;
  assign n449 = x29 & x157 ;
  assign n450 = x28 & x156 ;
  assign n451 = x28 | x156 ;
  assign n452 = n443 & n451 ;
  assign n453 = n442 & n451 ;
  assign n454 = ( n415 & n452 ) | ( n415 & n453 ) | ( n452 & n453 ) ;
  assign n455 = ( n414 & n452 ) | ( n414 & n453 ) | ( n452 & n453 ) ;
  assign n456 = ( n377 & n454 ) | ( n377 & n455 ) | ( n454 & n455 ) ;
  assign n457 = n450 | n456 ;
  assign n458 = ( ~n448 & n449 ) | ( ~n448 & n457 ) | ( n449 & n457 ) ;
  assign n459 = ( n448 & n449 ) | ( n448 & n457 ) | ( n449 & n457 ) ;
  assign n460 = ( n448 & n458 ) | ( n448 & ~n459 ) | ( n458 & ~n459 ) ;
  assign n461 = ( x30 & ~x158 ) | ( x30 & n459 ) | ( ~x158 & n459 ) ;
  assign n462 = ( ~x30 & x158 ) | ( ~x30 & n461 ) | ( x158 & n461 ) ;
  assign n463 = ( ~n459 & n461 ) | ( ~n459 & n462 ) | ( n461 & n462 ) ;
  assign n464 = x30 & x158 ;
  assign n465 = x30 | x158 ;
  assign n466 = ( n448 & n464 ) | ( n448 & n465 ) | ( n464 & n465 ) ;
  assign n467 = ( n450 & n464 ) | ( n450 & n466 ) | ( n464 & n466 ) ;
  assign n468 = ( n449 & n465 ) | ( n449 & n467 ) | ( n465 & n467 ) ;
  assign n469 = ( n456 & n466 ) | ( n456 & n468 ) | ( n466 & n468 ) ;
  assign n470 = ( x31 & ~x159 ) | ( x31 & n469 ) | ( ~x159 & n469 ) ;
  assign n471 = ( ~x31 & x159 ) | ( ~x31 & n470 ) | ( x159 & n470 ) ;
  assign n472 = ( ~n469 & n470 ) | ( ~n469 & n471 ) | ( n470 & n471 ) ;
  assign n473 = ( x31 & x159 ) | ( x31 & n468 ) | ( x159 & n468 ) ;
  assign n474 = ( x31 & x159 ) | ( x31 & n466 ) | ( x159 & n466 ) ;
  assign n475 = ( n456 & n473 ) | ( n456 & n474 ) | ( n473 & n474 ) ;
  assign n476 = ( x32 & ~x160 ) | ( x32 & n475 ) | ( ~x160 & n475 ) ;
  assign n477 = ( ~x32 & x160 ) | ( ~x32 & n476 ) | ( x160 & n476 ) ;
  assign n478 = ( ~n475 & n476 ) | ( ~n475 & n477 ) | ( n476 & n477 ) ;
  assign n479 = x32 & x160 ;
  assign n480 = x32 | x160 ;
  assign n481 = n474 & n480 ;
  assign n482 = n479 | n481 ;
  assign n483 = ( n473 & n479 ) | ( n473 & n480 ) | ( n479 & n480 ) ;
  assign n484 = ( n456 & n482 ) | ( n456 & n483 ) | ( n482 & n483 ) ;
  assign n485 = ( x33 & ~x161 ) | ( x33 & n484 ) | ( ~x161 & n484 ) ;
  assign n486 = ( ~x33 & x161 ) | ( ~x33 & n485 ) | ( x161 & n485 ) ;
  assign n487 = ( ~n484 & n485 ) | ( ~n484 & n486 ) | ( n485 & n486 ) ;
  assign n488 = ( x33 & x161 ) | ( x33 & n480 ) | ( x161 & n480 ) ;
  assign n489 = ( x33 & x161 ) | ( x33 & n479 ) | ( x161 & n479 ) ;
  assign n490 = ( n473 & n488 ) | ( n473 & n489 ) | ( n488 & n489 ) ;
  assign n491 = ( x33 & x161 ) | ( x33 & n482 ) | ( x161 & n482 ) ;
  assign n492 = ( n456 & n490 ) | ( n456 & n491 ) | ( n490 & n491 ) ;
  assign n493 = ( x34 & ~x162 ) | ( x34 & n492 ) | ( ~x162 & n492 ) ;
  assign n494 = ( ~x34 & x162 ) | ( ~x34 & n493 ) | ( x162 & n493 ) ;
  assign n495 = ( ~n492 & n493 ) | ( ~n492 & n494 ) | ( n493 & n494 ) ;
  assign n496 = x34 & x162 ;
  assign n497 = x34 | x162 ;
  assign n498 = n496 | n497 ;
  assign n499 = ( n492 & n496 ) | ( n492 & n498 ) | ( n496 & n498 ) ;
  assign n500 = ( x35 & ~x163 ) | ( x35 & n499 ) | ( ~x163 & n499 ) ;
  assign n501 = ( ~x35 & x163 ) | ( ~x35 & n500 ) | ( x163 & n500 ) ;
  assign n502 = ( ~n499 & n500 ) | ( ~n499 & n501 ) | ( n500 & n501 ) ;
  assign n503 = ( x35 & x163 ) | ( x35 & n496 ) | ( x163 & n496 ) ;
  assign n504 = ( x35 & x163 ) | ( x35 & n498 ) | ( x163 & n498 ) ;
  assign n505 = ( n492 & n503 ) | ( n492 & n504 ) | ( n503 & n504 ) ;
  assign n506 = ( x36 & ~x164 ) | ( x36 & n505 ) | ( ~x164 & n505 ) ;
  assign n507 = ( ~x36 & x164 ) | ( ~x36 & n506 ) | ( x164 & n506 ) ;
  assign n508 = ( ~n505 & n506 ) | ( ~n505 & n507 ) | ( n506 & n507 ) ;
  assign n509 = ( x36 & x164 ) | ( x36 & n503 ) | ( x164 & n503 ) ;
  assign n510 = x36 | x164 ;
  assign n511 = ( n504 & n509 ) | ( n504 & n510 ) | ( n509 & n510 ) ;
  assign n512 = ( n492 & n509 ) | ( n492 & n511 ) | ( n509 & n511 ) ;
  assign n513 = ( x37 & ~x165 ) | ( x37 & n512 ) | ( ~x165 & n512 ) ;
  assign n514 = ( ~x37 & x165 ) | ( ~x37 & n513 ) | ( x165 & n513 ) ;
  assign n515 = ( ~n512 & n513 ) | ( ~n512 & n514 ) | ( n513 & n514 ) ;
  assign n516 = x37 & x165 ;
  assign n517 = x37 | x165 ;
  assign n518 = n511 & n517 ;
  assign n519 = n516 | n518 ;
  assign n520 = ( x37 & x165 ) | ( x37 & n509 ) | ( x165 & n509 ) ;
  assign n521 = ( n492 & n519 ) | ( n492 & n520 ) | ( n519 & n520 ) ;
  assign n522 = ( x38 & ~x166 ) | ( x38 & n521 ) | ( ~x166 & n521 ) ;
  assign n523 = ( ~x38 & x166 ) | ( ~x38 & n522 ) | ( x166 & n522 ) ;
  assign n524 = ( ~n521 & n522 ) | ( ~n521 & n523 ) | ( n522 & n523 ) ;
  assign n525 = x38 & x166 ;
  assign n526 = x38 | x166 ;
  assign n527 = n525 | n526 ;
  assign n528 = ( n520 & n525 ) | ( n520 & n527 ) | ( n525 & n527 ) ;
  assign n529 = ( x38 & x166 ) | ( x38 & n519 ) | ( x166 & n519 ) ;
  assign n530 = ( n492 & n528 ) | ( n492 & n529 ) | ( n528 & n529 ) ;
  assign n531 = ( x39 & ~x167 ) | ( x39 & n530 ) | ( ~x167 & n530 ) ;
  assign n532 = ( ~x39 & x167 ) | ( ~x39 & n531 ) | ( x167 & n531 ) ;
  assign n533 = ( ~n530 & n531 ) | ( ~n530 & n532 ) | ( n531 & n532 ) ;
  assign n534 = x39 & x167 ;
  assign n535 = x39 | x167 ;
  assign n536 = n528 & n535 ;
  assign n537 = n534 | n536 ;
  assign n538 = ( x39 & x167 ) | ( x39 & n529 ) | ( x167 & n529 ) ;
  assign n539 = ( n492 & n537 ) | ( n492 & n538 ) | ( n537 & n538 ) ;
  assign n540 = ( x40 & ~x168 ) | ( x40 & n539 ) | ( ~x168 & n539 ) ;
  assign n541 = ( ~x40 & x168 ) | ( ~x40 & n540 ) | ( x168 & n540 ) ;
  assign n542 = ( ~n539 & n540 ) | ( ~n539 & n541 ) | ( n540 & n541 ) ;
  assign n543 = x40 & x168 ;
  assign n544 = x40 | x168 ;
  assign n545 = n543 | n544 ;
  assign n546 = ( n539 & n543 ) | ( n539 & n545 ) | ( n543 & n545 ) ;
  assign n547 = ( x41 & ~x169 ) | ( x41 & n546 ) | ( ~x169 & n546 ) ;
  assign n548 = ( ~x41 & x169 ) | ( ~x41 & n547 ) | ( x169 & n547 ) ;
  assign n549 = ( ~n546 & n547 ) | ( ~n546 & n548 ) | ( n547 & n548 ) ;
  assign n550 = ( x41 & x169 ) | ( x41 & n543 ) | ( x169 & n543 ) ;
  assign n551 = ( x41 & x169 ) | ( x41 & n545 ) | ( x169 & n545 ) ;
  assign n552 = ( n539 & n550 ) | ( n539 & n551 ) | ( n550 & n551 ) ;
  assign n553 = ( x42 & ~x170 ) | ( x42 & n552 ) | ( ~x170 & n552 ) ;
  assign n554 = ( ~x42 & x170 ) | ( ~x42 & n553 ) | ( x170 & n553 ) ;
  assign n555 = ( ~n552 & n553 ) | ( ~n552 & n554 ) | ( n553 & n554 ) ;
  assign n556 = ( x42 & x170 ) | ( x42 & n550 ) | ( x170 & n550 ) ;
  assign n557 = x42 | x170 ;
  assign n558 = ( n551 & n556 ) | ( n551 & n557 ) | ( n556 & n557 ) ;
  assign n559 = ( n539 & n556 ) | ( n539 & n558 ) | ( n556 & n558 ) ;
  assign n560 = ( x43 & ~x171 ) | ( x43 & n559 ) | ( ~x171 & n559 ) ;
  assign n561 = ( ~x43 & x171 ) | ( ~x43 & n560 ) | ( x171 & n560 ) ;
  assign n562 = ( ~n559 & n560 ) | ( ~n559 & n561 ) | ( n560 & n561 ) ;
  assign n563 = x43 & x171 ;
  assign n564 = x43 | x171 ;
  assign n565 = n558 & n564 ;
  assign n566 = n563 | n565 ;
  assign n567 = ( x43 & x171 ) | ( x43 & n556 ) | ( x171 & n556 ) ;
  assign n568 = ( n539 & n566 ) | ( n539 & n567 ) | ( n566 & n567 ) ;
  assign n569 = ( x44 & ~x172 ) | ( x44 & n568 ) | ( ~x172 & n568 ) ;
  assign n570 = ( ~x44 & x172 ) | ( ~x44 & n569 ) | ( x172 & n569 ) ;
  assign n571 = ( ~n568 & n569 ) | ( ~n568 & n570 ) | ( n569 & n570 ) ;
  assign n572 = x44 & x172 ;
  assign n573 = x44 | x172 ;
  assign n574 = n572 | n573 ;
  assign n575 = ( n567 & n572 ) | ( n567 & n574 ) | ( n572 & n574 ) ;
  assign n576 = ( x44 & x172 ) | ( x44 & n566 ) | ( x172 & n566 ) ;
  assign n577 = ( n539 & n575 ) | ( n539 & n576 ) | ( n575 & n576 ) ;
  assign n578 = ( x45 & ~x173 ) | ( x45 & n577 ) | ( ~x173 & n577 ) ;
  assign n579 = ( ~x45 & x173 ) | ( ~x45 & n578 ) | ( x173 & n578 ) ;
  assign n580 = ( ~n577 & n578 ) | ( ~n577 & n579 ) | ( n578 & n579 ) ;
  assign n581 = x45 & x173 ;
  assign n582 = x45 | x173 ;
  assign n583 = n575 & n582 ;
  assign n584 = n581 | n583 ;
  assign n585 = ( x45 & x173 ) | ( x45 & n576 ) | ( x173 & n576 ) ;
  assign n586 = ( n539 & n584 ) | ( n539 & n585 ) | ( n584 & n585 ) ;
  assign n587 = ( x46 & ~x174 ) | ( x46 & n586 ) | ( ~x174 & n586 ) ;
  assign n588 = ( ~x46 & x174 ) | ( ~x46 & n587 ) | ( x174 & n587 ) ;
  assign n589 = ( ~n586 & n587 ) | ( ~n586 & n588 ) | ( n587 & n588 ) ;
  assign n590 = x47 | x175 ;
  assign n591 = x47 & x175 ;
  assign n592 = x46 & x174 ;
  assign n593 = x46 | x174 ;
  assign n594 = n584 & n593 ;
  assign n595 = n585 & n593 ;
  assign n596 = ( n539 & n594 ) | ( n539 & n595 ) | ( n594 & n595 ) ;
  assign n597 = n592 | n596 ;
  assign n598 = ( ~n590 & n591 ) | ( ~n590 & n597 ) | ( n591 & n597 ) ;
  assign n599 = ( n590 & n591 ) | ( n590 & n597 ) | ( n591 & n597 ) ;
  assign n600 = ( n590 & n598 ) | ( n590 & ~n599 ) | ( n598 & ~n599 ) ;
  assign n601 = ( x48 & ~x176 ) | ( x48 & n599 ) | ( ~x176 & n599 ) ;
  assign n602 = ( ~x48 & x176 ) | ( ~x48 & n601 ) | ( x176 & n601 ) ;
  assign n603 = ( ~n599 & n601 ) | ( ~n599 & n602 ) | ( n601 & n602 ) ;
  assign n604 = x48 & x176 ;
  assign n605 = x48 | x176 ;
  assign n606 = ( n590 & n604 ) | ( n590 & n605 ) | ( n604 & n605 ) ;
  assign n607 = ( n592 & n604 ) | ( n592 & n606 ) | ( n604 & n606 ) ;
  assign n608 = ( n591 & n605 ) | ( n591 & n607 ) | ( n605 & n607 ) ;
  assign n609 = ( n596 & n606 ) | ( n596 & n608 ) | ( n606 & n608 ) ;
  assign n610 = ( x49 & ~x177 ) | ( x49 & n609 ) | ( ~x177 & n609 ) ;
  assign n611 = ( ~x49 & x177 ) | ( ~x49 & n610 ) | ( x177 & n610 ) ;
  assign n612 = ( ~n609 & n610 ) | ( ~n609 & n611 ) | ( n610 & n611 ) ;
  assign n613 = ( x49 & x177 ) | ( x49 & n608 ) | ( x177 & n608 ) ;
  assign n614 = ( x49 & x177 ) | ( x49 & n606 ) | ( x177 & n606 ) ;
  assign n615 = ( n596 & n613 ) | ( n596 & n614 ) | ( n613 & n614 ) ;
  assign n616 = ( x50 & ~x178 ) | ( x50 & n615 ) | ( ~x178 & n615 ) ;
  assign n617 = ( ~x50 & x178 ) | ( ~x50 & n616 ) | ( x178 & n616 ) ;
  assign n618 = ( ~n615 & n616 ) | ( ~n615 & n617 ) | ( n616 & n617 ) ;
  assign n619 = x50 & x178 ;
  assign n620 = x50 | x178 ;
  assign n621 = n614 & n620 ;
  assign n622 = n619 | n621 ;
  assign n623 = ( n613 & n619 ) | ( n613 & n620 ) | ( n619 & n620 ) ;
  assign n624 = ( n596 & n622 ) | ( n596 & n623 ) | ( n622 & n623 ) ;
  assign n625 = ( x51 & ~x179 ) | ( x51 & n624 ) | ( ~x179 & n624 ) ;
  assign n626 = ( ~x51 & x179 ) | ( ~x51 & n625 ) | ( x179 & n625 ) ;
  assign n627 = ( ~n624 & n625 ) | ( ~n624 & n626 ) | ( n625 & n626 ) ;
  assign n628 = ( x51 & x179 ) | ( x51 & n620 ) | ( x179 & n620 ) ;
  assign n629 = ( x51 & x179 ) | ( x51 & n619 ) | ( x179 & n619 ) ;
  assign n630 = ( n613 & n628 ) | ( n613 & n629 ) | ( n628 & n629 ) ;
  assign n631 = ( x51 & x179 ) | ( x51 & n622 ) | ( x179 & n622 ) ;
  assign n632 = ( n596 & n630 ) | ( n596 & n631 ) | ( n630 & n631 ) ;
  assign n633 = ( x52 & ~x180 ) | ( x52 & n632 ) | ( ~x180 & n632 ) ;
  assign n634 = ( ~x52 & x180 ) | ( ~x52 & n633 ) | ( x180 & n633 ) ;
  assign n635 = ( ~n632 & n633 ) | ( ~n632 & n634 ) | ( n633 & n634 ) ;
  assign n636 = x52 & x180 ;
  assign n637 = x52 | x180 ;
  assign n638 = n631 & n637 ;
  assign n639 = n636 | n638 ;
  assign n640 = ( n630 & n636 ) | ( n630 & n637 ) | ( n636 & n637 ) ;
  assign n641 = ( n596 & n639 ) | ( n596 & n640 ) | ( n639 & n640 ) ;
  assign n642 = ( x53 & ~x181 ) | ( x53 & n641 ) | ( ~x181 & n641 ) ;
  assign n643 = ( ~x53 & x181 ) | ( ~x53 & n642 ) | ( x181 & n642 ) ;
  assign n644 = ( ~n641 & n642 ) | ( ~n641 & n643 ) | ( n642 & n643 ) ;
  assign n645 = x54 | x182 ;
  assign n646 = x54 & x182 ;
  assign n647 = x53 & x181 ;
  assign n648 = x53 | x181 ;
  assign n649 = n640 & n648 ;
  assign n650 = n639 & n648 ;
  assign n651 = ( n596 & n649 ) | ( n596 & n650 ) | ( n649 & n650 ) ;
  assign n652 = n647 | n651 ;
  assign n653 = ( ~n645 & n646 ) | ( ~n645 & n652 ) | ( n646 & n652 ) ;
  assign n654 = ( n645 & n646 ) | ( n645 & n652 ) | ( n646 & n652 ) ;
  assign n655 = ( n645 & n653 ) | ( n645 & ~n654 ) | ( n653 & ~n654 ) ;
  assign n656 = ( x55 & ~x183 ) | ( x55 & n654 ) | ( ~x183 & n654 ) ;
  assign n657 = ( ~x55 & x183 ) | ( ~x55 & n656 ) | ( x183 & n656 ) ;
  assign n658 = ( ~n654 & n656 ) | ( ~n654 & n657 ) | ( n656 & n657 ) ;
  assign n659 = x55 & x183 ;
  assign n660 = x55 | x183 ;
  assign n661 = ( n645 & n659 ) | ( n645 & n660 ) | ( n659 & n660 ) ;
  assign n662 = ( n647 & n659 ) | ( n647 & n661 ) | ( n659 & n661 ) ;
  assign n663 = ( n646 & n660 ) | ( n646 & n662 ) | ( n660 & n662 ) ;
  assign n664 = ( n651 & n661 ) | ( n651 & n663 ) | ( n661 & n663 ) ;
  assign n665 = ( x56 & ~x184 ) | ( x56 & n664 ) | ( ~x184 & n664 ) ;
  assign n666 = ( ~x56 & x184 ) | ( ~x56 & n665 ) | ( x184 & n665 ) ;
  assign n667 = ( ~n664 & n665 ) | ( ~n664 & n666 ) | ( n665 & n666 ) ;
  assign n668 = ( x56 & x184 ) | ( x56 & n663 ) | ( x184 & n663 ) ;
  assign n669 = ( x56 & x184 ) | ( x56 & n661 ) | ( x184 & n661 ) ;
  assign n670 = ( n651 & n668 ) | ( n651 & n669 ) | ( n668 & n669 ) ;
  assign n671 = ( x57 & ~x185 ) | ( x57 & n670 ) | ( ~x185 & n670 ) ;
  assign n672 = ( ~x57 & x185 ) | ( ~x57 & n671 ) | ( x185 & n671 ) ;
  assign n673 = ( ~n670 & n671 ) | ( ~n670 & n672 ) | ( n671 & n672 ) ;
  assign n674 = x57 & x185 ;
  assign n675 = x57 | x185 ;
  assign n676 = n669 & n675 ;
  assign n677 = n674 | n676 ;
  assign n678 = ( n668 & n674 ) | ( n668 & n675 ) | ( n674 & n675 ) ;
  assign n679 = ( n651 & n677 ) | ( n651 & n678 ) | ( n677 & n678 ) ;
  assign n680 = ( x58 & ~x186 ) | ( x58 & n679 ) | ( ~x186 & n679 ) ;
  assign n681 = ( ~x58 & x186 ) | ( ~x58 & n680 ) | ( x186 & n680 ) ;
  assign n682 = ( ~n679 & n680 ) | ( ~n679 & n681 ) | ( n680 & n681 ) ;
  assign n683 = ( x58 & x186 ) | ( x58 & n675 ) | ( x186 & n675 ) ;
  assign n684 = ( x58 & x186 ) | ( x58 & n674 ) | ( x186 & n674 ) ;
  assign n685 = ( n668 & n683 ) | ( n668 & n684 ) | ( n683 & n684 ) ;
  assign n686 = ( x58 & x186 ) | ( x58 & n677 ) | ( x186 & n677 ) ;
  assign n687 = ( n651 & n685 ) | ( n651 & n686 ) | ( n685 & n686 ) ;
  assign n688 = ( x59 & ~x187 ) | ( x59 & n687 ) | ( ~x187 & n687 ) ;
  assign n689 = ( ~x59 & x187 ) | ( ~x59 & n688 ) | ( x187 & n688 ) ;
  assign n690 = ( ~n687 & n688 ) | ( ~n687 & n689 ) | ( n688 & n689 ) ;
  assign n691 = x59 & x187 ;
  assign n692 = x59 | x187 ;
  assign n693 = n686 & n692 ;
  assign n694 = n691 | n693 ;
  assign n695 = ( n685 & n691 ) | ( n685 & n692 ) | ( n691 & n692 ) ;
  assign n696 = ( n651 & n694 ) | ( n651 & n695 ) | ( n694 & n695 ) ;
  assign n697 = ( x60 & ~x188 ) | ( x60 & n696 ) | ( ~x188 & n696 ) ;
  assign n698 = ( ~x60 & x188 ) | ( ~x60 & n697 ) | ( x188 & n697 ) ;
  assign n699 = ( ~n696 & n697 ) | ( ~n696 & n698 ) | ( n697 & n698 ) ;
  assign n700 = ( x60 & x188 ) | ( x60 & n692 ) | ( x188 & n692 ) ;
  assign n701 = ( x60 & x188 ) | ( x60 & n691 ) | ( x188 & n691 ) ;
  assign n702 = ( n685 & n700 ) | ( n685 & n701 ) | ( n700 & n701 ) ;
  assign n703 = ( x60 & x188 ) | ( x60 & n694 ) | ( x188 & n694 ) ;
  assign n704 = ( n651 & n702 ) | ( n651 & n703 ) | ( n702 & n703 ) ;
  assign n705 = ( x61 & ~x189 ) | ( x61 & n704 ) | ( ~x189 & n704 ) ;
  assign n706 = ( ~x61 & x189 ) | ( ~x61 & n705 ) | ( x189 & n705 ) ;
  assign n707 = ( ~n704 & n705 ) | ( ~n704 & n706 ) | ( n705 & n706 ) ;
  assign n708 = x61 & x189 ;
  assign n709 = x61 | x189 ;
  assign n710 = n708 | n709 ;
  assign n711 = ( n704 & n708 ) | ( n704 & n710 ) | ( n708 & n710 ) ;
  assign n712 = ( x62 & ~x190 ) | ( x62 & n711 ) | ( ~x190 & n711 ) ;
  assign n713 = ( ~x62 & x190 ) | ( ~x62 & n712 ) | ( x190 & n712 ) ;
  assign n714 = ( ~n711 & n712 ) | ( ~n711 & n713 ) | ( n712 & n713 ) ;
  assign n715 = ( x62 & x190 ) | ( x62 & n708 ) | ( x190 & n708 ) ;
  assign n716 = ( x62 & x190 ) | ( x62 & n710 ) | ( x190 & n710 ) ;
  assign n717 = ( n704 & n715 ) | ( n704 & n716 ) | ( n715 & n716 ) ;
  assign n718 = ( x63 & ~x191 ) | ( x63 & n717 ) | ( ~x191 & n717 ) ;
  assign n719 = ( ~x63 & x191 ) | ( ~x63 & n718 ) | ( x191 & n718 ) ;
  assign n720 = ( ~n717 & n718 ) | ( ~n717 & n719 ) | ( n718 & n719 ) ;
  assign n721 = ( x63 & x191 ) | ( x63 & n715 ) | ( x191 & n715 ) ;
  assign n722 = x63 | x191 ;
  assign n723 = ( n716 & n721 ) | ( n716 & n722 ) | ( n721 & n722 ) ;
  assign n724 = ( n704 & n721 ) | ( n704 & n723 ) | ( n721 & n723 ) ;
  assign n725 = ( x64 & ~x192 ) | ( x64 & n724 ) | ( ~x192 & n724 ) ;
  assign n726 = ( ~x64 & x192 ) | ( ~x64 & n725 ) | ( x192 & n725 ) ;
  assign n727 = ( ~n724 & n725 ) | ( ~n724 & n726 ) | ( n725 & n726 ) ;
  assign n728 = x64 & x192 ;
  assign n729 = x64 | x192 ;
  assign n730 = n723 & n729 ;
  assign n731 = n728 | n730 ;
  assign n732 = ( x64 & x192 ) | ( x64 & n721 ) | ( x192 & n721 ) ;
  assign n733 = ( n704 & n731 ) | ( n704 & n732 ) | ( n731 & n732 ) ;
  assign n734 = ( x65 & ~x193 ) | ( x65 & n733 ) | ( ~x193 & n733 ) ;
  assign n735 = ( ~x65 & x193 ) | ( ~x65 & n734 ) | ( x193 & n734 ) ;
  assign n736 = ( ~n733 & n734 ) | ( ~n733 & n735 ) | ( n734 & n735 ) ;
  assign n737 = x65 & x193 ;
  assign n738 = x65 | x193 ;
  assign n739 = n737 | n738 ;
  assign n740 = ( n732 & n737 ) | ( n732 & n739 ) | ( n737 & n739 ) ;
  assign n741 = ( x65 & x193 ) | ( x65 & n731 ) | ( x193 & n731 ) ;
  assign n742 = ( n704 & n740 ) | ( n704 & n741 ) | ( n740 & n741 ) ;
  assign n743 = ( x66 & ~x194 ) | ( x66 & n742 ) | ( ~x194 & n742 ) ;
  assign n744 = ( ~x66 & x194 ) | ( ~x66 & n743 ) | ( x194 & n743 ) ;
  assign n745 = ( ~n742 & n743 ) | ( ~n742 & n744 ) | ( n743 & n744 ) ;
  assign n746 = x66 & x194 ;
  assign n747 = x66 | x194 ;
  assign n748 = n741 & n747 ;
  assign n749 = n746 | n748 ;
  assign n750 = n740 & n747 ;
  assign n751 = n746 | n750 ;
  assign n752 = ( n704 & n749 ) | ( n704 & n751 ) | ( n749 & n751 ) ;
  assign n753 = ( x67 & ~x195 ) | ( x67 & n752 ) | ( ~x195 & n752 ) ;
  assign n754 = ( ~x67 & x195 ) | ( ~x67 & n753 ) | ( x195 & n753 ) ;
  assign n755 = ( ~n752 & n753 ) | ( ~n752 & n754 ) | ( n753 & n754 ) ;
  assign n756 = x67 | x195 ;
  assign n757 = ( x67 & x195 ) | ( x67 & n746 ) | ( x195 & n746 ) ;
  assign n758 = ( n748 & n756 ) | ( n748 & n757 ) | ( n756 & n757 ) ;
  assign n759 = x67 & x195 ;
  assign n760 = ( n751 & n756 ) | ( n751 & n759 ) | ( n756 & n759 ) ;
  assign n761 = ( n704 & n758 ) | ( n704 & n760 ) | ( n758 & n760 ) ;
  assign n762 = ( x68 & ~x196 ) | ( x68 & n761 ) | ( ~x196 & n761 ) ;
  assign n763 = ( ~x68 & x196 ) | ( ~x68 & n762 ) | ( x196 & n762 ) ;
  assign n764 = ( ~n761 & n762 ) | ( ~n761 & n763 ) | ( n762 & n763 ) ;
  assign n765 = ( x68 & x196 ) | ( x68 & n757 ) | ( x196 & n757 ) ;
  assign n766 = ( x68 & x196 ) | ( x68 & n756 ) | ( x196 & n756 ) ;
  assign n767 = ( n748 & n765 ) | ( n748 & n766 ) | ( n765 & n766 ) ;
  assign n768 = ( x68 & x196 ) | ( x68 & n759 ) | ( x196 & n759 ) ;
  assign n769 = ( n751 & n766 ) | ( n751 & n768 ) | ( n766 & n768 ) ;
  assign n770 = ( n703 & n767 ) | ( n703 & n769 ) | ( n767 & n769 ) ;
  assign n771 = ( n702 & n767 ) | ( n702 & n769 ) | ( n767 & n769 ) ;
  assign n772 = ( n651 & n770 ) | ( n651 & n771 ) | ( n770 & n771 ) ;
  assign n773 = ( x69 & ~x197 ) | ( x69 & n772 ) | ( ~x197 & n772 ) ;
  assign n774 = ( ~x69 & x197 ) | ( ~x69 & n773 ) | ( x197 & n773 ) ;
  assign n775 = ( ~n772 & n773 ) | ( ~n772 & n774 ) | ( n773 & n774 ) ;
  assign n776 = x69 & x197 ;
  assign n777 = x69 | x197 ;
  assign n778 = n776 | n777 ;
  assign n779 = ( n772 & n776 ) | ( n772 & n778 ) | ( n776 & n778 ) ;
  assign n780 = ( x70 & ~x198 ) | ( x70 & n779 ) | ( ~x198 & n779 ) ;
  assign n781 = ( ~x70 & x198 ) | ( ~x70 & n780 ) | ( x198 & n780 ) ;
  assign n782 = ( ~n779 & n780 ) | ( ~n779 & n781 ) | ( n780 & n781 ) ;
  assign n783 = ( x70 & x198 ) | ( x70 & n776 ) | ( x198 & n776 ) ;
  assign n784 = ( x70 & x198 ) | ( x70 & n778 ) | ( x198 & n778 ) ;
  assign n785 = ( n772 & n783 ) | ( n772 & n784 ) | ( n783 & n784 ) ;
  assign n786 = ( x71 & ~x199 ) | ( x71 & n785 ) | ( ~x199 & n785 ) ;
  assign n787 = ( ~x71 & x199 ) | ( ~x71 & n786 ) | ( x199 & n786 ) ;
  assign n788 = ( ~n785 & n786 ) | ( ~n785 & n787 ) | ( n786 & n787 ) ;
  assign n789 = ( x71 & x199 ) | ( x71 & n783 ) | ( x199 & n783 ) ;
  assign n790 = x71 | x199 ;
  assign n791 = ( n784 & n789 ) | ( n784 & n790 ) | ( n789 & n790 ) ;
  assign n792 = ( n772 & n789 ) | ( n772 & n791 ) | ( n789 & n791 ) ;
  assign n793 = ( x72 & ~x200 ) | ( x72 & n792 ) | ( ~x200 & n792 ) ;
  assign n794 = ( ~x72 & x200 ) | ( ~x72 & n793 ) | ( x200 & n793 ) ;
  assign n795 = ( ~n792 & n793 ) | ( ~n792 & n794 ) | ( n793 & n794 ) ;
  assign n796 = x72 & x200 ;
  assign n797 = x72 | x200 ;
  assign n798 = n791 & n797 ;
  assign n799 = n796 | n798 ;
  assign n800 = ( x72 & x200 ) | ( x72 & n789 ) | ( x200 & n789 ) ;
  assign n801 = ( n772 & n799 ) | ( n772 & n800 ) | ( n799 & n800 ) ;
  assign n802 = ( x73 & ~x201 ) | ( x73 & n801 ) | ( ~x201 & n801 ) ;
  assign n803 = ( ~x73 & x201 ) | ( ~x73 & n802 ) | ( x201 & n802 ) ;
  assign n804 = ( ~n801 & n802 ) | ( ~n801 & n803 ) | ( n802 & n803 ) ;
  assign n805 = x73 & x201 ;
  assign n806 = x73 | x201 ;
  assign n807 = n805 | n806 ;
  assign n808 = ( n800 & n805 ) | ( n800 & n807 ) | ( n805 & n807 ) ;
  assign n809 = ( x73 & x201 ) | ( x73 & n799 ) | ( x201 & n799 ) ;
  assign n810 = ( n772 & n808 ) | ( n772 & n809 ) | ( n808 & n809 ) ;
  assign n811 = ( x74 & ~x202 ) | ( x74 & n810 ) | ( ~x202 & n810 ) ;
  assign n812 = ( ~x74 & x202 ) | ( ~x74 & n811 ) | ( x202 & n811 ) ;
  assign n813 = ( ~n810 & n811 ) | ( ~n810 & n812 ) | ( n811 & n812 ) ;
  assign n814 = x74 & x202 ;
  assign n815 = x74 | x202 ;
  assign n816 = n809 & n815 ;
  assign n817 = n814 | n816 ;
  assign n818 = n808 & n815 ;
  assign n819 = n814 | n818 ;
  assign n820 = ( n772 & n817 ) | ( n772 & n819 ) | ( n817 & n819 ) ;
  assign n821 = ( x75 & ~x203 ) | ( x75 & n820 ) | ( ~x203 & n820 ) ;
  assign n822 = ( ~x75 & x203 ) | ( ~x75 & n821 ) | ( x203 & n821 ) ;
  assign n823 = ( ~n820 & n821 ) | ( ~n820 & n822 ) | ( n821 & n822 ) ;
  assign n824 = x75 | x203 ;
  assign n825 = ( x75 & x203 ) | ( x75 & n814 ) | ( x203 & n814 ) ;
  assign n826 = ( n816 & n824 ) | ( n816 & n825 ) | ( n824 & n825 ) ;
  assign n827 = x75 & x203 ;
  assign n828 = ( n819 & n824 ) | ( n819 & n827 ) | ( n824 & n827 ) ;
  assign n829 = ( n772 & n826 ) | ( n772 & n828 ) | ( n826 & n828 ) ;
  assign n830 = ( x76 & ~x204 ) | ( x76 & n829 ) | ( ~x204 & n829 ) ;
  assign n831 = ( ~x76 & x204 ) | ( ~x76 & n830 ) | ( x204 & n830 ) ;
  assign n832 = ( ~n829 & n830 ) | ( ~n829 & n831 ) | ( n830 & n831 ) ;
  assign n833 = ( x76 & x204 ) | ( x76 & n825 ) | ( x204 & n825 ) ;
  assign n834 = ( x76 & x204 ) | ( x76 & n824 ) | ( x204 & n824 ) ;
  assign n835 = ( n816 & n833 ) | ( n816 & n834 ) | ( n833 & n834 ) ;
  assign n836 = ( x76 & x204 ) | ( x76 & n827 ) | ( x204 & n827 ) ;
  assign n837 = ( n819 & n834 ) | ( n819 & n836 ) | ( n834 & n836 ) ;
  assign n838 = ( n772 & n835 ) | ( n772 & n837 ) | ( n835 & n837 ) ;
  assign n839 = ( x77 & ~x205 ) | ( x77 & n838 ) | ( ~x205 & n838 ) ;
  assign n840 = ( ~x77 & x205 ) | ( ~x77 & n839 ) | ( x205 & n839 ) ;
  assign n841 = ( ~n838 & n839 ) | ( ~n838 & n840 ) | ( n839 & n840 ) ;
  assign n842 = x78 | x206 ;
  assign n843 = x78 & x206 ;
  assign n844 = x77 & x205 ;
  assign n845 = x77 | x205 ;
  assign n846 = n835 & n845 ;
  assign n847 = n837 & n845 ;
  assign n848 = ( n771 & n846 ) | ( n771 & n847 ) | ( n846 & n847 ) ;
  assign n849 = ( n770 & n846 ) | ( n770 & n847 ) | ( n846 & n847 ) ;
  assign n850 = ( n651 & n848 ) | ( n651 & n849 ) | ( n848 & n849 ) ;
  assign n851 = n844 | n850 ;
  assign n852 = ( ~n842 & n843 ) | ( ~n842 & n851 ) | ( n843 & n851 ) ;
  assign n853 = ( n842 & n843 ) | ( n842 & n851 ) | ( n843 & n851 ) ;
  assign n854 = ( n842 & n852 ) | ( n842 & ~n853 ) | ( n852 & ~n853 ) ;
  assign n855 = ( x79 & ~x207 ) | ( x79 & n853 ) | ( ~x207 & n853 ) ;
  assign n856 = ( ~x79 & x207 ) | ( ~x79 & n855 ) | ( x207 & n855 ) ;
  assign n857 = ( ~n853 & n855 ) | ( ~n853 & n856 ) | ( n855 & n856 ) ;
  assign n858 = x79 & x207 ;
  assign n859 = x79 | x207 ;
  assign n860 = ( n842 & n858 ) | ( n842 & n859 ) | ( n858 & n859 ) ;
  assign n861 = ( n844 & n858 ) | ( n844 & n860 ) | ( n858 & n860 ) ;
  assign n862 = ( n843 & n859 ) | ( n843 & n861 ) | ( n859 & n861 ) ;
  assign n863 = ( n850 & n860 ) | ( n850 & n862 ) | ( n860 & n862 ) ;
  assign n864 = ( x80 & ~x208 ) | ( x80 & n863 ) | ( ~x208 & n863 ) ;
  assign n865 = ( ~x80 & x208 ) | ( ~x80 & n864 ) | ( x208 & n864 ) ;
  assign n866 = ( ~n863 & n864 ) | ( ~n863 & n865 ) | ( n864 & n865 ) ;
  assign n867 = ( x80 & x208 ) | ( x80 & n862 ) | ( x208 & n862 ) ;
  assign n868 = ( x80 & x208 ) | ( x80 & n860 ) | ( x208 & n860 ) ;
  assign n869 = ( n850 & n867 ) | ( n850 & n868 ) | ( n867 & n868 ) ;
  assign n870 = ( x81 & ~x209 ) | ( x81 & n869 ) | ( ~x209 & n869 ) ;
  assign n871 = ( ~x81 & x209 ) | ( ~x81 & n870 ) | ( x209 & n870 ) ;
  assign n872 = ( ~n869 & n870 ) | ( ~n869 & n871 ) | ( n870 & n871 ) ;
  assign n873 = x81 & x209 ;
  assign n874 = x81 | x209 ;
  assign n875 = n868 & n874 ;
  assign n876 = n873 | n875 ;
  assign n877 = ( n867 & n873 ) | ( n867 & n874 ) | ( n873 & n874 ) ;
  assign n878 = ( n850 & n876 ) | ( n850 & n877 ) | ( n876 & n877 ) ;
  assign n879 = ( x82 & ~x210 ) | ( x82 & n878 ) | ( ~x210 & n878 ) ;
  assign n880 = ( ~x82 & x210 ) | ( ~x82 & n879 ) | ( x210 & n879 ) ;
  assign n881 = ( ~n878 & n879 ) | ( ~n878 & n880 ) | ( n879 & n880 ) ;
  assign n882 = ( x82 & x210 ) | ( x82 & n874 ) | ( x210 & n874 ) ;
  assign n883 = ( x82 & x210 ) | ( x82 & n873 ) | ( x210 & n873 ) ;
  assign n884 = ( n867 & n882 ) | ( n867 & n883 ) | ( n882 & n883 ) ;
  assign n885 = ( x82 & x210 ) | ( x82 & n876 ) | ( x210 & n876 ) ;
  assign n886 = ( n850 & n884 ) | ( n850 & n885 ) | ( n884 & n885 ) ;
  assign n887 = ( x83 & ~x211 ) | ( x83 & n886 ) | ( ~x211 & n886 ) ;
  assign n888 = ( ~x83 & x211 ) | ( ~x83 & n887 ) | ( x211 & n887 ) ;
  assign n889 = ( ~n886 & n887 ) | ( ~n886 & n888 ) | ( n887 & n888 ) ;
  assign n890 = x83 & x211 ;
  assign n891 = x83 | x211 ;
  assign n892 = n885 & n891 ;
  assign n893 = n890 | n892 ;
  assign n894 = ( n884 & n890 ) | ( n884 & n891 ) | ( n890 & n891 ) ;
  assign n895 = ( n850 & n893 ) | ( n850 & n894 ) | ( n893 & n894 ) ;
  assign n896 = ( x84 & ~x212 ) | ( x84 & n895 ) | ( ~x212 & n895 ) ;
  assign n897 = ( ~x84 & x212 ) | ( ~x84 & n896 ) | ( x212 & n896 ) ;
  assign n898 = ( ~n895 & n896 ) | ( ~n895 & n897 ) | ( n896 & n897 ) ;
  assign n899 = ( x84 & x212 ) | ( x84 & n891 ) | ( x212 & n891 ) ;
  assign n900 = ( x84 & x212 ) | ( x84 & n890 ) | ( x212 & n890 ) ;
  assign n901 = ( n884 & n899 ) | ( n884 & n900 ) | ( n899 & n900 ) ;
  assign n902 = x84 | x212 ;
  assign n903 = ( n892 & n900 ) | ( n892 & n902 ) | ( n900 & n902 ) ;
  assign n904 = ( n850 & n901 ) | ( n850 & n903 ) | ( n901 & n903 ) ;
  assign n905 = ( x85 & ~x213 ) | ( x85 & n904 ) | ( ~x213 & n904 ) ;
  assign n906 = ( ~x85 & x213 ) | ( ~x85 & n905 ) | ( x213 & n905 ) ;
  assign n907 = ( ~n904 & n905 ) | ( ~n904 & n906 ) | ( n905 & n906 ) ;
  assign n908 = x85 & x213 ;
  assign n909 = x85 | x213 ;
  assign n910 = n903 & n909 ;
  assign n911 = n908 | n910 ;
  assign n912 = ( x85 & x213 ) | ( x85 & n901 ) | ( x213 & n901 ) ;
  assign n913 = ( n850 & n911 ) | ( n850 & n912 ) | ( n911 & n912 ) ;
  assign n914 = ( x86 & ~x214 ) | ( x86 & n913 ) | ( ~x214 & n913 ) ;
  assign n915 = ( ~x86 & x214 ) | ( ~x86 & n914 ) | ( x214 & n914 ) ;
  assign n916 = ( ~n913 & n914 ) | ( ~n913 & n915 ) | ( n914 & n915 ) ;
  assign n917 = x87 | x215 ;
  assign n918 = x87 & x215 ;
  assign n919 = x86 & x214 ;
  assign n920 = x86 | x214 ;
  assign n921 = n911 & n920 ;
  assign n922 = n912 & n920 ;
  assign n923 = ( n849 & n921 ) | ( n849 & n922 ) | ( n921 & n922 ) ;
  assign n924 = ( n848 & n921 ) | ( n848 & n922 ) | ( n921 & n922 ) ;
  assign n925 = ( n651 & n923 ) | ( n651 & n924 ) | ( n923 & n924 ) ;
  assign n926 = n919 | n925 ;
  assign n927 = ( ~n917 & n918 ) | ( ~n917 & n926 ) | ( n918 & n926 ) ;
  assign n928 = ( n917 & n918 ) | ( n917 & n926 ) | ( n918 & n926 ) ;
  assign n929 = ( n917 & n927 ) | ( n917 & ~n928 ) | ( n927 & ~n928 ) ;
  assign n930 = ( x88 & ~x216 ) | ( x88 & n928 ) | ( ~x216 & n928 ) ;
  assign n931 = ( ~x88 & x216 ) | ( ~x88 & n930 ) | ( x216 & n930 ) ;
  assign n932 = ( ~n928 & n930 ) | ( ~n928 & n931 ) | ( n930 & n931 ) ;
  assign n933 = x88 & x216 ;
  assign n934 = x88 | x216 ;
  assign n935 = ( n917 & n933 ) | ( n917 & n934 ) | ( n933 & n934 ) ;
  assign n936 = ( n919 & n933 ) | ( n919 & n935 ) | ( n933 & n935 ) ;
  assign n937 = ( n918 & n934 ) | ( n918 & n936 ) | ( n934 & n936 ) ;
  assign n938 = ( n925 & n935 ) | ( n925 & n937 ) | ( n935 & n937 ) ;
  assign n939 = ( x89 & ~x217 ) | ( x89 & n938 ) | ( ~x217 & n938 ) ;
  assign n940 = ( ~x89 & x217 ) | ( ~x89 & n939 ) | ( x217 & n939 ) ;
  assign n941 = ( ~n938 & n939 ) | ( ~n938 & n940 ) | ( n939 & n940 ) ;
  assign n942 = ( x89 & x217 ) | ( x89 & n937 ) | ( x217 & n937 ) ;
  assign n943 = ( x89 & x217 ) | ( x89 & n935 ) | ( x217 & n935 ) ;
  assign n944 = ( n925 & n942 ) | ( n925 & n943 ) | ( n942 & n943 ) ;
  assign n945 = ( x90 & ~x218 ) | ( x90 & n944 ) | ( ~x218 & n944 ) ;
  assign n946 = ( ~x90 & x218 ) | ( ~x90 & n945 ) | ( x218 & n945 ) ;
  assign n947 = ( ~n944 & n945 ) | ( ~n944 & n946 ) | ( n945 & n946 ) ;
  assign n948 = x90 & x218 ;
  assign n949 = x90 | x218 ;
  assign n950 = n943 & n949 ;
  assign n951 = n948 | n950 ;
  assign n952 = ( n942 & n948 ) | ( n942 & n949 ) | ( n948 & n949 ) ;
  assign n953 = ( n925 & n951 ) | ( n925 & n952 ) | ( n951 & n952 ) ;
  assign n954 = ( x91 & ~x219 ) | ( x91 & n953 ) | ( ~x219 & n953 ) ;
  assign n955 = ( ~x91 & x219 ) | ( ~x91 & n954 ) | ( x219 & n954 ) ;
  assign n956 = ( ~n953 & n954 ) | ( ~n953 & n955 ) | ( n954 & n955 ) ;
  assign n957 = ( x91 & x219 ) | ( x91 & n949 ) | ( x219 & n949 ) ;
  assign n958 = ( x91 & x219 ) | ( x91 & n948 ) | ( x219 & n948 ) ;
  assign n959 = ( n942 & n957 ) | ( n942 & n958 ) | ( n957 & n958 ) ;
  assign n960 = ( x91 & x219 ) | ( x91 & n951 ) | ( x219 & n951 ) ;
  assign n961 = ( n925 & n959 ) | ( n925 & n960 ) | ( n959 & n960 ) ;
  assign n962 = ( x92 & ~x220 ) | ( x92 & n961 ) | ( ~x220 & n961 ) ;
  assign n963 = ( ~x92 & x220 ) | ( ~x92 & n962 ) | ( x220 & n962 ) ;
  assign n964 = ( ~n961 & n962 ) | ( ~n961 & n963 ) | ( n962 & n963 ) ;
  assign n965 = x92 & x220 ;
  assign n966 = x92 | x220 ;
  assign n967 = n960 & n966 ;
  assign n968 = n965 | n967 ;
  assign n969 = ( n959 & n965 ) | ( n959 & n966 ) | ( n965 & n966 ) ;
  assign n970 = ( n925 & n968 ) | ( n925 & n969 ) | ( n968 & n969 ) ;
  assign n971 = ( x93 & ~x221 ) | ( x93 & n970 ) | ( ~x221 & n970 ) ;
  assign n972 = ( ~x93 & x221 ) | ( ~x93 & n971 ) | ( x221 & n971 ) ;
  assign n973 = ( ~n970 & n971 ) | ( ~n970 & n972 ) | ( n971 & n972 ) ;
  assign n974 = ( x93 & x221 ) | ( x93 & n966 ) | ( x221 & n966 ) ;
  assign n975 = ( x93 & x221 ) | ( x93 & n965 ) | ( x221 & n965 ) ;
  assign n976 = ( n959 & n974 ) | ( n959 & n975 ) | ( n974 & n975 ) ;
  assign n977 = x93 | x221 ;
  assign n978 = ( n967 & n975 ) | ( n967 & n977 ) | ( n975 & n977 ) ;
  assign n979 = ( n925 & n976 ) | ( n925 & n978 ) | ( n976 & n978 ) ;
  assign n980 = ( x94 & ~x222 ) | ( x94 & n979 ) | ( ~x222 & n979 ) ;
  assign n981 = ( ~x94 & x222 ) | ( ~x94 & n980 ) | ( x222 & n980 ) ;
  assign n982 = ( ~n979 & n980 ) | ( ~n979 & n981 ) | ( n980 & n981 ) ;
  assign n983 = x94 & x222 ;
  assign n984 = x94 | x222 ;
  assign n985 = n978 & n984 ;
  assign n986 = n983 | n985 ;
  assign n987 = ( x94 & x222 ) | ( x94 & n976 ) | ( x222 & n976 ) ;
  assign n988 = ( n925 & n986 ) | ( n925 & n987 ) | ( n986 & n987 ) ;
  assign n989 = ( x95 & ~x223 ) | ( x95 & n988 ) | ( ~x223 & n988 ) ;
  assign n990 = ( ~x95 & x223 ) | ( ~x95 & n989 ) | ( x223 & n989 ) ;
  assign n991 = ( ~n988 & n989 ) | ( ~n988 & n990 ) | ( n989 & n990 ) ;
  assign n992 = x95 | x223 ;
  assign n993 = x95 & x223 ;
  assign n994 = ( n986 & n992 ) | ( n986 & n993 ) | ( n992 & n993 ) ;
  assign n995 = ( x95 & x223 ) | ( x95 & n987 ) | ( x223 & n987 ) ;
  assign n996 = ( n925 & n994 ) | ( n925 & n995 ) | ( n994 & n995 ) ;
  assign n997 = ( x96 & ~x224 ) | ( x96 & n996 ) | ( ~x224 & n996 ) ;
  assign n998 = ( ~x96 & x224 ) | ( ~x96 & n997 ) | ( x224 & n997 ) ;
  assign n999 = ( ~n996 & n997 ) | ( ~n996 & n998 ) | ( n997 & n998 ) ;
  assign n1000 = x96 & x224 ;
  assign n1001 = x96 | x224 ;
  assign n1002 = n1000 | n1001 ;
  assign n1003 = ( n996 & n1000 ) | ( n996 & n1002 ) | ( n1000 & n1002 ) ;
  assign n1004 = ( x97 & ~x225 ) | ( x97 & n1003 ) | ( ~x225 & n1003 ) ;
  assign n1005 = ( ~x97 & x225 ) | ( ~x97 & n1004 ) | ( x225 & n1004 ) ;
  assign n1006 = ( ~n1003 & n1004 ) | ( ~n1003 & n1005 ) | ( n1004 & n1005 ) ;
  assign n1007 = ( x97 & x225 ) | ( x97 & n1000 ) | ( x225 & n1000 ) ;
  assign n1008 = ( x97 & x225 ) | ( x97 & n1002 ) | ( x225 & n1002 ) ;
  assign n1009 = ( n996 & n1007 ) | ( n996 & n1008 ) | ( n1007 & n1008 ) ;
  assign n1010 = ( x98 & ~x226 ) | ( x98 & n1009 ) | ( ~x226 & n1009 ) ;
  assign n1011 = ( ~x98 & x226 ) | ( ~x98 & n1010 ) | ( x226 & n1010 ) ;
  assign n1012 = ( ~n1009 & n1010 ) | ( ~n1009 & n1011 ) | ( n1010 & n1011 ) ;
  assign n1013 = ( x98 & x226 ) | ( x98 & n1007 ) | ( x226 & n1007 ) ;
  assign n1014 = x98 | x226 ;
  assign n1015 = ( n1008 & n1013 ) | ( n1008 & n1014 ) | ( n1013 & n1014 ) ;
  assign n1016 = ( n996 & n1013 ) | ( n996 & n1015 ) | ( n1013 & n1015 ) ;
  assign n1017 = ( x99 & ~x227 ) | ( x99 & n1016 ) | ( ~x227 & n1016 ) ;
  assign n1018 = ( ~x99 & x227 ) | ( ~x99 & n1017 ) | ( x227 & n1017 ) ;
  assign n1019 = ( ~n1016 & n1017 ) | ( ~n1016 & n1018 ) | ( n1017 & n1018 ) ;
  assign n1020 = x99 & x227 ;
  assign n1021 = x99 | x227 ;
  assign n1022 = n1015 & n1021 ;
  assign n1023 = n1020 | n1022 ;
  assign n1024 = ( x99 & x227 ) | ( x99 & n1013 ) | ( x227 & n1013 ) ;
  assign n1025 = ( n996 & n1023 ) | ( n996 & n1024 ) | ( n1023 & n1024 ) ;
  assign n1026 = ( x100 & ~x228 ) | ( x100 & n1025 ) | ( ~x228 & n1025 ) ;
  assign n1027 = ( ~x100 & x228 ) | ( ~x100 & n1026 ) | ( x228 & n1026 ) ;
  assign n1028 = ( ~n1025 & n1026 ) | ( ~n1025 & n1027 ) | ( n1026 & n1027 ) ;
  assign n1029 = x100 & x228 ;
  assign n1030 = x100 | x228 ;
  assign n1031 = n1029 | n1030 ;
  assign n1032 = ( n1024 & n1029 ) | ( n1024 & n1031 ) | ( n1029 & n1031 ) ;
  assign n1033 = ( x100 & x228 ) | ( x100 & n1023 ) | ( x228 & n1023 ) ;
  assign n1034 = ( n996 & n1032 ) | ( n996 & n1033 ) | ( n1032 & n1033 ) ;
  assign n1035 = ( x101 & ~x229 ) | ( x101 & n1034 ) | ( ~x229 & n1034 ) ;
  assign n1036 = ( ~x101 & x229 ) | ( ~x101 & n1035 ) | ( x229 & n1035 ) ;
  assign n1037 = ( ~n1034 & n1035 ) | ( ~n1034 & n1036 ) | ( n1035 & n1036 ) ;
  assign n1038 = x101 & x229 ;
  assign n1039 = x101 | x229 ;
  assign n1040 = n1033 & n1039 ;
  assign n1041 = n1038 | n1040 ;
  assign n1042 = n1032 & n1039 ;
  assign n1043 = n1038 | n1042 ;
  assign n1044 = ( n996 & n1041 ) | ( n996 & n1043 ) | ( n1041 & n1043 ) ;
  assign n1045 = ( x102 & ~x230 ) | ( x102 & n1044 ) | ( ~x230 & n1044 ) ;
  assign n1046 = ( ~x102 & x230 ) | ( ~x102 & n1045 ) | ( x230 & n1045 ) ;
  assign n1047 = ( ~n1044 & n1045 ) | ( ~n1044 & n1046 ) | ( n1045 & n1046 ) ;
  assign n1048 = x102 | x230 ;
  assign n1049 = ( x102 & x230 ) | ( x102 & n1038 ) | ( x230 & n1038 ) ;
  assign n1050 = ( n1040 & n1048 ) | ( n1040 & n1049 ) | ( n1048 & n1049 ) ;
  assign n1051 = x102 & x230 ;
  assign n1052 = ( n1043 & n1048 ) | ( n1043 & n1051 ) | ( n1048 & n1051 ) ;
  assign n1053 = ( n996 & n1050 ) | ( n996 & n1052 ) | ( n1050 & n1052 ) ;
  assign n1054 = ( x103 & ~x231 ) | ( x103 & n1053 ) | ( ~x231 & n1053 ) ;
  assign n1055 = ( ~x103 & x231 ) | ( ~x103 & n1054 ) | ( x231 & n1054 ) ;
  assign n1056 = ( ~n1053 & n1054 ) | ( ~n1053 & n1055 ) | ( n1054 & n1055 ) ;
  assign n1057 = ( x103 & x231 ) | ( x103 & n1049 ) | ( x231 & n1049 ) ;
  assign n1058 = ( x103 & x231 ) | ( x103 & n1048 ) | ( x231 & n1048 ) ;
  assign n1059 = ( n1040 & n1057 ) | ( n1040 & n1058 ) | ( n1057 & n1058 ) ;
  assign n1060 = ( x103 & x231 ) | ( x103 & n1051 ) | ( x231 & n1051 ) ;
  assign n1061 = ( n1043 & n1058 ) | ( n1043 & n1060 ) | ( n1058 & n1060 ) ;
  assign n1062 = ( n996 & n1059 ) | ( n996 & n1061 ) | ( n1059 & n1061 ) ;
  assign n1063 = ( x104 & ~x232 ) | ( x104 & n1062 ) | ( ~x232 & n1062 ) ;
  assign n1064 = ( ~x104 & x232 ) | ( ~x104 & n1063 ) | ( x232 & n1063 ) ;
  assign n1065 = ( ~n1062 & n1063 ) | ( ~n1062 & n1064 ) | ( n1063 & n1064 ) ;
  assign n1066 = x104 & x232 ;
  assign n1067 = x104 | x232 ;
  assign n1068 = n1061 & n1067 ;
  assign n1069 = n1066 | n1068 ;
  assign n1070 = ( n1059 & n1066 ) | ( n1059 & n1067 ) | ( n1066 & n1067 ) ;
  assign n1071 = ( n996 & n1069 ) | ( n996 & n1070 ) | ( n1069 & n1070 ) ;
  assign n1072 = ( x105 & ~x233 ) | ( x105 & n1071 ) | ( ~x233 & n1071 ) ;
  assign n1073 = ( ~x105 & x233 ) | ( ~x105 & n1072 ) | ( x233 & n1072 ) ;
  assign n1074 = ( ~n1071 & n1072 ) | ( ~n1071 & n1073 ) | ( n1072 & n1073 ) ;
  assign n1075 = ( x105 & x233 ) | ( x105 & n1067 ) | ( x233 & n1067 ) ;
  assign n1076 = ( x105 & x233 ) | ( x105 & n1066 ) | ( x233 & n1066 ) ;
  assign n1077 = ( n1059 & n1075 ) | ( n1059 & n1076 ) | ( n1075 & n1076 ) ;
  assign n1078 = ( x105 & x233 ) | ( x105 & n1069 ) | ( x233 & n1069 ) ;
  assign n1079 = ( n994 & n1077 ) | ( n994 & n1078 ) | ( n1077 & n1078 ) ;
  assign n1080 = ( n995 & n1077 ) | ( n995 & n1078 ) | ( n1077 & n1078 ) ;
  assign n1081 = ( n925 & n1079 ) | ( n925 & n1080 ) | ( n1079 & n1080 ) ;
  assign n1082 = ( x106 & ~x234 ) | ( x106 & n1081 ) | ( ~x234 & n1081 ) ;
  assign n1083 = ( ~x106 & x234 ) | ( ~x106 & n1082 ) | ( x234 & n1082 ) ;
  assign n1084 = ( ~n1081 & n1082 ) | ( ~n1081 & n1083 ) | ( n1082 & n1083 ) ;
  assign n1085 = x106 & x234 ;
  assign n1086 = x106 | x234 ;
  assign n1087 = n1085 | n1086 ;
  assign n1088 = ( n1081 & n1085 ) | ( n1081 & n1087 ) | ( n1085 & n1087 ) ;
  assign n1089 = ( x107 & ~x235 ) | ( x107 & n1088 ) | ( ~x235 & n1088 ) ;
  assign n1090 = ( ~x107 & x235 ) | ( ~x107 & n1089 ) | ( x235 & n1089 ) ;
  assign n1091 = ( ~n1088 & n1089 ) | ( ~n1088 & n1090 ) | ( n1089 & n1090 ) ;
  assign n1092 = ( x107 & x235 ) | ( x107 & n1085 ) | ( x235 & n1085 ) ;
  assign n1093 = ( x107 & x235 ) | ( x107 & n1087 ) | ( x235 & n1087 ) ;
  assign n1094 = ( n1081 & n1092 ) | ( n1081 & n1093 ) | ( n1092 & n1093 ) ;
  assign n1095 = ( x108 & ~x236 ) | ( x108 & n1094 ) | ( ~x236 & n1094 ) ;
  assign n1096 = ( ~x108 & x236 ) | ( ~x108 & n1095 ) | ( x236 & n1095 ) ;
  assign n1097 = ( ~n1094 & n1095 ) | ( ~n1094 & n1096 ) | ( n1095 & n1096 ) ;
  assign n1098 = ( x108 & x236 ) | ( x108 & n1092 ) | ( x236 & n1092 ) ;
  assign n1099 = x108 | x236 ;
  assign n1100 = ( n1093 & n1098 ) | ( n1093 & n1099 ) | ( n1098 & n1099 ) ;
  assign n1101 = ( n1081 & n1098 ) | ( n1081 & n1100 ) | ( n1098 & n1100 ) ;
  assign n1102 = ( x109 & ~x237 ) | ( x109 & n1101 ) | ( ~x237 & n1101 ) ;
  assign n1103 = ( ~x109 & x237 ) | ( ~x109 & n1102 ) | ( x237 & n1102 ) ;
  assign n1104 = ( ~n1101 & n1102 ) | ( ~n1101 & n1103 ) | ( n1102 & n1103 ) ;
  assign n1105 = x109 & x237 ;
  assign n1106 = x109 | x237 ;
  assign n1107 = n1100 & n1106 ;
  assign n1108 = n1105 | n1107 ;
  assign n1109 = ( x109 & x237 ) | ( x109 & n1098 ) | ( x237 & n1098 ) ;
  assign n1110 = ( n1081 & n1108 ) | ( n1081 & n1109 ) | ( n1108 & n1109 ) ;
  assign n1111 = ( x110 & ~x238 ) | ( x110 & n1110 ) | ( ~x238 & n1110 ) ;
  assign n1112 = ( ~x110 & x238 ) | ( ~x110 & n1111 ) | ( x238 & n1111 ) ;
  assign n1113 = ( ~n1110 & n1111 ) | ( ~n1110 & n1112 ) | ( n1111 & n1112 ) ;
  assign n1114 = x110 & x238 ;
  assign n1115 = x110 | x238 ;
  assign n1116 = n1114 | n1115 ;
  assign n1117 = ( n1109 & n1114 ) | ( n1109 & n1116 ) | ( n1114 & n1116 ) ;
  assign n1118 = ( x110 & x238 ) | ( x110 & n1108 ) | ( x238 & n1108 ) ;
  assign n1119 = ( n1081 & n1117 ) | ( n1081 & n1118 ) | ( n1117 & n1118 ) ;
  assign n1120 = ( x111 & ~x239 ) | ( x111 & n1119 ) | ( ~x239 & n1119 ) ;
  assign n1121 = ( ~x111 & x239 ) | ( ~x111 & n1120 ) | ( x239 & n1120 ) ;
  assign n1122 = ( ~n1119 & n1120 ) | ( ~n1119 & n1121 ) | ( n1120 & n1121 ) ;
  assign n1123 = x111 & x239 ;
  assign n1124 = x111 | x239 ;
  assign n1125 = n1118 & n1124 ;
  assign n1126 = n1123 | n1125 ;
  assign n1127 = n1117 & n1124 ;
  assign n1128 = n1123 | n1127 ;
  assign n1129 = ( n1081 & n1126 ) | ( n1081 & n1128 ) | ( n1126 & n1128 ) ;
  assign n1130 = ( x112 & ~x240 ) | ( x112 & n1129 ) | ( ~x240 & n1129 ) ;
  assign n1131 = ( ~x112 & x240 ) | ( ~x112 & n1130 ) | ( x240 & n1130 ) ;
  assign n1132 = ( ~n1129 & n1130 ) | ( ~n1129 & n1131 ) | ( n1130 & n1131 ) ;
  assign n1133 = x112 | x240 ;
  assign n1134 = ( x112 & x240 ) | ( x112 & n1123 ) | ( x240 & n1123 ) ;
  assign n1135 = ( n1125 & n1133 ) | ( n1125 & n1134 ) | ( n1133 & n1134 ) ;
  assign n1136 = x112 & x240 ;
  assign n1137 = ( n1128 & n1133 ) | ( n1128 & n1136 ) | ( n1133 & n1136 ) ;
  assign n1138 = ( n1081 & n1135 ) | ( n1081 & n1137 ) | ( n1135 & n1137 ) ;
  assign n1139 = ( x113 & ~x241 ) | ( x113 & n1138 ) | ( ~x241 & n1138 ) ;
  assign n1140 = ( ~x113 & x241 ) | ( ~x113 & n1139 ) | ( x241 & n1139 ) ;
  assign n1141 = ( ~n1138 & n1139 ) | ( ~n1138 & n1140 ) | ( n1139 & n1140 ) ;
  assign n1142 = ( x113 & x241 ) | ( x113 & n1134 ) | ( x241 & n1134 ) ;
  assign n1143 = ( x113 & x241 ) | ( x113 & n1133 ) | ( x241 & n1133 ) ;
  assign n1144 = ( n1125 & n1142 ) | ( n1125 & n1143 ) | ( n1142 & n1143 ) ;
  assign n1145 = ( x113 & x241 ) | ( x113 & n1136 ) | ( x241 & n1136 ) ;
  assign n1146 = ( n1128 & n1143 ) | ( n1128 & n1145 ) | ( n1143 & n1145 ) ;
  assign n1147 = ( n1081 & n1144 ) | ( n1081 & n1146 ) | ( n1144 & n1146 ) ;
  assign n1148 = ( x114 & ~x242 ) | ( x114 & n1147 ) | ( ~x242 & n1147 ) ;
  assign n1149 = ( ~x114 & x242 ) | ( ~x114 & n1148 ) | ( x242 & n1148 ) ;
  assign n1150 = ( ~n1147 & n1148 ) | ( ~n1147 & n1149 ) | ( n1148 & n1149 ) ;
  assign n1151 = x114 & x242 ;
  assign n1152 = x114 | x242 ;
  assign n1153 = n1146 & n1152 ;
  assign n1154 = n1151 | n1153 ;
  assign n1155 = ( n1144 & n1151 ) | ( n1144 & n1152 ) | ( n1151 & n1152 ) ;
  assign n1156 = ( n1081 & n1154 ) | ( n1081 & n1155 ) | ( n1154 & n1155 ) ;
  assign n1157 = ( x115 & ~x243 ) | ( x115 & n1156 ) | ( ~x243 & n1156 ) ;
  assign n1158 = ( ~x115 & x243 ) | ( ~x115 & n1157 ) | ( x243 & n1157 ) ;
  assign n1159 = ( ~n1156 & n1157 ) | ( ~n1156 & n1158 ) | ( n1157 & n1158 ) ;
  assign n1160 = ( x115 & x243 ) | ( x115 & n1152 ) | ( x243 & n1152 ) ;
  assign n1161 = ( x115 & x243 ) | ( x115 & n1151 ) | ( x243 & n1151 ) ;
  assign n1162 = ( n1144 & n1160 ) | ( n1144 & n1161 ) | ( n1160 & n1161 ) ;
  assign n1163 = x115 | x243 ;
  assign n1164 = ( n1153 & n1161 ) | ( n1153 & n1163 ) | ( n1161 & n1163 ) ;
  assign n1165 = ( n1081 & n1162 ) | ( n1081 & n1164 ) | ( n1162 & n1164 ) ;
  assign n1166 = ( x116 & ~x244 ) | ( x116 & n1165 ) | ( ~x244 & n1165 ) ;
  assign n1167 = ( ~x116 & x244 ) | ( ~x116 & n1166 ) | ( x244 & n1166 ) ;
  assign n1168 = ( ~n1165 & n1166 ) | ( ~n1165 & n1167 ) | ( n1166 & n1167 ) ;
  assign n1169 = x117 | x245 ;
  assign n1170 = x117 & x245 ;
  assign n1171 = x116 & x244 ;
  assign n1172 = x116 | x244 ;
  assign n1173 = n1162 & n1172 ;
  assign n1174 = n1164 & n1172 ;
  assign n1175 = ( n1081 & n1173 ) | ( n1081 & n1174 ) | ( n1173 & n1174 ) ;
  assign n1176 = n1171 | n1175 ;
  assign n1177 = ( ~n1169 & n1170 ) | ( ~n1169 & n1176 ) | ( n1170 & n1176 ) ;
  assign n1178 = ( n1169 & n1170 ) | ( n1169 & n1176 ) | ( n1170 & n1176 ) ;
  assign n1179 = ( n1169 & n1177 ) | ( n1169 & ~n1178 ) | ( n1177 & ~n1178 ) ;
  assign n1180 = ( x118 & ~x246 ) | ( x118 & n1178 ) | ( ~x246 & n1178 ) ;
  assign n1181 = ( ~x118 & x246 ) | ( ~x118 & n1180 ) | ( x246 & n1180 ) ;
  assign n1182 = ( ~n1178 & n1180 ) | ( ~n1178 & n1181 ) | ( n1180 & n1181 ) ;
  assign n1183 = x118 & x246 ;
  assign n1184 = x118 | x246 ;
  assign n1185 = ( n1169 & n1183 ) | ( n1169 & n1184 ) | ( n1183 & n1184 ) ;
  assign n1186 = ( n1171 & n1183 ) | ( n1171 & n1185 ) | ( n1183 & n1185 ) ;
  assign n1187 = ( n1170 & n1184 ) | ( n1170 & n1186 ) | ( n1184 & n1186 ) ;
  assign n1188 = ( n1175 & n1185 ) | ( n1175 & n1187 ) | ( n1185 & n1187 ) ;
  assign n1189 = ( x119 & ~x247 ) | ( x119 & n1188 ) | ( ~x247 & n1188 ) ;
  assign n1190 = ( ~x119 & x247 ) | ( ~x119 & n1189 ) | ( x247 & n1189 ) ;
  assign n1191 = ( ~n1188 & n1189 ) | ( ~n1188 & n1190 ) | ( n1189 & n1190 ) ;
  assign n1192 = ( x119 & x247 ) | ( x119 & n1187 ) | ( x247 & n1187 ) ;
  assign n1193 = ( x119 & x247 ) | ( x119 & n1185 ) | ( x247 & n1185 ) ;
  assign n1194 = ( n1175 & n1192 ) | ( n1175 & n1193 ) | ( n1192 & n1193 ) ;
  assign n1195 = ( x120 & ~x248 ) | ( x120 & n1194 ) | ( ~x248 & n1194 ) ;
  assign n1196 = ( ~x120 & x248 ) | ( ~x120 & n1195 ) | ( x248 & n1195 ) ;
  assign n1197 = ( ~n1194 & n1195 ) | ( ~n1194 & n1196 ) | ( n1195 & n1196 ) ;
  assign n1198 = x120 & x248 ;
  assign n1199 = x120 | x248 ;
  assign n1200 = n1193 & n1199 ;
  assign n1201 = n1198 | n1200 ;
  assign n1202 = ( n1192 & n1198 ) | ( n1192 & n1199 ) | ( n1198 & n1199 ) ;
  assign n1203 = ( n1175 & n1201 ) | ( n1175 & n1202 ) | ( n1201 & n1202 ) ;
  assign n1204 = ( x121 & ~x249 ) | ( x121 & n1203 ) | ( ~x249 & n1203 ) ;
  assign n1205 = ( ~x121 & x249 ) | ( ~x121 & n1204 ) | ( x249 & n1204 ) ;
  assign n1206 = ( ~n1203 & n1204 ) | ( ~n1203 & n1205 ) | ( n1204 & n1205 ) ;
  assign n1207 = ( x121 & x249 ) | ( x121 & n1199 ) | ( x249 & n1199 ) ;
  assign n1208 = ( x121 & x249 ) | ( x121 & n1198 ) | ( x249 & n1198 ) ;
  assign n1209 = ( n1192 & n1207 ) | ( n1192 & n1208 ) | ( n1207 & n1208 ) ;
  assign n1210 = ( x121 & x249 ) | ( x121 & n1201 ) | ( x249 & n1201 ) ;
  assign n1211 = ( n1175 & n1209 ) | ( n1175 & n1210 ) | ( n1209 & n1210 ) ;
  assign n1212 = ( x122 & ~x250 ) | ( x122 & n1211 ) | ( ~x250 & n1211 ) ;
  assign n1213 = ( ~x122 & x250 ) | ( ~x122 & n1212 ) | ( x250 & n1212 ) ;
  assign n1214 = ( ~n1211 & n1212 ) | ( ~n1211 & n1213 ) | ( n1212 & n1213 ) ;
  assign n1215 = x122 & x250 ;
  assign n1216 = x122 | x250 ;
  assign n1217 = n1210 & n1216 ;
  assign n1218 = n1215 | n1217 ;
  assign n1219 = ( n1209 & n1215 ) | ( n1209 & n1216 ) | ( n1215 & n1216 ) ;
  assign n1220 = ( n1175 & n1218 ) | ( n1175 & n1219 ) | ( n1218 & n1219 ) ;
  assign n1221 = ( x123 & ~x251 ) | ( x123 & n1220 ) | ( ~x251 & n1220 ) ;
  assign n1222 = ( ~x123 & x251 ) | ( ~x123 & n1221 ) | ( x251 & n1221 ) ;
  assign n1223 = ( ~n1220 & n1221 ) | ( ~n1220 & n1222 ) | ( n1221 & n1222 ) ;
  assign n1224 = ( x123 & x251 ) | ( x123 & n1216 ) | ( x251 & n1216 ) ;
  assign n1225 = ( x123 & x251 ) | ( x123 & n1215 ) | ( x251 & n1215 ) ;
  assign n1226 = ( n1209 & n1224 ) | ( n1209 & n1225 ) | ( n1224 & n1225 ) ;
  assign n1227 = x123 | x251 ;
  assign n1228 = ( n1217 & n1225 ) | ( n1217 & n1227 ) | ( n1225 & n1227 ) ;
  assign n1229 = ( n1175 & n1226 ) | ( n1175 & n1228 ) | ( n1226 & n1228 ) ;
  assign n1230 = ( x124 & ~x252 ) | ( x124 & n1229 ) | ( ~x252 & n1229 ) ;
  assign n1231 = ( ~x124 & x252 ) | ( ~x124 & n1230 ) | ( x252 & n1230 ) ;
  assign n1232 = ( ~n1229 & n1230 ) | ( ~n1229 & n1231 ) | ( n1230 & n1231 ) ;
  assign n1233 = x124 & x252 ;
  assign n1234 = x124 | x252 ;
  assign n1235 = n1226 & n1234 ;
  assign n1236 = n1233 | n1235 ;
  assign n1237 = n1228 & n1234 ;
  assign n1238 = n1233 | n1237 ;
  assign n1239 = ( n1175 & n1236 ) | ( n1175 & n1238 ) | ( n1236 & n1238 ) ;
  assign n1240 = ( x125 & ~x253 ) | ( x125 & n1239 ) | ( ~x253 & n1239 ) ;
  assign n1241 = ( ~x125 & x253 ) | ( ~x125 & n1240 ) | ( x253 & n1240 ) ;
  assign n1242 = ( ~n1239 & n1240 ) | ( ~n1239 & n1241 ) | ( n1240 & n1241 ) ;
  assign n1243 = x125 | x253 ;
  assign n1244 = ( x125 & x253 ) | ( x125 & n1233 ) | ( x253 & n1233 ) ;
  assign n1245 = ( n1235 & n1243 ) | ( n1235 & n1244 ) | ( n1243 & n1244 ) ;
  assign n1246 = x125 & x253 ;
  assign n1247 = ( n1238 & n1243 ) | ( n1238 & n1246 ) | ( n1243 & n1246 ) ;
  assign n1248 = ( n1175 & n1245 ) | ( n1175 & n1247 ) | ( n1245 & n1247 ) ;
  assign n1249 = ( x126 & ~x254 ) | ( x126 & n1248 ) | ( ~x254 & n1248 ) ;
  assign n1250 = ( ~x126 & x254 ) | ( ~x126 & n1249 ) | ( x254 & n1249 ) ;
  assign n1251 = ( ~n1248 & n1249 ) | ( ~n1248 & n1250 ) | ( n1249 & n1250 ) ;
  assign n1252 = ( x126 & x254 ) | ( x126 & n1244 ) | ( x254 & n1244 ) ;
  assign n1253 = ( x126 & x254 ) | ( x126 & n1243 ) | ( x254 & n1243 ) ;
  assign n1254 = ( n1235 & n1252 ) | ( n1235 & n1253 ) | ( n1252 & n1253 ) ;
  assign n1255 = ( x126 & x254 ) | ( x126 & n1246 ) | ( x254 & n1246 ) ;
  assign n1256 = ( n1238 & n1253 ) | ( n1238 & n1255 ) | ( n1253 & n1255 ) ;
  assign n1257 = ( n1175 & n1254 ) | ( n1175 & n1256 ) | ( n1254 & n1256 ) ;
  assign n1258 = ( x127 & ~x255 ) | ( x127 & n1257 ) | ( ~x255 & n1257 ) ;
  assign n1259 = ( ~x127 & x255 ) | ( ~x127 & n1258 ) | ( x255 & n1258 ) ;
  assign n1260 = ( ~n1257 & n1258 ) | ( ~n1257 & n1259 ) | ( n1258 & n1259 ) ;
  assign n1261 = ( x127 & x255 ) | ( x127 & n1257 ) | ( x255 & n1257 ) ;
  assign y0 = n259 ;
  assign y1 = n263 ;
  assign y2 = n267 ;
  assign y3 = n271 ;
  assign y4 = n275 ;
  assign y5 = n282 ;
  assign y6 = n286 ;
  assign y7 = n293 ;
  assign y8 = n299 ;
  assign y9 = n310 ;
  assign y10 = n313 ;
  assign y11 = n322 ;
  assign y12 = n333 ;
  assign y13 = n336 ;
  assign y14 = n345 ;
  assign y15 = n351 ;
  assign y16 = n358 ;
  assign y17 = n364 ;
  assign y18 = n371 ;
  assign y19 = n380 ;
  assign y20 = n387 ;
  assign y21 = n393 ;
  assign y22 = n400 ;
  assign y23 = n409 ;
  assign y24 = n420 ;
  assign y25 = n423 ;
  assign y26 = n432 ;
  assign y27 = n438 ;
  assign y28 = n447 ;
  assign y29 = n460 ;
  assign y30 = n463 ;
  assign y31 = n472 ;
  assign y32 = n478 ;
  assign y33 = n487 ;
  assign y34 = n495 ;
  assign y35 = n502 ;
  assign y36 = n508 ;
  assign y37 = n515 ;
  assign y38 = n524 ;
  assign y39 = n533 ;
  assign y40 = n542 ;
  assign y41 = n549 ;
  assign y42 = n555 ;
  assign y43 = n562 ;
  assign y44 = n571 ;
  assign y45 = n580 ;
  assign y46 = n589 ;
  assign y47 = n600 ;
  assign y48 = n603 ;
  assign y49 = n612 ;
  assign y50 = n618 ;
  assign y51 = n627 ;
  assign y52 = n635 ;
  assign y53 = n644 ;
  assign y54 = n655 ;
  assign y55 = n658 ;
  assign y56 = n667 ;
  assign y57 = n673 ;
  assign y58 = n682 ;
  assign y59 = n690 ;
  assign y60 = n699 ;
  assign y61 = n707 ;
  assign y62 = n714 ;
  assign y63 = n720 ;
  assign y64 = n727 ;
  assign y65 = n736 ;
  assign y66 = n745 ;
  assign y67 = n755 ;
  assign y68 = n764 ;
  assign y69 = n775 ;
  assign y70 = n782 ;
  assign y71 = n788 ;
  assign y72 = n795 ;
  assign y73 = n804 ;
  assign y74 = n813 ;
  assign y75 = n823 ;
  assign y76 = n832 ;
  assign y77 = n841 ;
  assign y78 = n854 ;
  assign y79 = n857 ;
  assign y80 = n866 ;
  assign y81 = n872 ;
  assign y82 = n881 ;
  assign y83 = n889 ;
  assign y84 = n898 ;
  assign y85 = n907 ;
  assign y86 = n916 ;
  assign y87 = n929 ;
  assign y88 = n932 ;
  assign y89 = n941 ;
  assign y90 = n947 ;
  assign y91 = n956 ;
  assign y92 = n964 ;
  assign y93 = n973 ;
  assign y94 = n982 ;
  assign y95 = n991 ;
  assign y96 = n999 ;
  assign y97 = n1006 ;
  assign y98 = n1012 ;
  assign y99 = n1019 ;
  assign y100 = n1028 ;
  assign y101 = n1037 ;
  assign y102 = n1047 ;
  assign y103 = n1056 ;
  assign y104 = n1065 ;
  assign y105 = n1074 ;
  assign y106 = n1084 ;
  assign y107 = n1091 ;
  assign y108 = n1097 ;
  assign y109 = n1104 ;
  assign y110 = n1113 ;
  assign y111 = n1122 ;
  assign y112 = n1132 ;
  assign y113 = n1141 ;
  assign y114 = n1150 ;
  assign y115 = n1159 ;
  assign y116 = n1168 ;
  assign y117 = n1179 ;
  assign y118 = n1182 ;
  assign y119 = n1191 ;
  assign y120 = n1197 ;
  assign y121 = n1206 ;
  assign y122 = n1214 ;
  assign y123 = n1223 ;
  assign y124 = n1232 ;
  assign y125 = n1242 ;
  assign y126 = n1251 ;
  assign y127 = n1260 ;
  assign y128 = n1261 ;
endmodule
