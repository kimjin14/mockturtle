//Written by the Majority Logic Package Fri Nov 14 22:36:45 2014
module top (
            cin, a0, b0, b1, a1, b2, a2, b3, a3, b4, a4, b5, a5, b6, a6, b7, a7, b8, a8, b9, a9, b10, a10, b11, a11, b12, a12, b13, a13, b14, a14, b15, a15, b16, a16, b17, a17, b18, a18, b19, a19, b20, a20, b21, a21, b22, a22, b23, a23, b24, a24, b25, a25, b26, a26, b27, a27, b28, a28, b29, a29, b30, a30, a31, b31, 
            s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15, s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29, s30, s31, s32);
input cin, a0, b0, b1, a1, b2, a2, b3, a3, b4, a4, b5, a5, b6, a6, b7, a7, b8, a8, b9, a9, b10, a10, b11, a11, b12, a12, b13, a13, b14, a14, b15, a15, b16, a16, b17, a17, b18, a18, b19, a19, b20, a20, b21, a21, b22, a22, b23, a23, b24, a24, b25, a25, b26, a26, b27, a27, b28, a28, b29, a29, b30, a30, a31, b31;
output s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15, s16, s17, s18, s19, s20, s21, s22, s23, s24, s25, s26, s27, s28, s29, s30, s31, s32;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609;
assign w0 = a1 & ~w119;
assign w1 = w48 & w9;
assign w2 = ~w145 & ~w104;
assign w3 = (~w273 & w77) | (~w273 & w27) | (w77 & w27);
assign w4 = w496 & ~w14;
assign w5 = w198 & ~w601;
assign w6 = (~w560 & w81) | (~w560 & w80) | (w81 & w80);
assign w7 = w514 & w28;
assign w8 = b10 & a10;
assign w9 = (~w580 & w158) | (~w580 & w34) | (w158 & w34);
assign w10 = ~w14 & w434;
assign w11 = b22 & a22;
assign w12 = (~w137 & w475) | (~w137 & w431) | (w475 & w431);
assign w13 = ~w447 & ~w171;
assign w14 = w75 & w480;
assign w15 = (~w247 & w27) | (~w247 & w3) | (w27 & w3);
assign w16 = ~w500 & w184;
assign w17 = ~w264 & w289;
assign w18 = ~b23 & ~a23;
assign w19 = (~w75 & w360) | (~w75 & w419) | (w360 & w419);
assign w20 = (w290 & w388) | (w290 & ~w38) | (w388 & ~w38);
assign w21 = ~w592 & ~w515;
assign w22 = (~w478 & w6) | (~w478 & w44) | (w6 & w44);
assign w23 = (~w580 & w51) | (~w580 & w36) | (w51 & w36);
assign w24 = (w580 & w102) | (w580 & w5) | (w102 & w5);
assign w25 = ~w104 & ~w8;
assign w26 = b13 & a13;
assign w27 = ~w348 & w258;
assign w28 = w479 & ~w485;
assign w29 = ~w335 & ~w299;
assign w30 = ~w284 & ~w568;
assign w31 = (~w75 & w336) | (~w75 & w134) | (w336 & w134);
assign w32 = w26 & ~w398;
assign w33 = (w556 & w541) | (w556 & w88) | (w541 & w88);
assign w34 = (~w386 & w562) | (~w386 & w601) | (w562 & w601);
assign w35 = ~w307 & ~w46;
assign w36 = (~w317 & w463) | (~w317 & w601) | (w463 & w601);
assign w37 = ~w112 & ~w457;
assign w38 = ~w139 & w30;
assign w39 = ~w322 & w372;
assign w40 = a1 & ~w166;
assign w41 = (~w149 & w541) | (~w149 & w33) | (w541 & w33);
assign w42 = w511 & ~w172;
assign w43 = w48 & w158;
assign w44 = w310 & ~w478;
assign w45 = w125 | w118;
assign w46 = (w16 & w148) | (w16 & w400) | (w148 & w400);
assign w47 = w580 & w524;
assign w48 = ~w382 & ~w573;
assign w49 = (~w75 & w162) | (~w75 & w12) | (w162 & w12);
assign w50 = (w560 & w69) | (w560 & w420) | (w69 & w420);
assign w51 = (~w317 & w463) | (~w317 & w327) | (w463 & w327);
assign w52 = ~w100 & w409;
assign w53 = (w560 & w293) | (w560 & w205) | (w293 & w205);
assign w54 = b18 & a18;
assign w55 = ~b5 & ~a5;
assign w56 = (w118 & w125) | (w118 & ~w137) | (w125 & ~w137);
assign w57 = ~w227 & ~w464;
assign w58 = (~w318 & ~w111) | (~w318 & w490) | (~w111 & w490);
assign w59 = (~w75 & w369) | (~w75 & w305) | (w369 & w305);
assign w60 = w164 & ~b1;
assign w61 = w523 & ~w151;
assign w62 = (~w75 & w51) | (~w75 & w23) | (w51 & w23);
assign w63 = (w159 & w163) | (w159 & ~w601) | (w163 & ~w601);
assign w64 = ~w145 & w25;
assign w65 = ~w193 & ~w351;
assign w66 = ~w144 & ~w422;
assign w67 = ~w29 & ~w386;
assign w68 = ~w605 & w213;
assign w69 = ~w322 & w82;
assign w70 = w309 | ~w207;
assign w71 = w116 & w349;
assign w72 = w465 & ~w8;
assign w73 = w580 & w570;
assign w74 = ~w567 & ~w341;
assign w75 = ~w396 & ~w61;
assign w76 = ~w179 & w587;
assign w77 = ~w348 & ~w497;
assign w78 = ~w569 & ~w513;
assign w79 = (w534 & w340) | (w534 & w350) | (w340 & w350);
assign w80 = w455 & ~w379;
assign w81 = w455 & ~w245;
assign w82 = (w430 & ~w143) | (w430 & ~w38) | (~w143 & ~w38);
assign w83 = (w560 & w410) | (w560 & w443) | (w410 & w443);
assign w84 = ~b29 & ~a29;
assign w85 = w224 & ~w255;
assign w86 = ~w273 & ~w555;
assign w87 = w263 & ~w72;
assign w88 = ~w331 & ~w131;
assign w89 = ~w242 & ~w11;
assign w90 = (~w601 & w582) | (~w601 & w357) | (w582 & w357);
assign w91 = ~w255 & w92;
assign w92 = ~w142 & ~w157;
assign w93 = (w312 & w552) | (w312 & ~w75) | (w552 & ~w75);
assign w94 = ~w30 & ~w71;
assign w95 = w278 & ~w184;
assign w96 = (~w58 & ~w501) | (~w58 & w270) | (~w501 & w270);
assign w97 = ~w313 & w192;
assign w98 = ~w127 & ~w254;
assign w99 = w437 & w597;
assign w100 = (w256 & w149) | (w256 & w381) | (w149 & w381);
assign w101 = (~w568 & ~w139) | (~w568 & w384) | (~w139 & w384);
assign w102 = w198 & ~w327;
assign w103 = ~w437 & ~w597;
assign w104 = b9 & a9;
assign w105 = (~w11 & w131) | (~w11 & ~w556) | (w131 & ~w556);
assign w106 = ~w196 & ~w157;
assign w107 = w87 & ~w469;
assign w108 = ~w133 & ~w598;
assign w109 = (~w429 & w549) | (~w429 & ~w301) | (w549 & ~w301);
assign w110 = ~w354 & w252;
assign w111 = ~w55 & ~w318;
assign w112 = (w277 & w395) | (w277 & w472) | (w395 & w472);
assign w113 = ~w478 & ~w579;
assign w114 = w564 & w101;
assign w115 = w263 & w106;
assign w116 = ~w25 & w91;
assign w117 = w394 & ~w422;
assign w118 = (w286 & w289) | (w286 & w199) | (w289 & w199);
assign w119 = ~w110 & ~w166;
assign w120 = (w273 & w456) | (w273 & w393) | (w456 & w393);
assign w121 = (w590 & ~w75) | (w590 & w298) | (~w75 & w298);
assign w122 = ~w135 & ~w545;
assign w123 = ~w587 & ~w575;
assign w124 = (~w560 & w461) | (~w560 & w607) | (w461 & w607);
assign w125 = (w289 & w520) | (w289 & w17) | (w520 & w17);
assign w126 = (w314 & w313) | (w314 & w542) | (w313 & w542);
assign w127 = ~w148 & w521;
assign w128 = ~w225 & ~w249;
assign w129 = (w75 & w42) | (w75 & w499) | (w42 & w499);
assign w130 = w356 & ~w513;
assign w131 = w573 & ~w11;
assign w132 = ~w464 & ~w500;
assign w133 = ~w8 & ~w388;
assign w134 = (w186 & ~w585) | (w186 & ~w137) | (~w585 & ~w137);
assign w135 = (~w148 & w488) | (~w148 & w489) | (w488 & w489);
assign w136 = w465 & ~w176;
assign w137 = w580 & w531;
assign w138 = w110 & w259;
assign w139 = ~w568 & ~w141;
assign w140 = ~w311 & ~w226;
assign w141 = b7 & a7;
assign w142 = ~b11 & ~a11;
assign w143 = ~w142 & ~w539;
assign w144 = ~w18 & ~w529;
assign w145 = b8 & a8;
assign w146 = ~w322 & w290;
assign w147 = ~w389 & ~w141;
assign w148 = (w259 & w40) | (w259 & w138) | (w40 & w138);
assign w149 = ~w327 & w167;
assign w150 = ~w342 & ~w50;
assign w151 = (~w71 & ~w7) | (~w71 & w94) | (~w7 & w94);
assign w152 = w155 & ~w378;
assign w153 = b30 & a30;
assign w154 = w596 & ~w537;
assign w155 = ~w575 & w429;
assign w156 = ~w311 & ~w146;
assign w157 = ~b12 & ~a12;
assign w158 = (~w386 & w562) | (~w386 & w327) | (w562 & w327);
assign w159 = (w210 & w383) | (w210 & ~w562) | (w383 & ~w562);
assign w160 = ~w577 & w13;
assign w161 = ~w572 & w508;
assign w162 = (w520 & w70) | (w520 & w475) | (w70 & w475);
assign w163 = (w210 & w383) | (w210 & w386) | (w383 & w386);
assign w164 = ~a0 & ~b0;
assign w165 = w221 & w240;
assign w166 = (~b1 & w354) | (~b1 & w60) | (w354 & w60);
assign w167 = ~w268 & w589;
assign w168 = b15 & a15;
assign w169 = (~w534 & w360) | (~w534 & w452) | (w360 & w452);
assign w170 = (w111 & w544) | (w111 & w334) | (w544 & w334);
assign w171 = w193 & ~w282;
assign w172 = ~w171 & w218;
assign w173 = ~w460 & ~w19;
assign w174 = b28 & a28;
assign w175 = ~w129 & w407;
assign w176 = ~w255 & ~w8;
assign w177 = ~w264 & ~w84;
assign w178 = ~b26 & ~a26;
assign w179 = (~w257 & w66) | (~w257 & w279) | (w66 & w279);
assign w180 = (w507 & w551) | (w507 & w303) | (w551 & w303);
assign w181 = b4 & a4;
assign w182 = (w541 & ~w149) | (w541 & w406) | (~w149 & w406);
assign w183 = ~w255 & ~w72;
assign w184 = ~w581 & ~w181;
assign w185 = ~w577 & w327;
assign w186 = (~w190 & ~w338) | (~w190 & w453) | (~w338 & w453);
assign w187 = w385 & w351;
assign w188 = (w240 & w221) | (w240 & w137) | (w221 & w137);
assign w189 = (w580 & w340) | (w580 & w79) | (w340 & w79);
assign w190 = w144 & w117;
assign w191 = (~w556 & w387) | (~w556 & w212) | (w387 & w212);
assign w192 = ~w153 & ~w314;
assign w193 = ~b16 & ~a16;
assign w194 = w105 & w387;
assign w195 = w564 & w561;
assign w196 = b12 & a12;
assign w197 = ~b18 & ~a18;
assign w198 = w468 & w317;
assign w199 = w517 & w177;
assign w200 = (~w176 & w136) | (~w176 & w379) | (w136 & w379);
assign w201 = ~w550 & ~w602;
assign w202 = (w599 & ~w108) | (w599 & w379) | (~w108 & w379);
assign w203 = (~w75 & w182) | (~w75 & w404) | (w182 & w404);
assign w204 = (w286 & w319) | (w286 & w126) | (w319 & w126);
assign w205 = ~w564 & ~w101;
assign w206 = ~b25 & ~a25;
assign w207 = ~w253 & ~w84;
assign w208 = ~w225 & ~w141;
assign w209 = (w599 & ~w108) | (w599 & w245) | (~w108 & w245);
assign w210 = ~w382 & ~w89;
assign w211 = (~w75 & w292) | (~w75 & w326) | (w292 & w326);
assign w212 = w331 & w131;
assign w213 = (w595 & w149) | (w595 & w414) | (w149 & w414);
assign w214 = (w159 & w163) | (w159 & ~w327) | (w163 & ~w327);
assign w215 = ~w18 & w437;
assign w216 = (~w137 & w553) | (~w137 & w109) | (w553 & w109);
assign w217 = ~w314 & w373;
assign w218 = ~w447 & ~w197;
assign w219 = (w217 & w97) | (w217 & ~w286) | (w97 & ~w286);
assign w220 = (w277 & w316) | (w277 & w424) | (w316 & w424);
assign w221 = w338 & w99;
assign w222 = w432 & w96;
assign w223 = ~b28 & ~a28;
assign w224 = ~w465 & ~w104;
assign w225 = (~w141 & ~w116) | (~w141 & w147) | (~w116 & w147);
assign w226 = w388 & ~w322;
assign w227 = b2 & a2;
assign w228 = ~w40 & w260;
assign w229 = ~w164 & ~w354;
assign w230 = ~w432 & ~w111;
assign w231 = ~w32 & ~w484;
assign w232 = w273 & ~w231;
assign w233 = ~w429 & w575;
assign w234 = (~w84 & w177) | (~w84 & w286) | (w177 & w286);
assign w235 = ~w241 & ~w59;
assign w236 = ~w346 & w66;
assign w237 = ~w271 & ~w84;
assign w238 = ~b15 & ~a15;
assign w239 = w597 & w190;
assign w240 = (w338 & w239) | (w338 & w532) | (w239 & w532);
assign w241 = (w75 & w165) | (w75 & w188) | (w165 & w188);
assign w242 = ~b22 & ~a22;
assign w243 = ~w87 & ~w21;
assign w244 = ~w396 & w47;
assign w245 = w2 & ~w38;
assign w246 = ~w322 & w20;
assign w247 = (w560 & w246) | (w560 & w39) | (w246 & w39);
assign w248 = ~w335 & ~w565;
assign w249 = w284 & w141;
assign w250 = ~w380 & ~w62;
assign w251 = (w155 & w179) | (w155 & w509) | (w179 & w509);
assign w252 = ~w164 & b1;
assign w253 = b29 & a29;
assign w254 = (w132 & w148) | (w132 & w512) | (w148 & w512);
assign w255 = ~b10 & ~a10;
assign w256 = w155 & w261;
assign w257 = b25 & a25;
assign w258 = ~w497 & w26;
assign w259 = ~w294 & ~w227;
assign w260 = ~w110 & ~w259;
assign w261 = w394 & w557;
assign w262 = w196 & w8;
assign w263 = ~w255 & w143;
assign w264 = ~w174 & ~w253;
assign w265 = (w560 & w546) | (w560 & w154) | (w546 & w154);
assign w266 = ~w6 & w295;
assign w267 = w490 & ~w270;
assign w268 = w54 & w248;
assign w269 = w471 & w139;
assign w270 = ~w57 & w334;
assign w271 = ~b30 & ~a30;
assign w272 = w528 & ~w334;
assign w273 = w388 & ~w91;
assign w274 = (w61 & ~w371) | (w61 & w526) | (~w371 & w526);
assign w275 = (~w597 & ~w338) | (~w597 & w103) | (~w338 & w103);
assign w276 = a0 & b0;
assign w277 = (w334 & w148) | (w334 & w270) | (w148 & w270);
assign w278 = w500 & ~w184;
assign w279 = ~w346 & ~w257;
assign w280 = b6 & a6;
assign w281 = ~w53 & ~w339;
assign w282 = b17 & a17;
assign w283 = ~w597 & w453;
assign w284 = ~b8 & ~a8;
assign w285 = w386 & ~w382;
assign w286 = ~w251 & w325;
assign w287 = w115 & ~w355;
assign w288 = ~w111 & w330;
assign w289 = w517 & ~w84;
assign w290 = ~w224 & w388;
assign w291 = ~w78 & ~w297;
assign w292 = w520 | w286;
assign w293 = ~w564 & ~w561;
assign w294 = ~b2 & ~a2;
assign w295 = ~w310 & w478;
assign w296 = (~w75 & w576) | (~w75 & w337) | (w576 & w337);
assign w297 = w569 & w513;
assign w298 = ~w137 & w590;
assign w299 = b20 & a20;
assign w300 = ~w10 & ~w358;
assign w301 = (~w575 & ~w590) | (~w575 & w535) | (~w590 & w535);
assign w302 = (w580 & w533) | (w580 & w90) | (w533 & w90);
assign w303 = w86 & w156;
assign w304 = ~w124 & ~w265;
assign w305 = (w275 & w563) | (w275 & ~w137) | (w563 & ~w137);
assign w306 = ~a31 & ~b31;
assign w307 = (~w148 & w95) | (~w148 & w506) | (w95 & w506);
assign w308 = b16 & a16;
assign w309 = w174 & ~w207;
assign w310 = (w560 & w209) | (w560 & w202) | (w209 & w202);
assign w311 = w497 & w291;
assign w312 = ~w595 | ~w213;
assign w313 = ~w264 & w237;
assign w314 = ~w578 & ~w306;
assign w315 = ~w251 & w362;
assign w316 = (~w469 & ~w446) | (~w469 & ~w288) | (~w446 & ~w288);
assign w317 = ~w299 & ~w386;
assign w318 = b5 & a5;
assign w319 = w314 & ~w373;
assign w320 = ~w534 & ~w371;
assign w321 = ~w548 & ~w574;
assign w322 = ~w64 & w183;
assign w323 = ~w61 & w324;
assign w324 = ~w396 & w73;
assign w325 = w362 & ~w256;
assign w326 = (w286 & w520) | (w286 & ~w137) | (w520 & ~w137);
assign w327 = w248 & w172;
assign w328 = (w534 & w42) | (w534 & w377) | (w42 & w377);
assign w329 = (w387 & w149) | (w387 & w194) | (w149 & w194);
assign w330 = ~w318 & ~w280;
assign w331 = ~w504 & ~w18;
assign w332 = ~b27 & ~a27;
assign w333 = ~w605 & ~w312;
assign w334 = ~w500 & ~w581;
assign w335 = b19 & a19;
assign w336 = ~w585 | w186;
assign w337 = (~w137 & w234) | (~w137 & w435) | (w234 & w435);
assign w338 = (w508 & w149) | (w508 & w161) | (w149 & w161);
assign w339 = (~w560 & w114) | (~w560 & w195) | (w114 & w195);
assign w340 = ~w486 & ~w13;
assign w341 = (~w148 & w272) | (~w148 & w370) | (w272 & w370);
assign w342 = w87 & w220;
assign w343 = w397 | w495;
assign w344 = (~w58 & ~w501) | (~w58 & w334) | (~w501 & w334);
assign w345 = ~w54 & ~w335;
assign w346 = ~w257 & ~w206;
assign w347 = w97 & w217;
assign w348 = ~w356 & ~w569;
assign w349 = w389 & w568;
assign w350 = ~w486 & ~w160;
assign w351 = ~w282 & ~w447;
assign w352 = w587 & ~w261;
assign w353 = ~w449 & ~w423;
assign w354 = ~cin & ~w276;
assign w355 = ~w224 & ~w322;
assign w356 = ~b14 & ~a14;
assign w357 = ~w48 & ~w562;
assign w358 = (w438 & w14) | (w438 & w606) | (w14 & w606);
assign w359 = w145 & ~w224;
assign w360 = w486 & w13;
assign w361 = (~w520 & w347) | (~w520 & w219) | (w347 & w219);
assign w362 = ~w332 & w438;
assign w363 = w534 & w577;
assign w364 = (w560 & w405) | (w560 & w200) | (w405 & w200);
assign w365 = (w430 & ~w143) | (w430 & ~w537) | (~w143 & ~w537);
assign w366 = ~w15 & ~w390;
assign w367 = w61 & w65;
assign w368 = (~w75 & w109) | (~w75 & w216) | (w109 & w216);
assign w369 = w563 | w275;
assign w370 = w528 & ~w270;
assign w371 = ~w308 & ~w193;
assign w372 = (w290 & w388) | (w290 & ~w537) | (w388 & ~w537);
assign w373 = ~w153 & ~w237;
assign w374 = ~w471 & ~w139;
assign w375 = ~w577 & w172;
assign w376 = ~w403 & ~w421;
assign w377 = w511 & ~w375;
assign w378 = ~w179 & w352;
assign w379 = (w2 & ~w101) | (w2 & w433) | (~w101 & w433);
assign w380 = (w75 & w102) | (w75 & w24) | (w102 & w24);
assign w381 = ~w572 & w256;
assign w382 = b21 & a21;
assign w383 = ~w48 & w210;
assign w384 = ~w471 & ~w568;
assign w385 = w193 & w351;
assign w386 = ~b20 & ~a20;
assign w387 = w331 & ~w11;
assign w388 = (~w196 & ~w106) | (~w196 & w503) | (~w106 & w503);
assign w389 = ~w485 & w473;
assign w390 = (w247 & w393) | (w247 & w120) | (w393 & w120);
assign w391 = ~w49 & ~w608;
assign w392 = (w149 & w387) | (w149 & w191) | (w387 & w191);
assign w393 = w348 & ~w258;
assign w394 = ~w11 & ~w504;
assign w395 = w374 & ~w288;
assign w396 = ~w523 & w493;
assign w397 = ~w338 & w518;
assign w398 = ~w130 & ~w492;
assign w399 = (~w75 & w343) | (~w75 & w442) | (w343 & w442);
assign w400 = ~w57 & w16;
assign w401 = (w351 & w385) | (w351 & ~w61) | (w385 & ~w61);
assign w402 = ~w228 & ~w148;
assign w403 = ~w517 & ~w296;
assign w404 = (w541 & w41) | (w541 & ~w137) | (w41 & ~w137);
assign w405 = (~w176 & w136) | (~w176 & w245) | (w136 & w245);
assign w406 = w33 | w541;
assign w407 = (w75 & w519) | (w75 & w547) | (w519 & w547);
assign w408 = (w387 & w392) | (w387 & w137) | (w392 & w137);
assign w409 = ~w251 & ~w332;
assign w410 = ~w21 & ~w107;
assign w411 = ~w569 & ~w26;
assign w412 = ~cin & w164;
assign w413 = ~w83 & ~w440;
assign w414 = ~w572 & w595;
assign w415 = w389 & ~w564;
assign w416 = w4 & ~w368;
assign w417 = (w210 & w383) | (w210 & ~w158) | (w383 & ~w158);
assign w418 = w598 & w465;
assign w419 = (~w580 & w360) | (~w580 & w169) | (w360 & w169);
assign w420 = ~w322 & w365;
assign w421 = (~w75 & w45) | (~w75 & w56) | (w45 & w56);
assign w422 = b24 & a24;
assign w423 = (w75 & w333) | (w75 & w591) | (w333 & w591);
assign w424 = (~w469 & ~w446) | (~w469 & ~w554) | (~w446 & ~w554);
assign w425 = ~w597 & ~w190;
assign w426 = b27 & a27;
assign w427 = (w75 & w329) | (w75 & w408) | (w329 & w408);
assign w428 = ~w466 & ~w180;
assign w429 = ~w426 & ~w332;
assign w430 = ~w143 & ~w85;
assign w431 = (~w207 & w309) | (~w207 & w520) | (w309 & w520);
assign w432 = ~w471 & ~w280;
assign w433 = w284 & w2;
assign w434 = w52 & ~w438;
assign w435 = (~w84 & w177) | (~w84 & w520) | (w177 & w520);
assign w436 = ~w266 & ~w22;
assign w437 = ~w529 & ~w422;
assign w438 = ~w223 & ~w174;
assign w439 = w115 & w322;
assign w440 = (w507 & w439) | (w507 & w287) | (w439 & w287);
assign w441 = (w288 & w554) | (w288 & ~w334) | (w554 & ~w334);
assign w442 = (w495 & w397) | (w495 & ~w137) | (w397 & ~w137);
assign w443 = (~w21 & w446) | (~w21 & w243) | (w446 & w243);
assign w444 = ~w145 & ~w467;
assign w445 = w18 & ~w437;
assign w446 = w64 & ~w537;
assign w447 = ~b17 & ~a17;
assign w448 = (w111 & w544) | (w111 & w270) | (w544 & w270);
assign w449 = w605 & w93;
assign w450 = ~w427 & ~w203;
assign w451 = (~w560 & w525) | (~w560 & w482) | (w525 & w482);
assign w452 = w486 & w160;
assign w453 = (~w437 & ~w117) | (~w437 & w604) | (~w117 & w604);
assign w454 = ~a1 & w119;
assign w455 = ~w465 & ~w273;
assign w456 = w348 & w497;
assign w457 = (w139 & w269) | (w139 & w560) | (w269 & w560);
assign w458 = w490 & ~w334;
assign w459 = ~w389 & ~w168;
assign w460 = (w75 & w340) | (w75 & w189) | (w340 & w189);
assign w461 = (~w224 & w359) | (~w224 & w38) | (w359 & w38);
assign w462 = ~w121 & ~w483;
assign w463 = ~w468 & ~w317;
assign w464 = b3 & a3;
assign w465 = ~b9 & ~a9;
assign w466 = (~w231 & w247) | (~w231 & w232) | (w247 & w232);
assign w467 = w116 & w415;
assign w468 = (~w335 & ~w248) | (~w335 & w345) | (~w248 & w345);
assign w469 = w64 & ~w38;
assign w470 = ~w0 & ~w454;
assign w471 = ~b6 & ~a6;
assign w472 = w374 & ~w554;
assign w473 = ~w356 & ~w238;
assign w474 = w179 & ~w587;
assign w475 = (~w207 & w309) | (~w207 & w286) | (w309 & w286);
assign w476 = ~w432 & ~w318;
assign w477 = (w217 & w97) | (w217 & ~w520) | (w97 & ~w520);
assign w478 = ~w497 & ~w26;
assign w479 = w183 & w492;
assign w480 = w137 & w152;
assign w481 = w31 & ~w399;
assign w482 = w600 & ~w379;
assign w483 = (w75 & w417) | (w75 & w494) | (w417 & w494);
assign w484 = ~w26 & ~w291;
assign w485 = w497 & ~w569;
assign w486 = ~w54 & ~w197;
assign w487 = ~w605 & w595;
assign w488 = (w230 & w476) | (w230 & w458) | (w476 & w458);
assign w489 = (w230 & w476) | (w230 & w267) | (w476 & w267);
assign w490 = ~w181 & ~w318;
assign w491 = ~w451 & ~w364;
assign w492 = ~w356 & w513;
assign w493 = (w7 & w208) | (w7 & w128) | (w208 & w128);
assign w494 = (w580 & w214) | (w580 & w63) | (w214 & w63);
assign w495 = ~w338 & w571;
assign w496 = ~w251 & ~w100;
assign w497 = ~b13 & ~a13;
assign w498 = ~w268 & ~w601;
assign w499 = (w580 & w42) | (w580 & w328) | (w42 & w328);
assign w500 = ~b3 & ~a3;
assign w501 = ~w318 & ~w111;
assign w502 = (w288 & w554) | (w288 & ~w270) | (w554 & ~w270);
assign w503 = ~w539 & ~w196;
assign w504 = b23 & a23;
assign w505 = (w314 & w542) | (w314 & w237) | (w542 & w237);
assign w506 = (~w184 & w278) | (~w184 & w57) | (w278 & w57);
assign w507 = (~w560 & w38) | (~w560 & w537) | (w38 & w537);
assign w508 = ~w18 & w394;
assign w509 = ~w587 & w155;
assign w510 = ~w578 & ~w602;
assign w511 = ~w54 & ~w248;
assign w512 = w227 & w132;
assign w513 = ~w168 & ~w238;
assign w514 = ~w522 & ~w113;
assign w515 = ~w539 & ~w106;
assign w516 = (w244 & w187) | (w244 & w401) | (w187 & w401);
assign w517 = ~w153 & ~w271;
assign w518 = ~w445 & ~w215;
assign w519 = ~w268 & ~w327;
assign w520 = w315 & ~w100;
assign w521 = ~w227 & ~w132;
assign w522 = w478 & w579;
assign w523 = ~w471 & ~w560;
assign w524 = w534 & ~w308;
assign w525 = w600 & ~w245;
assign w526 = (~w371 & w593) | (~w371 & w396) | (w593 & w396);
assign w527 = w346 & ~w66;
assign w528 = ~w181 & ~w111;
assign w529 = ~b24 & ~a24;
assign w530 = w229 & ~w543;
assign w531 = w363 & ~w540;
assign w532 = w597 & ~w453;
assign w533 = ~w48 & ~w158;
assign w534 = (~w168 & w603) | (~w168 & w459) | (w603 & w459);
assign w535 = (~w575 & w179) | (~w575 & w123) | (w179 & w123);
assign w536 = (w204 & w559) | (w204 & ~w137) | (w559 & ~w137);
assign w537 = ~w284 & w101;
assign w538 = (w65 & ~w244) | (w65 & w367) | (~w244 & w367);
assign w539 = b11 & a11;
assign w540 = w572 & ~w167;
assign w541 = ~w331 & w11;
assign w542 = w153 & w314;
assign w543 = cin & w276;
assign w544 = w181 & w111;
assign w545 = (w148 & w584) | (w148 & w222) | (w584 & w222);
assign w546 = w596 & ~w38;
assign w547 = (w580 & w519) | (w580 & w498) | (w519 & w498);
assign w548 = (~w75 & w43) | (~w75 & w1) | (w43 & w1);
assign w549 = w378 & ~w429;
assign w550 = (w75 & w361) | (w75 & w609) | (w361 & w609);
assign w551 = w86 & w140;
assign w552 = (~w213 & ~w595) | (~w213 & ~w137) | (~w595 & ~w137);
assign w553 = (~w429 & w378) | (~w429 & w233) | (w378 & w233);
assign w554 = ~w280 & w58;
assign w555 = ~w497 & w398;
assign w556 = ~w285 & w89;
assign w557 = ~w422 & ~w257;
assign w558 = w144 & w346;
assign w559 = (w520 & w505) | (w520 & w126) | (w505 & w126);
assign w560 = (~w148 & w441) | (~w148 & w502) | (w441 & w502);
assign w561 = ~w568 & ~w139;
assign w562 = (~w386 & w268) | (~w386 & w67) | (w268 & w67);
assign w563 = (~w338 & w283) | (~w338 & w425) | (w283 & w425);
assign w564 = ~w284 & ~w145;
assign w565 = ~b19 & ~a19;
assign w566 = w559 | w204;
assign w567 = (w148 & w170) | (w148 & w448) | (w170 & w448);
assign w568 = ~b7 & ~a7;
assign w569 = b14 & a14;
assign w570 = w534 & w371;
assign w571 = w518 & ~w508;
assign w572 = ~w573 & w556;
assign w573 = ~b21 & ~a21;
assign w574 = (w75 & w533) | (w75 & w302) | (w533 & w302);
assign w575 = b26 & a26;
assign w576 = (w520 & ~w84) | (w520 & w234) | (~w84 & w234);
assign w577 = w371 & ~w282;
assign w578 = a31 & b31;
assign w579 = ~w196 & ~w92;
assign w580 = (~w467 & ~w7) | (~w467 & w444) | (~w7 & w444);
assign w581 = ~b4 & ~a4;
assign w582 = ~w48 & w386;
assign w583 = ~w174 & w207;
assign w584 = w432 & w344;
assign w585 = w437 & w338;
assign w586 = ~w323 & ~w274;
assign w587 = ~w575 & ~w178;
assign w588 = ~w412 & ~w530;
assign w589 = ~w382 & w29;
assign w590 = w572 & ~w149;
assign w591 = (w137 & w487) | (w137 & w68) | (w487 & w68);
assign w592 = w539 & w106;
assign w593 = (~w371 & ~w580) | (~w371 & w320) | (~w580 & w320);
assign w594 = ~w538 & ~w516;
assign w595 = w117 & w558;
assign w596 = ~w145 & w224;
assign w597 = ~w527 & ~w236;
assign w598 = (w8 & w92) | (w8 & w262) | (w92 & w262);
assign w599 = (w465 & w133) | (w465 & w418) | (w133 & w418);
assign w600 = ~w465 & w176;
assign w601 = (w327 & ~w534) | (w327 & w185) | (~w534 & w185);
assign w602 = (~w75 & w566) | (~w75 & w536) | (w566 & w536);
assign w603 = w388 & w411;
assign w604 = ~w144 & ~w437;
assign w605 = ~w76 & ~w474;
assign w606 = ~w52 & w438;
assign w607 = (~w224 & w359) | (~w224 & w537) | (w359 & w537);
assign w608 = ~w211 & w583;
assign w609 = (w137 & w219) | (w137 & w477) | (w219 & w477);
assign one = 1;
assign s0 = w588;// level 5
assign s1 = ~w470;// level 6
assign s2 = w402;// level 6
assign s3 = w98;// level 7
assign s4 = w35;// level 7
assign s5 = w74;// level 7
assign s6 = w122;// level 7
assign s7 = ~w37;// level 8
assign s8 = w281;// level 8
assign s9 = ~w304;// level 8
assign s10 = w491;// level 8
assign s11 = w150;// level 9
assign s12 = w413;// level 9
assign s13 = ~w436;// level 10
assign s14 = ~w366;// level 9
assign s15 = w428;// level 9
assign s16 = ~w586;// level 11
assign s17 = ~w594;// level 11
assign s18 = w173;// level 11
assign s19 = w175;// level 11
assign s20 = ~w250;// level 11
assign s21 = w321;// level 11
assign s22 = w462;// level 11
assign s23 = ~w450;// level 11
assign s24 = ~w481;// level 11
assign s25 = w235;// level 11
assign s26 = ~w353;// level 12
assign s27 = ~w416;// level 12
assign s28 = ~w300;// level 12
assign s29 = ~w391;// level 12
assign s30 = w376;// level 12
assign s31 = w201;// level 11
assign s32 = ~w510;// level 11
endmodule
