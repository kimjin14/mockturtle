module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 ;
  assign n129 = x0 & x64 ;
  assign n130 = x2 & ~n129 ;
  assign n131 = ~x0 & x1 ;
  assign n132 = x64 & n131 ;
  assign n133 = ~x1 & x2 ;
  assign n134 = x1 & ~x2 ;
  assign n135 = n133 | n134 ;
  assign n136 = x0 & x65 ;
  assign n137 = ~n135 & n136 ;
  assign n138 = n132 | n137 ;
  assign n139 = x0 & n135 ;
  assign n140 = x64 & ~x65 ;
  assign n141 = ~x64 & x65 ;
  assign n142 = n140 | n141 ;
  assign n143 = n139 & n142 ;
  assign n144 = n138 | n143 ;
  assign n145 = x2 & ~n144 ;
  assign n146 = ~x2 & n144 ;
  assign n147 = n145 | n146 ;
  assign n148 = n130 | n147 ;
  assign n149 = n130 & n147 ;
  assign n150 = n148 & ~n149 ;
  assign n151 = ~x66 & n141 ;
  assign n152 = x66 | n151 ;
  assign n153 = ( ~n141 & n151 ) | ( ~n141 & n152 ) | ( n151 & n152 ) ;
  assign n154 = n139 & n153 ;
  assign n155 = x65 & n131 ;
  assign n156 = x0 | x1 ;
  assign n157 = x64 & ~n156 ;
  assign n158 = ( n135 & n155 ) | ( n135 & n157 ) | ( n155 & n157 ) ;
  assign n159 = x0 & x66 ;
  assign n160 = ( ~n135 & n155 ) | ( ~n135 & n159 ) | ( n155 & n159 ) ;
  assign n161 = n158 | n160 ;
  assign n162 = n154 | n161 ;
  assign n163 = x2 & ~n162 ;
  assign n164 = ~x2 & n162 ;
  assign n165 = n163 | n164 ;
  assign n166 = n149 & n165 ;
  assign n167 = n149 | n165 ;
  assign n168 = ~n166 & n167 ;
  assign n169 = x2 & ~x3 ;
  assign n170 = ~x2 & x3 ;
  assign n171 = n169 | n170 ;
  assign n172 = x64 & n171 ;
  assign n173 = x66 | x67 ;
  assign n174 = x66 & x67 ;
  assign n175 = n173 & ~n174 ;
  assign n176 = ( x64 & n141 ) | ( x64 & ~n142 ) | ( n141 & ~n142 ) ;
  assign n177 = ( x65 & x66 ) | ( x65 & n176 ) | ( x66 & n176 ) ;
  assign n178 = n175 & n177 ;
  assign n179 = n175 | n177 ;
  assign n180 = ~n178 & n179 ;
  assign n181 = n139 & n180 ;
  assign n182 = x66 & n131 ;
  assign n183 = x65 & ~n156 ;
  assign n184 = ( n135 & n182 ) | ( n135 & n183 ) | ( n182 & n183 ) ;
  assign n185 = x0 & x67 ;
  assign n186 = ( ~n135 & n182 ) | ( ~n135 & n185 ) | ( n182 & n185 ) ;
  assign n187 = n184 | n186 ;
  assign n188 = n181 | n187 ;
  assign n189 = x2 | n188 ;
  assign n190 = ~x2 & n189 ;
  assign n191 = ( ~n188 & n189 ) | ( ~n188 & n190 ) | ( n189 & n190 ) ;
  assign n192 = n172 & n191 ;
  assign n193 = n172 | n191 ;
  assign n194 = ~n192 & n193 ;
  assign n195 = n166 & n194 ;
  assign n196 = n166 | n194 ;
  assign n197 = ~n195 & n196 ;
  assign n198 = ~x3 & x4 ;
  assign n199 = x3 & ~x4 ;
  assign n200 = n198 | n199 ;
  assign n201 = ~n171 & n200 ;
  assign n202 = x64 & n201 ;
  assign n203 = ~x4 & x5 ;
  assign n204 = x4 & ~x5 ;
  assign n205 = n203 | n204 ;
  assign n206 = n171 & ~n205 ;
  assign n207 = x65 & n206 ;
  assign n208 = n202 | n207 ;
  assign n209 = n171 & n205 ;
  assign n210 = n142 & n209 ;
  assign n211 = n208 | n210 ;
  assign n212 = x5 | n211 ;
  assign n213 = ~x5 & n212 ;
  assign n214 = ( ~n211 & n212 ) | ( ~n211 & n213 ) | ( n212 & n213 ) ;
  assign n215 = x5 & ~n172 ;
  assign n216 = n214 & n215 ;
  assign n217 = n214 | n215 ;
  assign n218 = ~n216 & n217 ;
  assign n219 = x67 & n131 ;
  assign n220 = x66 & ~n156 ;
  assign n221 = ( n135 & n219 ) | ( n135 & n220 ) | ( n219 & n220 ) ;
  assign n222 = x0 & x68 ;
  assign n223 = ( ~n135 & n219 ) | ( ~n135 & n222 ) | ( n219 & n222 ) ;
  assign n224 = n221 | n223 ;
  assign n225 = n139 | n224 ;
  assign n226 = n174 | n178 ;
  assign n227 = ( x67 & ~x68 ) | ( x67 & n226 ) | ( ~x68 & n226 ) ;
  assign n228 = ( ~x67 & x68 ) | ( ~x67 & n227 ) | ( x68 & n227 ) ;
  assign n229 = ( ~n226 & n227 ) | ( ~n226 & n228 ) | ( n227 & n228 ) ;
  assign n230 = ( n224 & n225 ) | ( n224 & n229 ) | ( n225 & n229 ) ;
  assign n231 = x2 & ~n230 ;
  assign n232 = ~x2 & n230 ;
  assign n233 = n231 | n232 ;
  assign n234 = n218 & n233 ;
  assign n235 = n218 & ~n234 ;
  assign n236 = n233 & ~n234 ;
  assign n237 = n235 | n236 ;
  assign n238 = n192 | n195 ;
  assign n239 = n237 & n238 ;
  assign n240 = n237 | n238 ;
  assign n241 = ~n239 & n240 ;
  assign n242 = x65 & n201 ;
  assign n243 = ~n171 & n205 ;
  assign n244 = x64 & ~n200 ;
  assign n245 = n243 & n244 ;
  assign n246 = n242 | n245 ;
  assign n247 = x66 & n206 ;
  assign n248 = n246 | n247 ;
  assign n249 = ( n153 & n209 ) | ( n153 & n248 ) | ( n209 & n248 ) ;
  assign n250 = n248 | n249 ;
  assign n251 = x5 & ~n250 ;
  assign n252 = ~x5 & n250 ;
  assign n253 = n251 | n252 ;
  assign n254 = n216 & n253 ;
  assign n255 = n216 | n253 ;
  assign n256 = ~n254 & n255 ;
  assign n257 = x68 | x69 ;
  assign n258 = x68 & x69 ;
  assign n259 = n257 & ~n258 ;
  assign n260 = x67 & x68 ;
  assign n261 = ( n226 & ~n229 ) | ( n226 & n260 ) | ( ~n229 & n260 ) ;
  assign n262 = n259 & n261 ;
  assign n263 = n259 | n261 ;
  assign n264 = ~n262 & n263 ;
  assign n265 = x68 & n131 ;
  assign n266 = x67 & ~n156 ;
  assign n267 = ( n135 & n265 ) | ( n135 & n266 ) | ( n265 & n266 ) ;
  assign n268 = x0 & x69 ;
  assign n269 = ( ~n135 & n265 ) | ( ~n135 & n268 ) | ( n265 & n268 ) ;
  assign n270 = n267 | n269 ;
  assign n271 = n139 | n270 ;
  assign n272 = ( n264 & n270 ) | ( n264 & n271 ) | ( n270 & n271 ) ;
  assign n273 = x2 & ~n272 ;
  assign n274 = ~x2 & n272 ;
  assign n275 = n273 | n274 ;
  assign n276 = n256 & n275 ;
  assign n277 = n256 & ~n276 ;
  assign n278 = ~n256 & n275 ;
  assign n279 = n277 | n278 ;
  assign n280 = n234 | n239 ;
  assign n281 = n279 & n280 ;
  assign n282 = n279 | n280 ;
  assign n283 = ~n281 & n282 ;
  assign n284 = n276 | n281 ;
  assign n285 = x67 & n206 ;
  assign n286 = x66 & n201 ;
  assign n287 = x65 & ~n200 ;
  assign n288 = n243 & n287 ;
  assign n289 = n286 | n288 ;
  assign n290 = n285 | n289 ;
  assign n291 = n180 & n209 ;
  assign n292 = n290 | n291 ;
  assign n293 = x5 & ~n292 ;
  assign n294 = ~x5 & n292 ;
  assign n295 = n293 | n294 ;
  assign n296 = x5 & ~x6 ;
  assign n297 = ~x5 & x6 ;
  assign n298 = n296 | n297 ;
  assign n299 = x64 & n298 ;
  assign n300 = ( n254 & n295 ) | ( n254 & ~n299 ) | ( n295 & ~n299 ) ;
  assign n301 = ( ~n254 & n299 ) | ( ~n254 & n300 ) | ( n299 & n300 ) ;
  assign n302 = ( ~n295 & n300 ) | ( ~n295 & n301 ) | ( n300 & n301 ) ;
  assign n303 = x69 | x70 ;
  assign n304 = x69 & x70 ;
  assign n305 = n303 & ~n304 ;
  assign n306 = n258 & n305 ;
  assign n307 = ( n262 & n305 ) | ( n262 & n306 ) | ( n305 & n306 ) ;
  assign n308 = n258 | n305 ;
  assign n309 = n262 | n308 ;
  assign n310 = ~n307 & n309 ;
  assign n311 = x69 & n131 ;
  assign n312 = x68 & ~n156 ;
  assign n313 = ( n135 & n311 ) | ( n135 & n312 ) | ( n311 & n312 ) ;
  assign n314 = x0 & x70 ;
  assign n315 = ( ~n135 & n311 ) | ( ~n135 & n314 ) | ( n311 & n314 ) ;
  assign n316 = n313 | n315 ;
  assign n317 = ( n139 & n310 ) | ( n139 & n316 ) | ( n310 & n316 ) ;
  assign n318 = ( x2 & ~n316 ) | ( x2 & n317 ) | ( ~n316 & n317 ) ;
  assign n319 = ~n317 & n318 ;
  assign n320 = n316 | n318 ;
  assign n321 = ( ~x2 & n319 ) | ( ~x2 & n320 ) | ( n319 & n320 ) ;
  assign n322 = n302 & n321 ;
  assign n323 = n302 | n321 ;
  assign n324 = ~n322 & n323 ;
  assign n325 = n284 & n324 ;
  assign n326 = n284 | n324 ;
  assign n327 = ~n325 & n326 ;
  assign n328 = n322 | n325 ;
  assign n329 = ~x6 & x7 ;
  assign n330 = x6 & ~x7 ;
  assign n331 = n329 | n330 ;
  assign n332 = ~n298 & n331 ;
  assign n333 = x64 & n332 ;
  assign n334 = ~x7 & x8 ;
  assign n335 = x7 & ~x8 ;
  assign n336 = n334 | n335 ;
  assign n337 = n298 & ~n336 ;
  assign n338 = x65 & n337 ;
  assign n339 = n333 | n338 ;
  assign n340 = n298 & n336 ;
  assign n341 = n142 & n340 ;
  assign n342 = n339 | n341 ;
  assign n343 = x8 | n342 ;
  assign n344 = ~x8 & n343 ;
  assign n345 = ( ~n342 & n343 ) | ( ~n342 & n344 ) | ( n343 & n344 ) ;
  assign n346 = x8 & ~n299 ;
  assign n347 = n345 & n346 ;
  assign n348 = n345 | n346 ;
  assign n349 = ~n347 & n348 ;
  assign n350 = n209 & n229 ;
  assign n351 = x68 & n206 ;
  assign n352 = x67 & n201 ;
  assign n353 = x66 & ~n200 ;
  assign n354 = n243 & n353 ;
  assign n355 = n352 | n354 ;
  assign n356 = n351 | n355 ;
  assign n357 = n350 | n356 ;
  assign n358 = x5 | n357 ;
  assign n359 = ~x5 & n358 ;
  assign n360 = ( ~n357 & n358 ) | ( ~n357 & n359 ) | ( n358 & n359 ) ;
  assign n361 = n349 & n360 ;
  assign n362 = n349 & ~n361 ;
  assign n363 = n360 & ~n361 ;
  assign n364 = n362 | n363 ;
  assign n365 = ( n254 & n295 ) | ( n254 & n299 ) | ( n295 & n299 ) ;
  assign n366 = n364 | n365 ;
  assign n367 = n364 & n365 ;
  assign n368 = n366 & ~n367 ;
  assign n369 = x70 | x71 ;
  assign n370 = x70 & x71 ;
  assign n371 = n369 & ~n370 ;
  assign n372 = n304 | n306 ;
  assign n373 = ( n262 & n303 ) | ( n262 & n372 ) | ( n303 & n372 ) ;
  assign n374 = n371 & n373 ;
  assign n375 = n371 | n373 ;
  assign n376 = ~n374 & n375 ;
  assign n377 = x70 & n131 ;
  assign n378 = x69 & ~n156 ;
  assign n379 = ( n135 & n377 ) | ( n135 & n378 ) | ( n377 & n378 ) ;
  assign n380 = x0 & x71 ;
  assign n381 = ( ~n135 & n377 ) | ( ~n135 & n380 ) | ( n377 & n380 ) ;
  assign n382 = n379 | n381 ;
  assign n383 = ( n139 & n376 ) | ( n139 & n382 ) | ( n376 & n382 ) ;
  assign n384 = ( x2 & ~n382 ) | ( x2 & n383 ) | ( ~n382 & n383 ) ;
  assign n385 = ~n383 & n384 ;
  assign n386 = n382 | n384 ;
  assign n387 = ( ~x2 & n385 ) | ( ~x2 & n386 ) | ( n385 & n386 ) ;
  assign n388 = n368 & n387 ;
  assign n389 = n368 | n387 ;
  assign n390 = ~n388 & n389 ;
  assign n391 = n328 & n390 ;
  assign n392 = n328 | n390 ;
  assign n393 = ~n391 & n392 ;
  assign n394 = x66 & n337 ;
  assign n395 = x65 & n332 ;
  assign n396 = ~n298 & n336 ;
  assign n397 = x64 & ~n331 ;
  assign n398 = n396 & n397 ;
  assign n399 = n395 | n398 ;
  assign n400 = n394 | n399 ;
  assign n401 = n153 & n340 ;
  assign n402 = n400 | n401 ;
  assign n403 = x8 | n402 ;
  assign n404 = ~x8 & n403 ;
  assign n405 = ( ~n402 & n403 ) | ( ~n402 & n404 ) | ( n403 & n404 ) ;
  assign n406 = n347 | n405 ;
  assign n407 = n347 & n405 ;
  assign n408 = n406 & ~n407 ;
  assign n409 = n209 & n264 ;
  assign n410 = x69 & n206 ;
  assign n411 = x68 & n201 ;
  assign n412 = x67 & ~n200 ;
  assign n413 = n243 & n412 ;
  assign n414 = n411 | n413 ;
  assign n415 = n410 | n414 ;
  assign n416 = n409 | n415 ;
  assign n417 = x5 | n416 ;
  assign n418 = ~x5 & n417 ;
  assign n419 = ( ~n416 & n417 ) | ( ~n416 & n418 ) | ( n417 & n418 ) ;
  assign n420 = n408 & n419 ;
  assign n421 = n408 & ~n420 ;
  assign n422 = ~n408 & n419 ;
  assign n423 = n421 | n422 ;
  assign n424 = n361 | n367 ;
  assign n425 = n423 | n424 ;
  assign n426 = n423 & n424 ;
  assign n427 = n425 & ~n426 ;
  assign n428 = x71 | x72 ;
  assign n429 = x71 & x72 ;
  assign n430 = n428 & ~n429 ;
  assign n431 = n370 & n430 ;
  assign n432 = ( n374 & n430 ) | ( n374 & n431 ) | ( n430 & n431 ) ;
  assign n433 = n370 | n430 ;
  assign n434 = n374 | n433 ;
  assign n435 = ~n432 & n434 ;
  assign n436 = x71 & n131 ;
  assign n437 = x70 & ~n156 ;
  assign n438 = ( n135 & n436 ) | ( n135 & n437 ) | ( n436 & n437 ) ;
  assign n439 = x0 & x72 ;
  assign n440 = ( ~n135 & n436 ) | ( ~n135 & n439 ) | ( n436 & n439 ) ;
  assign n441 = n438 | n440 ;
  assign n442 = n139 | n441 ;
  assign n443 = ( n435 & n441 ) | ( n435 & n442 ) | ( n441 & n442 ) ;
  assign n444 = x2 & n443 ;
  assign n445 = x2 & ~n444 ;
  assign n446 = ( n443 & ~n444 ) | ( n443 & n445 ) | ( ~n444 & n445 ) ;
  assign n447 = n427 & n446 ;
  assign n448 = n427 & ~n447 ;
  assign n449 = ~n427 & n446 ;
  assign n450 = n448 | n449 ;
  assign n451 = n388 | n391 ;
  assign n452 = n450 & n451 ;
  assign n453 = n450 | n451 ;
  assign n454 = ~n452 & n453 ;
  assign n455 = x8 & ~x9 ;
  assign n456 = ~x8 & x9 ;
  assign n457 = n455 | n456 ;
  assign n458 = x64 & n457 ;
  assign n459 = x67 & n337 ;
  assign n460 = x66 & n332 ;
  assign n461 = x65 & ~n331 ;
  assign n462 = n396 & n461 ;
  assign n463 = n460 | n462 ;
  assign n464 = n459 | n463 ;
  assign n465 = n180 & n340 ;
  assign n466 = n464 | n465 ;
  assign n467 = x8 & ~n466 ;
  assign n468 = ~x8 & n466 ;
  assign n469 = n467 | n468 ;
  assign n470 = ( n407 & n458 ) | ( n407 & n469 ) | ( n458 & n469 ) ;
  assign n471 = ( n407 & n469 ) | ( n407 & ~n470 ) | ( n469 & ~n470 ) ;
  assign n472 = ( n458 & ~n470 ) | ( n458 & n471 ) | ( ~n470 & n471 ) ;
  assign n473 = x70 & n206 ;
  assign n474 = x69 & n201 ;
  assign n475 = x68 & ~n200 ;
  assign n476 = n243 & n475 ;
  assign n477 = n474 | n476 ;
  assign n478 = n473 | n477 ;
  assign n479 = n209 | n478 ;
  assign n480 = ( n310 & n478 ) | ( n310 & n479 ) | ( n478 & n479 ) ;
  assign n481 = x5 & ~n480 ;
  assign n482 = ~x5 & n480 ;
  assign n483 = n481 | n482 ;
  assign n484 = n472 & n483 ;
  assign n485 = n472 & ~n484 ;
  assign n486 = ~n472 & n483 ;
  assign n487 = n485 | n486 ;
  assign n488 = n420 | n426 ;
  assign n489 = n487 | n488 ;
  assign n490 = n487 & n488 ;
  assign n491 = n489 & ~n490 ;
  assign n492 = x72 | x73 ;
  assign n493 = x72 & x73 ;
  assign n494 = n492 & ~n493 ;
  assign n495 = n429 | n431 ;
  assign n496 = ( n374 & n428 ) | ( n374 & n495 ) | ( n428 & n495 ) ;
  assign n497 = n494 | n496 ;
  assign n498 = n494 & n496 ;
  assign n499 = n497 & ~n498 ;
  assign n500 = x72 & n131 ;
  assign n501 = x71 & ~n156 ;
  assign n502 = ( n135 & n500 ) | ( n135 & n501 ) | ( n500 & n501 ) ;
  assign n503 = x0 & x73 ;
  assign n504 = ( ~n135 & n500 ) | ( ~n135 & n503 ) | ( n500 & n503 ) ;
  assign n505 = n502 | n504 ;
  assign n506 = n139 | n505 ;
  assign n507 = ( n499 & n505 ) | ( n499 & n506 ) | ( n505 & n506 ) ;
  assign n508 = x2 & n507 ;
  assign n509 = x2 & ~n508 ;
  assign n510 = ( n507 & ~n508 ) | ( n507 & n509 ) | ( ~n508 & n509 ) ;
  assign n511 = n491 & n510 ;
  assign n512 = n491 & ~n511 ;
  assign n513 = ~n491 & n510 ;
  assign n514 = n512 | n513 ;
  assign n515 = n447 | n452 ;
  assign n516 = n514 & n515 ;
  assign n517 = n514 | n515 ;
  assign n518 = ~n516 & n517 ;
  assign n519 = n511 | n516 ;
  assign n520 = ~x9 & x10 ;
  assign n521 = x9 & ~x10 ;
  assign n522 = n520 | n521 ;
  assign n523 = ~n457 & n522 ;
  assign n524 = x64 & n523 ;
  assign n525 = ~x10 & x11 ;
  assign n526 = x10 & ~x11 ;
  assign n527 = n525 | n526 ;
  assign n528 = n457 & ~n527 ;
  assign n529 = x65 & n528 ;
  assign n530 = n524 | n529 ;
  assign n531 = n457 & n527 ;
  assign n532 = n142 & n531 ;
  assign n533 = n530 | n532 ;
  assign n534 = x11 | n533 ;
  assign n535 = ~x11 & n534 ;
  assign n536 = ( ~n533 & n534 ) | ( ~n533 & n535 ) | ( n534 & n535 ) ;
  assign n537 = x11 & ~n458 ;
  assign n538 = n536 & n537 ;
  assign n539 = n536 | n537 ;
  assign n540 = ~n538 & n539 ;
  assign n541 = n229 & n340 ;
  assign n542 = x68 & n337 ;
  assign n543 = x67 & n332 ;
  assign n544 = x66 & ~n331 ;
  assign n545 = n396 & n544 ;
  assign n546 = n543 | n545 ;
  assign n547 = n542 | n546 ;
  assign n548 = n541 | n547 ;
  assign n549 = x8 | n548 ;
  assign n550 = ~x8 & n549 ;
  assign n551 = ( ~n548 & n549 ) | ( ~n548 & n550 ) | ( n549 & n550 ) ;
  assign n552 = n540 | n551 ;
  assign n553 = n540 & n551 ;
  assign n554 = n552 & ~n553 ;
  assign n555 = n470 | n554 ;
  assign n556 = n470 & n554 ;
  assign n557 = n555 & ~n556 ;
  assign n558 = x71 & n206 ;
  assign n559 = x70 & n201 ;
  assign n560 = x69 & ~n200 ;
  assign n561 = n243 & n560 ;
  assign n562 = n559 | n561 ;
  assign n563 = n558 | n562 ;
  assign n564 = n209 | n563 ;
  assign n565 = ( n376 & n563 ) | ( n376 & n564 ) | ( n563 & n564 ) ;
  assign n566 = x5 & ~n565 ;
  assign n567 = ~x5 & n565 ;
  assign n568 = n566 | n567 ;
  assign n569 = n557 & n568 ;
  assign n570 = n557 & ~n569 ;
  assign n571 = ~n557 & n568 ;
  assign n572 = n570 | n571 ;
  assign n573 = n484 | n490 ;
  assign n574 = n572 | n573 ;
  assign n575 = n572 & n573 ;
  assign n576 = n574 & ~n575 ;
  assign n577 = x73 & n131 ;
  assign n578 = x72 & ~n156 ;
  assign n579 = ( n135 & n577 ) | ( n135 & n578 ) | ( n577 & n578 ) ;
  assign n580 = x0 & x74 ;
  assign n581 = ( ~n135 & n577 ) | ( ~n135 & n580 ) | ( n577 & n580 ) ;
  assign n582 = n579 | n581 ;
  assign n583 = n139 | n582 ;
  assign n584 = n493 | n498 ;
  assign n585 = ( x73 & ~x74 ) | ( x73 & n584 ) | ( ~x74 & n584 ) ;
  assign n586 = ( ~x73 & x74 ) | ( ~x73 & n585 ) | ( x74 & n585 ) ;
  assign n587 = ( ~n584 & n585 ) | ( ~n584 & n586 ) | ( n585 & n586 ) ;
  assign n588 = ( n582 & n583 ) | ( n582 & n587 ) | ( n583 & n587 ) ;
  assign n589 = x2 & n588 ;
  assign n590 = x2 & ~n589 ;
  assign n591 = ( n588 & ~n589 ) | ( n588 & n590 ) | ( ~n589 & n590 ) ;
  assign n592 = n576 | n591 ;
  assign n593 = n576 & n591 ;
  assign n594 = n592 & ~n593 ;
  assign n595 = n519 | n594 ;
  assign n596 = n519 & n594 ;
  assign n597 = n595 & ~n596 ;
  assign n598 = n593 | n596 ;
  assign n599 = x73 | x74 ;
  assign n600 = x74 | x75 ;
  assign n601 = x74 & x75 ;
  assign n602 = n600 & ~n601 ;
  assign n603 = n599 & n602 ;
  assign n604 = x73 & x74 ;
  assign n605 = n602 & n604 ;
  assign n606 = ( n584 & n603 ) | ( n584 & n605 ) | ( n603 & n605 ) ;
  assign n607 = ( n584 & n599 ) | ( n584 & n604 ) | ( n599 & n604 ) ;
  assign n608 = n602 | n607 ;
  assign n609 = ~n606 & n608 ;
  assign n610 = x74 & n131 ;
  assign n611 = x73 & ~n156 ;
  assign n612 = ( n135 & n610 ) | ( n135 & n611 ) | ( n610 & n611 ) ;
  assign n613 = x0 & x75 ;
  assign n614 = ( ~n135 & n610 ) | ( ~n135 & n613 ) | ( n610 & n613 ) ;
  assign n615 = n612 | n614 ;
  assign n616 = n139 | n615 ;
  assign n617 = ( n609 & n615 ) | ( n609 & n616 ) | ( n615 & n616 ) ;
  assign n618 = x2 & n617 ;
  assign n619 = x2 & ~n618 ;
  assign n620 = ( n617 & ~n618 ) | ( n617 & n619 ) | ( ~n618 & n619 ) ;
  assign n621 = n569 | n575 ;
  assign n622 = x72 & n206 ;
  assign n623 = x71 & n201 ;
  assign n624 = x70 & ~n200 ;
  assign n625 = n243 & n624 ;
  assign n626 = n623 | n625 ;
  assign n627 = n622 | n626 ;
  assign n628 = n209 | n627 ;
  assign n629 = ( n435 & n627 ) | ( n435 & n628 ) | ( n627 & n628 ) ;
  assign n630 = x5 & n629 ;
  assign n631 = x5 | n629 ;
  assign n632 = ~n630 & n631 ;
  assign n633 = x66 & n528 ;
  assign n634 = x65 & n523 ;
  assign n635 = ~n457 & n527 ;
  assign n636 = x64 & ~n522 ;
  assign n637 = n635 & n636 ;
  assign n638 = n634 | n637 ;
  assign n639 = n633 | n638 ;
  assign n640 = n153 & n531 ;
  assign n641 = n639 | n640 ;
  assign n642 = x11 | n641 ;
  assign n643 = ~x11 & n642 ;
  assign n644 = ( ~n641 & n642 ) | ( ~n641 & n643 ) | ( n642 & n643 ) ;
  assign n645 = n538 | n644 ;
  assign n646 = n538 & n644 ;
  assign n647 = n645 & ~n646 ;
  assign n648 = n264 & n340 ;
  assign n649 = x69 & n337 ;
  assign n650 = x68 & n332 ;
  assign n651 = x67 & ~n331 ;
  assign n652 = n396 & n651 ;
  assign n653 = n650 | n652 ;
  assign n654 = n649 | n653 ;
  assign n655 = n648 | n654 ;
  assign n656 = x8 | n655 ;
  assign n657 = ~x8 & n656 ;
  assign n658 = ( ~n655 & n656 ) | ( ~n655 & n657 ) | ( n656 & n657 ) ;
  assign n659 = n647 & n658 ;
  assign n660 = n647 & ~n659 ;
  assign n661 = ~n647 & n658 ;
  assign n662 = n660 | n661 ;
  assign n663 = n553 | n556 ;
  assign n664 = n662 & n663 ;
  assign n665 = n662 | n663 ;
  assign n666 = ~n664 & n665 ;
  assign n667 = n632 & n666 ;
  assign n668 = n666 & ~n667 ;
  assign n669 = ( n632 & ~n667 ) | ( n632 & n668 ) | ( ~n667 & n668 ) ;
  assign n670 = ( n620 & n621 ) | ( n620 & ~n669 ) | ( n621 & ~n669 ) ;
  assign n671 = ( ~n621 & n669 ) | ( ~n621 & n670 ) | ( n669 & n670 ) ;
  assign n672 = ( ~n620 & n670 ) | ( ~n620 & n671 ) | ( n670 & n671 ) ;
  assign n673 = n598 & n672 ;
  assign n674 = n598 | n672 ;
  assign n675 = ~n673 & n674 ;
  assign n676 = x11 & ~x12 ;
  assign n677 = ~x11 & x12 ;
  assign n678 = n676 | n677 ;
  assign n679 = x64 & n678 ;
  assign n680 = x67 & n528 ;
  assign n681 = x66 & n523 ;
  assign n682 = x65 & ~n522 ;
  assign n683 = n635 & n682 ;
  assign n684 = n681 | n683 ;
  assign n685 = n680 | n684 ;
  assign n686 = n180 & n531 ;
  assign n687 = n685 | n686 ;
  assign n688 = x11 & ~n687 ;
  assign n689 = ~x11 & n687 ;
  assign n690 = n688 | n689 ;
  assign n691 = ( n646 & n679 ) | ( n646 & n690 ) | ( n679 & n690 ) ;
  assign n692 = ( n646 & n690 ) | ( n646 & ~n691 ) | ( n690 & ~n691 ) ;
  assign n693 = ( n679 & ~n691 ) | ( n679 & n692 ) | ( ~n691 & n692 ) ;
  assign n694 = x70 & n337 ;
  assign n695 = x69 & n332 ;
  assign n696 = x68 & ~n331 ;
  assign n697 = n396 & n696 ;
  assign n698 = n695 | n697 ;
  assign n699 = n694 | n698 ;
  assign n700 = n340 | n699 ;
  assign n701 = ( n310 & n699 ) | ( n310 & n700 ) | ( n699 & n700 ) ;
  assign n702 = x8 & ~n701 ;
  assign n703 = ~x8 & n701 ;
  assign n704 = n702 | n703 ;
  assign n705 = n693 & n704 ;
  assign n706 = n693 & ~n705 ;
  assign n707 = ~n693 & n704 ;
  assign n708 = n706 | n707 ;
  assign n709 = n659 | n664 ;
  assign n710 = n708 | n709 ;
  assign n711 = n708 & n709 ;
  assign n712 = n710 & ~n711 ;
  assign n713 = x73 & n206 ;
  assign n714 = x72 & n201 ;
  assign n715 = x71 & ~n200 ;
  assign n716 = n243 & n715 ;
  assign n717 = n714 | n716 ;
  assign n718 = n713 | n717 ;
  assign n719 = ( n209 & n499 ) | ( n209 & n718 ) | ( n499 & n718 ) ;
  assign n720 = ( x5 & ~n718 ) | ( x5 & n719 ) | ( ~n718 & n719 ) ;
  assign n721 = ~n719 & n720 ;
  assign n722 = n718 | n720 ;
  assign n723 = ( ~x5 & n721 ) | ( ~x5 & n722 ) | ( n721 & n722 ) ;
  assign n724 = n712 | n723 ;
  assign n725 = n712 & n723 ;
  assign n726 = n724 & ~n725 ;
  assign n727 = n621 & n669 ;
  assign n728 = n667 | n727 ;
  assign n729 = n726 & n728 ;
  assign n730 = n726 | n728 ;
  assign n731 = ~n729 & n730 ;
  assign n732 = x75 | x76 ;
  assign n733 = x75 & x76 ;
  assign n734 = n732 & ~n733 ;
  assign n735 = n601 | n603 ;
  assign n736 = n601 | n605 ;
  assign n737 = ( n584 & n735 ) | ( n584 & n736 ) | ( n735 & n736 ) ;
  assign n738 = n734 | n737 ;
  assign n739 = n734 & n737 ;
  assign n740 = n738 & ~n739 ;
  assign n741 = x75 & n131 ;
  assign n742 = x74 & ~n156 ;
  assign n743 = ( n135 & n741 ) | ( n135 & n742 ) | ( n741 & n742 ) ;
  assign n744 = x0 & x76 ;
  assign n745 = ( ~n135 & n741 ) | ( ~n135 & n744 ) | ( n741 & n744 ) ;
  assign n746 = n743 | n745 ;
  assign n747 = n139 | n746 ;
  assign n748 = ( n740 & n746 ) | ( n740 & n747 ) | ( n746 & n747 ) ;
  assign n749 = x2 & n748 ;
  assign n750 = x2 & ~n749 ;
  assign n751 = ( n748 & ~n749 ) | ( n748 & n750 ) | ( ~n749 & n750 ) ;
  assign n752 = n731 & n751 ;
  assign n753 = n731 & ~n752 ;
  assign n754 = ~n731 & n751 ;
  assign n755 = n753 | n754 ;
  assign n756 = ( n620 & n621 ) | ( n620 & n669 ) | ( n621 & n669 ) ;
  assign n757 = ( n673 & ~n727 ) | ( n673 & n756 ) | ( ~n727 & n756 ) ;
  assign n758 = n755 & n757 ;
  assign n759 = n755 | n757 ;
  assign n760 = ~n758 & n759 ;
  assign n761 = n752 | n758 ;
  assign n762 = n725 | n729 ;
  assign n763 = ~x12 & x13 ;
  assign n764 = x12 & ~x13 ;
  assign n765 = n763 | n764 ;
  assign n766 = ~n678 & n765 ;
  assign n767 = x64 & n766 ;
  assign n768 = ~x13 & x14 ;
  assign n769 = x13 & ~x14 ;
  assign n770 = n768 | n769 ;
  assign n771 = n678 & ~n770 ;
  assign n772 = x65 & n771 ;
  assign n773 = n767 | n772 ;
  assign n774 = n678 & n770 ;
  assign n775 = n142 & n774 ;
  assign n776 = n773 | n775 ;
  assign n777 = x14 | n776 ;
  assign n778 = ~x14 & n777 ;
  assign n779 = ( ~n776 & n777 ) | ( ~n776 & n778 ) | ( n777 & n778 ) ;
  assign n780 = x14 & ~n679 ;
  assign n781 = n779 & n780 ;
  assign n782 = n779 | n780 ;
  assign n783 = ~n781 & n782 ;
  assign n784 = n229 & n531 ;
  assign n785 = x68 & n528 ;
  assign n786 = x67 & n523 ;
  assign n787 = x66 & ~n522 ;
  assign n788 = n635 & n787 ;
  assign n789 = n786 | n788 ;
  assign n790 = n785 | n789 ;
  assign n791 = n784 | n790 ;
  assign n792 = x11 | n791 ;
  assign n793 = ~x11 & n792 ;
  assign n794 = ( ~n791 & n792 ) | ( ~n791 & n793 ) | ( n792 & n793 ) ;
  assign n795 = n783 | n794 ;
  assign n796 = n783 & n794 ;
  assign n797 = n795 & ~n796 ;
  assign n798 = n691 | n797 ;
  assign n799 = n691 & n797 ;
  assign n800 = n798 & ~n799 ;
  assign n801 = x71 & n337 ;
  assign n802 = x70 & n332 ;
  assign n803 = x69 & ~n331 ;
  assign n804 = n396 & n803 ;
  assign n805 = n802 | n804 ;
  assign n806 = n801 | n805 ;
  assign n807 = n340 | n806 ;
  assign n808 = ( n376 & n806 ) | ( n376 & n807 ) | ( n806 & n807 ) ;
  assign n809 = x8 & ~n808 ;
  assign n810 = ~x8 & n808 ;
  assign n811 = n809 | n810 ;
  assign n812 = n800 & n811 ;
  assign n813 = n800 & ~n812 ;
  assign n814 = ~n800 & n811 ;
  assign n815 = n813 | n814 ;
  assign n816 = n705 | n711 ;
  assign n817 = n815 | n816 ;
  assign n818 = n815 & n816 ;
  assign n819 = n817 & ~n818 ;
  assign n820 = x74 & n206 ;
  assign n821 = x73 & n201 ;
  assign n822 = x72 & ~n200 ;
  assign n823 = n243 & n822 ;
  assign n824 = n821 | n823 ;
  assign n825 = n820 | n824 ;
  assign n826 = n209 | n825 ;
  assign n827 = ( n587 & n825 ) | ( n587 & n826 ) | ( n825 & n826 ) ;
  assign n828 = x5 & n827 ;
  assign n829 = x5 & ~n828 ;
  assign n830 = ( n827 & ~n828 ) | ( n827 & n829 ) | ( ~n828 & n829 ) ;
  assign n831 = n819 | n830 ;
  assign n832 = n762 & n831 ;
  assign n833 = n819 & n830 ;
  assign n834 = n831 & ~n833 ;
  assign n835 = ~n832 & n834 ;
  assign n836 = x76 & n131 ;
  assign n837 = x75 & ~n156 ;
  assign n838 = ( n135 & n836 ) | ( n135 & n837 ) | ( n836 & n837 ) ;
  assign n839 = x0 & x77 ;
  assign n840 = ( ~n135 & n836 ) | ( ~n135 & n839 ) | ( n836 & n839 ) ;
  assign n841 = n838 | n840 ;
  assign n842 = n139 | n841 ;
  assign n843 = n733 | n739 ;
  assign n844 = ( x76 & ~x77 ) | ( x76 & n843 ) | ( ~x77 & n843 ) ;
  assign n845 = ( ~x76 & x77 ) | ( ~x76 & n844 ) | ( x77 & n844 ) ;
  assign n846 = ( ~n843 & n844 ) | ( ~n843 & n845 ) | ( n844 & n845 ) ;
  assign n847 = ( n841 & n842 ) | ( n841 & n846 ) | ( n842 & n846 ) ;
  assign n848 = x2 & n847 ;
  assign n849 = x2 & ~n848 ;
  assign n850 = ( n847 & ~n848 ) | ( n847 & n849 ) | ( ~n848 & n849 ) ;
  assign n851 = n762 & ~n834 ;
  assign n852 = ( n835 & ~n850 ) | ( n835 & n851 ) | ( ~n850 & n851 ) ;
  assign n853 = ( n850 & ~n851 ) | ( n850 & n852 ) | ( ~n851 & n852 ) ;
  assign n854 = ( ~n835 & n852 ) | ( ~n835 & n853 ) | ( n852 & n853 ) ;
  assign n855 = n761 & n854 ;
  assign n856 = n761 | n854 ;
  assign n857 = ~n855 & n856 ;
  assign n858 = x76 | x77 ;
  assign n859 = x77 | x78 ;
  assign n860 = x77 & x78 ;
  assign n861 = n859 & ~n860 ;
  assign n862 = n858 & n861 ;
  assign n863 = x76 & x77 ;
  assign n864 = n861 & n863 ;
  assign n865 = ( n843 & n862 ) | ( n843 & n864 ) | ( n862 & n864 ) ;
  assign n866 = ( n843 & n858 ) | ( n843 & n863 ) | ( n858 & n863 ) ;
  assign n867 = n861 | n866 ;
  assign n868 = ~n865 & n867 ;
  assign n869 = x77 & n131 ;
  assign n870 = x76 & ~n156 ;
  assign n871 = ( n135 & n869 ) | ( n135 & n870 ) | ( n869 & n870 ) ;
  assign n872 = x0 & x78 ;
  assign n873 = ( ~n135 & n869 ) | ( ~n135 & n872 ) | ( n869 & n872 ) ;
  assign n874 = n871 | n873 ;
  assign n875 = n139 | n874 ;
  assign n876 = ( n868 & n874 ) | ( n868 & n875 ) | ( n874 & n875 ) ;
  assign n877 = x2 & n876 ;
  assign n878 = x2 & ~n877 ;
  assign n879 = ( n876 & ~n877 ) | ( n876 & n878 ) | ( ~n877 & n878 ) ;
  assign n880 = n812 | n818 ;
  assign n881 = x72 & n337 ;
  assign n882 = x71 & n332 ;
  assign n883 = x70 & ~n331 ;
  assign n884 = n396 & n883 ;
  assign n885 = n882 | n884 ;
  assign n886 = n881 | n885 ;
  assign n887 = n340 | n886 ;
  assign n888 = ( n435 & n886 ) | ( n435 & n887 ) | ( n886 & n887 ) ;
  assign n889 = x8 & n888 ;
  assign n890 = x8 | n888 ;
  assign n891 = ~n889 & n890 ;
  assign n892 = n264 & n531 ;
  assign n893 = x69 & n528 ;
  assign n894 = x68 & n523 ;
  assign n895 = x67 & ~n522 ;
  assign n896 = n635 & n895 ;
  assign n897 = n894 | n896 ;
  assign n898 = n893 | n897 ;
  assign n899 = n892 | n898 ;
  assign n900 = x11 | n899 ;
  assign n901 = ~x11 & n900 ;
  assign n902 = ( ~n899 & n900 ) | ( ~n899 & n901 ) | ( n900 & n901 ) ;
  assign n903 = x66 & n771 ;
  assign n904 = x65 & n766 ;
  assign n905 = ~n678 & n770 ;
  assign n906 = x64 & ~n765 ;
  assign n907 = n905 & n906 ;
  assign n908 = n904 | n907 ;
  assign n909 = n903 | n908 ;
  assign n910 = n153 & n774 ;
  assign n911 = n909 | n910 ;
  assign n912 = x14 | n911 ;
  assign n913 = ~x14 & n912 ;
  assign n914 = ( ~n911 & n912 ) | ( ~n911 & n913 ) | ( n912 & n913 ) ;
  assign n915 = n781 | n914 ;
  assign n916 = n781 & n914 ;
  assign n917 = n915 & ~n916 ;
  assign n918 = n796 | n799 ;
  assign n919 = ( n902 & n917 ) | ( n902 & n918 ) | ( n917 & n918 ) ;
  assign n920 = ( n917 & n918 ) | ( n917 & ~n919 ) | ( n918 & ~n919 ) ;
  assign n921 = ( n902 & ~n919 ) | ( n902 & n920 ) | ( ~n919 & n920 ) ;
  assign n922 = n891 | n921 ;
  assign n923 = n891 & n921 ;
  assign n924 = n922 & ~n923 ;
  assign n925 = n880 & n924 ;
  assign n926 = n880 | n924 ;
  assign n927 = ~n925 & n926 ;
  assign n928 = x75 & n206 ;
  assign n929 = x74 & n201 ;
  assign n930 = x73 & ~n200 ;
  assign n931 = n243 & n930 ;
  assign n932 = n929 | n931 ;
  assign n933 = n928 | n932 ;
  assign n934 = n209 | n933 ;
  assign n935 = ( n609 & n933 ) | ( n609 & n934 ) | ( n933 & n934 ) ;
  assign n936 = x5 & n935 ;
  assign n937 = x5 & ~n936 ;
  assign n938 = ( n935 & ~n936 ) | ( n935 & n937 ) | ( ~n936 & n937 ) ;
  assign n939 = n927 | n938 ;
  assign n940 = n927 & n938 ;
  assign n941 = n939 & ~n940 ;
  assign n942 = n832 | n833 ;
  assign n943 = n941 & n942 ;
  assign n944 = n941 | n942 ;
  assign n945 = ~n943 & n944 ;
  assign n946 = n835 | n851 ;
  assign n947 = ( n761 & n850 ) | ( n761 & n946 ) | ( n850 & n946 ) ;
  assign n948 = ( n879 & n945 ) | ( n879 & n947 ) | ( n945 & n947 ) ;
  assign n949 = ( n945 & n947 ) | ( n945 & ~n948 ) | ( n947 & ~n948 ) ;
  assign n950 = ( n879 & ~n948 ) | ( n879 & n949 ) | ( ~n948 & n949 ) ;
  assign n951 = x78 | x79 ;
  assign n952 = x78 & x79 ;
  assign n953 = n951 & ~n952 ;
  assign n954 = n860 | n862 ;
  assign n955 = n953 & n954 ;
  assign n956 = n860 | n864 ;
  assign n957 = n953 & n956 ;
  assign n958 = ( n843 & n955 ) | ( n843 & n957 ) | ( n955 & n957 ) ;
  assign n959 = ( n843 & n954 ) | ( n843 & n956 ) | ( n954 & n956 ) ;
  assign n960 = n953 | n959 ;
  assign n961 = ~n958 & n960 ;
  assign n962 = x78 & n131 ;
  assign n963 = x77 & ~n156 ;
  assign n964 = ( n135 & n962 ) | ( n135 & n963 ) | ( n962 & n963 ) ;
  assign n965 = x0 & x79 ;
  assign n966 = ( ~n135 & n962 ) | ( ~n135 & n965 ) | ( n962 & n965 ) ;
  assign n967 = n964 | n966 ;
  assign n968 = n139 | n967 ;
  assign n969 = ( n961 & n967 ) | ( n961 & n968 ) | ( n967 & n968 ) ;
  assign n970 = x2 & n969 ;
  assign n971 = x2 & ~n970 ;
  assign n972 = ( n969 & ~n970 ) | ( n969 & n971 ) | ( ~n970 & n971 ) ;
  assign n973 = n940 | n943 ;
  assign n974 = n923 | n925 ;
  assign n975 = x73 & n337 ;
  assign n976 = x72 & n332 ;
  assign n977 = x71 & ~n331 ;
  assign n978 = n396 & n977 ;
  assign n979 = n976 | n978 ;
  assign n980 = n975 | n979 ;
  assign n981 = ( n340 & n499 ) | ( n340 & n980 ) | ( n499 & n980 ) ;
  assign n982 = ( x8 & ~n980 ) | ( x8 & n981 ) | ( ~n980 & n981 ) ;
  assign n983 = ~n981 & n982 ;
  assign n984 = n980 | n982 ;
  assign n985 = ( ~x8 & n983 ) | ( ~x8 & n984 ) | ( n983 & n984 ) ;
  assign n986 = x14 & ~x15 ;
  assign n987 = ~x14 & x15 ;
  assign n988 = n986 | n987 ;
  assign n989 = x64 & n988 ;
  assign n990 = x67 & n771 ;
  assign n991 = x66 & n766 ;
  assign n992 = x65 & ~n765 ;
  assign n993 = n905 & n992 ;
  assign n994 = n991 | n993 ;
  assign n995 = n990 | n994 ;
  assign n996 = n180 & n774 ;
  assign n997 = n995 | n996 ;
  assign n998 = x14 & ~n997 ;
  assign n999 = ~x14 & n997 ;
  assign n1000 = n998 | n999 ;
  assign n1001 = ( n916 & n989 ) | ( n916 & n1000 ) | ( n989 & n1000 ) ;
  assign n1002 = ( n916 & n1000 ) | ( n916 & ~n1001 ) | ( n1000 & ~n1001 ) ;
  assign n1003 = ( n989 & ~n1001 ) | ( n989 & n1002 ) | ( ~n1001 & n1002 ) ;
  assign n1004 = x70 & n528 ;
  assign n1005 = x69 & n523 ;
  assign n1006 = x68 & ~n522 ;
  assign n1007 = n635 & n1006 ;
  assign n1008 = n1005 | n1007 ;
  assign n1009 = n1004 | n1008 ;
  assign n1010 = n531 | n1009 ;
  assign n1011 = ( n310 & n1009 ) | ( n310 & n1010 ) | ( n1009 & n1010 ) ;
  assign n1012 = x11 & ~n1011 ;
  assign n1013 = ~x11 & n1011 ;
  assign n1014 = n1012 | n1013 ;
  assign n1015 = n1003 & n1014 ;
  assign n1016 = n1003 & ~n1015 ;
  assign n1017 = ~n1003 & n1014 ;
  assign n1018 = n919 | n1017 ;
  assign n1019 = n1016 | n1018 ;
  assign n1020 = ( n919 & n1016 ) | ( n919 & n1017 ) | ( n1016 & n1017 ) ;
  assign n1021 = n1019 & ~n1020 ;
  assign n1022 = n985 & n1021 ;
  assign n1023 = n1021 & ~n1022 ;
  assign n1024 = ( n985 & ~n1022 ) | ( n985 & n1023 ) | ( ~n1022 & n1023 ) ;
  assign n1025 = n974 & n1024 ;
  assign n1026 = n974 | n1024 ;
  assign n1027 = ~n1025 & n1026 ;
  assign n1028 = x76 & n206 ;
  assign n1029 = x75 & n201 ;
  assign n1030 = x74 & ~n200 ;
  assign n1031 = n243 & n1030 ;
  assign n1032 = n1029 | n1031 ;
  assign n1033 = n1028 | n1032 ;
  assign n1034 = n209 | n1033 ;
  assign n1035 = ( n740 & n1033 ) | ( n740 & n1034 ) | ( n1033 & n1034 ) ;
  assign n1036 = x5 & n1035 ;
  assign n1037 = x5 & ~n1036 ;
  assign n1038 = ( n1035 & ~n1036 ) | ( n1035 & n1037 ) | ( ~n1036 & n1037 ) ;
  assign n1039 = n1027 & n1038 ;
  assign n1040 = n1027 & ~n1039 ;
  assign n1041 = ~n1027 & n1038 ;
  assign n1042 = n1040 | n1041 ;
  assign n1043 = n973 & n1042 ;
  assign n1044 = n973 | n1042 ;
  assign n1045 = ~n1043 & n1044 ;
  assign n1046 = ( n948 & n972 ) | ( n948 & n1045 ) | ( n972 & n1045 ) ;
  assign n1047 = ( n948 & n1045 ) | ( n948 & ~n1046 ) | ( n1045 & ~n1046 ) ;
  assign n1048 = ( n972 & ~n1046 ) | ( n972 & n1047 ) | ( ~n1046 & n1047 ) ;
  assign n1049 = n1039 | n1043 ;
  assign n1050 = n1022 | n1025 ;
  assign n1051 = n1015 | n1020 ;
  assign n1052 = x71 & n528 ;
  assign n1053 = x70 & n523 ;
  assign n1054 = x69 & ~n522 ;
  assign n1055 = n635 & n1054 ;
  assign n1056 = n1053 | n1055 ;
  assign n1057 = n1052 | n1056 ;
  assign n1058 = n531 | n1057 ;
  assign n1059 = ( n376 & n1057 ) | ( n376 & n1058 ) | ( n1057 & n1058 ) ;
  assign n1060 = x11 & ~n1059 ;
  assign n1061 = ~x11 & n1059 ;
  assign n1062 = n1060 | n1061 ;
  assign n1063 = ~x15 & x16 ;
  assign n1064 = x15 & ~x16 ;
  assign n1065 = n1063 | n1064 ;
  assign n1066 = ~n988 & n1065 ;
  assign n1067 = x64 & n1066 ;
  assign n1068 = ~x16 & x17 ;
  assign n1069 = x16 & ~x17 ;
  assign n1070 = n1068 | n1069 ;
  assign n1071 = n988 & ~n1070 ;
  assign n1072 = x65 & n1071 ;
  assign n1073 = n1067 | n1072 ;
  assign n1074 = n988 & n1070 ;
  assign n1075 = n142 & n1074 ;
  assign n1076 = n1073 | n1075 ;
  assign n1077 = x17 | n1076 ;
  assign n1078 = ~x17 & n1077 ;
  assign n1079 = ( ~n1076 & n1077 ) | ( ~n1076 & n1078 ) | ( n1077 & n1078 ) ;
  assign n1080 = x17 & ~n989 ;
  assign n1081 = n1079 & n1080 ;
  assign n1082 = n1079 | n1080 ;
  assign n1083 = ~n1081 & n1082 ;
  assign n1084 = n229 & n774 ;
  assign n1085 = x68 & n771 ;
  assign n1086 = x67 & n766 ;
  assign n1087 = x66 & ~n765 ;
  assign n1088 = n905 & n1087 ;
  assign n1089 = n1086 | n1088 ;
  assign n1090 = n1085 | n1089 ;
  assign n1091 = n1084 | n1090 ;
  assign n1092 = x14 | n1091 ;
  assign n1093 = ~x14 & n1092 ;
  assign n1094 = ( ~n1091 & n1092 ) | ( ~n1091 & n1093 ) | ( n1092 & n1093 ) ;
  assign n1095 = n1083 | n1094 ;
  assign n1096 = n1083 & n1094 ;
  assign n1097 = n1095 & ~n1096 ;
  assign n1098 = n1001 | n1097 ;
  assign n1099 = n1001 & n1097 ;
  assign n1100 = n1098 & ~n1099 ;
  assign n1101 = n1062 | n1100 ;
  assign n1102 = n1062 & n1100 ;
  assign n1103 = n1101 & ~n1102 ;
  assign n1104 = n1051 & n1103 ;
  assign n1105 = n1051 | n1103 ;
  assign n1106 = ~n1104 & n1105 ;
  assign n1107 = x74 & n337 ;
  assign n1108 = x73 & n332 ;
  assign n1109 = x72 & ~n331 ;
  assign n1110 = n396 & n1109 ;
  assign n1111 = n1108 | n1110 ;
  assign n1112 = n1107 | n1111 ;
  assign n1113 = n340 | n1112 ;
  assign n1114 = ( n587 & n1112 ) | ( n587 & n1113 ) | ( n1112 & n1113 ) ;
  assign n1115 = x8 & n1114 ;
  assign n1116 = x8 & ~n1115 ;
  assign n1117 = ( n1114 & ~n1115 ) | ( n1114 & n1116 ) | ( ~n1115 & n1116 ) ;
  assign n1118 = n1106 | n1117 ;
  assign n1119 = n1106 & n1117 ;
  assign n1120 = n1118 & ~n1119 ;
  assign n1121 = n1050 & n1120 ;
  assign n1122 = n1050 | n1120 ;
  assign n1123 = ~n1121 & n1122 ;
  assign n1124 = x77 & n206 ;
  assign n1125 = x76 & n201 ;
  assign n1126 = x75 & ~n200 ;
  assign n1127 = n243 & n1126 ;
  assign n1128 = n1125 | n1127 ;
  assign n1129 = n1124 | n1128 ;
  assign n1130 = n209 | n1129 ;
  assign n1131 = ( n846 & n1129 ) | ( n846 & n1130 ) | ( n1129 & n1130 ) ;
  assign n1132 = x5 & n1131 ;
  assign n1133 = x5 & ~n1132 ;
  assign n1134 = ( n1131 & ~n1132 ) | ( n1131 & n1133 ) | ( ~n1132 & n1133 ) ;
  assign n1135 = n1123 | n1134 ;
  assign n1136 = n1123 & n1134 ;
  assign n1137 = n1135 & ~n1136 ;
  assign n1138 = n1049 & n1137 ;
  assign n1139 = n1049 | n1137 ;
  assign n1140 = ~n1138 & n1139 ;
  assign n1141 = x79 | x80 ;
  assign n1142 = x79 & x80 ;
  assign n1143 = n1141 & ~n1142 ;
  assign n1144 = n952 | n958 ;
  assign n1145 = n1143 & n1144 ;
  assign n1146 = n1143 | n1144 ;
  assign n1147 = ~n1145 & n1146 ;
  assign n1148 = x79 & n131 ;
  assign n1149 = x78 & ~n156 ;
  assign n1150 = ( n135 & n1148 ) | ( n135 & n1149 ) | ( n1148 & n1149 ) ;
  assign n1151 = x0 & x80 ;
  assign n1152 = ( ~n135 & n1148 ) | ( ~n135 & n1151 ) | ( n1148 & n1151 ) ;
  assign n1153 = n1150 | n1152 ;
  assign n1154 = n139 | n1153 ;
  assign n1155 = ( n1147 & n1153 ) | ( n1147 & n1154 ) | ( n1153 & n1154 ) ;
  assign n1156 = x2 & n1155 ;
  assign n1157 = x2 & ~n1156 ;
  assign n1158 = ( n1155 & ~n1156 ) | ( n1155 & n1157 ) | ( ~n1156 & n1157 ) ;
  assign n1159 = n1140 & n1158 ;
  assign n1160 = n1158 & ~n1159 ;
  assign n1161 = ( n1140 & ~n1159 ) | ( n1140 & n1160 ) | ( ~n1159 & n1160 ) ;
  assign n1162 = n1046 & n1161 ;
  assign n1163 = n1046 | n1161 ;
  assign n1164 = ~n1162 & n1163 ;
  assign n1165 = x72 & n528 ;
  assign n1166 = x71 & n523 ;
  assign n1167 = x70 & ~n522 ;
  assign n1168 = n635 & n1167 ;
  assign n1169 = n1166 | n1168 ;
  assign n1170 = n1165 | n1169 ;
  assign n1171 = ( n435 & n531 ) | ( n435 & n1170 ) | ( n531 & n1170 ) ;
  assign n1172 = ( x11 & ~n1170 ) | ( x11 & n1171 ) | ( ~n1170 & n1171 ) ;
  assign n1173 = ~n1171 & n1172 ;
  assign n1174 = n1170 | n1172 ;
  assign n1175 = ( ~x11 & n1173 ) | ( ~x11 & n1174 ) | ( n1173 & n1174 ) ;
  assign n1176 = n264 & n774 ;
  assign n1177 = x69 & n771 ;
  assign n1178 = x68 & n766 ;
  assign n1179 = x67 & ~n765 ;
  assign n1180 = n905 & n1179 ;
  assign n1181 = n1178 | n1180 ;
  assign n1182 = n1177 | n1181 ;
  assign n1183 = n1176 | n1182 ;
  assign n1184 = x14 | n1183 ;
  assign n1185 = ~x14 & n1184 ;
  assign n1186 = ( ~n1183 & n1184 ) | ( ~n1183 & n1185 ) | ( n1184 & n1185 ) ;
  assign n1187 = x66 & n1071 ;
  assign n1188 = x65 & n1066 ;
  assign n1189 = ~n988 & n1070 ;
  assign n1190 = x64 & ~n1065 ;
  assign n1191 = n1189 & n1190 ;
  assign n1192 = n1188 | n1191 ;
  assign n1193 = n1187 | n1192 ;
  assign n1194 = n153 & n1074 ;
  assign n1195 = n1193 | n1194 ;
  assign n1196 = x17 | n1195 ;
  assign n1197 = ~x17 & n1196 ;
  assign n1198 = ( ~n1195 & n1196 ) | ( ~n1195 & n1197 ) | ( n1196 & n1197 ) ;
  assign n1199 = n1081 | n1198 ;
  assign n1200 = n1081 & n1198 ;
  assign n1201 = n1199 & ~n1200 ;
  assign n1202 = n1096 | n1099 ;
  assign n1203 = ( n1186 & n1201 ) | ( n1186 & n1202 ) | ( n1201 & n1202 ) ;
  assign n1204 = ( n1201 & n1202 ) | ( n1201 & ~n1203 ) | ( n1202 & ~n1203 ) ;
  assign n1205 = ( n1186 & ~n1203 ) | ( n1186 & n1204 ) | ( ~n1203 & n1204 ) ;
  assign n1206 = n1175 | n1205 ;
  assign n1207 = n1175 & n1205 ;
  assign n1208 = n1206 & ~n1207 ;
  assign n1209 = n1102 | n1104 ;
  assign n1210 = n1208 & n1209 ;
  assign n1211 = n1208 | n1209 ;
  assign n1212 = ~n1210 & n1211 ;
  assign n1213 = x75 & n337 ;
  assign n1214 = x74 & n332 ;
  assign n1215 = x73 & ~n331 ;
  assign n1216 = n396 & n1215 ;
  assign n1217 = n1214 | n1216 ;
  assign n1218 = n1213 | n1217 ;
  assign n1219 = n340 | n1218 ;
  assign n1220 = ( n609 & n1218 ) | ( n609 & n1219 ) | ( n1218 & n1219 ) ;
  assign n1221 = x8 & n1220 ;
  assign n1222 = x8 & ~n1221 ;
  assign n1223 = ( n1220 & ~n1221 ) | ( n1220 & n1222 ) | ( ~n1221 & n1222 ) ;
  assign n1224 = n1212 | n1223 ;
  assign n1225 = n1212 & n1223 ;
  assign n1226 = n1224 & ~n1225 ;
  assign n1227 = n1119 | n1121 ;
  assign n1228 = n1226 & n1227 ;
  assign n1229 = n1226 | n1227 ;
  assign n1230 = ~n1228 & n1229 ;
  assign n1231 = x78 & n206 ;
  assign n1232 = x77 & n201 ;
  assign n1233 = x76 & ~n200 ;
  assign n1234 = n243 & n1233 ;
  assign n1235 = n1232 | n1234 ;
  assign n1236 = n1231 | n1235 ;
  assign n1237 = n209 | n1236 ;
  assign n1238 = ( n868 & n1236 ) | ( n868 & n1237 ) | ( n1236 & n1237 ) ;
  assign n1239 = x5 & n1238 ;
  assign n1240 = x5 & ~n1239 ;
  assign n1241 = ( n1238 & ~n1239 ) | ( n1238 & n1240 ) | ( ~n1239 & n1240 ) ;
  assign n1242 = n1230 | n1241 ;
  assign n1243 = n1230 & n1241 ;
  assign n1244 = n1242 & ~n1243 ;
  assign n1245 = n1136 | n1138 ;
  assign n1246 = n1244 & n1245 ;
  assign n1247 = n1244 | n1245 ;
  assign n1248 = ~n1246 & n1247 ;
  assign n1249 = x80 | x81 ;
  assign n1250 = x80 & x81 ;
  assign n1251 = n1249 & ~n1250 ;
  assign n1252 = n1142 & n1251 ;
  assign n1253 = ( n1145 & n1251 ) | ( n1145 & n1252 ) | ( n1251 & n1252 ) ;
  assign n1254 = n1142 | n1251 ;
  assign n1255 = n1145 | n1254 ;
  assign n1256 = ~n1253 & n1255 ;
  assign n1257 = x80 & n131 ;
  assign n1258 = x79 & ~n156 ;
  assign n1259 = ( n135 & n1257 ) | ( n135 & n1258 ) | ( n1257 & n1258 ) ;
  assign n1260 = x0 & x81 ;
  assign n1261 = ( ~n135 & n1257 ) | ( ~n135 & n1260 ) | ( n1257 & n1260 ) ;
  assign n1262 = n1259 | n1261 ;
  assign n1263 = n139 | n1262 ;
  assign n1264 = ( n1256 & n1262 ) | ( n1256 & n1263 ) | ( n1262 & n1263 ) ;
  assign n1265 = x2 & n1264 ;
  assign n1266 = x2 & ~n1265 ;
  assign n1267 = ( n1264 & ~n1265 ) | ( n1264 & n1266 ) | ( ~n1265 & n1266 ) ;
  assign n1268 = n1248 & n1267 ;
  assign n1269 = n1248 & ~n1268 ;
  assign n1270 = ~n1248 & n1267 ;
  assign n1271 = n1269 | n1270 ;
  assign n1272 = n1159 | n1162 ;
  assign n1273 = n1271 & n1272 ;
  assign n1274 = n1271 | n1272 ;
  assign n1275 = ~n1273 & n1274 ;
  assign n1276 = n1207 | n1210 ;
  assign n1277 = x70 & n771 ;
  assign n1278 = x69 & n766 ;
  assign n1279 = x68 & ~n765 ;
  assign n1280 = n905 & n1279 ;
  assign n1281 = n1278 | n1280 ;
  assign n1282 = n1277 | n1281 ;
  assign n1283 = n774 | n1282 ;
  assign n1284 = ( n310 & n1282 ) | ( n310 & n1283 ) | ( n1282 & n1283 ) ;
  assign n1285 = x14 & ~n1284 ;
  assign n1286 = ~x14 & n1284 ;
  assign n1287 = n1285 | n1286 ;
  assign n1288 = x17 & ~x18 ;
  assign n1289 = ~x17 & x18 ;
  assign n1290 = n1288 | n1289 ;
  assign n1291 = x64 & n1290 ;
  assign n1292 = x67 & n1071 ;
  assign n1293 = x66 & n1066 ;
  assign n1294 = x65 & ~n1065 ;
  assign n1295 = n1189 & n1294 ;
  assign n1296 = n1293 | n1295 ;
  assign n1297 = n1292 | n1296 ;
  assign n1298 = n180 & n1074 ;
  assign n1299 = n1297 | n1298 ;
  assign n1300 = x17 & ~n1299 ;
  assign n1301 = ~x17 & n1299 ;
  assign n1302 = n1300 | n1301 ;
  assign n1303 = ( n1200 & n1291 ) | ( n1200 & n1302 ) | ( n1291 & n1302 ) ;
  assign n1304 = ( n1200 & n1302 ) | ( n1200 & ~n1303 ) | ( n1302 & ~n1303 ) ;
  assign n1305 = ( n1291 & ~n1303 ) | ( n1291 & n1304 ) | ( ~n1303 & n1304 ) ;
  assign n1306 = ( n1203 & n1287 ) | ( n1203 & ~n1305 ) | ( n1287 & ~n1305 ) ;
  assign n1307 = ( ~n1203 & n1305 ) | ( ~n1203 & n1306 ) | ( n1305 & n1306 ) ;
  assign n1308 = ( ~n1287 & n1306 ) | ( ~n1287 & n1307 ) | ( n1306 & n1307 ) ;
  assign n1309 = x73 & n528 ;
  assign n1310 = x72 & n523 ;
  assign n1311 = x71 & ~n522 ;
  assign n1312 = n635 & n1311 ;
  assign n1313 = n1310 | n1312 ;
  assign n1314 = n1309 | n1313 ;
  assign n1315 = n531 | n1314 ;
  assign n1316 = ( n499 & n1314 ) | ( n499 & n1315 ) | ( n1314 & n1315 ) ;
  assign n1317 = x11 & n1316 ;
  assign n1318 = x11 | n1316 ;
  assign n1319 = ~n1317 & n1318 ;
  assign n1320 = n1308 & n1319 ;
  assign n1321 = n1308 | n1319 ;
  assign n1322 = ~n1320 & n1321 ;
  assign n1323 = n1276 & n1322 ;
  assign n1324 = n1276 | n1322 ;
  assign n1325 = ~n1323 & n1324 ;
  assign n1326 = x76 & n337 ;
  assign n1327 = x75 & n332 ;
  assign n1328 = x74 & ~n331 ;
  assign n1329 = n396 & n1328 ;
  assign n1330 = n1327 | n1329 ;
  assign n1331 = n1326 | n1330 ;
  assign n1332 = n340 | n1331 ;
  assign n1333 = ( n740 & n1331 ) | ( n740 & n1332 ) | ( n1331 & n1332 ) ;
  assign n1334 = x8 & n1333 ;
  assign n1335 = x8 & ~n1334 ;
  assign n1336 = ( n1333 & ~n1334 ) | ( n1333 & n1335 ) | ( ~n1334 & n1335 ) ;
  assign n1337 = n1325 | n1336 ;
  assign n1338 = n1325 & n1336 ;
  assign n1339 = n1337 & ~n1338 ;
  assign n1340 = n1225 | n1228 ;
  assign n1341 = n1339 & n1340 ;
  assign n1342 = n1339 | n1340 ;
  assign n1343 = ~n1341 & n1342 ;
  assign n1344 = x79 & n206 ;
  assign n1345 = x78 & n201 ;
  assign n1346 = x77 & ~n200 ;
  assign n1347 = n243 & n1346 ;
  assign n1348 = n1345 | n1347 ;
  assign n1349 = n1344 | n1348 ;
  assign n1350 = n209 | n1349 ;
  assign n1351 = ( n961 & n1349 ) | ( n961 & n1350 ) | ( n1349 & n1350 ) ;
  assign n1352 = x5 & n1351 ;
  assign n1353 = x5 & ~n1352 ;
  assign n1354 = ( n1351 & ~n1352 ) | ( n1351 & n1353 ) | ( ~n1352 & n1353 ) ;
  assign n1355 = n1343 & n1354 ;
  assign n1356 = n1343 | n1354 ;
  assign n1357 = ~n1355 & n1356 ;
  assign n1358 = n1243 | n1246 ;
  assign n1359 = n1357 & n1358 ;
  assign n1360 = n1357 | n1358 ;
  assign n1361 = ~n1359 & n1360 ;
  assign n1362 = x81 | x82 ;
  assign n1363 = x81 & x82 ;
  assign n1364 = n1362 & ~n1363 ;
  assign n1365 = n1250 | n1252 ;
  assign n1366 = n1364 & n1365 ;
  assign n1367 = n1249 & n1364 ;
  assign n1368 = ( n1145 & n1366 ) | ( n1145 & n1367 ) | ( n1366 & n1367 ) ;
  assign n1369 = ( n1145 & n1249 ) | ( n1145 & n1365 ) | ( n1249 & n1365 ) ;
  assign n1370 = n1364 | n1369 ;
  assign n1371 = ~n1368 & n1370 ;
  assign n1372 = x81 & n131 ;
  assign n1373 = x80 & ~n156 ;
  assign n1374 = ( n135 & n1372 ) | ( n135 & n1373 ) | ( n1372 & n1373 ) ;
  assign n1375 = x0 & x82 ;
  assign n1376 = ( ~n135 & n1372 ) | ( ~n135 & n1375 ) | ( n1372 & n1375 ) ;
  assign n1377 = n1374 | n1376 ;
  assign n1378 = n139 | n1377 ;
  assign n1379 = ( n1371 & n1377 ) | ( n1371 & n1378 ) | ( n1377 & n1378 ) ;
  assign n1380 = x2 & n1379 ;
  assign n1381 = x2 & ~n1380 ;
  assign n1382 = ( n1379 & ~n1380 ) | ( n1379 & n1381 ) | ( ~n1380 & n1381 ) ;
  assign n1383 = n1361 & n1382 ;
  assign n1384 = n1361 & ~n1383 ;
  assign n1385 = ~n1361 & n1382 ;
  assign n1386 = n1384 | n1385 ;
  assign n1387 = n1268 | n1273 ;
  assign n1388 = n1386 & n1387 ;
  assign n1389 = n1386 | n1387 ;
  assign n1390 = ~n1388 & n1389 ;
  assign n1391 = x71 & n771 ;
  assign n1392 = x70 & n766 ;
  assign n1393 = x69 & ~n765 ;
  assign n1394 = n905 & n1393 ;
  assign n1395 = n1392 | n1394 ;
  assign n1396 = n1391 | n1395 ;
  assign n1397 = n774 | n1396 ;
  assign n1398 = ( n376 & n1396 ) | ( n376 & n1397 ) | ( n1396 & n1397 ) ;
  assign n1399 = x14 & ~n1398 ;
  assign n1400 = ~x14 & n1398 ;
  assign n1401 = n1399 | n1400 ;
  assign n1402 = n229 & n1074 ;
  assign n1403 = x68 & n1071 ;
  assign n1404 = x67 & n1066 ;
  assign n1405 = x66 & ~n1065 ;
  assign n1406 = n1189 & n1405 ;
  assign n1407 = n1404 | n1406 ;
  assign n1408 = n1403 | n1407 ;
  assign n1409 = n1402 | n1408 ;
  assign n1410 = x17 | n1409 ;
  assign n1411 = ~x17 & n1410 ;
  assign n1412 = ( ~n1409 & n1410 ) | ( ~n1409 & n1411 ) | ( n1410 & n1411 ) ;
  assign n1413 = ~x18 & x19 ;
  assign n1414 = x18 & ~x19 ;
  assign n1415 = n1413 | n1414 ;
  assign n1416 = ~n1290 & n1415 ;
  assign n1417 = x64 & n1416 ;
  assign n1418 = ~x19 & x20 ;
  assign n1419 = x19 & ~x20 ;
  assign n1420 = n1418 | n1419 ;
  assign n1421 = n1290 & ~n1420 ;
  assign n1422 = x65 & n1421 ;
  assign n1423 = n1417 | n1422 ;
  assign n1424 = n1290 & n1420 ;
  assign n1425 = n142 & n1424 ;
  assign n1426 = n1423 | n1425 ;
  assign n1427 = x20 | n1426 ;
  assign n1428 = ~x20 & n1427 ;
  assign n1429 = ( ~n1426 & n1427 ) | ( ~n1426 & n1428 ) | ( n1427 & n1428 ) ;
  assign n1430 = x20 & ~n1291 ;
  assign n1431 = n1429 & n1430 ;
  assign n1432 = n1429 | n1430 ;
  assign n1433 = ~n1431 & n1432 ;
  assign n1434 = ( n1303 & n1412 ) | ( n1303 & n1433 ) | ( n1412 & n1433 ) ;
  assign n1435 = ( n1303 & n1433 ) | ( n1303 & ~n1434 ) | ( n1433 & ~n1434 ) ;
  assign n1436 = ( n1412 & ~n1434 ) | ( n1412 & n1435 ) | ( ~n1434 & n1435 ) ;
  assign n1437 = n1401 & n1436 ;
  assign n1438 = n1401 | n1436 ;
  assign n1439 = ~n1437 & n1438 ;
  assign n1440 = ( n1203 & n1287 ) | ( n1203 & n1305 ) | ( n1287 & n1305 ) ;
  assign n1441 = n1439 | n1440 ;
  assign n1442 = n1439 & n1440 ;
  assign n1443 = n1441 & ~n1442 ;
  assign n1444 = x74 & n528 ;
  assign n1445 = x73 & n523 ;
  assign n1446 = x72 & ~n522 ;
  assign n1447 = n635 & n1446 ;
  assign n1448 = n1445 | n1447 ;
  assign n1449 = n1444 | n1448 ;
  assign n1450 = n531 | n1449 ;
  assign n1451 = ( n587 & n1449 ) | ( n587 & n1450 ) | ( n1449 & n1450 ) ;
  assign n1452 = x11 & n1451 ;
  assign n1453 = x11 & ~n1452 ;
  assign n1454 = ( n1451 & ~n1452 ) | ( n1451 & n1453 ) | ( ~n1452 & n1453 ) ;
  assign n1455 = n1443 & n1454 ;
  assign n1456 = n1443 & ~n1455 ;
  assign n1457 = ~n1443 & n1454 ;
  assign n1458 = n1456 | n1457 ;
  assign n1459 = n1320 | n1323 ;
  assign n1460 = n1458 | n1459 ;
  assign n1461 = n1458 & n1459 ;
  assign n1462 = n1460 & ~n1461 ;
  assign n1463 = x77 & n337 ;
  assign n1464 = x76 & n332 ;
  assign n1465 = x75 & ~n331 ;
  assign n1466 = n396 & n1465 ;
  assign n1467 = n1464 | n1466 ;
  assign n1468 = n1463 | n1467 ;
  assign n1469 = n340 | n1468 ;
  assign n1470 = ( n846 & n1468 ) | ( n846 & n1469 ) | ( n1468 & n1469 ) ;
  assign n1471 = x8 & n1470 ;
  assign n1472 = x8 & ~n1471 ;
  assign n1473 = ( n1470 & ~n1471 ) | ( n1470 & n1472 ) | ( ~n1471 & n1472 ) ;
  assign n1474 = n1462 | n1473 ;
  assign n1475 = n1462 & n1473 ;
  assign n1476 = n1474 & ~n1475 ;
  assign n1477 = n1338 | n1341 ;
  assign n1478 = n1476 & n1477 ;
  assign n1479 = n1476 | n1477 ;
  assign n1480 = ~n1478 & n1479 ;
  assign n1481 = x80 & n206 ;
  assign n1482 = x79 & n201 ;
  assign n1483 = x78 & ~n200 ;
  assign n1484 = n243 & n1483 ;
  assign n1485 = n1482 | n1484 ;
  assign n1486 = n1481 | n1485 ;
  assign n1487 = n209 | n1486 ;
  assign n1488 = ( n1147 & n1486 ) | ( n1147 & n1487 ) | ( n1486 & n1487 ) ;
  assign n1489 = x5 & n1488 ;
  assign n1490 = x5 & ~n1489 ;
  assign n1491 = ( n1488 & ~n1489 ) | ( n1488 & n1490 ) | ( ~n1489 & n1490 ) ;
  assign n1492 = n1480 & n1491 ;
  assign n1493 = n1480 & ~n1492 ;
  assign n1494 = ~n1480 & n1491 ;
  assign n1495 = n1493 | n1494 ;
  assign n1496 = n1355 | n1359 ;
  assign n1497 = n1495 | n1496 ;
  assign n1498 = n1495 & n1496 ;
  assign n1499 = n1497 & ~n1498 ;
  assign n1500 = x82 | x83 ;
  assign n1501 = x82 & x83 ;
  assign n1502 = n1500 & ~n1501 ;
  assign n1503 = n1363 | n1366 ;
  assign n1504 = n1502 & n1503 ;
  assign n1505 = n1363 | n1367 ;
  assign n1506 = n1502 & n1505 ;
  assign n1507 = ( n1145 & n1504 ) | ( n1145 & n1506 ) | ( n1504 & n1506 ) ;
  assign n1508 = ( n1145 & n1503 ) | ( n1145 & n1505 ) | ( n1503 & n1505 ) ;
  assign n1509 = n1502 | n1508 ;
  assign n1510 = ~n1507 & n1509 ;
  assign n1511 = x82 & n131 ;
  assign n1512 = x81 & ~n156 ;
  assign n1513 = ( n135 & n1511 ) | ( n135 & n1512 ) | ( n1511 & n1512 ) ;
  assign n1514 = x0 & x83 ;
  assign n1515 = ( ~n135 & n1511 ) | ( ~n135 & n1514 ) | ( n1511 & n1514 ) ;
  assign n1516 = n1513 | n1515 ;
  assign n1517 = n139 | n1516 ;
  assign n1518 = ( n1510 & n1516 ) | ( n1510 & n1517 ) | ( n1516 & n1517 ) ;
  assign n1519 = x2 & n1518 ;
  assign n1520 = x2 & ~n1519 ;
  assign n1521 = ( n1518 & ~n1519 ) | ( n1518 & n1520 ) | ( ~n1519 & n1520 ) ;
  assign n1522 = n1499 & n1521 ;
  assign n1523 = n1499 & ~n1522 ;
  assign n1524 = ~n1499 & n1521 ;
  assign n1525 = n1523 | n1524 ;
  assign n1526 = n1383 | n1388 ;
  assign n1527 = n1525 & n1526 ;
  assign n1528 = n1525 | n1526 ;
  assign n1529 = ~n1527 & n1528 ;
  assign n1530 = n1522 | n1527 ;
  assign n1531 = x83 | x84 ;
  assign n1532 = x83 & x84 ;
  assign n1533 = n1531 & ~n1532 ;
  assign n1534 = n1501 | n1507 ;
  assign n1535 = n1533 & n1534 ;
  assign n1536 = n1533 | n1534 ;
  assign n1537 = ~n1535 & n1536 ;
  assign n1538 = x83 & n131 ;
  assign n1539 = x82 & ~n156 ;
  assign n1540 = ( n135 & n1538 ) | ( n135 & n1539 ) | ( n1538 & n1539 ) ;
  assign n1541 = x0 & x84 ;
  assign n1542 = ( ~n135 & n1538 ) | ( ~n135 & n1541 ) | ( n1538 & n1541 ) ;
  assign n1543 = n1540 | n1542 ;
  assign n1544 = n139 | n1543 ;
  assign n1545 = ( n1537 & n1543 ) | ( n1537 & n1544 ) | ( n1543 & n1544 ) ;
  assign n1546 = x2 & n1545 ;
  assign n1547 = x2 & ~n1546 ;
  assign n1548 = ( n1545 & ~n1546 ) | ( n1545 & n1547 ) | ( ~n1546 & n1547 ) ;
  assign n1549 = x81 & n206 ;
  assign n1550 = x80 & n201 ;
  assign n1551 = x79 & ~n200 ;
  assign n1552 = n243 & n1551 ;
  assign n1553 = n1550 | n1552 ;
  assign n1554 = n1549 | n1553 ;
  assign n1555 = n209 | n1554 ;
  assign n1556 = ( n1256 & n1554 ) | ( n1256 & n1555 ) | ( n1554 & n1555 ) ;
  assign n1557 = x5 & n1556 ;
  assign n1558 = x5 & ~n1557 ;
  assign n1559 = ( n1556 & ~n1557 ) | ( n1556 & n1558 ) | ( ~n1557 & n1558 ) ;
  assign n1560 = x72 & n771 ;
  assign n1561 = x71 & n766 ;
  assign n1562 = x70 & ~n765 ;
  assign n1563 = n905 & n1562 ;
  assign n1564 = n1561 | n1563 ;
  assign n1565 = n1560 | n1564 ;
  assign n1566 = ( n435 & n774 ) | ( n435 & n1565 ) | ( n774 & n1565 ) ;
  assign n1567 = ( x14 & ~n1565 ) | ( x14 & n1566 ) | ( ~n1565 & n1566 ) ;
  assign n1568 = ~n1566 & n1567 ;
  assign n1569 = n1565 | n1567 ;
  assign n1570 = ( ~x14 & n1568 ) | ( ~x14 & n1569 ) | ( n1568 & n1569 ) ;
  assign n1571 = n264 & n1074 ;
  assign n1572 = x69 & n1071 ;
  assign n1573 = x68 & n1066 ;
  assign n1574 = x67 & ~n1065 ;
  assign n1575 = n1189 & n1574 ;
  assign n1576 = n1573 | n1575 ;
  assign n1577 = n1572 | n1576 ;
  assign n1578 = n1571 | n1577 ;
  assign n1579 = x17 | n1578 ;
  assign n1580 = ~x17 & n1579 ;
  assign n1581 = ( ~n1578 & n1579 ) | ( ~n1578 & n1580 ) | ( n1579 & n1580 ) ;
  assign n1582 = x66 & n1421 ;
  assign n1583 = x65 & n1416 ;
  assign n1584 = ~n1290 & n1420 ;
  assign n1585 = x64 & ~n1415 ;
  assign n1586 = n1584 & n1585 ;
  assign n1587 = n1583 | n1586 ;
  assign n1588 = n1582 | n1587 ;
  assign n1589 = n153 & n1424 ;
  assign n1590 = n1588 | n1589 ;
  assign n1591 = x20 | n1590 ;
  assign n1592 = ~x20 & n1591 ;
  assign n1593 = ( ~n1590 & n1591 ) | ( ~n1590 & n1592 ) | ( n1591 & n1592 ) ;
  assign n1594 = n1431 | n1593 ;
  assign n1595 = n1431 & n1593 ;
  assign n1596 = n1594 & ~n1595 ;
  assign n1597 = ( n1434 & n1581 ) | ( n1434 & n1596 ) | ( n1581 & n1596 ) ;
  assign n1598 = ( n1434 & n1596 ) | ( n1434 & ~n1597 ) | ( n1596 & ~n1597 ) ;
  assign n1599 = ( n1581 & ~n1597 ) | ( n1581 & n1598 ) | ( ~n1597 & n1598 ) ;
  assign n1600 = n1570 | n1599 ;
  assign n1601 = n1570 & n1599 ;
  assign n1602 = n1600 & ~n1601 ;
  assign n1603 = n1437 | n1442 ;
  assign n1604 = n1602 & n1603 ;
  assign n1605 = n1602 | n1603 ;
  assign n1606 = ~n1604 & n1605 ;
  assign n1607 = x75 & n528 ;
  assign n1608 = x74 & n523 ;
  assign n1609 = x73 & ~n522 ;
  assign n1610 = n635 & n1609 ;
  assign n1611 = n1608 | n1610 ;
  assign n1612 = n1607 | n1611 ;
  assign n1613 = n531 | n1612 ;
  assign n1614 = ( n609 & n1612 ) | ( n609 & n1613 ) | ( n1612 & n1613 ) ;
  assign n1615 = x11 & n1614 ;
  assign n1616 = x11 & ~n1615 ;
  assign n1617 = ( n1614 & ~n1615 ) | ( n1614 & n1616 ) | ( ~n1615 & n1616 ) ;
  assign n1618 = n1606 | n1617 ;
  assign n1619 = n1606 & n1617 ;
  assign n1620 = n1618 & ~n1619 ;
  assign n1621 = n1455 | n1461 ;
  assign n1622 = n1620 & n1621 ;
  assign n1623 = n1620 | n1621 ;
  assign n1624 = ~n1622 & n1623 ;
  assign n1625 = x78 & n337 ;
  assign n1626 = x77 & n332 ;
  assign n1627 = x76 & ~n331 ;
  assign n1628 = n396 & n1627 ;
  assign n1629 = n1626 | n1628 ;
  assign n1630 = n1625 | n1629 ;
  assign n1631 = n340 | n1630 ;
  assign n1632 = ( n868 & n1630 ) | ( n868 & n1631 ) | ( n1630 & n1631 ) ;
  assign n1633 = x8 & n1632 ;
  assign n1634 = x8 & ~n1633 ;
  assign n1635 = ( n1632 & ~n1633 ) | ( n1632 & n1634 ) | ( ~n1633 & n1634 ) ;
  assign n1636 = n1624 & n1635 ;
  assign n1637 = n1624 & ~n1636 ;
  assign n1638 = ~n1624 & n1635 ;
  assign n1639 = n1637 | n1638 ;
  assign n1640 = n1475 | n1478 ;
  assign n1641 = n1639 & n1640 ;
  assign n1642 = n1639 | n1640 ;
  assign n1643 = ~n1641 & n1642 ;
  assign n1644 = n1492 | n1498 ;
  assign n1645 = ( n1559 & n1643 ) | ( n1559 & n1644 ) | ( n1643 & n1644 ) ;
  assign n1646 = ( n1643 & n1644 ) | ( n1643 & ~n1645 ) | ( n1644 & ~n1645 ) ;
  assign n1647 = ( n1559 & ~n1645 ) | ( n1559 & n1646 ) | ( ~n1645 & n1646 ) ;
  assign n1648 = n1548 & n1647 ;
  assign n1649 = n1548 | n1647 ;
  assign n1650 = ~n1648 & n1649 ;
  assign n1651 = n1530 & n1650 ;
  assign n1652 = n1530 | n1650 ;
  assign n1653 = ~n1651 & n1652 ;
  assign n1654 = n1601 | n1604 ;
  assign n1655 = x70 & n1071 ;
  assign n1656 = x69 & n1066 ;
  assign n1657 = x68 & ~n1065 ;
  assign n1658 = n1189 & n1657 ;
  assign n1659 = n1656 | n1658 ;
  assign n1660 = n1655 | n1659 ;
  assign n1661 = n1074 | n1660 ;
  assign n1662 = ( n310 & n1660 ) | ( n310 & n1661 ) | ( n1660 & n1661 ) ;
  assign n1663 = x17 & ~n1662 ;
  assign n1664 = ~x17 & n1662 ;
  assign n1665 = n1663 | n1664 ;
  assign n1666 = x20 & ~x21 ;
  assign n1667 = ~x20 & x21 ;
  assign n1668 = n1666 | n1667 ;
  assign n1669 = x64 & n1668 ;
  assign n1670 = x67 & n1421 ;
  assign n1671 = x66 & n1416 ;
  assign n1672 = x65 & ~n1415 ;
  assign n1673 = n1584 & n1672 ;
  assign n1674 = n1671 | n1673 ;
  assign n1675 = n1670 | n1674 ;
  assign n1676 = n180 & n1424 ;
  assign n1677 = n1675 | n1676 ;
  assign n1678 = x20 & ~n1677 ;
  assign n1679 = ~x20 & n1677 ;
  assign n1680 = n1678 | n1679 ;
  assign n1681 = ( n1595 & n1669 ) | ( n1595 & n1680 ) | ( n1669 & n1680 ) ;
  assign n1682 = ( n1595 & n1680 ) | ( n1595 & ~n1681 ) | ( n1680 & ~n1681 ) ;
  assign n1683 = ( n1669 & ~n1681 ) | ( n1669 & n1682 ) | ( ~n1681 & n1682 ) ;
  assign n1684 = ( n1597 & n1665 ) | ( n1597 & ~n1683 ) | ( n1665 & ~n1683 ) ;
  assign n1685 = ( ~n1597 & n1683 ) | ( ~n1597 & n1684 ) | ( n1683 & n1684 ) ;
  assign n1686 = ( ~n1665 & n1684 ) | ( ~n1665 & n1685 ) | ( n1684 & n1685 ) ;
  assign n1687 = x73 & n771 ;
  assign n1688 = x72 & n766 ;
  assign n1689 = x71 & ~n765 ;
  assign n1690 = n905 & n1689 ;
  assign n1691 = n1688 | n1690 ;
  assign n1692 = n1687 | n1691 ;
  assign n1693 = n774 | n1692 ;
  assign n1694 = ( n499 & n1692 ) | ( n499 & n1693 ) | ( n1692 & n1693 ) ;
  assign n1695 = x14 & n1694 ;
  assign n1696 = x14 | n1694 ;
  assign n1697 = ~n1695 & n1696 ;
  assign n1698 = n1686 & n1697 ;
  assign n1699 = n1686 | n1697 ;
  assign n1700 = ~n1698 & n1699 ;
  assign n1701 = n1654 & n1700 ;
  assign n1702 = n1654 | n1700 ;
  assign n1703 = ~n1701 & n1702 ;
  assign n1704 = x76 & n528 ;
  assign n1705 = x75 & n523 ;
  assign n1706 = x74 & ~n522 ;
  assign n1707 = n635 & n1706 ;
  assign n1708 = n1705 | n1707 ;
  assign n1709 = n1704 | n1708 ;
  assign n1710 = n531 | n1709 ;
  assign n1711 = ( n740 & n1709 ) | ( n740 & n1710 ) | ( n1709 & n1710 ) ;
  assign n1712 = x11 & n1711 ;
  assign n1713 = x11 & ~n1712 ;
  assign n1714 = ( n1711 & ~n1712 ) | ( n1711 & n1713 ) | ( ~n1712 & n1713 ) ;
  assign n1715 = n1703 | n1714 ;
  assign n1716 = n1703 & n1714 ;
  assign n1717 = n1715 & ~n1716 ;
  assign n1718 = n1619 | n1622 ;
  assign n1719 = n1717 & n1718 ;
  assign n1720 = n1717 | n1718 ;
  assign n1721 = ~n1719 & n1720 ;
  assign n1722 = x79 & n337 ;
  assign n1723 = x78 & n332 ;
  assign n1724 = x77 & ~n331 ;
  assign n1725 = n396 & n1724 ;
  assign n1726 = n1723 | n1725 ;
  assign n1727 = n1722 | n1726 ;
  assign n1728 = n340 | n1727 ;
  assign n1729 = ( n961 & n1727 ) | ( n961 & n1728 ) | ( n1727 & n1728 ) ;
  assign n1730 = x8 & n1729 ;
  assign n1731 = x8 & ~n1730 ;
  assign n1732 = ( n1729 & ~n1730 ) | ( n1729 & n1731 ) | ( ~n1730 & n1731 ) ;
  assign n1733 = n1721 & n1732 ;
  assign n1734 = n1721 | n1732 ;
  assign n1735 = ~n1733 & n1734 ;
  assign n1736 = n1636 | n1735 ;
  assign n1737 = n1641 | n1736 ;
  assign n1738 = ( n1636 & n1641 ) | ( n1636 & n1735 ) | ( n1641 & n1735 ) ;
  assign n1739 = n1737 & ~n1738 ;
  assign n1740 = x82 & n206 ;
  assign n1741 = x81 & n201 ;
  assign n1742 = x80 & ~n200 ;
  assign n1743 = n243 & n1742 ;
  assign n1744 = n1741 | n1743 ;
  assign n1745 = n1740 | n1744 ;
  assign n1746 = n209 | n1745 ;
  assign n1747 = ( n1371 & n1745 ) | ( n1371 & n1746 ) | ( n1745 & n1746 ) ;
  assign n1748 = x5 & n1747 ;
  assign n1749 = x5 & ~n1748 ;
  assign n1750 = ( n1747 & ~n1748 ) | ( n1747 & n1749 ) | ( ~n1748 & n1749 ) ;
  assign n1751 = n1739 & n1750 ;
  assign n1752 = n1739 & ~n1751 ;
  assign n1753 = ~n1739 & n1750 ;
  assign n1754 = n1752 | n1753 ;
  assign n1755 = n1645 | n1754 ;
  assign n1756 = n1645 & n1754 ;
  assign n1757 = n1755 & ~n1756 ;
  assign n1758 = x84 | x85 ;
  assign n1759 = x84 & x85 ;
  assign n1760 = n1758 & ~n1759 ;
  assign n1761 = n1532 & n1760 ;
  assign n1762 = ( n1535 & n1760 ) | ( n1535 & n1761 ) | ( n1760 & n1761 ) ;
  assign n1763 = n1532 | n1760 ;
  assign n1764 = n1535 | n1763 ;
  assign n1765 = ~n1762 & n1764 ;
  assign n1766 = x84 & n131 ;
  assign n1767 = x83 & ~n156 ;
  assign n1768 = ( n135 & n1766 ) | ( n135 & n1767 ) | ( n1766 & n1767 ) ;
  assign n1769 = x0 & x85 ;
  assign n1770 = ( ~n135 & n1766 ) | ( ~n135 & n1769 ) | ( n1766 & n1769 ) ;
  assign n1771 = n1768 | n1770 ;
  assign n1772 = n139 | n1771 ;
  assign n1773 = ( n1765 & n1771 ) | ( n1765 & n1772 ) | ( n1771 & n1772 ) ;
  assign n1774 = x2 & n1773 ;
  assign n1775 = x2 & ~n1774 ;
  assign n1776 = ( n1773 & ~n1774 ) | ( n1773 & n1775 ) | ( ~n1774 & n1775 ) ;
  assign n1777 = n1757 & n1776 ;
  assign n1778 = n1757 & ~n1777 ;
  assign n1779 = ~n1757 & n1776 ;
  assign n1780 = n1778 | n1779 ;
  assign n1781 = n1648 | n1651 ;
  assign n1782 = n1780 & n1781 ;
  assign n1783 = n1780 | n1781 ;
  assign n1784 = ~n1782 & n1783 ;
  assign n1785 = n1733 | n1738 ;
  assign n1786 = n1716 | n1719 ;
  assign n1787 = x71 & n1071 ;
  assign n1788 = x70 & n1066 ;
  assign n1789 = x69 & ~n1065 ;
  assign n1790 = n1189 & n1789 ;
  assign n1791 = n1788 | n1790 ;
  assign n1792 = n1787 | n1791 ;
  assign n1793 = n1074 | n1792 ;
  assign n1794 = ( n376 & n1792 ) | ( n376 & n1793 ) | ( n1792 & n1793 ) ;
  assign n1795 = x17 & ~n1794 ;
  assign n1796 = ~x17 & n1794 ;
  assign n1797 = n1795 | n1796 ;
  assign n1798 = n229 & n1424 ;
  assign n1799 = x68 & n1421 ;
  assign n1800 = x67 & n1416 ;
  assign n1801 = x66 & ~n1415 ;
  assign n1802 = n1584 & n1801 ;
  assign n1803 = n1800 | n1802 ;
  assign n1804 = n1799 | n1803 ;
  assign n1805 = n1798 | n1804 ;
  assign n1806 = x20 | n1805 ;
  assign n1807 = ~x20 & n1806 ;
  assign n1808 = ( ~n1805 & n1806 ) | ( ~n1805 & n1807 ) | ( n1806 & n1807 ) ;
  assign n1809 = ~x21 & x22 ;
  assign n1810 = x21 & ~x22 ;
  assign n1811 = n1809 | n1810 ;
  assign n1812 = ~n1668 & n1811 ;
  assign n1813 = x64 & n1812 ;
  assign n1814 = ~x22 & x23 ;
  assign n1815 = x22 & ~x23 ;
  assign n1816 = n1814 | n1815 ;
  assign n1817 = n1668 & ~n1816 ;
  assign n1818 = x65 & n1817 ;
  assign n1819 = n1813 | n1818 ;
  assign n1820 = n1668 & n1816 ;
  assign n1821 = n142 & n1820 ;
  assign n1822 = n1819 | n1821 ;
  assign n1823 = x23 | n1822 ;
  assign n1824 = ~x23 & n1823 ;
  assign n1825 = ( ~n1822 & n1823 ) | ( ~n1822 & n1824 ) | ( n1823 & n1824 ) ;
  assign n1826 = x23 & ~n1669 ;
  assign n1827 = n1825 & n1826 ;
  assign n1828 = n1825 | n1826 ;
  assign n1829 = ~n1827 & n1828 ;
  assign n1830 = ( n1681 & n1808 ) | ( n1681 & n1829 ) | ( n1808 & n1829 ) ;
  assign n1831 = ( n1681 & n1829 ) | ( n1681 & ~n1830 ) | ( n1829 & ~n1830 ) ;
  assign n1832 = ( n1808 & ~n1830 ) | ( n1808 & n1831 ) | ( ~n1830 & n1831 ) ;
  assign n1833 = n1797 & n1832 ;
  assign n1834 = n1797 | n1832 ;
  assign n1835 = ~n1833 & n1834 ;
  assign n1836 = ( n1597 & n1665 ) | ( n1597 & n1683 ) | ( n1665 & n1683 ) ;
  assign n1837 = n1835 | n1836 ;
  assign n1838 = n1835 & n1836 ;
  assign n1839 = n1837 & ~n1838 ;
  assign n1840 = x74 & n771 ;
  assign n1841 = x73 & n766 ;
  assign n1842 = x72 & ~n765 ;
  assign n1843 = n905 & n1842 ;
  assign n1844 = n1841 | n1843 ;
  assign n1845 = n1840 | n1844 ;
  assign n1846 = n774 | n1845 ;
  assign n1847 = ( n587 & n1845 ) | ( n587 & n1846 ) | ( n1845 & n1846 ) ;
  assign n1848 = x14 & n1847 ;
  assign n1849 = x14 & ~n1848 ;
  assign n1850 = ( n1847 & ~n1848 ) | ( n1847 & n1849 ) | ( ~n1848 & n1849 ) ;
  assign n1851 = n1839 & n1850 ;
  assign n1852 = n1839 & ~n1851 ;
  assign n1853 = ~n1839 & n1850 ;
  assign n1854 = n1852 | n1853 ;
  assign n1855 = n1698 | n1701 ;
  assign n1856 = n1854 | n1855 ;
  assign n1857 = n1854 & n1855 ;
  assign n1858 = n1856 & ~n1857 ;
  assign n1859 = x77 & n528 ;
  assign n1860 = x76 & n523 ;
  assign n1861 = x75 & ~n522 ;
  assign n1862 = n635 & n1861 ;
  assign n1863 = n1860 | n1862 ;
  assign n1864 = n1859 | n1863 ;
  assign n1865 = n531 | n1864 ;
  assign n1866 = ( n846 & n1864 ) | ( n846 & n1865 ) | ( n1864 & n1865 ) ;
  assign n1867 = x11 & n1866 ;
  assign n1868 = x11 & ~n1867 ;
  assign n1869 = ( n1866 & ~n1867 ) | ( n1866 & n1868 ) | ( ~n1867 & n1868 ) ;
  assign n1870 = n1858 | n1869 ;
  assign n1871 = n1858 & n1869 ;
  assign n1872 = n1870 & ~n1871 ;
  assign n1873 = n1786 & n1872 ;
  assign n1874 = n1786 | n1872 ;
  assign n1875 = ~n1873 & n1874 ;
  assign n1876 = x80 & n337 ;
  assign n1877 = x79 & n332 ;
  assign n1878 = x78 & ~n331 ;
  assign n1879 = n396 & n1878 ;
  assign n1880 = n1877 | n1879 ;
  assign n1881 = n1876 | n1880 ;
  assign n1882 = n340 | n1881 ;
  assign n1883 = ( n1147 & n1881 ) | ( n1147 & n1882 ) | ( n1881 & n1882 ) ;
  assign n1884 = x8 & n1883 ;
  assign n1885 = x8 & ~n1884 ;
  assign n1886 = ( n1883 & ~n1884 ) | ( n1883 & n1885 ) | ( ~n1884 & n1885 ) ;
  assign n1887 = n1875 & n1886 ;
  assign n1888 = n1875 | n1886 ;
  assign n1889 = ~n1887 & n1888 ;
  assign n1890 = n1785 & n1889 ;
  assign n1891 = n1785 | n1889 ;
  assign n1892 = ~n1890 & n1891 ;
  assign n1893 = x83 & n206 ;
  assign n1894 = x82 & n201 ;
  assign n1895 = x81 & ~n200 ;
  assign n1896 = n243 & n1895 ;
  assign n1897 = n1894 | n1896 ;
  assign n1898 = n1893 | n1897 ;
  assign n1899 = n209 | n1898 ;
  assign n1900 = ( n1510 & n1898 ) | ( n1510 & n1899 ) | ( n1898 & n1899 ) ;
  assign n1901 = x5 & n1900 ;
  assign n1902 = x5 & ~n1901 ;
  assign n1903 = ( n1900 & ~n1901 ) | ( n1900 & n1902 ) | ( ~n1901 & n1902 ) ;
  assign n1904 = n1892 & n1903 ;
  assign n1905 = n1892 & ~n1904 ;
  assign n1906 = ~n1892 & n1903 ;
  assign n1907 = n1905 | n1906 ;
  assign n1908 = n1751 | n1756 ;
  assign n1909 = n1907 | n1908 ;
  assign n1910 = n1907 & n1908 ;
  assign n1911 = n1909 & ~n1910 ;
  assign n1912 = x85 | x86 ;
  assign n1913 = x85 & x86 ;
  assign n1914 = n1912 & ~n1913 ;
  assign n1915 = n1759 | n1761 ;
  assign n1916 = n1914 & n1915 ;
  assign n1917 = n1758 & n1914 ;
  assign n1918 = ( n1535 & n1916 ) | ( n1535 & n1917 ) | ( n1916 & n1917 ) ;
  assign n1919 = ( n1535 & n1758 ) | ( n1535 & n1915 ) | ( n1758 & n1915 ) ;
  assign n1920 = n1914 | n1919 ;
  assign n1921 = ~n1918 & n1920 ;
  assign n1922 = x85 & n131 ;
  assign n1923 = x84 & ~n156 ;
  assign n1924 = ( n135 & n1922 ) | ( n135 & n1923 ) | ( n1922 & n1923 ) ;
  assign n1925 = x0 & x86 ;
  assign n1926 = ( ~n135 & n1922 ) | ( ~n135 & n1925 ) | ( n1922 & n1925 ) ;
  assign n1927 = n1924 | n1926 ;
  assign n1928 = n139 | n1927 ;
  assign n1929 = ( n1921 & n1927 ) | ( n1921 & n1928 ) | ( n1927 & n1928 ) ;
  assign n1930 = x2 & n1929 ;
  assign n1931 = x2 & ~n1930 ;
  assign n1932 = ( n1929 & ~n1930 ) | ( n1929 & n1931 ) | ( ~n1930 & n1931 ) ;
  assign n1933 = n1911 | n1932 ;
  assign n1934 = n1911 & n1932 ;
  assign n1935 = n1933 & ~n1934 ;
  assign n1936 = n1777 | n1782 ;
  assign n1937 = n1935 & n1936 ;
  assign n1938 = n1935 | n1936 ;
  assign n1939 = ~n1937 & n1938 ;
  assign n1940 = n1904 | n1910 ;
  assign n1941 = x84 & n206 ;
  assign n1942 = x83 & n201 ;
  assign n1943 = x82 & ~n200 ;
  assign n1944 = n243 & n1943 ;
  assign n1945 = n1942 | n1944 ;
  assign n1946 = n1941 | n1945 ;
  assign n1947 = n209 | n1946 ;
  assign n1948 = ( n1537 & n1946 ) | ( n1537 & n1947 ) | ( n1946 & n1947 ) ;
  assign n1949 = x5 & n1948 ;
  assign n1950 = x5 & ~n1949 ;
  assign n1951 = ( n1948 & ~n1949 ) | ( n1948 & n1950 ) | ( ~n1949 & n1950 ) ;
  assign n1952 = n1887 | n1890 ;
  assign n1953 = x72 & n1071 ;
  assign n1954 = x71 & n1066 ;
  assign n1955 = x70 & ~n1065 ;
  assign n1956 = n1189 & n1955 ;
  assign n1957 = n1954 | n1956 ;
  assign n1958 = n1953 | n1957 ;
  assign n1959 = ( n435 & n1074 ) | ( n435 & n1958 ) | ( n1074 & n1958 ) ;
  assign n1960 = ( x17 & ~n1958 ) | ( x17 & n1959 ) | ( ~n1958 & n1959 ) ;
  assign n1961 = ~n1959 & n1960 ;
  assign n1962 = n1958 | n1960 ;
  assign n1963 = ( ~x17 & n1961 ) | ( ~x17 & n1962 ) | ( n1961 & n1962 ) ;
  assign n1964 = n264 & n1424 ;
  assign n1965 = x69 & n1421 ;
  assign n1966 = x68 & n1416 ;
  assign n1967 = x67 & ~n1415 ;
  assign n1968 = n1584 & n1967 ;
  assign n1969 = n1966 | n1968 ;
  assign n1970 = n1965 | n1969 ;
  assign n1971 = n1964 | n1970 ;
  assign n1972 = x20 | n1971 ;
  assign n1973 = ~x20 & n1972 ;
  assign n1974 = ( ~n1971 & n1972 ) | ( ~n1971 & n1973 ) | ( n1972 & n1973 ) ;
  assign n1975 = x66 & n1817 ;
  assign n1976 = x65 & n1812 ;
  assign n1977 = ~n1668 & n1816 ;
  assign n1978 = x64 & ~n1811 ;
  assign n1979 = n1977 & n1978 ;
  assign n1980 = n1976 | n1979 ;
  assign n1981 = n1975 | n1980 ;
  assign n1982 = n153 & n1820 ;
  assign n1983 = n1981 | n1982 ;
  assign n1984 = x23 | n1983 ;
  assign n1985 = ~x23 & n1984 ;
  assign n1986 = ( ~n1983 & n1984 ) | ( ~n1983 & n1985 ) | ( n1984 & n1985 ) ;
  assign n1987 = n1827 | n1986 ;
  assign n1988 = n1827 & n1986 ;
  assign n1989 = n1987 & ~n1988 ;
  assign n1990 = ( n1830 & n1974 ) | ( n1830 & n1989 ) | ( n1974 & n1989 ) ;
  assign n1991 = ( n1830 & n1989 ) | ( n1830 & ~n1990 ) | ( n1989 & ~n1990 ) ;
  assign n1992 = ( n1974 & ~n1990 ) | ( n1974 & n1991 ) | ( ~n1990 & n1991 ) ;
  assign n1993 = n1963 | n1992 ;
  assign n1994 = n1963 & n1992 ;
  assign n1995 = n1993 & ~n1994 ;
  assign n1996 = n1833 | n1838 ;
  assign n1997 = n1995 & n1996 ;
  assign n1998 = n1995 | n1996 ;
  assign n1999 = ~n1997 & n1998 ;
  assign n2000 = x75 & n771 ;
  assign n2001 = x74 & n766 ;
  assign n2002 = x73 & ~n765 ;
  assign n2003 = n905 & n2002 ;
  assign n2004 = n2001 | n2003 ;
  assign n2005 = n2000 | n2004 ;
  assign n2006 = n774 | n2005 ;
  assign n2007 = ( n609 & n2005 ) | ( n609 & n2006 ) | ( n2005 & n2006 ) ;
  assign n2008 = x14 & n2007 ;
  assign n2009 = x14 & ~n2008 ;
  assign n2010 = ( n2007 & ~n2008 ) | ( n2007 & n2009 ) | ( ~n2008 & n2009 ) ;
  assign n2011 = n1999 | n2010 ;
  assign n2012 = n1999 & n2010 ;
  assign n2013 = n2011 & ~n2012 ;
  assign n2014 = n1851 | n1857 ;
  assign n2015 = n2013 & n2014 ;
  assign n2016 = n2013 | n2014 ;
  assign n2017 = ~n2015 & n2016 ;
  assign n2018 = x78 & n528 ;
  assign n2019 = x77 & n523 ;
  assign n2020 = x76 & ~n522 ;
  assign n2021 = n635 & n2020 ;
  assign n2022 = n2019 | n2021 ;
  assign n2023 = n2018 | n2022 ;
  assign n2024 = n531 | n2023 ;
  assign n2025 = ( n868 & n2023 ) | ( n868 & n2024 ) | ( n2023 & n2024 ) ;
  assign n2026 = x11 & n2025 ;
  assign n2027 = x11 & ~n2026 ;
  assign n2028 = ( n2025 & ~n2026 ) | ( n2025 & n2027 ) | ( ~n2026 & n2027 ) ;
  assign n2029 = n2017 & n2028 ;
  assign n2030 = n2017 & ~n2029 ;
  assign n2031 = ~n2017 & n2028 ;
  assign n2032 = n2030 | n2031 ;
  assign n2033 = n1871 | n1873 ;
  assign n2034 = n2032 & n2033 ;
  assign n2035 = n2032 | n2033 ;
  assign n2036 = ~n2034 & n2035 ;
  assign n2037 = x81 & n337 ;
  assign n2038 = x80 & n332 ;
  assign n2039 = x79 & ~n331 ;
  assign n2040 = n396 & n2039 ;
  assign n2041 = n2038 | n2040 ;
  assign n2042 = n2037 | n2041 ;
  assign n2043 = n340 | n2042 ;
  assign n2044 = ( n1256 & n2042 ) | ( n1256 & n2043 ) | ( n2042 & n2043 ) ;
  assign n2045 = x8 & n2044 ;
  assign n2046 = x8 & ~n2045 ;
  assign n2047 = ( n2044 & ~n2045 ) | ( n2044 & n2046 ) | ( ~n2045 & n2046 ) ;
  assign n2048 = ( n1952 & n2036 ) | ( n1952 & ~n2047 ) | ( n2036 & ~n2047 ) ;
  assign n2049 = ( ~n2036 & n2047 ) | ( ~n2036 & n2048 ) | ( n2047 & n2048 ) ;
  assign n2050 = ( ~n1952 & n2048 ) | ( ~n1952 & n2049 ) | ( n2048 & n2049 ) ;
  assign n2051 = n1951 & n2050 ;
  assign n2052 = n1951 | n2050 ;
  assign n2053 = ~n2051 & n2052 ;
  assign n2054 = n1940 | n2053 ;
  assign n2055 = n1940 & n2053 ;
  assign n2056 = n2054 & ~n2055 ;
  assign n2057 = x86 | x87 ;
  assign n2058 = x86 & x87 ;
  assign n2059 = n2057 & ~n2058 ;
  assign n2060 = n1913 | n1916 ;
  assign n2061 = n2059 & n2060 ;
  assign n2062 = n1913 | n1917 ;
  assign n2063 = n2059 & n2062 ;
  assign n2064 = ( n1535 & n2061 ) | ( n1535 & n2063 ) | ( n2061 & n2063 ) ;
  assign n2065 = ( n1535 & n2060 ) | ( n1535 & n2062 ) | ( n2060 & n2062 ) ;
  assign n2066 = n2059 | n2065 ;
  assign n2067 = ~n2064 & n2066 ;
  assign n2068 = x86 & n131 ;
  assign n2069 = x85 & ~n156 ;
  assign n2070 = ( n135 & n2068 ) | ( n135 & n2069 ) | ( n2068 & n2069 ) ;
  assign n2071 = x0 & x87 ;
  assign n2072 = ( ~n135 & n2068 ) | ( ~n135 & n2071 ) | ( n2068 & n2071 ) ;
  assign n2073 = n2070 | n2072 ;
  assign n2074 = n139 | n2073 ;
  assign n2075 = ( n2067 & n2073 ) | ( n2067 & n2074 ) | ( n2073 & n2074 ) ;
  assign n2076 = x2 & n2075 ;
  assign n2077 = x2 & ~n2076 ;
  assign n2078 = ( n2075 & ~n2076 ) | ( n2075 & n2077 ) | ( ~n2076 & n2077 ) ;
  assign n2079 = n2056 & n2078 ;
  assign n2080 = n2056 & ~n2079 ;
  assign n2081 = ~n2056 & n2078 ;
  assign n2082 = n2080 | n2081 ;
  assign n2083 = n1934 | n1937 ;
  assign n2084 = n2082 & n2083 ;
  assign n2085 = n2082 | n2083 ;
  assign n2086 = ~n2084 & n2085 ;
  assign n2087 = x87 | x88 ;
  assign n2088 = x87 & x88 ;
  assign n2089 = n2087 & ~n2088 ;
  assign n2090 = n2058 | n2061 ;
  assign n2091 = n2058 | n2063 ;
  assign n2092 = ( n1535 & n2090 ) | ( n1535 & n2091 ) | ( n2090 & n2091 ) ;
  assign n2093 = n2089 | n2092 ;
  assign n2094 = n2089 & n2092 ;
  assign n2095 = n2093 & ~n2094 ;
  assign n2096 = x87 & n131 ;
  assign n2097 = x86 & ~n156 ;
  assign n2098 = ( n135 & n2096 ) | ( n135 & n2097 ) | ( n2096 & n2097 ) ;
  assign n2099 = x0 & x88 ;
  assign n2100 = ( ~n135 & n2096 ) | ( ~n135 & n2099 ) | ( n2096 & n2099 ) ;
  assign n2101 = n2098 | n2100 ;
  assign n2102 = n139 | n2101 ;
  assign n2103 = ( n2095 & n2101 ) | ( n2095 & n2102 ) | ( n2101 & n2102 ) ;
  assign n2104 = x2 & n2103 ;
  assign n2105 = x2 & ~n2104 ;
  assign n2106 = ( n2103 & ~n2104 ) | ( n2103 & n2105 ) | ( ~n2104 & n2105 ) ;
  assign n2107 = x85 & n206 ;
  assign n2108 = x84 & n201 ;
  assign n2109 = x83 & ~n200 ;
  assign n2110 = n243 & n2109 ;
  assign n2111 = n2108 | n2110 ;
  assign n2112 = n2107 | n2111 ;
  assign n2113 = n209 | n2112 ;
  assign n2114 = ( n1765 & n2112 ) | ( n1765 & n2113 ) | ( n2112 & n2113 ) ;
  assign n2115 = x5 & n2114 ;
  assign n2116 = x5 & ~n2115 ;
  assign n2117 = ( n2114 & ~n2115 ) | ( n2114 & n2116 ) | ( ~n2115 & n2116 ) ;
  assign n2118 = n2051 | n2055 ;
  assign n2119 = n1994 | n1997 ;
  assign n2120 = x70 & n1421 ;
  assign n2121 = x69 & n1416 ;
  assign n2122 = x68 & ~n1415 ;
  assign n2123 = n1584 & n2122 ;
  assign n2124 = n2121 | n2123 ;
  assign n2125 = n2120 | n2124 ;
  assign n2126 = n1424 | n2125 ;
  assign n2127 = ( n310 & n2125 ) | ( n310 & n2126 ) | ( n2125 & n2126 ) ;
  assign n2128 = x20 & ~n2127 ;
  assign n2129 = ~x20 & n2127 ;
  assign n2130 = n2128 | n2129 ;
  assign n2131 = x23 & ~x24 ;
  assign n2132 = ~x23 & x24 ;
  assign n2133 = n2131 | n2132 ;
  assign n2134 = x64 & n2133 ;
  assign n2135 = x67 & n1817 ;
  assign n2136 = x66 & n1812 ;
  assign n2137 = x65 & ~n1811 ;
  assign n2138 = n1977 & n2137 ;
  assign n2139 = n2136 | n2138 ;
  assign n2140 = n2135 | n2139 ;
  assign n2141 = n180 & n1820 ;
  assign n2142 = n2140 | n2141 ;
  assign n2143 = x23 & ~n2142 ;
  assign n2144 = ~x23 & n2142 ;
  assign n2145 = n2143 | n2144 ;
  assign n2146 = ( n1988 & n2134 ) | ( n1988 & n2145 ) | ( n2134 & n2145 ) ;
  assign n2147 = ( n1988 & n2145 ) | ( n1988 & ~n2146 ) | ( n2145 & ~n2146 ) ;
  assign n2148 = ( n2134 & ~n2146 ) | ( n2134 & n2147 ) | ( ~n2146 & n2147 ) ;
  assign n2149 = ( n1990 & n2130 ) | ( n1990 & ~n2148 ) | ( n2130 & ~n2148 ) ;
  assign n2150 = ( ~n1990 & n2148 ) | ( ~n1990 & n2149 ) | ( n2148 & n2149 ) ;
  assign n2151 = ( ~n2130 & n2149 ) | ( ~n2130 & n2150 ) | ( n2149 & n2150 ) ;
  assign n2152 = x73 & n1071 ;
  assign n2153 = x72 & n1066 ;
  assign n2154 = x71 & ~n1065 ;
  assign n2155 = n1189 & n2154 ;
  assign n2156 = n2153 | n2155 ;
  assign n2157 = n2152 | n2156 ;
  assign n2158 = n1074 | n2157 ;
  assign n2159 = ( n499 & n2157 ) | ( n499 & n2158 ) | ( n2157 & n2158 ) ;
  assign n2160 = x17 & n2159 ;
  assign n2161 = x17 | n2159 ;
  assign n2162 = ~n2160 & n2161 ;
  assign n2163 = n2151 & n2162 ;
  assign n2164 = n2151 | n2162 ;
  assign n2165 = ~n2163 & n2164 ;
  assign n2166 = n2119 & n2165 ;
  assign n2167 = n2119 | n2165 ;
  assign n2168 = ~n2166 & n2167 ;
  assign n2169 = x76 & n771 ;
  assign n2170 = x75 & n766 ;
  assign n2171 = x74 & ~n765 ;
  assign n2172 = n905 & n2171 ;
  assign n2173 = n2170 | n2172 ;
  assign n2174 = n2169 | n2173 ;
  assign n2175 = n774 | n2174 ;
  assign n2176 = ( n740 & n2174 ) | ( n740 & n2175 ) | ( n2174 & n2175 ) ;
  assign n2177 = x14 & n2176 ;
  assign n2178 = x14 & ~n2177 ;
  assign n2179 = ( n2176 & ~n2177 ) | ( n2176 & n2178 ) | ( ~n2177 & n2178 ) ;
  assign n2180 = n2168 | n2179 ;
  assign n2181 = n2168 & n2179 ;
  assign n2182 = n2180 & ~n2181 ;
  assign n2183 = n2012 | n2015 ;
  assign n2184 = n2182 & n2183 ;
  assign n2185 = n2182 | n2183 ;
  assign n2186 = ~n2184 & n2185 ;
  assign n2187 = x79 & n528 ;
  assign n2188 = x78 & n523 ;
  assign n2189 = x77 & ~n522 ;
  assign n2190 = n635 & n2189 ;
  assign n2191 = n2188 | n2190 ;
  assign n2192 = n2187 | n2191 ;
  assign n2193 = n531 | n2192 ;
  assign n2194 = ( n961 & n2192 ) | ( n961 & n2193 ) | ( n2192 & n2193 ) ;
  assign n2195 = x11 & n2194 ;
  assign n2196 = x11 & ~n2195 ;
  assign n2197 = ( n2194 & ~n2195 ) | ( n2194 & n2196 ) | ( ~n2195 & n2196 ) ;
  assign n2198 = n2186 & n2197 ;
  assign n2199 = n2186 & ~n2198 ;
  assign n2200 = ~n2186 & n2197 ;
  assign n2201 = n2199 | n2200 ;
  assign n2202 = n2029 | n2034 ;
  assign n2203 = n2201 | n2202 ;
  assign n2204 = n2201 & n2202 ;
  assign n2205 = n2203 & ~n2204 ;
  assign n2206 = x82 & n337 ;
  assign n2207 = x81 & n332 ;
  assign n2208 = x80 & ~n331 ;
  assign n2209 = n396 & n2208 ;
  assign n2210 = n2207 | n2209 ;
  assign n2211 = n2206 | n2210 ;
  assign n2212 = n340 | n2211 ;
  assign n2213 = ( n1371 & n2211 ) | ( n1371 & n2212 ) | ( n2211 & n2212 ) ;
  assign n2214 = x8 & n2213 ;
  assign n2215 = x8 & ~n2214 ;
  assign n2216 = ( n2213 & ~n2214 ) | ( n2213 & n2215 ) | ( ~n2214 & n2215 ) ;
  assign n2217 = n2205 | n2216 ;
  assign n2218 = n2205 & n2216 ;
  assign n2219 = n2217 & ~n2218 ;
  assign n2220 = ( n1952 & n2036 ) | ( n1952 & n2047 ) | ( n2036 & n2047 ) ;
  assign n2221 = n2219 & n2220 ;
  assign n2222 = n2219 | n2220 ;
  assign n2223 = ~n2221 & n2222 ;
  assign n2224 = ( n2117 & n2118 ) | ( n2117 & ~n2223 ) | ( n2118 & ~n2223 ) ;
  assign n2225 = ( ~n2118 & n2223 ) | ( ~n2118 & n2224 ) | ( n2223 & n2224 ) ;
  assign n2226 = ( ~n2117 & n2224 ) | ( ~n2117 & n2225 ) | ( n2224 & n2225 ) ;
  assign n2227 = n2106 & n2226 ;
  assign n2228 = n2106 | n2226 ;
  assign n2229 = ~n2227 & n2228 ;
  assign n2230 = n2079 | n2084 ;
  assign n2231 = n2229 & n2230 ;
  assign n2232 = n2229 | n2230 ;
  assign n2233 = ~n2231 & n2232 ;
  assign n2234 = x88 & n131 ;
  assign n2235 = x87 & ~n156 ;
  assign n2236 = ( n135 & n2234 ) | ( n135 & n2235 ) | ( n2234 & n2235 ) ;
  assign n2237 = x0 & x89 ;
  assign n2238 = ( ~n135 & n2234 ) | ( ~n135 & n2237 ) | ( n2234 & n2237 ) ;
  assign n2239 = n2236 | n2238 ;
  assign n2240 = n139 | n2239 ;
  assign n2241 = n2088 | n2094 ;
  assign n2242 = ( x88 & ~x89 ) | ( x88 & n2241 ) | ( ~x89 & n2241 ) ;
  assign n2243 = ( ~x88 & x89 ) | ( ~x88 & n2242 ) | ( x89 & n2242 ) ;
  assign n2244 = ( ~n2241 & n2242 ) | ( ~n2241 & n2243 ) | ( n2242 & n2243 ) ;
  assign n2245 = ( n2239 & n2240 ) | ( n2239 & n2244 ) | ( n2240 & n2244 ) ;
  assign n2246 = x2 & n2245 ;
  assign n2247 = x2 & ~n2246 ;
  assign n2248 = ( n2245 & ~n2246 ) | ( n2245 & n2247 ) | ( ~n2246 & n2247 ) ;
  assign n2249 = ( n2117 & n2118 ) | ( n2117 & n2223 ) | ( n2118 & n2223 ) ;
  assign n2250 = x71 & n1421 ;
  assign n2251 = x70 & n1416 ;
  assign n2252 = x69 & ~n1415 ;
  assign n2253 = n1584 & n2252 ;
  assign n2254 = n2251 | n2253 ;
  assign n2255 = n2250 | n2254 ;
  assign n2256 = n1424 | n2255 ;
  assign n2257 = ( n376 & n2255 ) | ( n376 & n2256 ) | ( n2255 & n2256 ) ;
  assign n2258 = x20 & ~n2257 ;
  assign n2259 = ~x20 & n2257 ;
  assign n2260 = n2258 | n2259 ;
  assign n2261 = n229 & n1820 ;
  assign n2262 = x68 & n1817 ;
  assign n2263 = x67 & n1812 ;
  assign n2264 = x66 & ~n1811 ;
  assign n2265 = n1977 & n2264 ;
  assign n2266 = n2263 | n2265 ;
  assign n2267 = n2262 | n2266 ;
  assign n2268 = n2261 | n2267 ;
  assign n2269 = x23 | n2268 ;
  assign n2270 = ~x23 & n2269 ;
  assign n2271 = ( ~n2268 & n2269 ) | ( ~n2268 & n2270 ) | ( n2269 & n2270 ) ;
  assign n2272 = ~x24 & x25 ;
  assign n2273 = x24 & ~x25 ;
  assign n2274 = n2272 | n2273 ;
  assign n2275 = ~n2133 & n2274 ;
  assign n2276 = x64 & n2275 ;
  assign n2277 = ~x25 & x26 ;
  assign n2278 = x25 & ~x26 ;
  assign n2279 = n2277 | n2278 ;
  assign n2280 = n2133 & ~n2279 ;
  assign n2281 = x65 & n2280 ;
  assign n2282 = n2276 | n2281 ;
  assign n2283 = n2133 & n2279 ;
  assign n2284 = n142 & n2283 ;
  assign n2285 = n2282 | n2284 ;
  assign n2286 = x26 | n2285 ;
  assign n2287 = ~x26 & n2286 ;
  assign n2288 = ( ~n2285 & n2286 ) | ( ~n2285 & n2287 ) | ( n2286 & n2287 ) ;
  assign n2289 = x26 & ~n2134 ;
  assign n2290 = n2288 & n2289 ;
  assign n2291 = n2288 | n2289 ;
  assign n2292 = ~n2290 & n2291 ;
  assign n2293 = ( n2146 & n2271 ) | ( n2146 & n2292 ) | ( n2271 & n2292 ) ;
  assign n2294 = ( n2146 & n2292 ) | ( n2146 & ~n2293 ) | ( n2292 & ~n2293 ) ;
  assign n2295 = ( n2271 & ~n2293 ) | ( n2271 & n2294 ) | ( ~n2293 & n2294 ) ;
  assign n2296 = n2260 & n2295 ;
  assign n2297 = n2260 | n2295 ;
  assign n2298 = ~n2296 & n2297 ;
  assign n2299 = ( n1990 & n2130 ) | ( n1990 & n2148 ) | ( n2130 & n2148 ) ;
  assign n2300 = n2298 | n2299 ;
  assign n2301 = n2298 & n2299 ;
  assign n2302 = n2300 & ~n2301 ;
  assign n2303 = x74 & n1071 ;
  assign n2304 = x73 & n1066 ;
  assign n2305 = x72 & ~n1065 ;
  assign n2306 = n1189 & n2305 ;
  assign n2307 = n2304 | n2306 ;
  assign n2308 = n2303 | n2307 ;
  assign n2309 = n1074 | n2308 ;
  assign n2310 = ( n587 & n2308 ) | ( n587 & n2309 ) | ( n2308 & n2309 ) ;
  assign n2311 = x17 & n2310 ;
  assign n2312 = x17 & ~n2311 ;
  assign n2313 = ( n2310 & ~n2311 ) | ( n2310 & n2312 ) | ( ~n2311 & n2312 ) ;
  assign n2314 = n2302 & n2313 ;
  assign n2315 = n2302 & ~n2314 ;
  assign n2316 = ~n2302 & n2313 ;
  assign n2317 = n2315 | n2316 ;
  assign n2318 = n2163 | n2166 ;
  assign n2319 = n2317 | n2318 ;
  assign n2320 = n2317 & n2318 ;
  assign n2321 = n2319 & ~n2320 ;
  assign n2322 = x77 & n771 ;
  assign n2323 = x76 & n766 ;
  assign n2324 = x75 & ~n765 ;
  assign n2325 = n905 & n2324 ;
  assign n2326 = n2323 | n2325 ;
  assign n2327 = n2322 | n2326 ;
  assign n2328 = n774 | n2327 ;
  assign n2329 = ( n846 & n2327 ) | ( n846 & n2328 ) | ( n2327 & n2328 ) ;
  assign n2330 = x14 & n2329 ;
  assign n2331 = x14 & ~n2330 ;
  assign n2332 = ( n2329 & ~n2330 ) | ( n2329 & n2331 ) | ( ~n2330 & n2331 ) ;
  assign n2333 = n2321 | n2332 ;
  assign n2334 = n2321 & n2332 ;
  assign n2335 = n2333 & ~n2334 ;
  assign n2336 = n2181 | n2184 ;
  assign n2337 = n2335 & n2336 ;
  assign n2338 = n2335 | n2336 ;
  assign n2339 = ~n2337 & n2338 ;
  assign n2340 = x80 & n528 ;
  assign n2341 = x79 & n523 ;
  assign n2342 = x78 & ~n522 ;
  assign n2343 = n635 & n2342 ;
  assign n2344 = n2341 | n2343 ;
  assign n2345 = n2340 | n2344 ;
  assign n2346 = n531 | n2345 ;
  assign n2347 = ( n1147 & n2345 ) | ( n1147 & n2346 ) | ( n2345 & n2346 ) ;
  assign n2348 = x11 & n2347 ;
  assign n2349 = x11 & ~n2348 ;
  assign n2350 = ( n2347 & ~n2348 ) | ( n2347 & n2349 ) | ( ~n2348 & n2349 ) ;
  assign n2351 = n2339 & n2350 ;
  assign n2352 = n2339 & ~n2351 ;
  assign n2353 = ~n2339 & n2350 ;
  assign n2354 = n2352 | n2353 ;
  assign n2355 = n2198 | n2204 ;
  assign n2356 = n2354 | n2355 ;
  assign n2357 = n2354 & n2355 ;
  assign n2358 = n2356 & ~n2357 ;
  assign n2359 = x83 & n337 ;
  assign n2360 = x82 & n332 ;
  assign n2361 = x81 & ~n331 ;
  assign n2362 = n396 & n2361 ;
  assign n2363 = n2360 | n2362 ;
  assign n2364 = n2359 | n2363 ;
  assign n2365 = n340 | n2364 ;
  assign n2366 = ( n1510 & n2364 ) | ( n1510 & n2365 ) | ( n2364 & n2365 ) ;
  assign n2367 = x8 & n2366 ;
  assign n2368 = x8 & ~n2367 ;
  assign n2369 = ( n2366 & ~n2367 ) | ( n2366 & n2368 ) | ( ~n2367 & n2368 ) ;
  assign n2370 = n2358 & n2369 ;
  assign n2371 = n2358 & ~n2370 ;
  assign n2372 = ~n2358 & n2369 ;
  assign n2373 = n2371 | n2372 ;
  assign n2374 = n2218 | n2221 ;
  assign n2375 = n2373 & n2374 ;
  assign n2376 = n2373 & ~n2375 ;
  assign n2377 = n2374 & ~n2375 ;
  assign n2378 = n2376 | n2377 ;
  assign n2379 = x86 & n206 ;
  assign n2380 = x85 & n201 ;
  assign n2381 = x84 & ~n200 ;
  assign n2382 = n243 & n2381 ;
  assign n2383 = n2380 | n2382 ;
  assign n2384 = n2379 | n2383 ;
  assign n2385 = n209 | n2384 ;
  assign n2386 = ( n1921 & n2384 ) | ( n1921 & n2385 ) | ( n2384 & n2385 ) ;
  assign n2387 = x5 & n2386 ;
  assign n2388 = x5 & ~n2387 ;
  assign n2389 = ( n2386 & ~n2387 ) | ( n2386 & n2388 ) | ( ~n2387 & n2388 ) ;
  assign n2390 = ( n2249 & n2378 ) | ( n2249 & ~n2389 ) | ( n2378 & ~n2389 ) ;
  assign n2391 = ( ~n2378 & n2389 ) | ( ~n2378 & n2390 ) | ( n2389 & n2390 ) ;
  assign n2392 = ( ~n2249 & n2390 ) | ( ~n2249 & n2391 ) | ( n2390 & n2391 ) ;
  assign n2393 = n2248 & n2392 ;
  assign n2394 = n2248 | n2392 ;
  assign n2395 = ~n2393 & n2394 ;
  assign n2396 = n2227 | n2231 ;
  assign n2397 = n2395 & n2396 ;
  assign n2398 = n2395 | n2396 ;
  assign n2399 = ~n2397 & n2398 ;
  assign n2400 = x88 | x89 ;
  assign n2401 = x89 | x90 ;
  assign n2402 = x89 & x90 ;
  assign n2403 = n2401 & ~n2402 ;
  assign n2404 = n2400 & n2403 ;
  assign n2405 = x88 & x89 ;
  assign n2406 = n2403 & n2405 ;
  assign n2407 = ( n2241 & n2404 ) | ( n2241 & n2406 ) | ( n2404 & n2406 ) ;
  assign n2408 = ( n2241 & n2400 ) | ( n2241 & n2405 ) | ( n2400 & n2405 ) ;
  assign n2409 = n2403 | n2408 ;
  assign n2410 = ~n2407 & n2409 ;
  assign n2411 = x89 & n131 ;
  assign n2412 = x88 & ~n156 ;
  assign n2413 = ( n135 & n2411 ) | ( n135 & n2412 ) | ( n2411 & n2412 ) ;
  assign n2414 = x0 & x90 ;
  assign n2415 = ( ~n135 & n2411 ) | ( ~n135 & n2414 ) | ( n2411 & n2414 ) ;
  assign n2416 = n2413 | n2415 ;
  assign n2417 = n139 | n2416 ;
  assign n2418 = ( n2410 & n2416 ) | ( n2410 & n2417 ) | ( n2416 & n2417 ) ;
  assign n2419 = x2 & n2418 ;
  assign n2420 = x2 & ~n2419 ;
  assign n2421 = ( n2418 & ~n2419 ) | ( n2418 & n2420 ) | ( ~n2419 & n2420 ) ;
  assign n2422 = x87 & n206 ;
  assign n2423 = x86 & n201 ;
  assign n2424 = x85 & ~n200 ;
  assign n2425 = n243 & n2424 ;
  assign n2426 = n2423 | n2425 ;
  assign n2427 = n2422 | n2426 ;
  assign n2428 = n209 | n2427 ;
  assign n2429 = ( n2067 & n2427 ) | ( n2067 & n2428 ) | ( n2427 & n2428 ) ;
  assign n2430 = x5 & n2429 ;
  assign n2431 = x5 & ~n2430 ;
  assign n2432 = ( n2429 & ~n2430 ) | ( n2429 & n2431 ) | ( ~n2430 & n2431 ) ;
  assign n2433 = n2351 | n2357 ;
  assign n2434 = x81 & n528 ;
  assign n2435 = x80 & n523 ;
  assign n2436 = x79 & ~n522 ;
  assign n2437 = n635 & n2436 ;
  assign n2438 = n2435 | n2437 ;
  assign n2439 = n2434 | n2438 ;
  assign n2440 = n531 | n2439 ;
  assign n2441 = ( n1256 & n2439 ) | ( n1256 & n2440 ) | ( n2439 & n2440 ) ;
  assign n2442 = x11 & n2441 ;
  assign n2443 = x11 & ~n2442 ;
  assign n2444 = ( n2441 & ~n2442 ) | ( n2441 & n2443 ) | ( ~n2442 & n2443 ) ;
  assign n2445 = x78 & n771 ;
  assign n2446 = x77 & n766 ;
  assign n2447 = x76 & ~n765 ;
  assign n2448 = n905 & n2447 ;
  assign n2449 = n2446 | n2448 ;
  assign n2450 = n2445 | n2449 ;
  assign n2451 = n774 | n2450 ;
  assign n2452 = ( n868 & n2450 ) | ( n868 & n2451 ) | ( n2450 & n2451 ) ;
  assign n2453 = x14 & n2452 ;
  assign n2454 = x14 & ~n2453 ;
  assign n2455 = ( n2452 & ~n2453 ) | ( n2452 & n2454 ) | ( ~n2453 & n2454 ) ;
  assign n2456 = n2334 | n2337 ;
  assign n2457 = x72 & n1421 ;
  assign n2458 = x71 & n1416 ;
  assign n2459 = x70 & ~n1415 ;
  assign n2460 = n1584 & n2459 ;
  assign n2461 = n2458 | n2460 ;
  assign n2462 = n2457 | n2461 ;
  assign n2463 = ( n435 & n1424 ) | ( n435 & n2462 ) | ( n1424 & n2462 ) ;
  assign n2464 = ( x20 & ~n2462 ) | ( x20 & n2463 ) | ( ~n2462 & n2463 ) ;
  assign n2465 = ~n2463 & n2464 ;
  assign n2466 = n2462 | n2464 ;
  assign n2467 = ( ~x20 & n2465 ) | ( ~x20 & n2466 ) | ( n2465 & n2466 ) ;
  assign n2468 = n264 & n1820 ;
  assign n2469 = x69 & n1817 ;
  assign n2470 = x68 & n1812 ;
  assign n2471 = x67 & ~n1811 ;
  assign n2472 = n1977 & n2471 ;
  assign n2473 = n2470 | n2472 ;
  assign n2474 = n2469 | n2473 ;
  assign n2475 = n2468 | n2474 ;
  assign n2476 = x23 | n2475 ;
  assign n2477 = ~x23 & n2476 ;
  assign n2478 = ( ~n2475 & n2476 ) | ( ~n2475 & n2477 ) | ( n2476 & n2477 ) ;
  assign n2479 = x66 & n2280 ;
  assign n2480 = x65 & n2275 ;
  assign n2481 = ~n2133 & n2279 ;
  assign n2482 = x64 & ~n2274 ;
  assign n2483 = n2481 & n2482 ;
  assign n2484 = n2480 | n2483 ;
  assign n2485 = n2479 | n2484 ;
  assign n2486 = n153 & n2283 ;
  assign n2487 = n2485 | n2486 ;
  assign n2488 = x26 | n2487 ;
  assign n2489 = ~x26 & n2488 ;
  assign n2490 = ( ~n2487 & n2488 ) | ( ~n2487 & n2489 ) | ( n2488 & n2489 ) ;
  assign n2491 = n2290 | n2490 ;
  assign n2492 = n2290 & n2490 ;
  assign n2493 = n2491 & ~n2492 ;
  assign n2494 = ( n2293 & n2478 ) | ( n2293 & n2493 ) | ( n2478 & n2493 ) ;
  assign n2495 = ( n2293 & n2493 ) | ( n2293 & ~n2494 ) | ( n2493 & ~n2494 ) ;
  assign n2496 = ( n2478 & ~n2494 ) | ( n2478 & n2495 ) | ( ~n2494 & n2495 ) ;
  assign n2497 = n2467 | n2496 ;
  assign n2498 = n2467 & n2496 ;
  assign n2499 = n2497 & ~n2498 ;
  assign n2500 = n2296 | n2301 ;
  assign n2501 = n2499 & n2500 ;
  assign n2502 = n2499 | n2500 ;
  assign n2503 = ~n2501 & n2502 ;
  assign n2504 = x75 & n1071 ;
  assign n2505 = x74 & n1066 ;
  assign n2506 = x73 & ~n1065 ;
  assign n2507 = n1189 & n2506 ;
  assign n2508 = n2505 | n2507 ;
  assign n2509 = n2504 | n2508 ;
  assign n2510 = n1074 | n2509 ;
  assign n2511 = ( n609 & n2509 ) | ( n609 & n2510 ) | ( n2509 & n2510 ) ;
  assign n2512 = x17 & n2511 ;
  assign n2513 = x17 & ~n2512 ;
  assign n2514 = ( n2511 & ~n2512 ) | ( n2511 & n2513 ) | ( ~n2512 & n2513 ) ;
  assign n2515 = n2503 | n2514 ;
  assign n2516 = n2503 & n2514 ;
  assign n2517 = n2515 & ~n2516 ;
  assign n2518 = n2314 | n2320 ;
  assign n2519 = n2517 & n2518 ;
  assign n2520 = n2517 | n2518 ;
  assign n2521 = ~n2519 & n2520 ;
  assign n2522 = ( n2455 & n2456 ) | ( n2455 & ~n2521 ) | ( n2456 & ~n2521 ) ;
  assign n2523 = ( ~n2456 & n2521 ) | ( ~n2456 & n2522 ) | ( n2521 & n2522 ) ;
  assign n2524 = ( ~n2455 & n2522 ) | ( ~n2455 & n2523 ) | ( n2522 & n2523 ) ;
  assign n2525 = n2444 & n2524 ;
  assign n2526 = n2444 | n2524 ;
  assign n2527 = ~n2525 & n2526 ;
  assign n2528 = n2433 | n2527 ;
  assign n2529 = n2433 & n2527 ;
  assign n2530 = n2528 & ~n2529 ;
  assign n2531 = x84 & n337 ;
  assign n2532 = x83 & n332 ;
  assign n2533 = x82 & ~n331 ;
  assign n2534 = n396 & n2533 ;
  assign n2535 = n2532 | n2534 ;
  assign n2536 = n2531 | n2535 ;
  assign n2537 = n340 | n2536 ;
  assign n2538 = ( n1537 & n2536 ) | ( n1537 & n2537 ) | ( n2536 & n2537 ) ;
  assign n2539 = x8 & n2538 ;
  assign n2540 = x8 & ~n2539 ;
  assign n2541 = ( n2538 & ~n2539 ) | ( n2538 & n2540 ) | ( ~n2539 & n2540 ) ;
  assign n2542 = n2530 & n2541 ;
  assign n2543 = n2530 & ~n2542 ;
  assign n2544 = ~n2530 & n2541 ;
  assign n2545 = n2543 | n2544 ;
  assign n2546 = n2370 | n2375 ;
  assign n2547 = n2545 | n2546 ;
  assign n2548 = n2545 & n2546 ;
  assign n2549 = n2547 & ~n2548 ;
  assign n2550 = ( n2249 & n2378 ) | ( n2249 & n2389 ) | ( n2378 & n2389 ) ;
  assign n2551 = ( n2432 & n2549 ) | ( n2432 & n2550 ) | ( n2549 & n2550 ) ;
  assign n2552 = ( n2549 & n2550 ) | ( n2549 & ~n2551 ) | ( n2550 & ~n2551 ) ;
  assign n2553 = ( n2432 & ~n2551 ) | ( n2432 & n2552 ) | ( ~n2551 & n2552 ) ;
  assign n2554 = n2421 & n2553 ;
  assign n2555 = n2421 | n2553 ;
  assign n2556 = ~n2554 & n2555 ;
  assign n2557 = n2393 | n2397 ;
  assign n2558 = n2556 & n2557 ;
  assign n2559 = n2556 | n2557 ;
  assign n2560 = ~n2558 & n2559 ;
  assign n2561 = n2554 | n2558 ;
  assign n2562 = n2498 | n2501 ;
  assign n2563 = x73 & n1421 ;
  assign n2564 = x72 & n1416 ;
  assign n2565 = x71 & ~n1415 ;
  assign n2566 = n1584 & n2565 ;
  assign n2567 = n2564 | n2566 ;
  assign n2568 = n2563 | n2567 ;
  assign n2569 = n1424 | n2568 ;
  assign n2570 = ( n499 & n2568 ) | ( n499 & n2569 ) | ( n2568 & n2569 ) ;
  assign n2571 = x20 & n2570 ;
  assign n2572 = x20 | n2570 ;
  assign n2573 = ~n2571 & n2572 ;
  assign n2574 = x70 & n1817 ;
  assign n2575 = x69 & n1812 ;
  assign n2576 = x68 & ~n1811 ;
  assign n2577 = n1977 & n2576 ;
  assign n2578 = n2575 | n2577 ;
  assign n2579 = n2574 | n2578 ;
  assign n2580 = n1820 | n2579 ;
  assign n2581 = ( n310 & n2579 ) | ( n310 & n2580 ) | ( n2579 & n2580 ) ;
  assign n2582 = x23 & ~n2581 ;
  assign n2583 = ~x23 & n2581 ;
  assign n2584 = n2582 | n2583 ;
  assign n2585 = x26 & ~x27 ;
  assign n2586 = ~x26 & x27 ;
  assign n2587 = n2585 | n2586 ;
  assign n2588 = x64 & n2587 ;
  assign n2589 = x67 & n2280 ;
  assign n2590 = x66 & n2275 ;
  assign n2591 = x65 & ~n2274 ;
  assign n2592 = n2481 & n2591 ;
  assign n2593 = n2590 | n2592 ;
  assign n2594 = n2589 | n2593 ;
  assign n2595 = n180 & n2283 ;
  assign n2596 = n2594 | n2595 ;
  assign n2597 = x26 & ~n2596 ;
  assign n2598 = ~x26 & n2596 ;
  assign n2599 = n2597 | n2598 ;
  assign n2600 = ( n2492 & n2588 ) | ( n2492 & n2599 ) | ( n2588 & n2599 ) ;
  assign n2601 = ( n2492 & n2599 ) | ( n2492 & ~n2600 ) | ( n2599 & ~n2600 ) ;
  assign n2602 = ( n2588 & ~n2600 ) | ( n2588 & n2601 ) | ( ~n2600 & n2601 ) ;
  assign n2603 = ( n2494 & n2584 ) | ( n2494 & ~n2602 ) | ( n2584 & ~n2602 ) ;
  assign n2604 = ( ~n2494 & n2602 ) | ( ~n2494 & n2603 ) | ( n2602 & n2603 ) ;
  assign n2605 = ( ~n2584 & n2603 ) | ( ~n2584 & n2604 ) | ( n2603 & n2604 ) ;
  assign n2606 = n2573 & n2605 ;
  assign n2607 = n2573 | n2605 ;
  assign n2608 = ~n2606 & n2607 ;
  assign n2609 = n2562 & n2608 ;
  assign n2610 = n2562 | n2608 ;
  assign n2611 = ~n2609 & n2610 ;
  assign n2612 = x76 & n1071 ;
  assign n2613 = x75 & n1066 ;
  assign n2614 = x74 & ~n1065 ;
  assign n2615 = n1189 & n2614 ;
  assign n2616 = n2613 | n2615 ;
  assign n2617 = n2612 | n2616 ;
  assign n2618 = n1074 | n2617 ;
  assign n2619 = ( n740 & n2617 ) | ( n740 & n2618 ) | ( n2617 & n2618 ) ;
  assign n2620 = x17 & n2619 ;
  assign n2621 = x17 & ~n2620 ;
  assign n2622 = ( n2619 & ~n2620 ) | ( n2619 & n2621 ) | ( ~n2620 & n2621 ) ;
  assign n2623 = n2611 | n2622 ;
  assign n2624 = n2611 & n2622 ;
  assign n2625 = n2623 & ~n2624 ;
  assign n2626 = n2516 | n2519 ;
  assign n2627 = n2625 & n2626 ;
  assign n2628 = n2625 | n2626 ;
  assign n2629 = ~n2627 & n2628 ;
  assign n2630 = x79 & n771 ;
  assign n2631 = x78 & n766 ;
  assign n2632 = x77 & ~n765 ;
  assign n2633 = n905 & n2632 ;
  assign n2634 = n2631 | n2633 ;
  assign n2635 = n2630 | n2634 ;
  assign n2636 = n774 | n2635 ;
  assign n2637 = ( n961 & n2635 ) | ( n961 & n2636 ) | ( n2635 & n2636 ) ;
  assign n2638 = x14 & n2637 ;
  assign n2639 = x14 & ~n2638 ;
  assign n2640 = ( n2637 & ~n2638 ) | ( n2637 & n2639 ) | ( ~n2638 & n2639 ) ;
  assign n2641 = n2629 & n2640 ;
  assign n2642 = n2629 & ~n2641 ;
  assign n2643 = ~n2629 & n2640 ;
  assign n2644 = n2642 | n2643 ;
  assign n2645 = ( n2455 & n2456 ) | ( n2455 & n2521 ) | ( n2456 & n2521 ) ;
  assign n2646 = n2644 | n2645 ;
  assign n2647 = n2644 & n2645 ;
  assign n2648 = n2646 & ~n2647 ;
  assign n2649 = x82 & n528 ;
  assign n2650 = x81 & n523 ;
  assign n2651 = x80 & ~n522 ;
  assign n2652 = n635 & n2651 ;
  assign n2653 = n2650 | n2652 ;
  assign n2654 = n2649 | n2653 ;
  assign n2655 = n531 | n2654 ;
  assign n2656 = ( n1371 & n2654 ) | ( n1371 & n2655 ) | ( n2654 & n2655 ) ;
  assign n2657 = x11 & n2656 ;
  assign n2658 = x11 & ~n2657 ;
  assign n2659 = ( n2656 & ~n2657 ) | ( n2656 & n2658 ) | ( ~n2657 & n2658 ) ;
  assign n2660 = n2648 & n2659 ;
  assign n2661 = n2648 & ~n2660 ;
  assign n2662 = ~n2648 & n2659 ;
  assign n2663 = n2661 | n2662 ;
  assign n2664 = n2525 | n2529 ;
  assign n2665 = n2663 | n2664 ;
  assign n2666 = n2663 & n2664 ;
  assign n2667 = n2665 & ~n2666 ;
  assign n2668 = x85 & n337 ;
  assign n2669 = x84 & n332 ;
  assign n2670 = x83 & ~n331 ;
  assign n2671 = n396 & n2670 ;
  assign n2672 = n2669 | n2671 ;
  assign n2673 = n2668 | n2672 ;
  assign n2674 = n340 | n2673 ;
  assign n2675 = ( n1765 & n2673 ) | ( n1765 & n2674 ) | ( n2673 & n2674 ) ;
  assign n2676 = x8 & n2675 ;
  assign n2677 = x8 & ~n2676 ;
  assign n2678 = ( n2675 & ~n2676 ) | ( n2675 & n2677 ) | ( ~n2676 & n2677 ) ;
  assign n2679 = n2667 | n2678 ;
  assign n2680 = n2667 & n2678 ;
  assign n2681 = n2679 & ~n2680 ;
  assign n2682 = n2542 | n2548 ;
  assign n2683 = n2681 & n2682 ;
  assign n2684 = n2681 | n2682 ;
  assign n2685 = ~n2683 & n2684 ;
  assign n2686 = x88 & n206 ;
  assign n2687 = x87 & n201 ;
  assign n2688 = x86 & ~n200 ;
  assign n2689 = n243 & n2688 ;
  assign n2690 = n2687 | n2689 ;
  assign n2691 = n2686 | n2690 ;
  assign n2692 = n209 | n2691 ;
  assign n2693 = ( n2095 & n2691 ) | ( n2095 & n2692 ) | ( n2691 & n2692 ) ;
  assign n2694 = x5 & n2693 ;
  assign n2695 = x5 & ~n2694 ;
  assign n2696 = ( n2693 & ~n2694 ) | ( n2693 & n2695 ) | ( ~n2694 & n2695 ) ;
  assign n2697 = n2685 & n2696 ;
  assign n2698 = n2685 & ~n2697 ;
  assign n2699 = ~n2685 & n2696 ;
  assign n2700 = n2698 | n2699 ;
  assign n2701 = n2551 | n2700 ;
  assign n2702 = n2551 & n2700 ;
  assign n2703 = n2701 & ~n2702 ;
  assign n2704 = x90 | x91 ;
  assign n2705 = x90 & x91 ;
  assign n2706 = n2704 & ~n2705 ;
  assign n2707 = n2402 | n2404 ;
  assign n2708 = n2706 & n2707 ;
  assign n2709 = n2402 | n2406 ;
  assign n2710 = n2706 & n2709 ;
  assign n2711 = ( n2241 & n2708 ) | ( n2241 & n2710 ) | ( n2708 & n2710 ) ;
  assign n2712 = ( n2241 & n2707 ) | ( n2241 & n2709 ) | ( n2707 & n2709 ) ;
  assign n2713 = n2706 | n2712 ;
  assign n2714 = ~n2711 & n2713 ;
  assign n2715 = x90 & n131 ;
  assign n2716 = x89 & ~n156 ;
  assign n2717 = ( n135 & n2715 ) | ( n135 & n2716 ) | ( n2715 & n2716 ) ;
  assign n2718 = x0 & x91 ;
  assign n2719 = ( ~n135 & n2715 ) | ( ~n135 & n2718 ) | ( n2715 & n2718 ) ;
  assign n2720 = n2717 | n2719 ;
  assign n2721 = n139 | n2720 ;
  assign n2722 = ( n2714 & n2720 ) | ( n2714 & n2721 ) | ( n2720 & n2721 ) ;
  assign n2723 = x2 & n2722 ;
  assign n2724 = x2 & ~n2723 ;
  assign n2725 = ( n2722 & ~n2723 ) | ( n2722 & n2724 ) | ( ~n2723 & n2724 ) ;
  assign n2726 = n2703 | n2725 ;
  assign n2727 = n2703 & n2725 ;
  assign n2728 = n2726 & ~n2727 ;
  assign n2729 = n2561 & n2728 ;
  assign n2730 = n2561 | n2728 ;
  assign n2731 = ~n2729 & n2730 ;
  assign n2732 = n2727 | n2729 ;
  assign n2733 = x80 & n771 ;
  assign n2734 = x79 & n766 ;
  assign n2735 = x78 & ~n765 ;
  assign n2736 = n905 & n2735 ;
  assign n2737 = n2734 | n2736 ;
  assign n2738 = n2733 | n2737 ;
  assign n2739 = n774 | n2738 ;
  assign n2740 = ( n1147 & n2738 ) | ( n1147 & n2739 ) | ( n2738 & n2739 ) ;
  assign n2741 = x14 & n2740 ;
  assign n2742 = x14 & ~n2741 ;
  assign n2743 = ( n2740 & ~n2741 ) | ( n2740 & n2742 ) | ( ~n2741 & n2742 ) ;
  assign n2744 = n2624 | n2627 ;
  assign n2745 = x71 & n1817 ;
  assign n2746 = x70 & n1812 ;
  assign n2747 = x69 & ~n1811 ;
  assign n2748 = n1977 & n2747 ;
  assign n2749 = n2746 | n2748 ;
  assign n2750 = n2745 | n2749 ;
  assign n2751 = n1820 | n2750 ;
  assign n2752 = ( n376 & n2750 ) | ( n376 & n2751 ) | ( n2750 & n2751 ) ;
  assign n2753 = x23 & ~n2752 ;
  assign n2754 = ~x23 & n2752 ;
  assign n2755 = n2753 | n2754 ;
  assign n2756 = n229 & n2283 ;
  assign n2757 = x68 & n2280 ;
  assign n2758 = x67 & n2275 ;
  assign n2759 = x66 & ~n2274 ;
  assign n2760 = n2481 & n2759 ;
  assign n2761 = n2758 | n2760 ;
  assign n2762 = n2757 | n2761 ;
  assign n2763 = n2756 | n2762 ;
  assign n2764 = x26 | n2763 ;
  assign n2765 = ~x26 & n2764 ;
  assign n2766 = ( ~n2763 & n2764 ) | ( ~n2763 & n2765 ) | ( n2764 & n2765 ) ;
  assign n2767 = ~x27 & x28 ;
  assign n2768 = x27 & ~x28 ;
  assign n2769 = n2767 | n2768 ;
  assign n2770 = ~n2587 & n2769 ;
  assign n2771 = x64 & n2770 ;
  assign n2772 = ~x28 & x29 ;
  assign n2773 = x28 & ~x29 ;
  assign n2774 = n2772 | n2773 ;
  assign n2775 = n2587 & ~n2774 ;
  assign n2776 = x65 & n2775 ;
  assign n2777 = n2771 | n2776 ;
  assign n2778 = n2587 & n2774 ;
  assign n2779 = n142 & n2778 ;
  assign n2780 = n2777 | n2779 ;
  assign n2781 = x29 | n2780 ;
  assign n2782 = ~x29 & n2781 ;
  assign n2783 = ( ~n2780 & n2781 ) | ( ~n2780 & n2782 ) | ( n2781 & n2782 ) ;
  assign n2784 = x29 & ~n2588 ;
  assign n2785 = n2783 & n2784 ;
  assign n2786 = n2783 | n2784 ;
  assign n2787 = ~n2785 & n2786 ;
  assign n2788 = ( n2600 & n2766 ) | ( n2600 & n2787 ) | ( n2766 & n2787 ) ;
  assign n2789 = ( n2600 & n2787 ) | ( n2600 & ~n2788 ) | ( n2787 & ~n2788 ) ;
  assign n2790 = ( n2766 & ~n2788 ) | ( n2766 & n2789 ) | ( ~n2788 & n2789 ) ;
  assign n2791 = n2755 & n2790 ;
  assign n2792 = n2755 | n2790 ;
  assign n2793 = ~n2791 & n2792 ;
  assign n2794 = ( n2494 & n2584 ) | ( n2494 & ~n2605 ) | ( n2584 & ~n2605 ) ;
  assign n2795 = n2793 & n2794 ;
  assign n2796 = n2793 | n2794 ;
  assign n2797 = ~n2795 & n2796 ;
  assign n2798 = x74 & n1421 ;
  assign n2799 = x73 & n1416 ;
  assign n2800 = x72 & ~n1415 ;
  assign n2801 = n1584 & n2800 ;
  assign n2802 = n2799 | n2801 ;
  assign n2803 = n2798 | n2802 ;
  assign n2804 = n1424 | n2803 ;
  assign n2805 = ( n587 & n2803 ) | ( n587 & n2804 ) | ( n2803 & n2804 ) ;
  assign n2806 = x20 & n2805 ;
  assign n2807 = x20 & ~n2806 ;
  assign n2808 = ( n2805 & ~n2806 ) | ( n2805 & n2807 ) | ( ~n2806 & n2807 ) ;
  assign n2809 = n2797 & n2808 ;
  assign n2810 = n2797 & ~n2809 ;
  assign n2811 = ~n2797 & n2808 ;
  assign n2812 = n2810 | n2811 ;
  assign n2813 = n2606 | n2609 ;
  assign n2814 = n2812 | n2813 ;
  assign n2815 = n2812 & n2813 ;
  assign n2816 = n2814 & ~n2815 ;
  assign n2817 = x77 & n1071 ;
  assign n2818 = x76 & n1066 ;
  assign n2819 = x75 & ~n1065 ;
  assign n2820 = n1189 & n2819 ;
  assign n2821 = n2818 | n2820 ;
  assign n2822 = n2817 | n2821 ;
  assign n2823 = n1074 | n2822 ;
  assign n2824 = ( n846 & n2822 ) | ( n846 & n2823 ) | ( n2822 & n2823 ) ;
  assign n2825 = x17 & n2824 ;
  assign n2826 = x17 & ~n2825 ;
  assign n2827 = ( n2824 & ~n2825 ) | ( n2824 & n2826 ) | ( ~n2825 & n2826 ) ;
  assign n2828 = ( n2744 & n2816 ) | ( n2744 & ~n2827 ) | ( n2816 & ~n2827 ) ;
  assign n2829 = ( ~n2816 & n2827 ) | ( ~n2816 & n2828 ) | ( n2827 & n2828 ) ;
  assign n2830 = ( ~n2744 & n2828 ) | ( ~n2744 & n2829 ) | ( n2828 & n2829 ) ;
  assign n2831 = n2743 & n2830 ;
  assign n2832 = n2743 | n2830 ;
  assign n2833 = ~n2831 & n2832 ;
  assign n2834 = n2641 | n2647 ;
  assign n2835 = n2833 | n2834 ;
  assign n2836 = n2833 & n2834 ;
  assign n2837 = n2835 & ~n2836 ;
  assign n2838 = x83 & n528 ;
  assign n2839 = x82 & n523 ;
  assign n2840 = x81 & ~n522 ;
  assign n2841 = n635 & n2840 ;
  assign n2842 = n2839 | n2841 ;
  assign n2843 = n2838 | n2842 ;
  assign n2844 = n531 | n2843 ;
  assign n2845 = ( n1510 & n2843 ) | ( n1510 & n2844 ) | ( n2843 & n2844 ) ;
  assign n2846 = x11 & n2845 ;
  assign n2847 = x11 & ~n2846 ;
  assign n2848 = ( n2845 & ~n2846 ) | ( n2845 & n2847 ) | ( ~n2846 & n2847 ) ;
  assign n2849 = n2837 & n2848 ;
  assign n2850 = n2837 & ~n2849 ;
  assign n2851 = ~n2837 & n2848 ;
  assign n2852 = n2850 | n2851 ;
  assign n2853 = n2660 | n2666 ;
  assign n2854 = n2852 | n2853 ;
  assign n2855 = n2852 & n2853 ;
  assign n2856 = n2854 & ~n2855 ;
  assign n2857 = x86 & n337 ;
  assign n2858 = x85 & n332 ;
  assign n2859 = x84 & ~n331 ;
  assign n2860 = n396 & n2859 ;
  assign n2861 = n2858 | n2860 ;
  assign n2862 = n2857 | n2861 ;
  assign n2863 = n340 | n2862 ;
  assign n2864 = ( n1921 & n2862 ) | ( n1921 & n2863 ) | ( n2862 & n2863 ) ;
  assign n2865 = x8 & n2864 ;
  assign n2866 = x8 & ~n2865 ;
  assign n2867 = ( n2864 & ~n2865 ) | ( n2864 & n2866 ) | ( ~n2865 & n2866 ) ;
  assign n2868 = n2856 | n2867 ;
  assign n2869 = n2856 & n2867 ;
  assign n2870 = n2868 & ~n2869 ;
  assign n2871 = n2680 | n2683 ;
  assign n2872 = n2870 & n2871 ;
  assign n2873 = n2870 | n2871 ;
  assign n2874 = ~n2872 & n2873 ;
  assign n2875 = x89 & n206 ;
  assign n2876 = x88 & n201 ;
  assign n2877 = x87 & ~n200 ;
  assign n2878 = n243 & n2877 ;
  assign n2879 = n2876 | n2878 ;
  assign n2880 = n2875 | n2879 ;
  assign n2881 = n209 | n2880 ;
  assign n2882 = ( n2244 & n2880 ) | ( n2244 & n2881 ) | ( n2880 & n2881 ) ;
  assign n2883 = x5 & n2882 ;
  assign n2884 = x5 & ~n2883 ;
  assign n2885 = ( n2882 & ~n2883 ) | ( n2882 & n2884 ) | ( ~n2883 & n2884 ) ;
  assign n2886 = n2874 & n2885 ;
  assign n2887 = n2874 & ~n2886 ;
  assign n2888 = ~n2874 & n2885 ;
  assign n2889 = n2887 | n2888 ;
  assign n2890 = n2697 | n2702 ;
  assign n2891 = n2889 | n2890 ;
  assign n2892 = n2889 & n2890 ;
  assign n2893 = n2891 & ~n2892 ;
  assign n2894 = x91 | x92 ;
  assign n2895 = x91 & x92 ;
  assign n2896 = n2894 & ~n2895 ;
  assign n2897 = n2705 | n2708 ;
  assign n2898 = n2896 & n2897 ;
  assign n2899 = n2705 | n2710 ;
  assign n2900 = n2896 & n2899 ;
  assign n2901 = ( n2241 & n2898 ) | ( n2241 & n2900 ) | ( n2898 & n2900 ) ;
  assign n2902 = ( n2241 & n2897 ) | ( n2241 & n2899 ) | ( n2897 & n2899 ) ;
  assign n2903 = n2896 | n2902 ;
  assign n2904 = ~n2901 & n2903 ;
  assign n2905 = x91 & n131 ;
  assign n2906 = x90 & ~n156 ;
  assign n2907 = ( n135 & n2905 ) | ( n135 & n2906 ) | ( n2905 & n2906 ) ;
  assign n2908 = x0 & x92 ;
  assign n2909 = ( ~n135 & n2905 ) | ( ~n135 & n2908 ) | ( n2905 & n2908 ) ;
  assign n2910 = n2907 | n2909 ;
  assign n2911 = n139 | n2910 ;
  assign n2912 = ( n2904 & n2910 ) | ( n2904 & n2911 ) | ( n2910 & n2911 ) ;
  assign n2913 = x2 & n2912 ;
  assign n2914 = x2 & ~n2913 ;
  assign n2915 = ( n2912 & ~n2913 ) | ( n2912 & n2914 ) | ( ~n2913 & n2914 ) ;
  assign n2916 = n2893 | n2915 ;
  assign n2917 = n2893 & n2915 ;
  assign n2918 = n2916 & ~n2917 ;
  assign n2919 = n2732 & n2918 ;
  assign n2920 = n2732 | n2918 ;
  assign n2921 = ~n2919 & n2920 ;
  assign n2922 = n2917 | n2919 ;
  assign n2923 = x92 | x93 ;
  assign n2924 = x92 & x93 ;
  assign n2925 = n2923 & ~n2924 ;
  assign n2926 = n2895 | n2898 ;
  assign n2927 = n2895 | n2900 ;
  assign n2928 = ( n2241 & n2926 ) | ( n2241 & n2927 ) | ( n2926 & n2927 ) ;
  assign n2929 = n2925 | n2928 ;
  assign n2930 = n2925 & n2928 ;
  assign n2931 = n2929 & ~n2930 ;
  assign n2932 = x92 & n131 ;
  assign n2933 = x91 & ~n156 ;
  assign n2934 = ( n135 & n2932 ) | ( n135 & n2933 ) | ( n2932 & n2933 ) ;
  assign n2935 = x0 & x93 ;
  assign n2936 = ( ~n135 & n2932 ) | ( ~n135 & n2935 ) | ( n2932 & n2935 ) ;
  assign n2937 = n2934 | n2936 ;
  assign n2938 = n139 | n2937 ;
  assign n2939 = ( n2931 & n2937 ) | ( n2931 & n2938 ) | ( n2937 & n2938 ) ;
  assign n2940 = x2 & n2939 ;
  assign n2941 = x2 & ~n2940 ;
  assign n2942 = ( n2939 & ~n2940 ) | ( n2939 & n2941 ) | ( ~n2940 & n2941 ) ;
  assign n2943 = x90 & n206 ;
  assign n2944 = x89 & n201 ;
  assign n2945 = x88 & ~n200 ;
  assign n2946 = n243 & n2945 ;
  assign n2947 = n2944 | n2946 ;
  assign n2948 = n2943 | n2947 ;
  assign n2949 = n209 | n2948 ;
  assign n2950 = ( n2410 & n2948 ) | ( n2410 & n2949 ) | ( n2948 & n2949 ) ;
  assign n2951 = x5 & n2950 ;
  assign n2952 = x5 & ~n2951 ;
  assign n2953 = ( n2950 & ~n2951 ) | ( n2950 & n2952 ) | ( ~n2951 & n2952 ) ;
  assign n2954 = x72 & n1817 ;
  assign n2955 = x71 & n1812 ;
  assign n2956 = x70 & ~n1811 ;
  assign n2957 = n1977 & n2956 ;
  assign n2958 = n2955 | n2957 ;
  assign n2959 = n2954 | n2958 ;
  assign n2960 = ( n435 & n1820 ) | ( n435 & n2959 ) | ( n1820 & n2959 ) ;
  assign n2961 = ( x23 & ~n2959 ) | ( x23 & n2960 ) | ( ~n2959 & n2960 ) ;
  assign n2962 = ~n2960 & n2961 ;
  assign n2963 = n2959 | n2961 ;
  assign n2964 = ( ~x23 & n2962 ) | ( ~x23 & n2963 ) | ( n2962 & n2963 ) ;
  assign n2965 = n264 & n2283 ;
  assign n2966 = x69 & n2280 ;
  assign n2967 = x68 & n2275 ;
  assign n2968 = x67 & ~n2274 ;
  assign n2969 = n2481 & n2968 ;
  assign n2970 = n2967 | n2969 ;
  assign n2971 = n2966 | n2970 ;
  assign n2972 = n2965 | n2971 ;
  assign n2973 = x26 | n2972 ;
  assign n2974 = ~x26 & n2973 ;
  assign n2975 = ( ~n2972 & n2973 ) | ( ~n2972 & n2974 ) | ( n2973 & n2974 ) ;
  assign n2976 = x66 & n2775 ;
  assign n2977 = x65 & n2770 ;
  assign n2978 = ~n2587 & n2774 ;
  assign n2979 = x64 & ~n2769 ;
  assign n2980 = n2978 & n2979 ;
  assign n2981 = n2977 | n2980 ;
  assign n2982 = n2976 | n2981 ;
  assign n2983 = n153 & n2778 ;
  assign n2984 = n2982 | n2983 ;
  assign n2985 = x29 | n2984 ;
  assign n2986 = ~x29 & n2985 ;
  assign n2987 = ( ~n2984 & n2985 ) | ( ~n2984 & n2986 ) | ( n2985 & n2986 ) ;
  assign n2988 = n2785 | n2987 ;
  assign n2989 = n2785 & n2987 ;
  assign n2990 = n2988 & ~n2989 ;
  assign n2991 = ( n2788 & n2975 ) | ( n2788 & n2990 ) | ( n2975 & n2990 ) ;
  assign n2992 = ( n2788 & n2990 ) | ( n2788 & ~n2991 ) | ( n2990 & ~n2991 ) ;
  assign n2993 = ( n2975 & ~n2991 ) | ( n2975 & n2992 ) | ( ~n2991 & n2992 ) ;
  assign n2994 = n2964 | n2993 ;
  assign n2995 = n2964 & n2993 ;
  assign n2996 = n2994 & ~n2995 ;
  assign n2997 = n2791 | n2795 ;
  assign n2998 = n2996 & n2997 ;
  assign n2999 = n2996 | n2997 ;
  assign n3000 = ~n2998 & n2999 ;
  assign n3001 = x75 & n1421 ;
  assign n3002 = x74 & n1416 ;
  assign n3003 = x73 & ~n1415 ;
  assign n3004 = n1584 & n3003 ;
  assign n3005 = n3002 | n3004 ;
  assign n3006 = n3001 | n3005 ;
  assign n3007 = n1424 | n3006 ;
  assign n3008 = ( n609 & n3006 ) | ( n609 & n3007 ) | ( n3006 & n3007 ) ;
  assign n3009 = x20 & n3008 ;
  assign n3010 = x20 & ~n3009 ;
  assign n3011 = ( n3008 & ~n3009 ) | ( n3008 & n3010 ) | ( ~n3009 & n3010 ) ;
  assign n3012 = n3000 | n3011 ;
  assign n3013 = n3000 & n3011 ;
  assign n3014 = n3012 & ~n3013 ;
  assign n3015 = n2809 | n2815 ;
  assign n3016 = n3014 & n3015 ;
  assign n3017 = n3014 | n3015 ;
  assign n3018 = ~n3016 & n3017 ;
  assign n3019 = x78 & n1071 ;
  assign n3020 = x77 & n1066 ;
  assign n3021 = x76 & ~n1065 ;
  assign n3022 = n1189 & n3021 ;
  assign n3023 = n3020 | n3022 ;
  assign n3024 = n3019 | n3023 ;
  assign n3025 = n1074 | n3024 ;
  assign n3026 = ( n868 & n3024 ) | ( n868 & n3025 ) | ( n3024 & n3025 ) ;
  assign n3027 = x17 & n3026 ;
  assign n3028 = x17 & ~n3027 ;
  assign n3029 = ( n3026 & ~n3027 ) | ( n3026 & n3028 ) | ( ~n3027 & n3028 ) ;
  assign n3030 = n3018 & n3029 ;
  assign n3031 = n3018 & ~n3030 ;
  assign n3032 = ~n3018 & n3029 ;
  assign n3033 = n3031 | n3032 ;
  assign n3034 = ( n2744 & n2816 ) | ( n2744 & n2827 ) | ( n2816 & n2827 ) ;
  assign n3035 = n3033 | n3034 ;
  assign n3036 = n3033 & n3034 ;
  assign n3037 = n3035 & ~n3036 ;
  assign n3038 = x81 & n771 ;
  assign n3039 = x80 & n766 ;
  assign n3040 = x79 & ~n765 ;
  assign n3041 = n905 & n3040 ;
  assign n3042 = n3039 | n3041 ;
  assign n3043 = n3038 | n3042 ;
  assign n3044 = n774 | n3043 ;
  assign n3045 = ( n1256 & n3043 ) | ( n1256 & n3044 ) | ( n3043 & n3044 ) ;
  assign n3046 = x14 & n3045 ;
  assign n3047 = x14 & ~n3046 ;
  assign n3048 = ( n3045 & ~n3046 ) | ( n3045 & n3047 ) | ( ~n3046 & n3047 ) ;
  assign n3049 = n3037 & n3048 ;
  assign n3050 = n3037 & ~n3049 ;
  assign n3051 = ~n3037 & n3048 ;
  assign n3052 = n3050 | n3051 ;
  assign n3053 = n2831 | n2836 ;
  assign n3054 = n3052 | n3053 ;
  assign n3055 = n3052 & n3053 ;
  assign n3056 = n3054 & ~n3055 ;
  assign n3057 = x84 & n528 ;
  assign n3058 = x83 & n523 ;
  assign n3059 = x82 & ~n522 ;
  assign n3060 = n635 & n3059 ;
  assign n3061 = n3058 | n3060 ;
  assign n3062 = n3057 | n3061 ;
  assign n3063 = n531 | n3062 ;
  assign n3064 = ( n1537 & n3062 ) | ( n1537 & n3063 ) | ( n3062 & n3063 ) ;
  assign n3065 = x11 & n3064 ;
  assign n3066 = x11 & ~n3065 ;
  assign n3067 = ( n3064 & ~n3065 ) | ( n3064 & n3066 ) | ( ~n3065 & n3066 ) ;
  assign n3068 = n3056 | n3067 ;
  assign n3069 = n2849 | n2855 ;
  assign n3070 = ( n3056 & n3067 ) | ( n3056 & n3069 ) | ( n3067 & n3069 ) ;
  assign n3071 = n3068 & ~n3070 ;
  assign n3072 = n3056 & n3067 ;
  assign n3073 = n3068 & ~n3072 ;
  assign n3074 = n3069 & ~n3073 ;
  assign n3075 = n3071 | n3074 ;
  assign n3076 = x87 & n337 ;
  assign n3077 = x86 & n332 ;
  assign n3078 = x85 & ~n331 ;
  assign n3079 = n396 & n3078 ;
  assign n3080 = n3077 | n3079 ;
  assign n3081 = n3076 | n3080 ;
  assign n3082 = n340 | n3081 ;
  assign n3083 = ( n2067 & n3081 ) | ( n2067 & n3082 ) | ( n3081 & n3082 ) ;
  assign n3084 = x8 & n3083 ;
  assign n3085 = x8 & ~n3084 ;
  assign n3086 = ( n3083 & ~n3084 ) | ( n3083 & n3085 ) | ( ~n3084 & n3085 ) ;
  assign n3087 = n3075 & n3086 ;
  assign n3088 = n3075 & ~n3087 ;
  assign n3089 = ~n3075 & n3086 ;
  assign n3090 = n3088 | n3089 ;
  assign n3091 = n2869 | n2872 ;
  assign n3092 = n3090 & n3091 ;
  assign n3093 = n3090 | n3091 ;
  assign n3094 = ~n3092 & n3093 ;
  assign n3095 = n2886 | n2892 ;
  assign n3096 = ( n2953 & n3094 ) | ( n2953 & n3095 ) | ( n3094 & n3095 ) ;
  assign n3097 = ( n3094 & n3095 ) | ( n3094 & ~n3096 ) | ( n3095 & ~n3096 ) ;
  assign n3098 = ( n2953 & ~n3096 ) | ( n2953 & n3097 ) | ( ~n3096 & n3097 ) ;
  assign n3099 = n2942 & n3098 ;
  assign n3100 = n2942 | n3098 ;
  assign n3101 = ~n3099 & n3100 ;
  assign n3102 = n2922 & n3101 ;
  assign n3103 = n2922 | n3101 ;
  assign n3104 = ~n3102 & n3103 ;
  assign n3105 = x88 & n337 ;
  assign n3106 = x87 & n332 ;
  assign n3107 = x86 & ~n331 ;
  assign n3108 = n396 & n3107 ;
  assign n3109 = n3106 | n3108 ;
  assign n3110 = n3105 | n3109 ;
  assign n3111 = n340 | n3110 ;
  assign n3112 = ( n2095 & n3110 ) | ( n2095 & n3111 ) | ( n3110 & n3111 ) ;
  assign n3113 = x8 & n3112 ;
  assign n3114 = x8 & ~n3113 ;
  assign n3115 = ( n3112 & ~n3113 ) | ( n3112 & n3114 ) | ( ~n3113 & n3114 ) ;
  assign n3116 = x85 & n528 ;
  assign n3117 = x84 & n523 ;
  assign n3118 = x83 & ~n522 ;
  assign n3119 = n635 & n3118 ;
  assign n3120 = n3117 | n3119 ;
  assign n3121 = n3116 | n3120 ;
  assign n3122 = n531 | n3121 ;
  assign n3123 = ( n1765 & n3121 ) | ( n1765 & n3122 ) | ( n3121 & n3122 ) ;
  assign n3124 = x11 & n3123 ;
  assign n3125 = x11 & ~n3124 ;
  assign n3126 = ( n3123 & ~n3124 ) | ( n3123 & n3125 ) | ( ~n3124 & n3125 ) ;
  assign n3127 = n2995 | n2998 ;
  assign n3128 = x70 & n2280 ;
  assign n3129 = x69 & n2275 ;
  assign n3130 = x68 & ~n2274 ;
  assign n3131 = n2481 & n3130 ;
  assign n3132 = n3129 | n3131 ;
  assign n3133 = n3128 | n3132 ;
  assign n3134 = n2283 | n3133 ;
  assign n3135 = ( n310 & n3133 ) | ( n310 & n3134 ) | ( n3133 & n3134 ) ;
  assign n3136 = x26 & ~n3135 ;
  assign n3137 = ~x26 & n3135 ;
  assign n3138 = n3136 | n3137 ;
  assign n3139 = x29 & ~x30 ;
  assign n3140 = ~x29 & x30 ;
  assign n3141 = n3139 | n3140 ;
  assign n3142 = x64 & n3141 ;
  assign n3143 = x67 & n2775 ;
  assign n3144 = x66 & n2770 ;
  assign n3145 = x65 & ~n2769 ;
  assign n3146 = n2978 & n3145 ;
  assign n3147 = n3144 | n3146 ;
  assign n3148 = n3143 | n3147 ;
  assign n3149 = n180 & n2778 ;
  assign n3150 = n3148 | n3149 ;
  assign n3151 = x29 & ~n3150 ;
  assign n3152 = ~x29 & n3150 ;
  assign n3153 = n3151 | n3152 ;
  assign n3154 = ( n2989 & n3142 ) | ( n2989 & n3153 ) | ( n3142 & n3153 ) ;
  assign n3155 = ( n2989 & n3153 ) | ( n2989 & ~n3154 ) | ( n3153 & ~n3154 ) ;
  assign n3156 = ( n3142 & ~n3154 ) | ( n3142 & n3155 ) | ( ~n3154 & n3155 ) ;
  assign n3157 = ( n2991 & n3138 ) | ( n2991 & ~n3156 ) | ( n3138 & ~n3156 ) ;
  assign n3158 = ( ~n2991 & n3156 ) | ( ~n2991 & n3157 ) | ( n3156 & n3157 ) ;
  assign n3159 = ( ~n3138 & n3157 ) | ( ~n3138 & n3158 ) | ( n3157 & n3158 ) ;
  assign n3160 = x73 & n1817 ;
  assign n3161 = x72 & n1812 ;
  assign n3162 = x71 & ~n1811 ;
  assign n3163 = n1977 & n3162 ;
  assign n3164 = n3161 | n3163 ;
  assign n3165 = n3160 | n3164 ;
  assign n3166 = ( n499 & n1820 ) | ( n499 & n3165 ) | ( n1820 & n3165 ) ;
  assign n3167 = ( x23 & ~n3165 ) | ( x23 & n3166 ) | ( ~n3165 & n3166 ) ;
  assign n3168 = ~n3166 & n3167 ;
  assign n3169 = n3165 | n3167 ;
  assign n3170 = ( ~x23 & n3168 ) | ( ~x23 & n3169 ) | ( n3168 & n3169 ) ;
  assign n3171 = n3159 & n3170 ;
  assign n3172 = n3159 | n3170 ;
  assign n3173 = ~n3171 & n3172 ;
  assign n3174 = n3127 & n3173 ;
  assign n3175 = n3127 | n3173 ;
  assign n3176 = ~n3174 & n3175 ;
  assign n3177 = x76 & n1421 ;
  assign n3178 = x75 & n1416 ;
  assign n3179 = x74 & ~n1415 ;
  assign n3180 = n1584 & n3179 ;
  assign n3181 = n3178 | n3180 ;
  assign n3182 = n3177 | n3181 ;
  assign n3183 = n1424 | n3182 ;
  assign n3184 = ( n740 & n3182 ) | ( n740 & n3183 ) | ( n3182 & n3183 ) ;
  assign n3185 = x20 & n3184 ;
  assign n3186 = x20 & ~n3185 ;
  assign n3187 = ( n3184 & ~n3185 ) | ( n3184 & n3186 ) | ( ~n3185 & n3186 ) ;
  assign n3188 = n3176 | n3187 ;
  assign n3189 = n3176 & n3187 ;
  assign n3190 = n3188 & ~n3189 ;
  assign n3191 = n3013 | n3016 ;
  assign n3192 = n3190 & n3191 ;
  assign n3193 = n3190 | n3191 ;
  assign n3194 = ~n3192 & n3193 ;
  assign n3195 = x79 & n1071 ;
  assign n3196 = x78 & n1066 ;
  assign n3197 = x77 & ~n1065 ;
  assign n3198 = n1189 & n3197 ;
  assign n3199 = n3196 | n3198 ;
  assign n3200 = n3195 | n3199 ;
  assign n3201 = n1074 | n3200 ;
  assign n3202 = ( n961 & n3200 ) | ( n961 & n3201 ) | ( n3200 & n3201 ) ;
  assign n3203 = x17 & n3202 ;
  assign n3204 = x17 & ~n3203 ;
  assign n3205 = ( n3202 & ~n3203 ) | ( n3202 & n3204 ) | ( ~n3203 & n3204 ) ;
  assign n3206 = n3194 & n3205 ;
  assign n3207 = n3194 & ~n3206 ;
  assign n3208 = ~n3194 & n3205 ;
  assign n3209 = n3207 | n3208 ;
  assign n3210 = n3030 | n3036 ;
  assign n3211 = n3209 | n3210 ;
  assign n3212 = n3209 & n3210 ;
  assign n3213 = n3211 & ~n3212 ;
  assign n3214 = x82 & n771 ;
  assign n3215 = x81 & n766 ;
  assign n3216 = x80 & ~n765 ;
  assign n3217 = n905 & n3216 ;
  assign n3218 = n3215 | n3217 ;
  assign n3219 = n3214 | n3218 ;
  assign n3220 = n774 | n3219 ;
  assign n3221 = ( n1371 & n3219 ) | ( n1371 & n3220 ) | ( n3219 & n3220 ) ;
  assign n3222 = x14 & n3221 ;
  assign n3223 = x14 & ~n3222 ;
  assign n3224 = ( n3221 & ~n3222 ) | ( n3221 & n3223 ) | ( ~n3222 & n3223 ) ;
  assign n3225 = n3213 & n3224 ;
  assign n3226 = n3213 & ~n3225 ;
  assign n3227 = ~n3213 & n3224 ;
  assign n3228 = n3226 | n3227 ;
  assign n3229 = n3049 | n3055 ;
  assign n3230 = n3228 | n3229 ;
  assign n3231 = n3228 & n3229 ;
  assign n3232 = n3230 & ~n3231 ;
  assign n3233 = ( n3070 & n3126 ) | ( n3070 & ~n3232 ) | ( n3126 & ~n3232 ) ;
  assign n3234 = ( ~n3070 & n3232 ) | ( ~n3070 & n3233 ) | ( n3232 & n3233 ) ;
  assign n3235 = ( ~n3126 & n3233 ) | ( ~n3126 & n3234 ) | ( n3233 & n3234 ) ;
  assign n3236 = n3115 & n3235 ;
  assign n3237 = n3115 | n3235 ;
  assign n3238 = ~n3236 & n3237 ;
  assign n3239 = n3087 | n3092 ;
  assign n3240 = n3238 | n3239 ;
  assign n3241 = n3238 & n3239 ;
  assign n3242 = n3240 & ~n3241 ;
  assign n3243 = x91 & n206 ;
  assign n3244 = x90 & n201 ;
  assign n3245 = x89 & ~n200 ;
  assign n3246 = n243 & n3245 ;
  assign n3247 = n3244 | n3246 ;
  assign n3248 = n3243 | n3247 ;
  assign n3249 = n209 | n3248 ;
  assign n3250 = ( n2714 & n3248 ) | ( n2714 & n3249 ) | ( n3248 & n3249 ) ;
  assign n3251 = x5 & n3250 ;
  assign n3252 = x5 & ~n3251 ;
  assign n3253 = ( n3250 & ~n3251 ) | ( n3250 & n3252 ) | ( ~n3251 & n3252 ) ;
  assign n3254 = n3242 & n3253 ;
  assign n3255 = n3242 & ~n3254 ;
  assign n3256 = ~n3242 & n3253 ;
  assign n3257 = n3255 | n3256 ;
  assign n3258 = n3096 | n3257 ;
  assign n3259 = n3096 & n3257 ;
  assign n3260 = n3258 & ~n3259 ;
  assign n3261 = x93 & n131 ;
  assign n3262 = x92 & ~n156 ;
  assign n3263 = ( n135 & n3261 ) | ( n135 & n3262 ) | ( n3261 & n3262 ) ;
  assign n3264 = x0 & x94 ;
  assign n3265 = ( ~n135 & n3261 ) | ( ~n135 & n3264 ) | ( n3261 & n3264 ) ;
  assign n3266 = n3263 | n3265 ;
  assign n3267 = n139 | n3266 ;
  assign n3268 = n2924 | n2930 ;
  assign n3269 = ( x93 & ~x94 ) | ( x93 & n3268 ) | ( ~x94 & n3268 ) ;
  assign n3270 = ( ~x93 & x94 ) | ( ~x93 & n3269 ) | ( x94 & n3269 ) ;
  assign n3271 = ( ~n3268 & n3269 ) | ( ~n3268 & n3270 ) | ( n3269 & n3270 ) ;
  assign n3272 = ( n3266 & n3267 ) | ( n3266 & n3271 ) | ( n3267 & n3271 ) ;
  assign n3273 = x2 & n3272 ;
  assign n3274 = x2 & ~n3273 ;
  assign n3275 = ( n3272 & ~n3273 ) | ( n3272 & n3274 ) | ( ~n3273 & n3274 ) ;
  assign n3276 = n3260 & n3275 ;
  assign n3277 = n3260 & ~n3276 ;
  assign n3278 = ~n3260 & n3275 ;
  assign n3279 = n3277 | n3278 ;
  assign n3280 = n3099 | n3102 ;
  assign n3281 = n3279 & n3280 ;
  assign n3282 = n3279 | n3280 ;
  assign n3283 = ~n3281 & n3282 ;
  assign n3284 = x71 & n2280 ;
  assign n3285 = x70 & n2275 ;
  assign n3286 = x69 & ~n2274 ;
  assign n3287 = n2481 & n3286 ;
  assign n3288 = n3285 | n3287 ;
  assign n3289 = n3284 | n3288 ;
  assign n3290 = n2283 | n3289 ;
  assign n3291 = ( n376 & n3289 ) | ( n376 & n3290 ) | ( n3289 & n3290 ) ;
  assign n3292 = x26 & ~n3291 ;
  assign n3293 = ~x26 & n3291 ;
  assign n3294 = n3292 | n3293 ;
  assign n3295 = n229 & n2778 ;
  assign n3296 = x68 & n2775 ;
  assign n3297 = x67 & n2770 ;
  assign n3298 = x66 & ~n2769 ;
  assign n3299 = n2978 & n3298 ;
  assign n3300 = n3297 | n3299 ;
  assign n3301 = n3296 | n3300 ;
  assign n3302 = n3295 | n3301 ;
  assign n3303 = x29 | n3302 ;
  assign n3304 = ~x29 & n3303 ;
  assign n3305 = ( ~n3302 & n3303 ) | ( ~n3302 & n3304 ) | ( n3303 & n3304 ) ;
  assign n3306 = ~x30 & x31 ;
  assign n3307 = x30 & ~x31 ;
  assign n3308 = n3306 | n3307 ;
  assign n3309 = ~n3141 & n3308 ;
  assign n3310 = x64 & n3309 ;
  assign n3311 = ~x31 & x32 ;
  assign n3312 = x31 & ~x32 ;
  assign n3313 = n3311 | n3312 ;
  assign n3314 = n3141 & ~n3313 ;
  assign n3315 = x65 & n3314 ;
  assign n3316 = n3310 | n3315 ;
  assign n3317 = n3141 & n3313 ;
  assign n3318 = n142 & n3317 ;
  assign n3319 = n3316 | n3318 ;
  assign n3320 = x32 | n3319 ;
  assign n3321 = ~x32 & n3320 ;
  assign n3322 = ( ~n3319 & n3320 ) | ( ~n3319 & n3321 ) | ( n3320 & n3321 ) ;
  assign n3323 = x32 & ~n3142 ;
  assign n3324 = n3322 & n3323 ;
  assign n3325 = n3322 | n3323 ;
  assign n3326 = ~n3324 & n3325 ;
  assign n3327 = ( n3154 & n3305 ) | ( n3154 & n3326 ) | ( n3305 & n3326 ) ;
  assign n3328 = ( n3154 & n3326 ) | ( n3154 & ~n3327 ) | ( n3326 & ~n3327 ) ;
  assign n3329 = ( n3305 & ~n3327 ) | ( n3305 & n3328 ) | ( ~n3327 & n3328 ) ;
  assign n3330 = n3294 & n3329 ;
  assign n3331 = n3294 | n3329 ;
  assign n3332 = ~n3330 & n3331 ;
  assign n3333 = ( n2991 & n3138 ) | ( n2991 & n3156 ) | ( n3138 & n3156 ) ;
  assign n3334 = n3332 | n3333 ;
  assign n3335 = n3332 & n3333 ;
  assign n3336 = n3334 & ~n3335 ;
  assign n3337 = x74 & n1817 ;
  assign n3338 = x73 & n1812 ;
  assign n3339 = x72 & ~n1811 ;
  assign n3340 = n1977 & n3339 ;
  assign n3341 = n3338 | n3340 ;
  assign n3342 = n3337 | n3341 ;
  assign n3343 = n1820 | n3342 ;
  assign n3344 = ( n587 & n3342 ) | ( n587 & n3343 ) | ( n3342 & n3343 ) ;
  assign n3345 = x23 & n3344 ;
  assign n3346 = x23 & ~n3345 ;
  assign n3347 = ( n3344 & ~n3345 ) | ( n3344 & n3346 ) | ( ~n3345 & n3346 ) ;
  assign n3348 = n3336 & n3347 ;
  assign n3349 = n3336 & ~n3348 ;
  assign n3350 = ~n3336 & n3347 ;
  assign n3351 = n3349 | n3350 ;
  assign n3352 = n3171 | n3174 ;
  assign n3353 = n3351 | n3352 ;
  assign n3354 = n3351 & n3352 ;
  assign n3355 = n3353 & ~n3354 ;
  assign n3356 = x77 & n1421 ;
  assign n3357 = x76 & n1416 ;
  assign n3358 = x75 & ~n1415 ;
  assign n3359 = n1584 & n3358 ;
  assign n3360 = n3357 | n3359 ;
  assign n3361 = n3356 | n3360 ;
  assign n3362 = n1424 | n3361 ;
  assign n3363 = ( n846 & n3361 ) | ( n846 & n3362 ) | ( n3361 & n3362 ) ;
  assign n3364 = x20 & n3363 ;
  assign n3365 = x20 & ~n3364 ;
  assign n3366 = ( n3363 & ~n3364 ) | ( n3363 & n3365 ) | ( ~n3364 & n3365 ) ;
  assign n3367 = n3355 | n3366 ;
  assign n3368 = n3355 & n3366 ;
  assign n3369 = n3367 & ~n3368 ;
  assign n3370 = n3189 | n3192 ;
  assign n3371 = n3369 & n3370 ;
  assign n3372 = n3369 | n3370 ;
  assign n3373 = ~n3371 & n3372 ;
  assign n3374 = x80 & n1071 ;
  assign n3375 = x79 & n1066 ;
  assign n3376 = x78 & ~n1065 ;
  assign n3377 = n1189 & n3376 ;
  assign n3378 = n3375 | n3377 ;
  assign n3379 = n3374 | n3378 ;
  assign n3380 = n1074 | n3379 ;
  assign n3381 = ( n1147 & n3379 ) | ( n1147 & n3380 ) | ( n3379 & n3380 ) ;
  assign n3382 = x17 & n3381 ;
  assign n3383 = x17 & ~n3382 ;
  assign n3384 = ( n3381 & ~n3382 ) | ( n3381 & n3383 ) | ( ~n3382 & n3383 ) ;
  assign n3385 = n3373 & n3384 ;
  assign n3386 = n3373 & ~n3385 ;
  assign n3387 = ~n3373 & n3384 ;
  assign n3388 = n3386 | n3387 ;
  assign n3389 = n3206 | n3212 ;
  assign n3390 = n3388 | n3389 ;
  assign n3391 = n3388 & n3389 ;
  assign n3392 = n3390 & ~n3391 ;
  assign n3393 = x83 & n771 ;
  assign n3394 = x82 & n766 ;
  assign n3395 = x81 & ~n765 ;
  assign n3396 = n905 & n3395 ;
  assign n3397 = n3394 | n3396 ;
  assign n3398 = n3393 | n3397 ;
  assign n3399 = n774 | n3398 ;
  assign n3400 = ( n1510 & n3398 ) | ( n1510 & n3399 ) | ( n3398 & n3399 ) ;
  assign n3401 = x14 & n3400 ;
  assign n3402 = x14 & ~n3401 ;
  assign n3403 = ( n3400 & ~n3401 ) | ( n3400 & n3402 ) | ( ~n3401 & n3402 ) ;
  assign n3404 = n3392 & n3403 ;
  assign n3405 = n3392 & ~n3404 ;
  assign n3406 = ~n3392 & n3403 ;
  assign n3407 = n3405 | n3406 ;
  assign n3408 = n3225 | n3231 ;
  assign n3409 = n3407 | n3408 ;
  assign n3410 = n3407 & n3408 ;
  assign n3411 = n3409 & ~n3410 ;
  assign n3412 = x86 & n528 ;
  assign n3413 = x85 & n523 ;
  assign n3414 = x84 & ~n522 ;
  assign n3415 = n635 & n3414 ;
  assign n3416 = n3413 | n3415 ;
  assign n3417 = n3412 | n3416 ;
  assign n3418 = n531 | n3417 ;
  assign n3419 = ( n1921 & n3417 ) | ( n1921 & n3418 ) | ( n3417 & n3418 ) ;
  assign n3420 = x11 & n3419 ;
  assign n3421 = x11 & ~n3420 ;
  assign n3422 = ( n3419 & ~n3420 ) | ( n3419 & n3421 ) | ( ~n3420 & n3421 ) ;
  assign n3423 = n3411 & n3422 ;
  assign n3424 = n3411 & ~n3423 ;
  assign n3425 = ~n3411 & n3422 ;
  assign n3426 = n3424 | n3425 ;
  assign n3427 = ( n3070 & n3126 ) | ( n3070 & n3232 ) | ( n3126 & n3232 ) ;
  assign n3428 = n3426 | n3427 ;
  assign n3429 = n3426 & n3427 ;
  assign n3430 = n3428 & ~n3429 ;
  assign n3431 = x89 & n337 ;
  assign n3432 = x88 & n332 ;
  assign n3433 = x87 & ~n331 ;
  assign n3434 = n396 & n3433 ;
  assign n3435 = n3432 | n3434 ;
  assign n3436 = n3431 | n3435 ;
  assign n3437 = n340 | n3436 ;
  assign n3438 = ( n2244 & n3436 ) | ( n2244 & n3437 ) | ( n3436 & n3437 ) ;
  assign n3439 = x8 & n3438 ;
  assign n3440 = x8 & ~n3439 ;
  assign n3441 = ( n3438 & ~n3439 ) | ( n3438 & n3440 ) | ( ~n3439 & n3440 ) ;
  assign n3442 = n3430 & n3441 ;
  assign n3443 = n3430 & ~n3442 ;
  assign n3444 = ~n3430 & n3441 ;
  assign n3445 = n3443 | n3444 ;
  assign n3446 = n3236 | n3241 ;
  assign n3447 = n3445 | n3446 ;
  assign n3448 = n3445 & n3446 ;
  assign n3449 = n3447 & ~n3448 ;
  assign n3450 = x92 & n206 ;
  assign n3451 = x91 & n201 ;
  assign n3452 = x90 & ~n200 ;
  assign n3453 = n243 & n3452 ;
  assign n3454 = n3451 | n3453 ;
  assign n3455 = n3450 | n3454 ;
  assign n3456 = n209 | n3455 ;
  assign n3457 = ( n2904 & n3455 ) | ( n2904 & n3456 ) | ( n3455 & n3456 ) ;
  assign n3458 = x5 & n3457 ;
  assign n3459 = x5 & ~n3458 ;
  assign n3460 = ( n3457 & ~n3458 ) | ( n3457 & n3459 ) | ( ~n3458 & n3459 ) ;
  assign n3461 = n3449 & n3460 ;
  assign n3462 = n3449 & ~n3461 ;
  assign n3463 = ~n3449 & n3460 ;
  assign n3464 = n3462 | n3463 ;
  assign n3465 = n3254 | n3259 ;
  assign n3466 = n3464 | n3465 ;
  assign n3467 = n3464 & n3465 ;
  assign n3468 = n3466 & ~n3467 ;
  assign n3469 = x93 | x94 ;
  assign n3470 = x94 | x95 ;
  assign n3471 = x94 & x95 ;
  assign n3472 = n3470 & ~n3471 ;
  assign n3473 = n3469 & n3472 ;
  assign n3474 = x93 & x94 ;
  assign n3475 = n3472 & n3474 ;
  assign n3476 = ( n3268 & n3473 ) | ( n3268 & n3475 ) | ( n3473 & n3475 ) ;
  assign n3477 = ( n3268 & n3469 ) | ( n3268 & n3474 ) | ( n3469 & n3474 ) ;
  assign n3478 = n3472 | n3477 ;
  assign n3479 = ~n3476 & n3478 ;
  assign n3480 = x94 & n131 ;
  assign n3481 = x93 & ~n156 ;
  assign n3482 = ( n135 & n3480 ) | ( n135 & n3481 ) | ( n3480 & n3481 ) ;
  assign n3483 = x0 & x95 ;
  assign n3484 = ( ~n135 & n3480 ) | ( ~n135 & n3483 ) | ( n3480 & n3483 ) ;
  assign n3485 = n3482 | n3484 ;
  assign n3486 = n139 | n3485 ;
  assign n3487 = ( n3479 & n3485 ) | ( n3479 & n3486 ) | ( n3485 & n3486 ) ;
  assign n3488 = x2 & n3487 ;
  assign n3489 = x2 & ~n3488 ;
  assign n3490 = ( n3487 & ~n3488 ) | ( n3487 & n3489 ) | ( ~n3488 & n3489 ) ;
  assign n3491 = n3468 & n3490 ;
  assign n3492 = n3468 & ~n3491 ;
  assign n3493 = ~n3468 & n3490 ;
  assign n3494 = n3492 | n3493 ;
  assign n3495 = n3276 | n3281 ;
  assign n3496 = n3494 & n3495 ;
  assign n3497 = n3494 | n3495 ;
  assign n3498 = ~n3496 & n3497 ;
  assign n3499 = x95 | x96 ;
  assign n3500 = x95 & x96 ;
  assign n3501 = n3499 & ~n3500 ;
  assign n3502 = n3471 | n3473 ;
  assign n3503 = n3501 & n3502 ;
  assign n3504 = n3471 | n3475 ;
  assign n3505 = n3501 & n3504 ;
  assign n3506 = ( n3268 & n3503 ) | ( n3268 & n3505 ) | ( n3503 & n3505 ) ;
  assign n3507 = ( n3268 & n3502 ) | ( n3268 & n3504 ) | ( n3502 & n3504 ) ;
  assign n3508 = n3501 | n3507 ;
  assign n3509 = ~n3506 & n3508 ;
  assign n3510 = x95 & n131 ;
  assign n3511 = x94 & ~n156 ;
  assign n3512 = ( n135 & n3510 ) | ( n135 & n3511 ) | ( n3510 & n3511 ) ;
  assign n3513 = x0 & x96 ;
  assign n3514 = ( ~n135 & n3510 ) | ( ~n135 & n3513 ) | ( n3510 & n3513 ) ;
  assign n3515 = n3512 | n3514 ;
  assign n3516 = n139 | n3515 ;
  assign n3517 = ( n3509 & n3515 ) | ( n3509 & n3516 ) | ( n3515 & n3516 ) ;
  assign n3518 = x2 & n3517 ;
  assign n3519 = x2 & ~n3518 ;
  assign n3520 = ( n3517 & ~n3518 ) | ( n3517 & n3519 ) | ( ~n3518 & n3519 ) ;
  assign n3521 = n3491 | n3496 ;
  assign n3522 = x87 & n528 ;
  assign n3523 = x86 & n523 ;
  assign n3524 = x85 & ~n522 ;
  assign n3525 = n635 & n3524 ;
  assign n3526 = n3523 | n3525 ;
  assign n3527 = n3522 | n3526 ;
  assign n3528 = n531 | n3527 ;
  assign n3529 = ( n2067 & n3527 ) | ( n2067 & n3528 ) | ( n3527 & n3528 ) ;
  assign n3530 = x11 & n3529 ;
  assign n3531 = x11 & ~n3530 ;
  assign n3532 = ( n3529 & ~n3530 ) | ( n3529 & n3531 ) | ( ~n3530 & n3531 ) ;
  assign n3533 = x84 & n771 ;
  assign n3534 = x83 & n766 ;
  assign n3535 = x82 & ~n765 ;
  assign n3536 = n905 & n3535 ;
  assign n3537 = n3534 | n3536 ;
  assign n3538 = n3533 | n3537 ;
  assign n3539 = n774 | n3538 ;
  assign n3540 = ( n1537 & n3538 ) | ( n1537 & n3539 ) | ( n3538 & n3539 ) ;
  assign n3541 = x14 & n3540 ;
  assign n3542 = x14 & ~n3541 ;
  assign n3543 = ( n3540 & ~n3541 ) | ( n3540 & n3542 ) | ( ~n3541 & n3542 ) ;
  assign n3544 = n3368 | n3371 ;
  assign n3545 = n3330 | n3335 ;
  assign n3546 = x72 & n2280 ;
  assign n3547 = x71 & n2275 ;
  assign n3548 = x70 & ~n2274 ;
  assign n3549 = n2481 & n3548 ;
  assign n3550 = n3547 | n3549 ;
  assign n3551 = n3546 | n3550 ;
  assign n3552 = ( n435 & n2283 ) | ( n435 & n3551 ) | ( n2283 & n3551 ) ;
  assign n3553 = ( x26 & ~n3551 ) | ( x26 & n3552 ) | ( ~n3551 & n3552 ) ;
  assign n3554 = ~n3552 & n3553 ;
  assign n3555 = n3551 | n3553 ;
  assign n3556 = ( ~x26 & n3554 ) | ( ~x26 & n3555 ) | ( n3554 & n3555 ) ;
  assign n3557 = n264 & n2778 ;
  assign n3558 = x69 & n2775 ;
  assign n3559 = x68 & n2770 ;
  assign n3560 = x67 & ~n2769 ;
  assign n3561 = n2978 & n3560 ;
  assign n3562 = n3559 | n3561 ;
  assign n3563 = n3558 | n3562 ;
  assign n3564 = n3557 | n3563 ;
  assign n3565 = x29 | n3564 ;
  assign n3566 = ~x29 & n3565 ;
  assign n3567 = ( ~n3564 & n3565 ) | ( ~n3564 & n3566 ) | ( n3565 & n3566 ) ;
  assign n3568 = x66 & n3314 ;
  assign n3569 = x65 & n3309 ;
  assign n3570 = ~n3141 & n3313 ;
  assign n3571 = x64 & ~n3308 ;
  assign n3572 = n3570 & n3571 ;
  assign n3573 = n3569 | n3572 ;
  assign n3574 = n3568 | n3573 ;
  assign n3575 = n153 & n3317 ;
  assign n3576 = n3574 | n3575 ;
  assign n3577 = x32 | n3576 ;
  assign n3578 = ~x32 & n3577 ;
  assign n3579 = ( ~n3576 & n3577 ) | ( ~n3576 & n3578 ) | ( n3577 & n3578 ) ;
  assign n3580 = n3324 | n3579 ;
  assign n3581 = n3324 & n3579 ;
  assign n3582 = n3580 & ~n3581 ;
  assign n3583 = ( n3327 & n3567 ) | ( n3327 & n3582 ) | ( n3567 & n3582 ) ;
  assign n3584 = ( n3327 & n3582 ) | ( n3327 & ~n3583 ) | ( n3582 & ~n3583 ) ;
  assign n3585 = ( n3567 & ~n3583 ) | ( n3567 & n3584 ) | ( ~n3583 & n3584 ) ;
  assign n3586 = n3556 & n3585 ;
  assign n3587 = n3585 & ~n3586 ;
  assign n3588 = ( n3556 & ~n3586 ) | ( n3556 & n3587 ) | ( ~n3586 & n3587 ) ;
  assign n3589 = n3545 | n3588 ;
  assign n3590 = n3545 & n3588 ;
  assign n3591 = n3589 & ~n3590 ;
  assign n3592 = x75 & n1817 ;
  assign n3593 = x74 & n1812 ;
  assign n3594 = x73 & ~n1811 ;
  assign n3595 = n1977 & n3594 ;
  assign n3596 = n3593 | n3595 ;
  assign n3597 = n3592 | n3596 ;
  assign n3598 = n1820 | n3597 ;
  assign n3599 = ( n609 & n3597 ) | ( n609 & n3598 ) | ( n3597 & n3598 ) ;
  assign n3600 = x23 & n3599 ;
  assign n3601 = x23 & ~n3600 ;
  assign n3602 = ( n3599 & ~n3600 ) | ( n3599 & n3601 ) | ( ~n3600 & n3601 ) ;
  assign n3603 = n3591 & n3602 ;
  assign n3604 = n3591 | n3602 ;
  assign n3605 = ~n3603 & n3604 ;
  assign n3606 = n3348 | n3354 ;
  assign n3607 = n3605 & n3606 ;
  assign n3608 = n3606 & ~n3607 ;
  assign n3609 = ( n3605 & ~n3607 ) | ( n3605 & n3608 ) | ( ~n3607 & n3608 ) ;
  assign n3610 = x78 & n1421 ;
  assign n3611 = x77 & n1416 ;
  assign n3612 = x76 & ~n1415 ;
  assign n3613 = n1584 & n3612 ;
  assign n3614 = n3611 | n3613 ;
  assign n3615 = n3610 | n3614 ;
  assign n3616 = n1424 | n3615 ;
  assign n3617 = ( n868 & n3615 ) | ( n868 & n3616 ) | ( n3615 & n3616 ) ;
  assign n3618 = x20 & n3617 ;
  assign n3619 = x20 & ~n3618 ;
  assign n3620 = ( n3617 & ~n3618 ) | ( n3617 & n3619 ) | ( ~n3618 & n3619 ) ;
  assign n3621 = n3609 | n3620 ;
  assign n3622 = n3609 & n3620 ;
  assign n3623 = n3621 & ~n3622 ;
  assign n3624 = n3544 & n3623 ;
  assign n3625 = n3544 | n3623 ;
  assign n3626 = ~n3624 & n3625 ;
  assign n3627 = x81 & n1071 ;
  assign n3628 = x80 & n1066 ;
  assign n3629 = x79 & ~n1065 ;
  assign n3630 = n1189 & n3629 ;
  assign n3631 = n3628 | n3630 ;
  assign n3632 = n3627 | n3631 ;
  assign n3633 = n1074 | n3632 ;
  assign n3634 = ( n1256 & n3632 ) | ( n1256 & n3633 ) | ( n3632 & n3633 ) ;
  assign n3635 = x17 & n3634 ;
  assign n3636 = x17 & ~n3635 ;
  assign n3637 = ( n3634 & ~n3635 ) | ( n3634 & n3636 ) | ( ~n3635 & n3636 ) ;
  assign n3638 = n3626 & n3637 ;
  assign n3639 = n3626 & ~n3638 ;
  assign n3640 = ~n3626 & n3637 ;
  assign n3641 = n3639 | n3640 ;
  assign n3642 = n3385 | n3391 ;
  assign n3643 = n3641 | n3642 ;
  assign n3644 = n3641 & n3642 ;
  assign n3645 = n3643 & ~n3644 ;
  assign n3646 = n3404 | n3410 ;
  assign n3647 = ( n3543 & n3645 ) | ( n3543 & n3646 ) | ( n3645 & n3646 ) ;
  assign n3648 = ( n3645 & n3646 ) | ( n3645 & ~n3647 ) | ( n3646 & ~n3647 ) ;
  assign n3649 = ( n3543 & ~n3647 ) | ( n3543 & n3648 ) | ( ~n3647 & n3648 ) ;
  assign n3650 = n3532 | n3649 ;
  assign n3651 = n3532 & n3649 ;
  assign n3652 = n3650 & ~n3651 ;
  assign n3653 = n3423 | n3429 ;
  assign n3654 = n3652 & n3653 ;
  assign n3655 = n3652 | n3653 ;
  assign n3656 = ~n3654 & n3655 ;
  assign n3657 = x90 & n337 ;
  assign n3658 = x89 & n332 ;
  assign n3659 = x88 & ~n331 ;
  assign n3660 = n396 & n3659 ;
  assign n3661 = n3658 | n3660 ;
  assign n3662 = n3657 | n3661 ;
  assign n3663 = n340 | n3662 ;
  assign n3664 = ( n2410 & n3662 ) | ( n2410 & n3663 ) | ( n3662 & n3663 ) ;
  assign n3665 = x8 & n3664 ;
  assign n3666 = x8 & ~n3665 ;
  assign n3667 = ( n3664 & ~n3665 ) | ( n3664 & n3666 ) | ( ~n3665 & n3666 ) ;
  assign n3668 = n3656 & n3667 ;
  assign n3669 = n3656 & ~n3668 ;
  assign n3670 = ~n3656 & n3667 ;
  assign n3671 = n3669 | n3670 ;
  assign n3672 = n3442 | n3448 ;
  assign n3673 = n3671 | n3672 ;
  assign n3674 = n3671 & n3672 ;
  assign n3675 = n3673 & ~n3674 ;
  assign n3676 = x93 & n206 ;
  assign n3677 = x92 & n201 ;
  assign n3678 = x91 & ~n200 ;
  assign n3679 = n243 & n3678 ;
  assign n3680 = n3677 | n3679 ;
  assign n3681 = n3676 | n3680 ;
  assign n3682 = n209 | n3681 ;
  assign n3683 = ( n2931 & n3681 ) | ( n2931 & n3682 ) | ( n3681 & n3682 ) ;
  assign n3684 = x5 & n3683 ;
  assign n3685 = x5 & ~n3684 ;
  assign n3686 = ( n3683 & ~n3684 ) | ( n3683 & n3685 ) | ( ~n3684 & n3685 ) ;
  assign n3687 = n3675 & n3686 ;
  assign n3688 = n3675 | n3686 ;
  assign n3689 = ~n3687 & n3688 ;
  assign n3690 = n3461 | n3467 ;
  assign n3691 = n3689 | n3690 ;
  assign n3692 = ( n3461 & n3467 ) | ( n3461 & n3689 ) | ( n3467 & n3689 ) ;
  assign n3693 = n3691 & ~n3692 ;
  assign n3694 = ( n3520 & n3521 ) | ( n3520 & ~n3693 ) | ( n3521 & ~n3693 ) ;
  assign n3695 = ( ~n3521 & n3693 ) | ( ~n3521 & n3694 ) | ( n3693 & n3694 ) ;
  assign n3696 = ( ~n3520 & n3694 ) | ( ~n3520 & n3695 ) | ( n3694 & n3695 ) ;
  assign n3697 = x96 | x97 ;
  assign n3698 = x96 & x97 ;
  assign n3699 = n3697 & ~n3698 ;
  assign n3700 = n3500 | n3503 ;
  assign n3701 = n3699 & n3700 ;
  assign n3702 = n3500 | n3505 ;
  assign n3703 = n3699 & n3702 ;
  assign n3704 = ( n3268 & n3701 ) | ( n3268 & n3703 ) | ( n3701 & n3703 ) ;
  assign n3705 = ( n3268 & n3700 ) | ( n3268 & n3702 ) | ( n3700 & n3702 ) ;
  assign n3706 = n3699 | n3705 ;
  assign n3707 = ~n3704 & n3706 ;
  assign n3708 = x96 & n131 ;
  assign n3709 = x95 & ~n156 ;
  assign n3710 = ( n135 & n3708 ) | ( n135 & n3709 ) | ( n3708 & n3709 ) ;
  assign n3711 = x0 & x97 ;
  assign n3712 = ( ~n135 & n3708 ) | ( ~n135 & n3711 ) | ( n3708 & n3711 ) ;
  assign n3713 = n3710 | n3712 ;
  assign n3714 = n139 | n3713 ;
  assign n3715 = ( n3707 & n3713 ) | ( n3707 & n3714 ) | ( n3713 & n3714 ) ;
  assign n3716 = x2 & n3715 ;
  assign n3717 = x2 & ~n3716 ;
  assign n3718 = ( n3715 & ~n3716 ) | ( n3715 & n3717 ) | ( ~n3716 & n3717 ) ;
  assign n3719 = x94 & n206 ;
  assign n3720 = x93 & n201 ;
  assign n3721 = x92 & ~n200 ;
  assign n3722 = n243 & n3721 ;
  assign n3723 = n3720 | n3722 ;
  assign n3724 = n3719 | n3723 ;
  assign n3725 = n209 | n3724 ;
  assign n3726 = ( n3271 & n3724 ) | ( n3271 & n3725 ) | ( n3724 & n3725 ) ;
  assign n3727 = x5 & n3726 ;
  assign n3728 = x5 & ~n3727 ;
  assign n3729 = ( n3726 & ~n3727 ) | ( n3726 & n3728 ) | ( ~n3727 & n3728 ) ;
  assign n3730 = n3687 | n3692 ;
  assign n3731 = n3651 | n3654 ;
  assign n3732 = x88 & n528 ;
  assign n3733 = x87 & n523 ;
  assign n3734 = x86 & ~n522 ;
  assign n3735 = n635 & n3734 ;
  assign n3736 = n3733 | n3735 ;
  assign n3737 = n3732 | n3736 ;
  assign n3738 = n531 | n3737 ;
  assign n3739 = ( n2095 & n3737 ) | ( n2095 & n3738 ) | ( n3737 & n3738 ) ;
  assign n3740 = x11 & n3739 ;
  assign n3741 = x11 & ~n3740 ;
  assign n3742 = ( n3739 & ~n3740 ) | ( n3739 & n3741 ) | ( ~n3740 & n3741 ) ;
  assign n3743 = x85 & n771 ;
  assign n3744 = x84 & n766 ;
  assign n3745 = x83 & ~n765 ;
  assign n3746 = n905 & n3745 ;
  assign n3747 = n3744 | n3746 ;
  assign n3748 = n3743 | n3747 ;
  assign n3749 = n774 | n3748 ;
  assign n3750 = ( n1765 & n3748 ) | ( n1765 & n3749 ) | ( n3748 & n3749 ) ;
  assign n3751 = x14 & n3750 ;
  assign n3752 = x14 & ~n3751 ;
  assign n3753 = ( n3750 & ~n3751 ) | ( n3750 & n3752 ) | ( ~n3751 & n3752 ) ;
  assign n3754 = n3638 | n3644 ;
  assign n3755 = x82 & n1071 ;
  assign n3756 = x81 & n1066 ;
  assign n3757 = x80 & ~n1065 ;
  assign n3758 = n1189 & n3757 ;
  assign n3759 = n3756 | n3758 ;
  assign n3760 = n3755 | n3759 ;
  assign n3761 = n1074 | n3760 ;
  assign n3762 = ( n1371 & n3760 ) | ( n1371 & n3761 ) | ( n3760 & n3761 ) ;
  assign n3763 = x17 & n3762 ;
  assign n3764 = x17 & ~n3763 ;
  assign n3765 = ( n3762 & ~n3763 ) | ( n3762 & n3764 ) | ( ~n3763 & n3764 ) ;
  assign n3766 = x79 & n1421 ;
  assign n3767 = x78 & n1416 ;
  assign n3768 = x77 & ~n1415 ;
  assign n3769 = n1584 & n3768 ;
  assign n3770 = n3767 | n3769 ;
  assign n3771 = n3766 | n3770 ;
  assign n3772 = n1424 | n3771 ;
  assign n3773 = ( n961 & n3771 ) | ( n961 & n3772 ) | ( n3771 & n3772 ) ;
  assign n3774 = x20 & n3773 ;
  assign n3775 = x20 & ~n3774 ;
  assign n3776 = ( n3773 & ~n3774 ) | ( n3773 & n3775 ) | ( ~n3774 & n3775 ) ;
  assign n3777 = n3622 | n3624 ;
  assign n3778 = n3603 | n3607 ;
  assign n3779 = x70 & n2775 ;
  assign n3780 = x69 & n2770 ;
  assign n3781 = x68 & ~n2769 ;
  assign n3782 = n2978 & n3781 ;
  assign n3783 = n3780 | n3782 ;
  assign n3784 = n3779 | n3783 ;
  assign n3785 = n2778 | n3784 ;
  assign n3786 = ( n310 & n3784 ) | ( n310 & n3785 ) | ( n3784 & n3785 ) ;
  assign n3787 = x29 & ~n3786 ;
  assign n3788 = ~x29 & n3786 ;
  assign n3789 = n3787 | n3788 ;
  assign n3790 = x32 & ~x33 ;
  assign n3791 = ~x32 & x33 ;
  assign n3792 = n3790 | n3791 ;
  assign n3793 = x64 & n3792 ;
  assign n3794 = x67 & n3314 ;
  assign n3795 = x66 & n3309 ;
  assign n3796 = x65 & ~n3308 ;
  assign n3797 = n3570 & n3796 ;
  assign n3798 = n3795 | n3797 ;
  assign n3799 = n3794 | n3798 ;
  assign n3800 = n180 & n3317 ;
  assign n3801 = n3799 | n3800 ;
  assign n3802 = x32 & ~n3801 ;
  assign n3803 = ~x32 & n3801 ;
  assign n3804 = n3802 | n3803 ;
  assign n3805 = ( n3581 & n3793 ) | ( n3581 & n3804 ) | ( n3793 & n3804 ) ;
  assign n3806 = ( n3581 & n3804 ) | ( n3581 & ~n3805 ) | ( n3804 & ~n3805 ) ;
  assign n3807 = ( n3793 & ~n3805 ) | ( n3793 & n3806 ) | ( ~n3805 & n3806 ) ;
  assign n3808 = ( n3583 & n3789 ) | ( n3583 & ~n3807 ) | ( n3789 & ~n3807 ) ;
  assign n3809 = ( ~n3583 & n3807 ) | ( ~n3583 & n3808 ) | ( n3807 & n3808 ) ;
  assign n3810 = ( ~n3789 & n3808 ) | ( ~n3789 & n3809 ) | ( n3808 & n3809 ) ;
  assign n3811 = x73 & n2280 ;
  assign n3812 = x72 & n2275 ;
  assign n3813 = x71 & ~n2274 ;
  assign n3814 = n2481 & n3813 ;
  assign n3815 = n3812 | n3814 ;
  assign n3816 = n3811 | n3815 ;
  assign n3817 = ( n499 & n2283 ) | ( n499 & n3816 ) | ( n2283 & n3816 ) ;
  assign n3818 = ( x26 & ~n3816 ) | ( x26 & n3817 ) | ( ~n3816 & n3817 ) ;
  assign n3819 = ~n3817 & n3818 ;
  assign n3820 = n3816 | n3818 ;
  assign n3821 = ( ~x26 & n3819 ) | ( ~x26 & n3820 ) | ( n3819 & n3820 ) ;
  assign n3822 = n3810 & n3821 ;
  assign n3823 = n3810 | n3821 ;
  assign n3824 = ~n3822 & n3823 ;
  assign n3825 = n3586 | n3590 ;
  assign n3826 = n3824 | n3825 ;
  assign n3827 = n3824 & n3825 ;
  assign n3828 = n3826 & ~n3827 ;
  assign n3829 = x76 & n1817 ;
  assign n3830 = x75 & n1812 ;
  assign n3831 = x74 & ~n1811 ;
  assign n3832 = n1977 & n3831 ;
  assign n3833 = n3830 | n3832 ;
  assign n3834 = n3829 | n3833 ;
  assign n3835 = n1820 | n3834 ;
  assign n3836 = ( n740 & n3834 ) | ( n740 & n3835 ) | ( n3834 & n3835 ) ;
  assign n3837 = x23 & n3836 ;
  assign n3838 = x23 & ~n3837 ;
  assign n3839 = ( n3836 & ~n3837 ) | ( n3836 & n3838 ) | ( ~n3837 & n3838 ) ;
  assign n3840 = n3828 | n3839 ;
  assign n3841 = n3828 & n3839 ;
  assign n3842 = n3840 & ~n3841 ;
  assign n3843 = n3778 & n3842 ;
  assign n3844 = n3778 | n3842 ;
  assign n3845 = ~n3843 & n3844 ;
  assign n3846 = ( n3776 & n3777 ) | ( n3776 & ~n3845 ) | ( n3777 & ~n3845 ) ;
  assign n3847 = ( ~n3777 & n3845 ) | ( ~n3777 & n3846 ) | ( n3845 & n3846 ) ;
  assign n3848 = ( ~n3776 & n3846 ) | ( ~n3776 & n3847 ) | ( n3846 & n3847 ) ;
  assign n3849 = n3765 & n3848 ;
  assign n3850 = n3765 | n3848 ;
  assign n3851 = ~n3849 & n3850 ;
  assign n3852 = n3754 | n3851 ;
  assign n3853 = n3754 & n3851 ;
  assign n3854 = n3852 & ~n3853 ;
  assign n3855 = ( n3647 & n3753 ) | ( n3647 & ~n3854 ) | ( n3753 & ~n3854 ) ;
  assign n3856 = ( ~n3647 & n3854 ) | ( ~n3647 & n3855 ) | ( n3854 & n3855 ) ;
  assign n3857 = ( ~n3753 & n3855 ) | ( ~n3753 & n3856 ) | ( n3855 & n3856 ) ;
  assign n3858 = n3742 | n3857 ;
  assign n3859 = n3742 & n3857 ;
  assign n3860 = n3858 & ~n3859 ;
  assign n3861 = n3731 & n3860 ;
  assign n3862 = n3731 | n3860 ;
  assign n3863 = ~n3861 & n3862 ;
  assign n3864 = x91 & n337 ;
  assign n3865 = x90 & n332 ;
  assign n3866 = x89 & ~n331 ;
  assign n3867 = n396 & n3866 ;
  assign n3868 = n3865 | n3867 ;
  assign n3869 = n3864 | n3868 ;
  assign n3870 = n340 | n3869 ;
  assign n3871 = ( n2714 & n3869 ) | ( n2714 & n3870 ) | ( n3869 & n3870 ) ;
  assign n3872 = x8 & n3871 ;
  assign n3873 = x8 & ~n3872 ;
  assign n3874 = ( n3871 & ~n3872 ) | ( n3871 & n3873 ) | ( ~n3872 & n3873 ) ;
  assign n3875 = n3863 & n3874 ;
  assign n3876 = n3863 & ~n3875 ;
  assign n3877 = ~n3863 & n3874 ;
  assign n3878 = n3876 | n3877 ;
  assign n3879 = n3668 | n3674 ;
  assign n3880 = n3878 | n3879 ;
  assign n3881 = n3878 & n3879 ;
  assign n3882 = n3880 & ~n3881 ;
  assign n3883 = ( n3729 & n3730 ) | ( n3729 & ~n3882 ) | ( n3730 & ~n3882 ) ;
  assign n3884 = ( ~n3730 & n3882 ) | ( ~n3730 & n3883 ) | ( n3882 & n3883 ) ;
  assign n3885 = ( ~n3729 & n3883 ) | ( ~n3729 & n3884 ) | ( n3883 & n3884 ) ;
  assign n3886 = n3718 & n3885 ;
  assign n3887 = n3718 | n3885 ;
  assign n3888 = ~n3886 & n3887 ;
  assign n3889 = ( n3520 & n3521 ) | ( n3520 & n3693 ) | ( n3521 & n3693 ) ;
  assign n3890 = n3888 | n3889 ;
  assign n3891 = n3888 & n3889 ;
  assign n3892 = n3890 & ~n3891 ;
  assign n3893 = ( n3729 & n3730 ) | ( n3729 & n3882 ) | ( n3730 & n3882 ) ;
  assign n3894 = x71 & n2775 ;
  assign n3895 = x70 & n2770 ;
  assign n3896 = x69 & ~n2769 ;
  assign n3897 = n2978 & n3896 ;
  assign n3898 = n3895 | n3897 ;
  assign n3899 = n3894 | n3898 ;
  assign n3900 = n2778 | n3899 ;
  assign n3901 = ( n376 & n3899 ) | ( n376 & n3900 ) | ( n3899 & n3900 ) ;
  assign n3902 = x29 & ~n3901 ;
  assign n3903 = ~x29 & n3901 ;
  assign n3904 = n3902 | n3903 ;
  assign n3905 = ~x33 & x34 ;
  assign n3906 = x33 & ~x34 ;
  assign n3907 = n3905 | n3906 ;
  assign n3908 = ~n3792 & n3907 ;
  assign n3909 = x64 & n3908 ;
  assign n3910 = ~x34 & x35 ;
  assign n3911 = x34 & ~x35 ;
  assign n3912 = n3910 | n3911 ;
  assign n3913 = n3792 & ~n3912 ;
  assign n3914 = x65 & n3913 ;
  assign n3915 = n3909 | n3914 ;
  assign n3916 = n3792 & n3912 ;
  assign n3917 = n142 & n3916 ;
  assign n3918 = n3915 | n3917 ;
  assign n3919 = x35 | n3918 ;
  assign n3920 = ~x35 & n3919 ;
  assign n3921 = ( ~n3918 & n3919 ) | ( ~n3918 & n3920 ) | ( n3919 & n3920 ) ;
  assign n3922 = x35 & ~n3793 ;
  assign n3923 = n3921 & n3922 ;
  assign n3924 = n3921 | n3922 ;
  assign n3925 = ~n3923 & n3924 ;
  assign n3926 = n229 & n3317 ;
  assign n3927 = x68 & n3314 ;
  assign n3928 = x67 & n3309 ;
  assign n3929 = x66 & ~n3308 ;
  assign n3930 = n3570 & n3929 ;
  assign n3931 = n3928 | n3930 ;
  assign n3932 = n3927 | n3931 ;
  assign n3933 = n3926 | n3932 ;
  assign n3934 = x32 | n3933 ;
  assign n3935 = ~x32 & n3934 ;
  assign n3936 = ( ~n3933 & n3934 ) | ( ~n3933 & n3935 ) | ( n3934 & n3935 ) ;
  assign n3937 = n3925 | n3936 ;
  assign n3938 = n3925 & n3936 ;
  assign n3939 = n3937 & ~n3938 ;
  assign n3940 = n3805 | n3939 ;
  assign n3941 = n3805 & n3939 ;
  assign n3942 = n3940 & ~n3941 ;
  assign n3943 = n3904 | n3942 ;
  assign n3944 = n3904 & n3942 ;
  assign n3945 = n3943 & ~n3944 ;
  assign n3946 = ( n3583 & n3789 ) | ( n3583 & n3807 ) | ( n3789 & n3807 ) ;
  assign n3947 = n3945 | n3946 ;
  assign n3948 = n3945 & n3946 ;
  assign n3949 = n3947 & ~n3948 ;
  assign n3950 = x74 & n2280 ;
  assign n3951 = x73 & n2275 ;
  assign n3952 = x72 & ~n2274 ;
  assign n3953 = n2481 & n3952 ;
  assign n3954 = n3951 | n3953 ;
  assign n3955 = n3950 | n3954 ;
  assign n3956 = n2283 | n3955 ;
  assign n3957 = ( n587 & n3955 ) | ( n587 & n3956 ) | ( n3955 & n3956 ) ;
  assign n3958 = x26 & n3957 ;
  assign n3959 = x26 & ~n3958 ;
  assign n3960 = ( n3957 & ~n3958 ) | ( n3957 & n3959 ) | ( ~n3958 & n3959 ) ;
  assign n3961 = n3949 & n3960 ;
  assign n3962 = n3949 & ~n3961 ;
  assign n3963 = ~n3949 & n3960 ;
  assign n3964 = n3962 | n3963 ;
  assign n3965 = n3822 | n3827 ;
  assign n3966 = n3964 | n3965 ;
  assign n3967 = n3964 & n3965 ;
  assign n3968 = n3966 & ~n3967 ;
  assign n3969 = x77 & n1817 ;
  assign n3970 = x76 & n1812 ;
  assign n3971 = x75 & ~n1811 ;
  assign n3972 = n1977 & n3971 ;
  assign n3973 = n3970 | n3972 ;
  assign n3974 = n3969 | n3973 ;
  assign n3975 = n1820 | n3974 ;
  assign n3976 = ( n846 & n3974 ) | ( n846 & n3975 ) | ( n3974 & n3975 ) ;
  assign n3977 = x23 & n3976 ;
  assign n3978 = x23 & ~n3977 ;
  assign n3979 = ( n3976 & ~n3977 ) | ( n3976 & n3978 ) | ( ~n3977 & n3978 ) ;
  assign n3980 = n3968 & n3979 ;
  assign n3981 = n3968 | n3979 ;
  assign n3982 = ~n3980 & n3981 ;
  assign n3983 = n3841 | n3843 ;
  assign n3984 = n3982 & n3983 ;
  assign n3985 = n3983 & ~n3984 ;
  assign n3986 = ( n3982 & ~n3984 ) | ( n3982 & n3985 ) | ( ~n3984 & n3985 ) ;
  assign n3987 = x80 & n1421 ;
  assign n3988 = x79 & n1416 ;
  assign n3989 = x78 & ~n1415 ;
  assign n3990 = n1584 & n3989 ;
  assign n3991 = n3988 | n3990 ;
  assign n3992 = n3987 | n3991 ;
  assign n3993 = n1424 | n3992 ;
  assign n3994 = ( n1147 & n3992 ) | ( n1147 & n3993 ) | ( n3992 & n3993 ) ;
  assign n3995 = x20 & n3994 ;
  assign n3996 = x20 & ~n3995 ;
  assign n3997 = ( n3994 & ~n3995 ) | ( n3994 & n3996 ) | ( ~n3995 & n3996 ) ;
  assign n3998 = n3986 & n3997 ;
  assign n3999 = n3986 & ~n3998 ;
  assign n4000 = ~n3986 & n3997 ;
  assign n4001 = n3999 | n4000 ;
  assign n4002 = ( n3776 & n3777 ) | ( n3776 & n3845 ) | ( n3777 & n3845 ) ;
  assign n4003 = n4001 | n4002 ;
  assign n4004 = n4001 & n4002 ;
  assign n4005 = n4003 & ~n4004 ;
  assign n4006 = x83 & n1071 ;
  assign n4007 = x82 & n1066 ;
  assign n4008 = x81 & ~n1065 ;
  assign n4009 = n1189 & n4008 ;
  assign n4010 = n4007 | n4009 ;
  assign n4011 = n4006 | n4010 ;
  assign n4012 = n1074 | n4011 ;
  assign n4013 = ( n1510 & n4011 ) | ( n1510 & n4012 ) | ( n4011 & n4012 ) ;
  assign n4014 = x17 & n4013 ;
  assign n4015 = x17 & ~n4014 ;
  assign n4016 = ( n4013 & ~n4014 ) | ( n4013 & n4015 ) | ( ~n4014 & n4015 ) ;
  assign n4017 = n4005 & n4016 ;
  assign n4018 = n4005 & ~n4017 ;
  assign n4019 = ~n4005 & n4016 ;
  assign n4020 = n4018 | n4019 ;
  assign n4021 = n3849 | n3853 ;
  assign n4022 = n4020 | n4021 ;
  assign n4023 = n4020 & n4021 ;
  assign n4024 = n4022 & ~n4023 ;
  assign n4025 = x86 & n771 ;
  assign n4026 = x85 & n766 ;
  assign n4027 = x84 & ~n765 ;
  assign n4028 = n905 & n4027 ;
  assign n4029 = n4026 | n4028 ;
  assign n4030 = n4025 | n4029 ;
  assign n4031 = n774 | n4030 ;
  assign n4032 = ( n1921 & n4030 ) | ( n1921 & n4031 ) | ( n4030 & n4031 ) ;
  assign n4033 = x14 & n4032 ;
  assign n4034 = x14 & ~n4033 ;
  assign n4035 = ( n4032 & ~n4033 ) | ( n4032 & n4034 ) | ( ~n4033 & n4034 ) ;
  assign n4036 = n4024 & n4035 ;
  assign n4037 = n4024 & ~n4036 ;
  assign n4038 = ~n4024 & n4035 ;
  assign n4039 = n4037 | n4038 ;
  assign n4040 = ( n3647 & n3753 ) | ( n3647 & n3854 ) | ( n3753 & n3854 ) ;
  assign n4041 = n4039 | n4040 ;
  assign n4042 = n4039 & n4040 ;
  assign n4043 = n4041 & ~n4042 ;
  assign n4044 = x89 & n528 ;
  assign n4045 = x88 & n523 ;
  assign n4046 = x87 & ~n522 ;
  assign n4047 = n635 & n4046 ;
  assign n4048 = n4045 | n4047 ;
  assign n4049 = n4044 | n4048 ;
  assign n4050 = n531 | n4049 ;
  assign n4051 = ( n2244 & n4049 ) | ( n2244 & n4050 ) | ( n4049 & n4050 ) ;
  assign n4052 = x11 & n4051 ;
  assign n4053 = x11 & ~n4052 ;
  assign n4054 = ( n4051 & ~n4052 ) | ( n4051 & n4053 ) | ( ~n4052 & n4053 ) ;
  assign n4055 = n4043 & n4054 ;
  assign n4056 = n4043 | n4054 ;
  assign n4057 = ~n4055 & n4056 ;
  assign n4058 = n3859 | n3861 ;
  assign n4059 = n4057 & n4058 ;
  assign n4060 = n4058 & ~n4059 ;
  assign n4061 = ( n4057 & ~n4059 ) | ( n4057 & n4060 ) | ( ~n4059 & n4060 ) ;
  assign n4062 = x92 & n337 ;
  assign n4063 = x91 & n332 ;
  assign n4064 = x90 & ~n331 ;
  assign n4065 = n396 & n4064 ;
  assign n4066 = n4063 | n4065 ;
  assign n4067 = n4062 | n4066 ;
  assign n4068 = n340 | n4067 ;
  assign n4069 = ( n2904 & n4067 ) | ( n2904 & n4068 ) | ( n4067 & n4068 ) ;
  assign n4070 = x8 & n4069 ;
  assign n4071 = x8 & ~n4070 ;
  assign n4072 = ( n4069 & ~n4070 ) | ( n4069 & n4071 ) | ( ~n4070 & n4071 ) ;
  assign n4073 = n4061 & n4072 ;
  assign n4074 = n4061 & ~n4073 ;
  assign n4075 = ~n4061 & n4072 ;
  assign n4076 = n4074 | n4075 ;
  assign n4077 = n3875 | n3881 ;
  assign n4078 = n4076 | n4077 ;
  assign n4079 = n4076 & n4077 ;
  assign n4080 = n4078 & ~n4079 ;
  assign n4081 = x95 & n206 ;
  assign n4082 = x94 & n201 ;
  assign n4083 = x93 & ~n200 ;
  assign n4084 = n243 & n4083 ;
  assign n4085 = n4082 | n4084 ;
  assign n4086 = n4081 | n4085 ;
  assign n4087 = n209 | n4086 ;
  assign n4088 = ( n3479 & n4086 ) | ( n3479 & n4087 ) | ( n4086 & n4087 ) ;
  assign n4089 = x5 & n4088 ;
  assign n4090 = x5 & ~n4089 ;
  assign n4091 = ( n4088 & ~n4089 ) | ( n4088 & n4090 ) | ( ~n4089 & n4090 ) ;
  assign n4092 = ( n3893 & n4080 ) | ( n3893 & ~n4091 ) | ( n4080 & ~n4091 ) ;
  assign n4093 = ( ~n4080 & n4091 ) | ( ~n4080 & n4092 ) | ( n4091 & n4092 ) ;
  assign n4094 = ( ~n3893 & n4092 ) | ( ~n3893 & n4093 ) | ( n4092 & n4093 ) ;
  assign n4095 = x97 | x98 ;
  assign n4096 = x97 & x98 ;
  assign n4097 = n4095 & ~n4096 ;
  assign n4098 = n3698 | n3701 ;
  assign n4099 = n4097 & n4098 ;
  assign n4100 = n3698 | n3703 ;
  assign n4101 = n4097 & n4100 ;
  assign n4102 = ( n3268 & n4099 ) | ( n3268 & n4101 ) | ( n4099 & n4101 ) ;
  assign n4103 = ( n3268 & n4098 ) | ( n3268 & n4100 ) | ( n4098 & n4100 ) ;
  assign n4104 = n4097 | n4103 ;
  assign n4105 = ~n4102 & n4104 ;
  assign n4106 = x97 & n131 ;
  assign n4107 = x96 & ~n156 ;
  assign n4108 = ( n135 & n4106 ) | ( n135 & n4107 ) | ( n4106 & n4107 ) ;
  assign n4109 = x0 & x98 ;
  assign n4110 = ( ~n135 & n4106 ) | ( ~n135 & n4109 ) | ( n4106 & n4109 ) ;
  assign n4111 = n4108 | n4110 ;
  assign n4112 = n139 | n4111 ;
  assign n4113 = ( n4105 & n4111 ) | ( n4105 & n4112 ) | ( n4111 & n4112 ) ;
  assign n4114 = x2 & n4113 ;
  assign n4115 = x2 & ~n4114 ;
  assign n4116 = ( n4113 & ~n4114 ) | ( n4113 & n4115 ) | ( ~n4114 & n4115 ) ;
  assign n4117 = n4094 | n4116 ;
  assign n4118 = ~n4116 & n4117 ;
  assign n4119 = ( ~n4094 & n4117 ) | ( ~n4094 & n4118 ) | ( n4117 & n4118 ) ;
  assign n4120 = n3886 | n3891 ;
  assign n4121 = n4119 & n4120 ;
  assign n4122 = n4119 | n4120 ;
  assign n4123 = ~n4121 & n4122 ;
  assign n4124 = ( n4094 & n4116 ) | ( n4094 & n4121 ) | ( n4116 & n4121 ) ;
  assign n4125 = n4055 | n4059 ;
  assign n4126 = n3980 | n3984 ;
  assign n4127 = n3944 | n3948 ;
  assign n4128 = x72 & n2775 ;
  assign n4129 = x71 & n2770 ;
  assign n4130 = x70 & ~n2769 ;
  assign n4131 = n2978 & n4130 ;
  assign n4132 = n4129 | n4131 ;
  assign n4133 = n4128 | n4132 ;
  assign n4134 = ( n435 & n2778 ) | ( n435 & n4133 ) | ( n2778 & n4133 ) ;
  assign n4135 = ( x29 & ~n4133 ) | ( x29 & n4134 ) | ( ~n4133 & n4134 ) ;
  assign n4136 = ~n4134 & n4135 ;
  assign n4137 = n4133 | n4135 ;
  assign n4138 = ( ~x29 & n4136 ) | ( ~x29 & n4137 ) | ( n4136 & n4137 ) ;
  assign n4139 = n264 & n3317 ;
  assign n4140 = x69 & n3314 ;
  assign n4141 = x68 & n3309 ;
  assign n4142 = x67 & ~n3308 ;
  assign n4143 = n3570 & n4142 ;
  assign n4144 = n4141 | n4143 ;
  assign n4145 = n4140 | n4144 ;
  assign n4146 = n4139 | n4145 ;
  assign n4147 = x32 | n4146 ;
  assign n4148 = ~x32 & n4147 ;
  assign n4149 = ( ~n4146 & n4147 ) | ( ~n4146 & n4148 ) | ( n4147 & n4148 ) ;
  assign n4150 = x66 & n3913 ;
  assign n4151 = x65 & n3908 ;
  assign n4152 = ~n3792 & n3912 ;
  assign n4153 = x64 & ~n3907 ;
  assign n4154 = n4152 & n4153 ;
  assign n4155 = n4151 | n4154 ;
  assign n4156 = n4150 | n4155 ;
  assign n4157 = n153 & n3916 ;
  assign n4158 = n4156 | n4157 ;
  assign n4159 = x35 | n4158 ;
  assign n4160 = ~x35 & n4159 ;
  assign n4161 = ( ~n4158 & n4159 ) | ( ~n4158 & n4160 ) | ( n4159 & n4160 ) ;
  assign n4162 = n3923 | n4161 ;
  assign n4163 = n3923 & n4161 ;
  assign n4164 = n4162 & ~n4163 ;
  assign n4165 = n3938 | n3941 ;
  assign n4166 = ( n4149 & n4164 ) | ( n4149 & n4165 ) | ( n4164 & n4165 ) ;
  assign n4167 = ( n4164 & n4165 ) | ( n4164 & ~n4166 ) | ( n4165 & ~n4166 ) ;
  assign n4168 = ( n4149 & ~n4166 ) | ( n4149 & n4167 ) | ( ~n4166 & n4167 ) ;
  assign n4169 = n4138 & n4168 ;
  assign n4170 = n4168 & ~n4169 ;
  assign n4171 = ( n4138 & ~n4169 ) | ( n4138 & n4170 ) | ( ~n4169 & n4170 ) ;
  assign n4172 = n4127 & n4171 ;
  assign n4173 = n4127 | n4171 ;
  assign n4174 = ~n4172 & n4173 ;
  assign n4175 = x75 & n2280 ;
  assign n4176 = x74 & n2275 ;
  assign n4177 = x73 & ~n2274 ;
  assign n4178 = n2481 & n4177 ;
  assign n4179 = n4176 | n4178 ;
  assign n4180 = n4175 | n4179 ;
  assign n4181 = n2283 | n4180 ;
  assign n4182 = ( n609 & n4180 ) | ( n609 & n4181 ) | ( n4180 & n4181 ) ;
  assign n4183 = x26 & n4182 ;
  assign n4184 = x26 & ~n4183 ;
  assign n4185 = ( n4182 & ~n4183 ) | ( n4182 & n4184 ) | ( ~n4183 & n4184 ) ;
  assign n4186 = ~n4174 & n4185 ;
  assign n4187 = n4174 & ~n4185 ;
  assign n4188 = n4186 | n4187 ;
  assign n4189 = n3961 | n3967 ;
  assign n4190 = n4188 & ~n4189 ;
  assign n4191 = ~n4188 & n4189 ;
  assign n4192 = x78 & n1817 ;
  assign n4193 = x77 & n1812 ;
  assign n4194 = x76 & ~n1811 ;
  assign n4195 = n1977 & n4194 ;
  assign n4196 = n4193 | n4195 ;
  assign n4197 = n4192 | n4196 ;
  assign n4198 = n1820 | n4197 ;
  assign n4199 = ( n868 & n4197 ) | ( n868 & n4198 ) | ( n4197 & n4198 ) ;
  assign n4200 = x23 & n4199 ;
  assign n4201 = x23 & ~n4200 ;
  assign n4202 = ( n4199 & ~n4200 ) | ( n4199 & n4201 ) | ( ~n4200 & n4201 ) ;
  assign n4203 = n4191 | n4202 ;
  assign n4204 = n4190 | n4203 ;
  assign n4205 = ( n4190 & n4191 ) | ( n4190 & n4202 ) | ( n4191 & n4202 ) ;
  assign n4206 = n4204 & ~n4205 ;
  assign n4207 = n4126 & n4206 ;
  assign n4208 = n4126 | n4206 ;
  assign n4209 = ~n4207 & n4208 ;
  assign n4210 = x81 & n1421 ;
  assign n4211 = x80 & n1416 ;
  assign n4212 = x79 & ~n1415 ;
  assign n4213 = n1584 & n4212 ;
  assign n4214 = n4211 | n4213 ;
  assign n4215 = n4210 | n4214 ;
  assign n4216 = n1424 | n4215 ;
  assign n4217 = ( n1256 & n4215 ) | ( n1256 & n4216 ) | ( n4215 & n4216 ) ;
  assign n4218 = x20 & n4217 ;
  assign n4219 = x20 & ~n4218 ;
  assign n4220 = ( n4217 & ~n4218 ) | ( n4217 & n4219 ) | ( ~n4218 & n4219 ) ;
  assign n4221 = n4209 & n4220 ;
  assign n4222 = n4209 & ~n4221 ;
  assign n4223 = ~n4209 & n4220 ;
  assign n4224 = n4222 | n4223 ;
  assign n4225 = n3998 | n4004 ;
  assign n4226 = n4224 | n4225 ;
  assign n4227 = n4224 & n4225 ;
  assign n4228 = n4226 & ~n4227 ;
  assign n4229 = x84 & n1071 ;
  assign n4230 = x83 & n1066 ;
  assign n4231 = x82 & ~n1065 ;
  assign n4232 = n1189 & n4231 ;
  assign n4233 = n4230 | n4232 ;
  assign n4234 = n4229 | n4233 ;
  assign n4235 = n1074 | n4234 ;
  assign n4236 = ( n1537 & n4234 ) | ( n1537 & n4235 ) | ( n4234 & n4235 ) ;
  assign n4237 = x17 & n4236 ;
  assign n4238 = x17 & ~n4237 ;
  assign n4239 = ( n4236 & ~n4237 ) | ( n4236 & n4238 ) | ( ~n4237 & n4238 ) ;
  assign n4240 = n4228 & n4239 ;
  assign n4241 = n4228 | n4239 ;
  assign n4242 = ~n4240 & n4241 ;
  assign n4243 = n4017 | n4023 ;
  assign n4244 = n4242 & n4243 ;
  assign n4245 = n4243 & ~n4244 ;
  assign n4246 = ( n4242 & ~n4244 ) | ( n4242 & n4245 ) | ( ~n4244 & n4245 ) ;
  assign n4247 = x87 & n771 ;
  assign n4248 = x86 & n766 ;
  assign n4249 = x85 & ~n765 ;
  assign n4250 = n905 & n4249 ;
  assign n4251 = n4248 | n4250 ;
  assign n4252 = n4247 | n4251 ;
  assign n4253 = n774 | n4252 ;
  assign n4254 = ( n2067 & n4252 ) | ( n2067 & n4253 ) | ( n4252 & n4253 ) ;
  assign n4255 = x14 & n4254 ;
  assign n4256 = x14 & ~n4255 ;
  assign n4257 = ( n4254 & ~n4255 ) | ( n4254 & n4256 ) | ( ~n4255 & n4256 ) ;
  assign n4258 = n4246 | n4257 ;
  assign n4259 = n4246 & n4257 ;
  assign n4260 = n4258 & ~n4259 ;
  assign n4261 = n4036 | n4042 ;
  assign n4262 = n4260 & n4261 ;
  assign n4263 = n4260 | n4261 ;
  assign n4264 = ~n4262 & n4263 ;
  assign n4265 = x90 & n528 ;
  assign n4266 = x89 & n523 ;
  assign n4267 = x88 & ~n522 ;
  assign n4268 = n635 & n4267 ;
  assign n4269 = n4266 | n4268 ;
  assign n4270 = n4265 | n4269 ;
  assign n4271 = n531 | n4270 ;
  assign n4272 = ( n2410 & n4270 ) | ( n2410 & n4271 ) | ( n4270 & n4271 ) ;
  assign n4273 = x11 & n4272 ;
  assign n4274 = x11 & ~n4273 ;
  assign n4275 = ( n4272 & ~n4273 ) | ( n4272 & n4274 ) | ( ~n4273 & n4274 ) ;
  assign n4276 = n4264 | n4275 ;
  assign n4277 = n4264 & n4275 ;
  assign n4278 = n4276 & ~n4277 ;
  assign n4279 = n4125 & n4278 ;
  assign n4280 = n4125 | n4278 ;
  assign n4281 = ~n4279 & n4280 ;
  assign n4282 = x93 & n337 ;
  assign n4283 = x92 & n332 ;
  assign n4284 = x91 & ~n331 ;
  assign n4285 = n396 & n4284 ;
  assign n4286 = n4283 | n4285 ;
  assign n4287 = n4282 | n4286 ;
  assign n4288 = n340 | n4287 ;
  assign n4289 = ( n2931 & n4287 ) | ( n2931 & n4288 ) | ( n4287 & n4288 ) ;
  assign n4290 = x8 & n4289 ;
  assign n4291 = x8 & ~n4290 ;
  assign n4292 = ( n4289 & ~n4290 ) | ( n4289 & n4291 ) | ( ~n4290 & n4291 ) ;
  assign n4293 = n4281 & n4292 ;
  assign n4294 = n4281 & ~n4293 ;
  assign n4295 = ~n4281 & n4292 ;
  assign n4296 = n4294 | n4295 ;
  assign n4297 = n4073 | n4079 ;
  assign n4298 = n4296 | n4297 ;
  assign n4299 = n4296 & n4297 ;
  assign n4300 = n4298 & ~n4299 ;
  assign n4301 = x96 & n206 ;
  assign n4302 = x95 & n201 ;
  assign n4303 = x94 & ~n200 ;
  assign n4304 = n243 & n4303 ;
  assign n4305 = n4302 | n4304 ;
  assign n4306 = n4301 | n4305 ;
  assign n4307 = n209 | n4306 ;
  assign n4308 = ( n3509 & n4306 ) | ( n3509 & n4307 ) | ( n4306 & n4307 ) ;
  assign n4309 = x5 & n4308 ;
  assign n4310 = x5 & ~n4309 ;
  assign n4311 = ( n4308 & ~n4309 ) | ( n4308 & n4310 ) | ( ~n4309 & n4310 ) ;
  assign n4312 = n4300 & n4311 ;
  assign n4313 = n4300 | n4311 ;
  assign n4314 = ~n4312 & n4313 ;
  assign n4315 = ( n3893 & n4080 ) | ( n3893 & n4091 ) | ( n4080 & n4091 ) ;
  assign n4316 = n4314 & n4315 ;
  assign n4317 = n4315 & ~n4316 ;
  assign n4318 = ( n4314 & ~n4316 ) | ( n4314 & n4317 ) | ( ~n4316 & n4317 ) ;
  assign n4319 = x98 | x99 ;
  assign n4320 = x98 & x99 ;
  assign n4321 = n4319 & ~n4320 ;
  assign n4322 = n4096 | n4102 ;
  assign n4323 = n4321 & n4322 ;
  assign n4324 = n4321 | n4322 ;
  assign n4325 = ~n4323 & n4324 ;
  assign n4326 = x98 & n131 ;
  assign n4327 = x97 & ~n156 ;
  assign n4328 = ( n135 & n4326 ) | ( n135 & n4327 ) | ( n4326 & n4327 ) ;
  assign n4329 = x0 & x99 ;
  assign n4330 = ( ~n135 & n4326 ) | ( ~n135 & n4329 ) | ( n4326 & n4329 ) ;
  assign n4331 = n4328 | n4330 ;
  assign n4332 = n139 | n4331 ;
  assign n4333 = ( n4325 & n4331 ) | ( n4325 & n4332 ) | ( n4331 & n4332 ) ;
  assign n4334 = x2 & n4333 ;
  assign n4335 = x2 & ~n4334 ;
  assign n4336 = ( n4333 & ~n4334 ) | ( n4333 & n4335 ) | ( ~n4334 & n4335 ) ;
  assign n4337 = ( n4124 & n4318 ) | ( n4124 & ~n4336 ) | ( n4318 & ~n4336 ) ;
  assign n4338 = ( ~n4318 & n4336 ) | ( ~n4318 & n4337 ) | ( n4336 & n4337 ) ;
  assign n4339 = ( ~n4124 & n4337 ) | ( ~n4124 & n4338 ) | ( n4337 & n4338 ) ;
  assign n4340 = n4312 | n4316 ;
  assign n4341 = x94 & n337 ;
  assign n4342 = x93 & n332 ;
  assign n4343 = x92 & ~n331 ;
  assign n4344 = n396 & n4343 ;
  assign n4345 = n4342 | n4344 ;
  assign n4346 = n4341 | n4345 ;
  assign n4347 = n340 | n4346 ;
  assign n4348 = ( n3271 & n4346 ) | ( n3271 & n4347 ) | ( n4346 & n4347 ) ;
  assign n4349 = x8 & n4348 ;
  assign n4350 = x8 & ~n4349 ;
  assign n4351 = ( n4348 & ~n4349 ) | ( n4348 & n4350 ) | ( ~n4349 & n4350 ) ;
  assign n4352 = x91 & n528 ;
  assign n4353 = x90 & n523 ;
  assign n4354 = x89 & ~n522 ;
  assign n4355 = n635 & n4354 ;
  assign n4356 = n4353 | n4355 ;
  assign n4357 = n4352 | n4356 ;
  assign n4358 = n531 | n4357 ;
  assign n4359 = ( n2714 & n4357 ) | ( n2714 & n4358 ) | ( n4357 & n4358 ) ;
  assign n4360 = x11 & n4359 ;
  assign n4361 = x11 & ~n4360 ;
  assign n4362 = ( n4359 & ~n4360 ) | ( n4359 & n4361 ) | ( ~n4360 & n4361 ) ;
  assign n4363 = n4259 | n4262 ;
  assign n4364 = x88 & n771 ;
  assign n4365 = x87 & n766 ;
  assign n4366 = x86 & ~n765 ;
  assign n4367 = n905 & n4366 ;
  assign n4368 = n4365 | n4367 ;
  assign n4369 = n4364 | n4368 ;
  assign n4370 = n774 | n4369 ;
  assign n4371 = ( n2095 & n4369 ) | ( n2095 & n4370 ) | ( n4369 & n4370 ) ;
  assign n4372 = x14 & n4371 ;
  assign n4373 = x14 & ~n4372 ;
  assign n4374 = ( n4371 & ~n4372 ) | ( n4371 & n4373 ) | ( ~n4372 & n4373 ) ;
  assign n4375 = x85 & n1071 ;
  assign n4376 = x84 & n1066 ;
  assign n4377 = x83 & ~n1065 ;
  assign n4378 = n1189 & n4377 ;
  assign n4379 = n4376 | n4378 ;
  assign n4380 = n4375 | n4379 ;
  assign n4381 = n1074 | n4380 ;
  assign n4382 = ( n1765 & n4380 ) | ( n1765 & n4381 ) | ( n4380 & n4381 ) ;
  assign n4383 = x17 & n4382 ;
  assign n4384 = x17 & ~n4383 ;
  assign n4385 = ( n4382 & ~n4383 ) | ( n4382 & n4384 ) | ( ~n4383 & n4384 ) ;
  assign n4386 = n4240 | n4244 ;
  assign n4387 = x82 & n1421 ;
  assign n4388 = x81 & n1416 ;
  assign n4389 = x80 & ~n1415 ;
  assign n4390 = n1584 & n4389 ;
  assign n4391 = n4388 | n4390 ;
  assign n4392 = n4387 | n4391 ;
  assign n4393 = n1424 | n4392 ;
  assign n4394 = ( n1371 & n4392 ) | ( n1371 & n4393 ) | ( n4392 & n4393 ) ;
  assign n4395 = x20 & n4394 ;
  assign n4396 = x20 & ~n4395 ;
  assign n4397 = ( n4394 & ~n4395 ) | ( n4394 & n4396 ) | ( ~n4395 & n4396 ) ;
  assign n4398 = x79 & n1817 ;
  assign n4399 = x78 & n1812 ;
  assign n4400 = x77 & ~n1811 ;
  assign n4401 = n1977 & n4400 ;
  assign n4402 = n4399 | n4401 ;
  assign n4403 = n4398 | n4402 ;
  assign n4404 = n1820 | n4403 ;
  assign n4405 = ( n961 & n4403 ) | ( n961 & n4404 ) | ( n4403 & n4404 ) ;
  assign n4406 = x23 & n4405 ;
  assign n4407 = x23 & ~n4406 ;
  assign n4408 = ( n4405 & ~n4406 ) | ( n4405 & n4407 ) | ( ~n4406 & n4407 ) ;
  assign n4409 = n4205 | n4207 ;
  assign n4410 = x70 & n3314 ;
  assign n4411 = x69 & n3309 ;
  assign n4412 = x68 & ~n3308 ;
  assign n4413 = n3570 & n4412 ;
  assign n4414 = n4411 | n4413 ;
  assign n4415 = n4410 | n4414 ;
  assign n4416 = n3317 | n4415 ;
  assign n4417 = ( n310 & n4415 ) | ( n310 & n4416 ) | ( n4415 & n4416 ) ;
  assign n4418 = x32 & ~n4417 ;
  assign n4419 = ~x32 & n4417 ;
  assign n4420 = n4418 | n4419 ;
  assign n4421 = x35 & ~x36 ;
  assign n4422 = ~x35 & x36 ;
  assign n4423 = n4421 | n4422 ;
  assign n4424 = x64 & n4423 ;
  assign n4425 = x67 & n3913 ;
  assign n4426 = x66 & n3908 ;
  assign n4427 = x65 & ~n3907 ;
  assign n4428 = n4152 & n4427 ;
  assign n4429 = n4426 | n4428 ;
  assign n4430 = n4425 | n4429 ;
  assign n4431 = n180 & n3916 ;
  assign n4432 = n4430 | n4431 ;
  assign n4433 = x35 & ~n4432 ;
  assign n4434 = ~x35 & n4432 ;
  assign n4435 = n4433 | n4434 ;
  assign n4436 = ( n4163 & n4424 ) | ( n4163 & n4435 ) | ( n4424 & n4435 ) ;
  assign n4437 = ( n4163 & n4435 ) | ( n4163 & ~n4436 ) | ( n4435 & ~n4436 ) ;
  assign n4438 = ( n4424 & ~n4436 ) | ( n4424 & n4437 ) | ( ~n4436 & n4437 ) ;
  assign n4439 = ( n4166 & n4420 ) | ( n4166 & ~n4438 ) | ( n4420 & ~n4438 ) ;
  assign n4440 = ( ~n4166 & n4438 ) | ( ~n4166 & n4439 ) | ( n4438 & n4439 ) ;
  assign n4441 = ( ~n4420 & n4439 ) | ( ~n4420 & n4440 ) | ( n4439 & n4440 ) ;
  assign n4442 = x73 & n2775 ;
  assign n4443 = x72 & n2770 ;
  assign n4444 = x71 & ~n2769 ;
  assign n4445 = n2978 & n4444 ;
  assign n4446 = n4443 | n4445 ;
  assign n4447 = n4442 | n4446 ;
  assign n4448 = ( n499 & n2778 ) | ( n499 & n4447 ) | ( n2778 & n4447 ) ;
  assign n4449 = ( x29 & ~n4447 ) | ( x29 & n4448 ) | ( ~n4447 & n4448 ) ;
  assign n4450 = ~n4448 & n4449 ;
  assign n4451 = n4447 | n4449 ;
  assign n4452 = ( ~x29 & n4450 ) | ( ~x29 & n4451 ) | ( n4450 & n4451 ) ;
  assign n4453 = n4441 & n4452 ;
  assign n4454 = n4441 | n4452 ;
  assign n4455 = ~n4453 & n4454 ;
  assign n4456 = n4169 | n4172 ;
  assign n4457 = n4455 | n4456 ;
  assign n4458 = n4455 & n4456 ;
  assign n4459 = n4457 & ~n4458 ;
  assign n4460 = x76 & n2280 ;
  assign n4461 = x75 & n2275 ;
  assign n4462 = x74 & ~n2274 ;
  assign n4463 = n2481 & n4462 ;
  assign n4464 = n4461 | n4463 ;
  assign n4465 = n4460 | n4464 ;
  assign n4466 = n2283 | n4465 ;
  assign n4467 = ( n740 & n4465 ) | ( n740 & n4466 ) | ( n4465 & n4466 ) ;
  assign n4468 = x26 & n4467 ;
  assign n4469 = x26 & ~n4468 ;
  assign n4470 = ( n4467 & ~n4468 ) | ( n4467 & n4469 ) | ( ~n4468 & n4469 ) ;
  assign n4471 = n4459 | n4470 ;
  assign n4472 = n4459 & n4470 ;
  assign n4473 = n4471 & ~n4472 ;
  assign n4474 = ( n4174 & n4185 ) | ( n4174 & n4189 ) | ( n4185 & n4189 ) ;
  assign n4475 = n4473 & n4474 ;
  assign n4476 = n4473 | n4474 ;
  assign n4477 = ~n4475 & n4476 ;
  assign n4478 = ( n4408 & n4409 ) | ( n4408 & ~n4477 ) | ( n4409 & ~n4477 ) ;
  assign n4479 = ( ~n4409 & n4477 ) | ( ~n4409 & n4478 ) | ( n4477 & n4478 ) ;
  assign n4480 = ( ~n4408 & n4478 ) | ( ~n4408 & n4479 ) | ( n4478 & n4479 ) ;
  assign n4481 = n4397 & n4480 ;
  assign n4482 = n4397 | n4480 ;
  assign n4483 = ~n4481 & n4482 ;
  assign n4484 = n4221 | n4227 ;
  assign n4485 = n4483 | n4484 ;
  assign n4486 = n4483 & n4484 ;
  assign n4487 = n4485 & ~n4486 ;
  assign n4488 = ( n4385 & n4386 ) | ( n4385 & ~n4487 ) | ( n4386 & ~n4487 ) ;
  assign n4489 = ( ~n4386 & n4487 ) | ( ~n4386 & n4488 ) | ( n4487 & n4488 ) ;
  assign n4490 = ( ~n4385 & n4488 ) | ( ~n4385 & n4489 ) | ( n4488 & n4489 ) ;
  assign n4491 = n4374 | n4490 ;
  assign n4492 = n4374 & n4490 ;
  assign n4493 = n4491 & ~n4492 ;
  assign n4494 = n4363 & n4493 ;
  assign n4495 = n4363 | n4493 ;
  assign n4496 = ~n4494 & n4495 ;
  assign n4497 = n4277 | n4279 ;
  assign n4498 = ( n4362 & n4496 ) | ( n4362 & n4497 ) | ( n4496 & n4497 ) ;
  assign n4499 = ( n4496 & n4497 ) | ( n4496 & ~n4498 ) | ( n4497 & ~n4498 ) ;
  assign n4500 = ( n4362 & ~n4498 ) | ( n4362 & n4499 ) | ( ~n4498 & n4499 ) ;
  assign n4501 = n4351 | n4500 ;
  assign n4502 = n4351 & n4500 ;
  assign n4503 = n4501 & ~n4502 ;
  assign n4504 = n4293 | n4299 ;
  assign n4505 = n4503 & n4504 ;
  assign n4506 = n4503 | n4504 ;
  assign n4507 = ~n4505 & n4506 ;
  assign n4508 = x97 & n206 ;
  assign n4509 = x96 & n201 ;
  assign n4510 = x95 & ~n200 ;
  assign n4511 = n243 & n4510 ;
  assign n4512 = n4509 | n4511 ;
  assign n4513 = n4508 | n4512 ;
  assign n4514 = n209 | n4513 ;
  assign n4515 = ( n3707 & n4513 ) | ( n3707 & n4514 ) | ( n4513 & n4514 ) ;
  assign n4516 = x5 & n4515 ;
  assign n4517 = x5 & ~n4516 ;
  assign n4518 = ( n4515 & ~n4516 ) | ( n4515 & n4517 ) | ( ~n4516 & n4517 ) ;
  assign n4519 = n4507 & n4518 ;
  assign n4520 = n4507 | n4518 ;
  assign n4521 = ~n4519 & n4520 ;
  assign n4522 = n4340 & n4521 ;
  assign n4523 = n4340 | n4521 ;
  assign n4524 = ~n4522 & n4523 ;
  assign n4525 = x99 | x100 ;
  assign n4526 = x99 & x100 ;
  assign n4527 = n4525 & ~n4526 ;
  assign n4528 = n4320 & n4527 ;
  assign n4529 = ( n4323 & n4527 ) | ( n4323 & n4528 ) | ( n4527 & n4528 ) ;
  assign n4530 = n4320 | n4527 ;
  assign n4531 = n4323 | n4530 ;
  assign n4532 = ~n4529 & n4531 ;
  assign n4533 = x99 & n131 ;
  assign n4534 = x98 & ~n156 ;
  assign n4535 = ( n135 & n4533 ) | ( n135 & n4534 ) | ( n4533 & n4534 ) ;
  assign n4536 = x0 & x100 ;
  assign n4537 = ( ~n135 & n4533 ) | ( ~n135 & n4536 ) | ( n4533 & n4536 ) ;
  assign n4538 = n4535 | n4537 ;
  assign n4539 = n139 | n4538 ;
  assign n4540 = ( n4532 & n4538 ) | ( n4532 & n4539 ) | ( n4538 & n4539 ) ;
  assign n4541 = x2 & n4540 ;
  assign n4542 = x2 & ~n4541 ;
  assign n4543 = ( n4540 & ~n4541 ) | ( n4540 & n4542 ) | ( ~n4541 & n4542 ) ;
  assign n4544 = n4524 & n4543 ;
  assign n4545 = n4524 & ~n4544 ;
  assign n4546 = ~n4524 & n4543 ;
  assign n4547 = n4545 | n4546 ;
  assign n4548 = ( n4124 & n4318 ) | ( n4124 & n4336 ) | ( n4318 & n4336 ) ;
  assign n4549 = n4547 | n4548 ;
  assign n4550 = n4547 & n4548 ;
  assign n4551 = n4549 & ~n4550 ;
  assign n4552 = n4544 | n4550 ;
  assign n4553 = x71 & n3314 ;
  assign n4554 = x70 & n3309 ;
  assign n4555 = x69 & ~n3308 ;
  assign n4556 = n3570 & n4555 ;
  assign n4557 = n4554 | n4556 ;
  assign n4558 = n4553 | n4557 ;
  assign n4559 = n3317 | n4558 ;
  assign n4560 = ( n376 & n4558 ) | ( n376 & n4559 ) | ( n4558 & n4559 ) ;
  assign n4561 = x32 & ~n4560 ;
  assign n4562 = ~x32 & n4560 ;
  assign n4563 = n4561 | n4562 ;
  assign n4564 = ~x36 & x37 ;
  assign n4565 = x36 & ~x37 ;
  assign n4566 = n4564 | n4565 ;
  assign n4567 = ~n4423 & n4566 ;
  assign n4568 = x64 & n4567 ;
  assign n4569 = ~x37 & x38 ;
  assign n4570 = x37 & ~x38 ;
  assign n4571 = n4569 | n4570 ;
  assign n4572 = n4423 & ~n4571 ;
  assign n4573 = x65 & n4572 ;
  assign n4574 = n4568 | n4573 ;
  assign n4575 = n4423 & n4571 ;
  assign n4576 = n142 & n4575 ;
  assign n4577 = n4574 | n4576 ;
  assign n4578 = x38 | n4577 ;
  assign n4579 = ~x38 & n4578 ;
  assign n4580 = ( ~n4577 & n4578 ) | ( ~n4577 & n4579 ) | ( n4578 & n4579 ) ;
  assign n4581 = x38 & ~n4424 ;
  assign n4582 = n4580 & n4581 ;
  assign n4583 = n4580 | n4581 ;
  assign n4584 = ~n4582 & n4583 ;
  assign n4585 = n229 & n3916 ;
  assign n4586 = x68 & n3913 ;
  assign n4587 = x67 & n3908 ;
  assign n4588 = x66 & ~n3907 ;
  assign n4589 = n4152 & n4588 ;
  assign n4590 = n4587 | n4589 ;
  assign n4591 = n4586 | n4590 ;
  assign n4592 = n4585 | n4591 ;
  assign n4593 = x35 | n4592 ;
  assign n4594 = ~x35 & n4593 ;
  assign n4595 = ( ~n4592 & n4593 ) | ( ~n4592 & n4594 ) | ( n4593 & n4594 ) ;
  assign n4596 = n4584 | n4595 ;
  assign n4597 = n4584 & n4595 ;
  assign n4598 = n4596 & ~n4597 ;
  assign n4599 = n4436 | n4598 ;
  assign n4600 = n4436 & n4598 ;
  assign n4601 = n4599 & ~n4600 ;
  assign n4602 = n4563 | n4601 ;
  assign n4603 = n4563 & n4601 ;
  assign n4604 = n4602 & ~n4603 ;
  assign n4605 = ( n4166 & n4420 ) | ( n4166 & n4438 ) | ( n4420 & n4438 ) ;
  assign n4606 = n4604 | n4605 ;
  assign n4607 = n4604 & n4605 ;
  assign n4608 = n4606 & ~n4607 ;
  assign n4609 = x74 & n2775 ;
  assign n4610 = x73 & n2770 ;
  assign n4611 = x72 & ~n2769 ;
  assign n4612 = n2978 & n4611 ;
  assign n4613 = n4610 | n4612 ;
  assign n4614 = n4609 | n4613 ;
  assign n4615 = n2778 | n4614 ;
  assign n4616 = ( n587 & n4614 ) | ( n587 & n4615 ) | ( n4614 & n4615 ) ;
  assign n4617 = x29 & n4616 ;
  assign n4618 = x29 & ~n4617 ;
  assign n4619 = ( n4616 & ~n4617 ) | ( n4616 & n4618 ) | ( ~n4617 & n4618 ) ;
  assign n4620 = n4608 | n4619 ;
  assign n4621 = n4608 & n4619 ;
  assign n4622 = n4620 & ~n4621 ;
  assign n4623 = n4453 | n4458 ;
  assign n4624 = n4622 & n4623 ;
  assign n4625 = n4622 | n4623 ;
  assign n4626 = ~n4624 & n4625 ;
  assign n4627 = x77 & n2280 ;
  assign n4628 = x76 & n2275 ;
  assign n4629 = x75 & ~n2274 ;
  assign n4630 = n2481 & n4629 ;
  assign n4631 = n4628 | n4630 ;
  assign n4632 = n4627 | n4631 ;
  assign n4633 = n2283 | n4632 ;
  assign n4634 = ( n846 & n4632 ) | ( n846 & n4633 ) | ( n4632 & n4633 ) ;
  assign n4635 = x26 & n4634 ;
  assign n4636 = x26 & ~n4635 ;
  assign n4637 = ( n4634 & ~n4635 ) | ( n4634 & n4636 ) | ( ~n4635 & n4636 ) ;
  assign n4638 = n4626 | n4637 ;
  assign n4639 = n4626 & n4637 ;
  assign n4640 = n4638 & ~n4639 ;
  assign n4641 = n4472 | n4475 ;
  assign n4642 = n4640 & n4641 ;
  assign n4643 = n4640 | n4641 ;
  assign n4644 = ~n4642 & n4643 ;
  assign n4645 = x80 & n1817 ;
  assign n4646 = x79 & n1812 ;
  assign n4647 = x78 & ~n1811 ;
  assign n4648 = n1977 & n4647 ;
  assign n4649 = n4646 | n4648 ;
  assign n4650 = n4645 | n4649 ;
  assign n4651 = n1820 | n4650 ;
  assign n4652 = ( n1147 & n4650 ) | ( n1147 & n4651 ) | ( n4650 & n4651 ) ;
  assign n4653 = x23 & n4652 ;
  assign n4654 = x23 & ~n4653 ;
  assign n4655 = ( n4652 & ~n4653 ) | ( n4652 & n4654 ) | ( ~n4653 & n4654 ) ;
  assign n4656 = n4644 & n4655 ;
  assign n4657 = n4644 & ~n4656 ;
  assign n4658 = ~n4644 & n4655 ;
  assign n4659 = n4657 | n4658 ;
  assign n4660 = ( n4408 & n4409 ) | ( n4408 & n4477 ) | ( n4409 & n4477 ) ;
  assign n4661 = n4659 | n4660 ;
  assign n4662 = n4659 & n4660 ;
  assign n4663 = n4661 & ~n4662 ;
  assign n4664 = x83 & n1421 ;
  assign n4665 = x82 & n1416 ;
  assign n4666 = x81 & ~n1415 ;
  assign n4667 = n1584 & n4666 ;
  assign n4668 = n4665 | n4667 ;
  assign n4669 = n4664 | n4668 ;
  assign n4670 = n1424 | n4669 ;
  assign n4671 = ( n1510 & n4669 ) | ( n1510 & n4670 ) | ( n4669 & n4670 ) ;
  assign n4672 = x20 & n4671 ;
  assign n4673 = x20 & ~n4672 ;
  assign n4674 = ( n4671 & ~n4672 ) | ( n4671 & n4673 ) | ( ~n4672 & n4673 ) ;
  assign n4675 = n4663 & n4674 ;
  assign n4676 = n4663 & ~n4675 ;
  assign n4677 = ~n4663 & n4674 ;
  assign n4678 = n4676 | n4677 ;
  assign n4679 = n4481 | n4486 ;
  assign n4680 = n4678 | n4679 ;
  assign n4681 = n4678 & n4679 ;
  assign n4682 = n4680 & ~n4681 ;
  assign n4683 = x86 & n1071 ;
  assign n4684 = x85 & n1066 ;
  assign n4685 = x84 & ~n1065 ;
  assign n4686 = n1189 & n4685 ;
  assign n4687 = n4684 | n4686 ;
  assign n4688 = n4683 | n4687 ;
  assign n4689 = n1074 | n4688 ;
  assign n4690 = ( n1921 & n4688 ) | ( n1921 & n4689 ) | ( n4688 & n4689 ) ;
  assign n4691 = x17 & n4690 ;
  assign n4692 = x17 & ~n4691 ;
  assign n4693 = ( n4690 & ~n4691 ) | ( n4690 & n4692 ) | ( ~n4691 & n4692 ) ;
  assign n4694 = n4682 & n4693 ;
  assign n4695 = n4682 & ~n4694 ;
  assign n4696 = ~n4682 & n4693 ;
  assign n4697 = n4695 | n4696 ;
  assign n4698 = ( n4385 & n4386 ) | ( n4385 & n4487 ) | ( n4386 & n4487 ) ;
  assign n4699 = n4697 | n4698 ;
  assign n4700 = n4697 & n4698 ;
  assign n4701 = n4699 & ~n4700 ;
  assign n4702 = x89 & n771 ;
  assign n4703 = x88 & n766 ;
  assign n4704 = x87 & ~n765 ;
  assign n4705 = n905 & n4704 ;
  assign n4706 = n4703 | n4705 ;
  assign n4707 = n4702 | n4706 ;
  assign n4708 = n774 | n4707 ;
  assign n4709 = ( n2244 & n4707 ) | ( n2244 & n4708 ) | ( n4707 & n4708 ) ;
  assign n4710 = x14 & n4709 ;
  assign n4711 = x14 & ~n4710 ;
  assign n4712 = ( n4709 & ~n4710 ) | ( n4709 & n4711 ) | ( ~n4710 & n4711 ) ;
  assign n4713 = n4701 & n4712 ;
  assign n4714 = n4701 | n4712 ;
  assign n4715 = ~n4713 & n4714 ;
  assign n4716 = n4492 | n4494 ;
  assign n4717 = n4715 & n4716 ;
  assign n4718 = n4716 & ~n4717 ;
  assign n4719 = ( n4715 & ~n4717 ) | ( n4715 & n4718 ) | ( ~n4717 & n4718 ) ;
  assign n4720 = x92 & n528 ;
  assign n4721 = x91 & n523 ;
  assign n4722 = x90 & ~n522 ;
  assign n4723 = n635 & n4722 ;
  assign n4724 = n4721 | n4723 ;
  assign n4725 = n4720 | n4724 ;
  assign n4726 = n531 | n4725 ;
  assign n4727 = ( n2904 & n4725 ) | ( n2904 & n4726 ) | ( n4725 & n4726 ) ;
  assign n4728 = x11 & n4727 ;
  assign n4729 = x11 & ~n4728 ;
  assign n4730 = ( n4727 & ~n4728 ) | ( n4727 & n4729 ) | ( ~n4728 & n4729 ) ;
  assign n4731 = n4719 | n4730 ;
  assign n4732 = n4719 & n4730 ;
  assign n4733 = n4731 & ~n4732 ;
  assign n4734 = n4498 | n4733 ;
  assign n4735 = n4498 & n4733 ;
  assign n4736 = n4734 & ~n4735 ;
  assign n4737 = x95 & n337 ;
  assign n4738 = x94 & n332 ;
  assign n4739 = x93 & ~n331 ;
  assign n4740 = n396 & n4739 ;
  assign n4741 = n4738 | n4740 ;
  assign n4742 = n4737 | n4741 ;
  assign n4743 = n340 | n4742 ;
  assign n4744 = ( n3479 & n4742 ) | ( n3479 & n4743 ) | ( n4742 & n4743 ) ;
  assign n4745 = x8 & n4744 ;
  assign n4746 = x8 & ~n4745 ;
  assign n4747 = ( n4744 & ~n4745 ) | ( n4744 & n4746 ) | ( ~n4745 & n4746 ) ;
  assign n4748 = n4736 | n4747 ;
  assign n4749 = n4736 & n4747 ;
  assign n4750 = n4748 & ~n4749 ;
  assign n4751 = n4502 | n4505 ;
  assign n4752 = n4750 & n4751 ;
  assign n4753 = n4750 | n4751 ;
  assign n4754 = ~n4752 & n4753 ;
  assign n4755 = x98 & n206 ;
  assign n4756 = x97 & n201 ;
  assign n4757 = x96 & ~n200 ;
  assign n4758 = n243 & n4757 ;
  assign n4759 = n4756 | n4758 ;
  assign n4760 = n4755 | n4759 ;
  assign n4761 = n209 | n4760 ;
  assign n4762 = ( n4105 & n4760 ) | ( n4105 & n4761 ) | ( n4760 & n4761 ) ;
  assign n4763 = x5 & n4762 ;
  assign n4764 = x5 & ~n4763 ;
  assign n4765 = ( n4762 & ~n4763 ) | ( n4762 & n4764 ) | ( ~n4763 & n4764 ) ;
  assign n4766 = n4754 & n4765 ;
  assign n4767 = n4754 & ~n4766 ;
  assign n4768 = ~n4754 & n4765 ;
  assign n4769 = n4767 | n4768 ;
  assign n4770 = n4519 | n4522 ;
  assign n4771 = n4769 | n4770 ;
  assign n4772 = n4769 & n4770 ;
  assign n4773 = n4771 & ~n4772 ;
  assign n4774 = x100 | x101 ;
  assign n4775 = x100 & x101 ;
  assign n4776 = n4774 & ~n4775 ;
  assign n4777 = n4526 | n4528 ;
  assign n4778 = n4776 & n4777 ;
  assign n4779 = n4525 & n4776 ;
  assign n4780 = ( n4323 & n4778 ) | ( n4323 & n4779 ) | ( n4778 & n4779 ) ;
  assign n4781 = ( n4323 & n4525 ) | ( n4323 & n4777 ) | ( n4525 & n4777 ) ;
  assign n4782 = n4776 | n4781 ;
  assign n4783 = ~n4780 & n4782 ;
  assign n4784 = x100 & n131 ;
  assign n4785 = x99 & ~n156 ;
  assign n4786 = ( n135 & n4784 ) | ( n135 & n4785 ) | ( n4784 & n4785 ) ;
  assign n4787 = x0 & x101 ;
  assign n4788 = ( ~n135 & n4784 ) | ( ~n135 & n4787 ) | ( n4784 & n4787 ) ;
  assign n4789 = n4786 | n4788 ;
  assign n4790 = n139 | n4789 ;
  assign n4791 = ( n4783 & n4789 ) | ( n4783 & n4790 ) | ( n4789 & n4790 ) ;
  assign n4792 = x2 & n4791 ;
  assign n4793 = x2 & ~n4792 ;
  assign n4794 = ( n4791 & ~n4792 ) | ( n4791 & n4793 ) | ( ~n4792 & n4793 ) ;
  assign n4795 = n4773 | n4794 ;
  assign n4796 = n4773 & n4794 ;
  assign n4797 = n4795 & ~n4796 ;
  assign n4798 = n4552 | n4797 ;
  assign n4799 = n4552 & n4797 ;
  assign n4800 = n4798 & ~n4799 ;
  assign n4801 = n4732 | n4735 ;
  assign n4802 = n4713 | n4717 ;
  assign n4803 = n4621 | n4624 ;
  assign n4804 = x72 & n3314 ;
  assign n4805 = x71 & n3309 ;
  assign n4806 = x70 & ~n3308 ;
  assign n4807 = n3570 & n4806 ;
  assign n4808 = n4805 | n4807 ;
  assign n4809 = n4804 | n4808 ;
  assign n4810 = ( n435 & n3317 ) | ( n435 & n4809 ) | ( n3317 & n4809 ) ;
  assign n4811 = ( x32 & ~n4809 ) | ( x32 & n4810 ) | ( ~n4809 & n4810 ) ;
  assign n4812 = ~n4810 & n4811 ;
  assign n4813 = n4809 | n4811 ;
  assign n4814 = ( ~x32 & n4812 ) | ( ~x32 & n4813 ) | ( n4812 & n4813 ) ;
  assign n4815 = n264 & n3916 ;
  assign n4816 = x69 & n3913 ;
  assign n4817 = x68 & n3908 ;
  assign n4818 = x67 & ~n3907 ;
  assign n4819 = n4152 & n4818 ;
  assign n4820 = n4817 | n4819 ;
  assign n4821 = n4816 | n4820 ;
  assign n4822 = n4815 | n4821 ;
  assign n4823 = x35 | n4822 ;
  assign n4824 = ~x35 & n4823 ;
  assign n4825 = ( ~n4822 & n4823 ) | ( ~n4822 & n4824 ) | ( n4823 & n4824 ) ;
  assign n4826 = x66 & n4572 ;
  assign n4827 = x65 & n4567 ;
  assign n4828 = ~n4423 & n4571 ;
  assign n4829 = x64 & ~n4566 ;
  assign n4830 = n4828 & n4829 ;
  assign n4831 = n4827 | n4830 ;
  assign n4832 = n4826 | n4831 ;
  assign n4833 = n153 & n4575 ;
  assign n4834 = n4832 | n4833 ;
  assign n4835 = x38 | n4834 ;
  assign n4836 = ~x38 & n4835 ;
  assign n4837 = ( ~n4834 & n4835 ) | ( ~n4834 & n4836 ) | ( n4835 & n4836 ) ;
  assign n4838 = n4582 | n4837 ;
  assign n4839 = n4582 & n4837 ;
  assign n4840 = n4838 & ~n4839 ;
  assign n4841 = n4597 | n4600 ;
  assign n4842 = ( n4825 & n4840 ) | ( n4825 & n4841 ) | ( n4840 & n4841 ) ;
  assign n4843 = ( n4840 & n4841 ) | ( n4840 & ~n4842 ) | ( n4841 & ~n4842 ) ;
  assign n4844 = ( n4825 & ~n4842 ) | ( n4825 & n4843 ) | ( ~n4842 & n4843 ) ;
  assign n4845 = n4814 & n4844 ;
  assign n4846 = n4814 | n4844 ;
  assign n4847 = ~n4845 & n4846 ;
  assign n4848 = n4603 | n4607 ;
  assign n4849 = n4847 & n4848 ;
  assign n4850 = n4847 | n4848 ;
  assign n4851 = ~n4849 & n4850 ;
  assign n4852 = x75 & n2775 ;
  assign n4853 = x74 & n2770 ;
  assign n4854 = x73 & ~n2769 ;
  assign n4855 = n2978 & n4854 ;
  assign n4856 = n4853 | n4855 ;
  assign n4857 = n4852 | n4856 ;
  assign n4858 = n2778 | n4857 ;
  assign n4859 = ( n609 & n4857 ) | ( n609 & n4858 ) | ( n4857 & n4858 ) ;
  assign n4860 = x29 & n4859 ;
  assign n4861 = x29 & ~n4860 ;
  assign n4862 = ( n4859 & ~n4860 ) | ( n4859 & n4861 ) | ( ~n4860 & n4861 ) ;
  assign n4863 = n4851 & n4862 ;
  assign n4864 = n4851 & ~n4863 ;
  assign n4865 = ~n4851 & n4862 ;
  assign n4866 = n4864 | n4865 ;
  assign n4867 = n4803 & n4866 ;
  assign n4868 = n4803 & ~n4867 ;
  assign n4869 = n4866 & ~n4867 ;
  assign n4870 = n4868 | n4869 ;
  assign n4871 = x78 & n2280 ;
  assign n4872 = x77 & n2275 ;
  assign n4873 = x76 & ~n2274 ;
  assign n4874 = n2481 & n4873 ;
  assign n4875 = n4872 | n4874 ;
  assign n4876 = n4871 | n4875 ;
  assign n4877 = n2283 | n4876 ;
  assign n4878 = ( n868 & n4876 ) | ( n868 & n4877 ) | ( n4876 & n4877 ) ;
  assign n4879 = x26 & n4878 ;
  assign n4880 = x26 & ~n4879 ;
  assign n4881 = ( n4878 & ~n4879 ) | ( n4878 & n4880 ) | ( ~n4879 & n4880 ) ;
  assign n4882 = n4870 | n4881 ;
  assign n4883 = n4870 & n4881 ;
  assign n4884 = n4882 & ~n4883 ;
  assign n4885 = n4639 | n4642 ;
  assign n4886 = n4884 & n4885 ;
  assign n4887 = n4884 | n4885 ;
  assign n4888 = ~n4886 & n4887 ;
  assign n4889 = x81 & n1817 ;
  assign n4890 = x80 & n1812 ;
  assign n4891 = x79 & ~n1811 ;
  assign n4892 = n1977 & n4891 ;
  assign n4893 = n4890 | n4892 ;
  assign n4894 = n4889 | n4893 ;
  assign n4895 = n1820 | n4894 ;
  assign n4896 = ( n1256 & n4894 ) | ( n1256 & n4895 ) | ( n4894 & n4895 ) ;
  assign n4897 = x23 & n4896 ;
  assign n4898 = x23 & ~n4897 ;
  assign n4899 = ( n4896 & ~n4897 ) | ( n4896 & n4898 ) | ( ~n4897 & n4898 ) ;
  assign n4900 = n4888 & n4899 ;
  assign n4901 = n4888 & ~n4900 ;
  assign n4902 = ~n4888 & n4899 ;
  assign n4903 = n4901 | n4902 ;
  assign n4904 = n4656 | n4662 ;
  assign n4905 = n4903 | n4904 ;
  assign n4906 = n4903 & n4904 ;
  assign n4907 = n4905 & ~n4906 ;
  assign n4908 = x84 & n1421 ;
  assign n4909 = x83 & n1416 ;
  assign n4910 = x82 & ~n1415 ;
  assign n4911 = n1584 & n4910 ;
  assign n4912 = n4909 | n4911 ;
  assign n4913 = n4908 | n4912 ;
  assign n4914 = n1424 | n4913 ;
  assign n4915 = ( n1537 & n4913 ) | ( n1537 & n4914 ) | ( n4913 & n4914 ) ;
  assign n4916 = x20 & n4915 ;
  assign n4917 = x20 & ~n4916 ;
  assign n4918 = ( n4915 & ~n4916 ) | ( n4915 & n4917 ) | ( ~n4916 & n4917 ) ;
  assign n4919 = n4907 & n4918 ;
  assign n4920 = n4907 & ~n4919 ;
  assign n4921 = ~n4907 & n4918 ;
  assign n4922 = n4920 | n4921 ;
  assign n4923 = n4675 | n4681 ;
  assign n4924 = n4922 | n4923 ;
  assign n4925 = n4922 & n4923 ;
  assign n4926 = n4924 & ~n4925 ;
  assign n4927 = x87 & n1071 ;
  assign n4928 = x86 & n1066 ;
  assign n4929 = x85 & ~n1065 ;
  assign n4930 = n1189 & n4929 ;
  assign n4931 = n4928 | n4930 ;
  assign n4932 = n4927 | n4931 ;
  assign n4933 = n1074 | n4932 ;
  assign n4934 = ( n2067 & n4932 ) | ( n2067 & n4933 ) | ( n4932 & n4933 ) ;
  assign n4935 = x17 & n4934 ;
  assign n4936 = x17 & ~n4935 ;
  assign n4937 = ( n4934 & ~n4935 ) | ( n4934 & n4936 ) | ( ~n4935 & n4936 ) ;
  assign n4938 = n4926 & n4937 ;
  assign n4939 = n4926 | n4937 ;
  assign n4940 = ~n4938 & n4939 ;
  assign n4941 = n4694 | n4700 ;
  assign n4942 = n4940 | n4941 ;
  assign n4943 = ( n4694 & n4700 ) | ( n4694 & n4940 ) | ( n4700 & n4940 ) ;
  assign n4944 = n4942 & ~n4943 ;
  assign n4945 = x90 & n771 ;
  assign n4946 = x89 & n766 ;
  assign n4947 = x88 & ~n765 ;
  assign n4948 = n905 & n4947 ;
  assign n4949 = n4946 | n4948 ;
  assign n4950 = n4945 | n4949 ;
  assign n4951 = n774 | n4950 ;
  assign n4952 = ( n2410 & n4950 ) | ( n2410 & n4951 ) | ( n4950 & n4951 ) ;
  assign n4953 = x14 & n4952 ;
  assign n4954 = x14 & ~n4953 ;
  assign n4955 = ( n4952 & ~n4953 ) | ( n4952 & n4954 ) | ( ~n4953 & n4954 ) ;
  assign n4956 = n4944 | n4955 ;
  assign n4957 = n4944 & n4955 ;
  assign n4958 = n4956 & ~n4957 ;
  assign n4959 = n4802 & n4958 ;
  assign n4960 = n4802 | n4958 ;
  assign n4961 = ~n4959 & n4960 ;
  assign n4962 = x93 & n528 ;
  assign n4963 = x92 & n523 ;
  assign n4964 = x91 & ~n522 ;
  assign n4965 = n635 & n4964 ;
  assign n4966 = n4963 | n4965 ;
  assign n4967 = n4962 | n4966 ;
  assign n4968 = n531 | n4967 ;
  assign n4969 = ( n2931 & n4967 ) | ( n2931 & n4968 ) | ( n4967 & n4968 ) ;
  assign n4970 = x11 & n4969 ;
  assign n4971 = x11 & ~n4970 ;
  assign n4972 = ( n4969 & ~n4970 ) | ( n4969 & n4971 ) | ( ~n4970 & n4971 ) ;
  assign n4973 = n4961 | n4972 ;
  assign n4974 = n4961 & n4972 ;
  assign n4975 = n4973 & ~n4974 ;
  assign n4976 = n4801 & n4975 ;
  assign n4977 = n4801 | n4975 ;
  assign n4978 = ~n4976 & n4977 ;
  assign n4979 = x96 & n337 ;
  assign n4980 = x95 & n332 ;
  assign n4981 = x94 & ~n331 ;
  assign n4982 = n396 & n4981 ;
  assign n4983 = n4980 | n4982 ;
  assign n4984 = n4979 | n4983 ;
  assign n4985 = n340 | n4984 ;
  assign n4986 = ( n3509 & n4984 ) | ( n3509 & n4985 ) | ( n4984 & n4985 ) ;
  assign n4987 = x8 & n4986 ;
  assign n4988 = x8 & ~n4987 ;
  assign n4989 = ( n4986 & ~n4987 ) | ( n4986 & n4988 ) | ( ~n4987 & n4988 ) ;
  assign n4990 = n4978 | n4989 ;
  assign n4991 = n4978 & n4989 ;
  assign n4992 = n4990 & ~n4991 ;
  assign n4993 = n4749 | n4752 ;
  assign n4994 = n4992 & n4993 ;
  assign n4995 = n4992 | n4993 ;
  assign n4996 = ~n4994 & n4995 ;
  assign n4997 = x99 & n206 ;
  assign n4998 = x98 & n201 ;
  assign n4999 = x97 & ~n200 ;
  assign n5000 = n243 & n4999 ;
  assign n5001 = n4998 | n5000 ;
  assign n5002 = n4997 | n5001 ;
  assign n5003 = n209 | n5002 ;
  assign n5004 = ( n4325 & n5002 ) | ( n4325 & n5003 ) | ( n5002 & n5003 ) ;
  assign n5005 = x5 & n5004 ;
  assign n5006 = x5 & ~n5005 ;
  assign n5007 = ( n5004 & ~n5005 ) | ( n5004 & n5006 ) | ( ~n5005 & n5006 ) ;
  assign n5008 = n4996 | n5007 ;
  assign n5009 = n4996 & n5007 ;
  assign n5010 = n5008 & ~n5009 ;
  assign n5011 = n4766 | n5010 ;
  assign n5012 = n4772 | n5011 ;
  assign n5013 = ( n4766 & n4772 ) | ( n4766 & n5010 ) | ( n4772 & n5010 ) ;
  assign n5014 = n5012 & ~n5013 ;
  assign n5015 = x101 | x102 ;
  assign n5016 = x101 & x102 ;
  assign n5017 = n5015 & ~n5016 ;
  assign n5018 = n4775 | n4778 ;
  assign n5019 = n5017 & n5018 ;
  assign n5020 = n4775 | n4779 ;
  assign n5021 = n5017 & n5020 ;
  assign n5022 = ( n4323 & n5019 ) | ( n4323 & n5021 ) | ( n5019 & n5021 ) ;
  assign n5023 = ( n4323 & n5018 ) | ( n4323 & n5020 ) | ( n5018 & n5020 ) ;
  assign n5024 = n5017 | n5023 ;
  assign n5025 = ~n5022 & n5024 ;
  assign n5026 = x101 & n131 ;
  assign n5027 = x100 & ~n156 ;
  assign n5028 = ( n135 & n5026 ) | ( n135 & n5027 ) | ( n5026 & n5027 ) ;
  assign n5029 = x0 & x102 ;
  assign n5030 = ( ~n135 & n5026 ) | ( ~n135 & n5029 ) | ( n5026 & n5029 ) ;
  assign n5031 = n5028 | n5030 ;
  assign n5032 = n139 | n5031 ;
  assign n5033 = ( n5025 & n5031 ) | ( n5025 & n5032 ) | ( n5031 & n5032 ) ;
  assign n5034 = x2 & n5033 ;
  assign n5035 = x2 & ~n5034 ;
  assign n5036 = ( n5033 & ~n5034 ) | ( n5033 & n5035 ) | ( ~n5034 & n5035 ) ;
  assign n5037 = n5014 & n5036 ;
  assign n5038 = n5014 & ~n5037 ;
  assign n5039 = ~n5014 & n5036 ;
  assign n5040 = n5038 | n5039 ;
  assign n5041 = n4796 | n4799 ;
  assign n5042 = n5040 & n5041 ;
  assign n5043 = n5040 | n5041 ;
  assign n5044 = ~n5042 & n5043 ;
  assign n5045 = n5009 | n5013 ;
  assign n5046 = x100 & n206 ;
  assign n5047 = x99 & n201 ;
  assign n5048 = x98 & ~n200 ;
  assign n5049 = n243 & n5048 ;
  assign n5050 = n5047 | n5049 ;
  assign n5051 = n5046 | n5050 ;
  assign n5052 = n209 | n5051 ;
  assign n5053 = ( n4532 & n5051 ) | ( n4532 & n5052 ) | ( n5051 & n5052 ) ;
  assign n5054 = x5 & n5053 ;
  assign n5055 = x5 & ~n5054 ;
  assign n5056 = ( n5053 & ~n5054 ) | ( n5053 & n5055 ) | ( ~n5054 & n5055 ) ;
  assign n5057 = x97 & n337 ;
  assign n5058 = x96 & n332 ;
  assign n5059 = x95 & ~n331 ;
  assign n5060 = n396 & n5059 ;
  assign n5061 = n5058 | n5060 ;
  assign n5062 = n5057 | n5061 ;
  assign n5063 = n340 | n5062 ;
  assign n5064 = ( n3707 & n5062 ) | ( n3707 & n5063 ) | ( n5062 & n5063 ) ;
  assign n5065 = x8 & n5064 ;
  assign n5066 = x8 & ~n5065 ;
  assign n5067 = ( n5064 & ~n5065 ) | ( n5064 & n5066 ) | ( ~n5065 & n5066 ) ;
  assign n5068 = n4991 | n4994 ;
  assign n5069 = x94 & n528 ;
  assign n5070 = x93 & n523 ;
  assign n5071 = x92 & ~n522 ;
  assign n5072 = n635 & n5071 ;
  assign n5073 = n5070 | n5072 ;
  assign n5074 = n5069 | n5073 ;
  assign n5075 = n531 | n5074 ;
  assign n5076 = ( n3271 & n5074 ) | ( n3271 & n5075 ) | ( n5074 & n5075 ) ;
  assign n5077 = x11 & n5076 ;
  assign n5078 = x11 & ~n5077 ;
  assign n5079 = ( n5076 & ~n5077 ) | ( n5076 & n5078 ) | ( ~n5077 & n5078 ) ;
  assign n5080 = x91 & n771 ;
  assign n5081 = x90 & n766 ;
  assign n5082 = x89 & ~n765 ;
  assign n5083 = n905 & n5082 ;
  assign n5084 = n5081 | n5083 ;
  assign n5085 = n5080 | n5084 ;
  assign n5086 = n774 | n5085 ;
  assign n5087 = ( n2714 & n5085 ) | ( n2714 & n5086 ) | ( n5085 & n5086 ) ;
  assign n5088 = x14 & n5087 ;
  assign n5089 = x14 & ~n5088 ;
  assign n5090 = ( n5087 & ~n5088 ) | ( n5087 & n5089 ) | ( ~n5088 & n5089 ) ;
  assign n5091 = n4957 | n4959 ;
  assign n5092 = n4938 | n4943 ;
  assign n5093 = n4900 | n4906 ;
  assign n5094 = x82 & n1817 ;
  assign n5095 = x81 & n1812 ;
  assign n5096 = x80 & ~n1811 ;
  assign n5097 = n1977 & n5096 ;
  assign n5098 = n5095 | n5097 ;
  assign n5099 = n5094 | n5098 ;
  assign n5100 = n1820 | n5099 ;
  assign n5101 = ( n1371 & n5099 ) | ( n1371 & n5100 ) | ( n5099 & n5100 ) ;
  assign n5102 = x23 & n5101 ;
  assign n5103 = x23 & ~n5102 ;
  assign n5104 = ( n5101 & ~n5102 ) | ( n5101 & n5103 ) | ( ~n5102 & n5103 ) ;
  assign n5105 = x79 & n2280 ;
  assign n5106 = x78 & n2275 ;
  assign n5107 = x77 & ~n2274 ;
  assign n5108 = n2481 & n5107 ;
  assign n5109 = n5106 | n5108 ;
  assign n5110 = n5105 | n5109 ;
  assign n5111 = n2283 | n5110 ;
  assign n5112 = ( n961 & n5110 ) | ( n961 & n5111 ) | ( n5110 & n5111 ) ;
  assign n5113 = x26 & n5112 ;
  assign n5114 = x26 & ~n5113 ;
  assign n5115 = ( n5112 & ~n5113 ) | ( n5112 & n5114 ) | ( ~n5113 & n5114 ) ;
  assign n5116 = x38 & ~x39 ;
  assign n5117 = ~x38 & x39 ;
  assign n5118 = n5116 | n5117 ;
  assign n5119 = x64 & n5118 ;
  assign n5120 = x67 & n4572 ;
  assign n5121 = x66 & n4567 ;
  assign n5122 = x65 & ~n4566 ;
  assign n5123 = n4828 & n5122 ;
  assign n5124 = n5121 | n5123 ;
  assign n5125 = n5120 | n5124 ;
  assign n5126 = n180 & n4575 ;
  assign n5127 = n5125 | n5126 ;
  assign n5128 = x38 & ~n5127 ;
  assign n5129 = ~x38 & n5127 ;
  assign n5130 = n5128 | n5129 ;
  assign n5131 = ( n4839 & n5119 ) | ( n4839 & n5130 ) | ( n5119 & n5130 ) ;
  assign n5132 = ( n4839 & n5130 ) | ( n4839 & ~n5131 ) | ( n5130 & ~n5131 ) ;
  assign n5133 = ( n5119 & ~n5131 ) | ( n5119 & n5132 ) | ( ~n5131 & n5132 ) ;
  assign n5134 = x70 & n3913 ;
  assign n5135 = x69 & n3908 ;
  assign n5136 = x68 & ~n3907 ;
  assign n5137 = n4152 & n5136 ;
  assign n5138 = n5135 | n5137 ;
  assign n5139 = n5134 | n5138 ;
  assign n5140 = n3916 | n5139 ;
  assign n5141 = ( n310 & n5139 ) | ( n310 & n5140 ) | ( n5139 & n5140 ) ;
  assign n5142 = x35 & ~n5141 ;
  assign n5143 = ~x35 & n5141 ;
  assign n5144 = n5142 | n5143 ;
  assign n5145 = n5133 & n5144 ;
  assign n5146 = n5133 & ~n5145 ;
  assign n5147 = ~n5133 & n5144 ;
  assign n5148 = n5146 | n5147 ;
  assign n5149 = n4842 | n5148 ;
  assign n5150 = n4842 & n5148 ;
  assign n5151 = n5149 & ~n5150 ;
  assign n5152 = x73 & n3314 ;
  assign n5153 = x72 & n3309 ;
  assign n5154 = x71 & ~n3308 ;
  assign n5155 = n3570 & n5154 ;
  assign n5156 = n5153 | n5155 ;
  assign n5157 = n5152 | n5156 ;
  assign n5158 = ( n499 & n3317 ) | ( n499 & n5157 ) | ( n3317 & n5157 ) ;
  assign n5159 = ( x32 & ~n5157 ) | ( x32 & n5158 ) | ( ~n5157 & n5158 ) ;
  assign n5160 = ~n5158 & n5159 ;
  assign n5161 = n5157 | n5159 ;
  assign n5162 = ( ~x32 & n5160 ) | ( ~x32 & n5161 ) | ( n5160 & n5161 ) ;
  assign n5163 = n5151 & n5162 ;
  assign n5164 = n5151 & ~n5163 ;
  assign n5165 = ~n5151 & n5162 ;
  assign n5166 = n4845 | n4849 ;
  assign n5167 = n5165 | n5166 ;
  assign n5168 = n5164 | n5167 ;
  assign n5169 = ( n5164 & n5165 ) | ( n5164 & n5166 ) | ( n5165 & n5166 ) ;
  assign n5170 = n5168 & ~n5169 ;
  assign n5171 = x76 & n2775 ;
  assign n5172 = x75 & n2770 ;
  assign n5173 = x74 & ~n2769 ;
  assign n5174 = n2978 & n5173 ;
  assign n5175 = n5172 | n5174 ;
  assign n5176 = n5171 | n5175 ;
  assign n5177 = n2778 | n5176 ;
  assign n5178 = ( n740 & n5176 ) | ( n740 & n5177 ) | ( n5176 & n5177 ) ;
  assign n5179 = x29 & n5178 ;
  assign n5180 = x29 & ~n5179 ;
  assign n5181 = ( n5178 & ~n5179 ) | ( n5178 & n5180 ) | ( ~n5179 & n5180 ) ;
  assign n5182 = n5170 | n5181 ;
  assign n5183 = n5170 & n5181 ;
  assign n5184 = n5182 & ~n5183 ;
  assign n5185 = n4863 | n4867 ;
  assign n5186 = n5184 & n5185 ;
  assign n5187 = n5184 | n5185 ;
  assign n5188 = ~n5186 & n5187 ;
  assign n5189 = n4883 | n4886 ;
  assign n5190 = ( n5115 & n5188 ) | ( n5115 & n5189 ) | ( n5188 & n5189 ) ;
  assign n5191 = ( n5188 & n5189 ) | ( n5188 & ~n5190 ) | ( n5189 & ~n5190 ) ;
  assign n5192 = ( n5115 & ~n5190 ) | ( n5115 & n5191 ) | ( ~n5190 & n5191 ) ;
  assign n5193 = n5104 & n5192 ;
  assign n5194 = n5104 | n5192 ;
  assign n5195 = ~n5193 & n5194 ;
  assign n5196 = n5093 | n5195 ;
  assign n5197 = n5093 & n5195 ;
  assign n5198 = n5196 & ~n5197 ;
  assign n5199 = x85 & n1421 ;
  assign n5200 = x84 & n1416 ;
  assign n5201 = x83 & ~n1415 ;
  assign n5202 = n1584 & n5201 ;
  assign n5203 = n5200 | n5202 ;
  assign n5204 = n5199 | n5203 ;
  assign n5205 = n1424 | n5204 ;
  assign n5206 = ( n1765 & n5204 ) | ( n1765 & n5205 ) | ( n5204 & n5205 ) ;
  assign n5207 = x20 & n5206 ;
  assign n5208 = x20 & ~n5207 ;
  assign n5209 = ( n5206 & ~n5207 ) | ( n5206 & n5208 ) | ( ~n5207 & n5208 ) ;
  assign n5210 = n5198 & n5209 ;
  assign n5211 = n5198 & ~n5210 ;
  assign n5212 = ~n5198 & n5209 ;
  assign n5213 = n5211 | n5212 ;
  assign n5214 = n4919 | n4925 ;
  assign n5215 = n5213 | n5214 ;
  assign n5216 = n5213 & n5214 ;
  assign n5217 = n5215 & ~n5216 ;
  assign n5218 = x88 & n1071 ;
  assign n5219 = x87 & n1066 ;
  assign n5220 = x86 & ~n1065 ;
  assign n5221 = n1189 & n5220 ;
  assign n5222 = n5219 | n5221 ;
  assign n5223 = n5218 | n5222 ;
  assign n5224 = n1074 | n5223 ;
  assign n5225 = ( n2095 & n5223 ) | ( n2095 & n5224 ) | ( n5223 & n5224 ) ;
  assign n5226 = x17 & n5225 ;
  assign n5227 = x17 & ~n5226 ;
  assign n5228 = ( n5225 & ~n5226 ) | ( n5225 & n5227 ) | ( ~n5226 & n5227 ) ;
  assign n5229 = n5217 | n5228 ;
  assign n5230 = n5217 & n5228 ;
  assign n5231 = n5229 & ~n5230 ;
  assign n5232 = n5092 & n5231 ;
  assign n5233 = n5092 | n5231 ;
  assign n5234 = ~n5232 & n5233 ;
  assign n5235 = ( n5090 & n5091 ) | ( n5090 & ~n5234 ) | ( n5091 & ~n5234 ) ;
  assign n5236 = ( ~n5091 & n5234 ) | ( ~n5091 & n5235 ) | ( n5234 & n5235 ) ;
  assign n5237 = ( ~n5090 & n5235 ) | ( ~n5090 & n5236 ) | ( n5235 & n5236 ) ;
  assign n5238 = n5079 & n5237 ;
  assign n5239 = n5079 | n5237 ;
  assign n5240 = ~n5238 & n5239 ;
  assign n5241 = n4974 | n4976 ;
  assign n5242 = n5240 & n5241 ;
  assign n5243 = n5240 | n5241 ;
  assign n5244 = ~n5242 & n5243 ;
  assign n5245 = ( n5067 & n5068 ) | ( n5067 & ~n5244 ) | ( n5068 & ~n5244 ) ;
  assign n5246 = ( ~n5068 & n5244 ) | ( ~n5068 & n5245 ) | ( n5244 & n5245 ) ;
  assign n5247 = ( ~n5067 & n5245 ) | ( ~n5067 & n5246 ) | ( n5245 & n5246 ) ;
  assign n5248 = n5056 | n5247 ;
  assign n5249 = n5056 & n5247 ;
  assign n5250 = n5248 & ~n5249 ;
  assign n5251 = n5045 & n5250 ;
  assign n5252 = n5045 | n5250 ;
  assign n5253 = ~n5251 & n5252 ;
  assign n5254 = x102 | x103 ;
  assign n5255 = x102 & x103 ;
  assign n5256 = n5254 & ~n5255 ;
  assign n5257 = n5016 | n5019 ;
  assign n5258 = n5256 & n5257 ;
  assign n5259 = n5016 | n5021 ;
  assign n5260 = n5256 & n5259 ;
  assign n5261 = ( n4323 & n5258 ) | ( n4323 & n5260 ) | ( n5258 & n5260 ) ;
  assign n5262 = ( n4323 & n5257 ) | ( n4323 & n5259 ) | ( n5257 & n5259 ) ;
  assign n5263 = n5256 | n5262 ;
  assign n5264 = ~n5261 & n5263 ;
  assign n5265 = x102 & n131 ;
  assign n5266 = x101 & ~n156 ;
  assign n5267 = ( n135 & n5265 ) | ( n135 & n5266 ) | ( n5265 & n5266 ) ;
  assign n5268 = x0 & x103 ;
  assign n5269 = ( ~n135 & n5265 ) | ( ~n135 & n5268 ) | ( n5265 & n5268 ) ;
  assign n5270 = n5267 | n5269 ;
  assign n5271 = n139 | n5270 ;
  assign n5272 = ( n5264 & n5270 ) | ( n5264 & n5271 ) | ( n5270 & n5271 ) ;
  assign n5273 = x2 & n5272 ;
  assign n5274 = x2 & ~n5273 ;
  assign n5275 = ( n5272 & ~n5273 ) | ( n5272 & n5274 ) | ( ~n5273 & n5274 ) ;
  assign n5276 = n5253 & n5275 ;
  assign n5277 = n5253 & ~n5276 ;
  assign n5278 = ~n5253 & n5275 ;
  assign n5279 = n5277 | n5278 ;
  assign n5280 = n5037 | n5042 ;
  assign n5281 = n5279 & n5280 ;
  assign n5282 = n5279 | n5280 ;
  assign n5283 = ~n5281 & n5282 ;
  assign n5284 = n5276 | n5281 ;
  assign n5285 = x103 | x104 ;
  assign n5286 = x103 & x104 ;
  assign n5287 = n5285 & ~n5286 ;
  assign n5288 = n5255 | n5258 ;
  assign n5289 = n5287 & n5288 ;
  assign n5290 = n5255 | n5260 ;
  assign n5291 = n5287 & n5290 ;
  assign n5292 = ( n4323 & n5289 ) | ( n4323 & n5291 ) | ( n5289 & n5291 ) ;
  assign n5293 = ( n4323 & n5288 ) | ( n4323 & n5290 ) | ( n5288 & n5290 ) ;
  assign n5294 = n5287 | n5293 ;
  assign n5295 = ~n5292 & n5294 ;
  assign n5296 = x103 & n131 ;
  assign n5297 = x102 & ~n156 ;
  assign n5298 = ( n135 & n5296 ) | ( n135 & n5297 ) | ( n5296 & n5297 ) ;
  assign n5299 = x0 & x104 ;
  assign n5300 = ( ~n135 & n5296 ) | ( ~n135 & n5299 ) | ( n5296 & n5299 ) ;
  assign n5301 = n5298 | n5300 ;
  assign n5302 = n139 | n5301 ;
  assign n5303 = ( n5295 & n5301 ) | ( n5295 & n5302 ) | ( n5301 & n5302 ) ;
  assign n5304 = x2 & n5303 ;
  assign n5305 = x2 & ~n5304 ;
  assign n5306 = ( n5303 & ~n5304 ) | ( n5303 & n5305 ) | ( ~n5304 & n5305 ) ;
  assign n5307 = x101 & n206 ;
  assign n5308 = x100 & n201 ;
  assign n5309 = x99 & ~n200 ;
  assign n5310 = n243 & n5309 ;
  assign n5311 = n5308 | n5310 ;
  assign n5312 = n5307 | n5311 ;
  assign n5313 = n209 | n5312 ;
  assign n5314 = ( n4783 & n5312 ) | ( n4783 & n5313 ) | ( n5312 & n5313 ) ;
  assign n5315 = x5 & n5314 ;
  assign n5316 = x5 & ~n5315 ;
  assign n5317 = ( n5314 & ~n5315 ) | ( n5314 & n5316 ) | ( ~n5315 & n5316 ) ;
  assign n5318 = n5238 | n5242 ;
  assign n5319 = x95 & n528 ;
  assign n5320 = x94 & n523 ;
  assign n5321 = x93 & ~n522 ;
  assign n5322 = n635 & n5321 ;
  assign n5323 = n5320 | n5322 ;
  assign n5324 = n5319 | n5323 ;
  assign n5325 = n531 | n5324 ;
  assign n5326 = ( n3479 & n5324 ) | ( n3479 & n5325 ) | ( n5324 & n5325 ) ;
  assign n5327 = x11 & n5326 ;
  assign n5328 = x11 & ~n5327 ;
  assign n5329 = ( n5326 & ~n5327 ) | ( n5326 & n5328 ) | ( ~n5327 & n5328 ) ;
  assign n5330 = ( n5090 & n5091 ) | ( n5090 & n5234 ) | ( n5091 & n5234 ) ;
  assign n5331 = n5163 | n5169 ;
  assign n5332 = ~x39 & x40 ;
  assign n5333 = x39 & ~x40 ;
  assign n5334 = n5332 | n5333 ;
  assign n5335 = ~n5118 & n5334 ;
  assign n5336 = x64 & n5335 ;
  assign n5337 = ~x40 & x41 ;
  assign n5338 = x40 & ~x41 ;
  assign n5339 = n5337 | n5338 ;
  assign n5340 = n5118 & ~n5339 ;
  assign n5341 = x65 & n5340 ;
  assign n5342 = n5336 | n5341 ;
  assign n5343 = n5118 & n5339 ;
  assign n5344 = n142 & n5343 ;
  assign n5345 = n5342 | n5344 ;
  assign n5346 = x41 | n5345 ;
  assign n5347 = ~x41 & n5346 ;
  assign n5348 = ( ~n5345 & n5346 ) | ( ~n5345 & n5347 ) | ( n5346 & n5347 ) ;
  assign n5349 = x41 & ~n5119 ;
  assign n5350 = n5348 & n5349 ;
  assign n5351 = n5348 | n5349 ;
  assign n5352 = ~n5350 & n5351 ;
  assign n5353 = n229 & n4575 ;
  assign n5354 = x68 & n4572 ;
  assign n5355 = x67 & n4567 ;
  assign n5356 = x66 & ~n4566 ;
  assign n5357 = n4828 & n5356 ;
  assign n5358 = n5355 | n5357 ;
  assign n5359 = n5354 | n5358 ;
  assign n5360 = n5353 | n5359 ;
  assign n5361 = x38 | n5360 ;
  assign n5362 = ~x38 & n5361 ;
  assign n5363 = ( ~n5360 & n5361 ) | ( ~n5360 & n5362 ) | ( n5361 & n5362 ) ;
  assign n5364 = n5352 | n5363 ;
  assign n5365 = n5352 & n5363 ;
  assign n5366 = n5364 & ~n5365 ;
  assign n5367 = n5131 | n5366 ;
  assign n5368 = n5131 & n5366 ;
  assign n5369 = n5367 & ~n5368 ;
  assign n5370 = x71 & n3913 ;
  assign n5371 = x70 & n3908 ;
  assign n5372 = x69 & ~n3907 ;
  assign n5373 = n4152 & n5372 ;
  assign n5374 = n5371 | n5373 ;
  assign n5375 = n5370 | n5374 ;
  assign n5376 = n3916 | n5375 ;
  assign n5377 = ( n376 & n5375 ) | ( n376 & n5376 ) | ( n5375 & n5376 ) ;
  assign n5378 = x35 & ~n5377 ;
  assign n5379 = ~x35 & n5377 ;
  assign n5380 = n5378 | n5379 ;
  assign n5381 = n5369 & n5380 ;
  assign n5382 = n5369 & ~n5381 ;
  assign n5383 = ~n5369 & n5380 ;
  assign n5384 = n5382 | n5383 ;
  assign n5385 = n5145 | n5150 ;
  assign n5386 = n5384 | n5385 ;
  assign n5387 = n5384 & n5385 ;
  assign n5388 = n5386 & ~n5387 ;
  assign n5389 = x74 & n3314 ;
  assign n5390 = x73 & n3309 ;
  assign n5391 = x72 & ~n3308 ;
  assign n5392 = n3570 & n5391 ;
  assign n5393 = n5390 | n5392 ;
  assign n5394 = n5389 | n5393 ;
  assign n5395 = n3317 | n5394 ;
  assign n5396 = ( n587 & n5394 ) | ( n587 & n5395 ) | ( n5394 & n5395 ) ;
  assign n5397 = x32 & n5396 ;
  assign n5398 = x32 & ~n5397 ;
  assign n5399 = ( n5396 & ~n5397 ) | ( n5396 & n5398 ) | ( ~n5397 & n5398 ) ;
  assign n5400 = n5388 | n5399 ;
  assign n5401 = n5331 & n5400 ;
  assign n5402 = n5388 & n5399 ;
  assign n5403 = n5400 & ~n5402 ;
  assign n5404 = ~n5401 & n5403 ;
  assign n5405 = x77 & n2775 ;
  assign n5406 = x76 & n2770 ;
  assign n5407 = x75 & ~n2769 ;
  assign n5408 = n2978 & n5407 ;
  assign n5409 = n5406 | n5408 ;
  assign n5410 = n5405 | n5409 ;
  assign n5411 = n2778 | n5410 ;
  assign n5412 = ( n846 & n5410 ) | ( n846 & n5411 ) | ( n5410 & n5411 ) ;
  assign n5413 = x29 & n5412 ;
  assign n5414 = x29 & ~n5413 ;
  assign n5415 = ( n5412 & ~n5413 ) | ( n5412 & n5414 ) | ( ~n5413 & n5414 ) ;
  assign n5416 = n5404 | n5415 ;
  assign n5417 = n5331 & ~n5403 ;
  assign n5418 = n5416 | n5417 ;
  assign n5419 = ( n5404 & n5415 ) | ( n5404 & n5417 ) | ( n5415 & n5417 ) ;
  assign n5420 = n5418 & ~n5419 ;
  assign n5421 = n5183 | n5186 ;
  assign n5422 = n5420 & n5421 ;
  assign n5423 = n5420 | n5421 ;
  assign n5424 = ~n5422 & n5423 ;
  assign n5425 = x80 & n2280 ;
  assign n5426 = x79 & n2275 ;
  assign n5427 = x78 & ~n2274 ;
  assign n5428 = n2481 & n5427 ;
  assign n5429 = n5426 | n5428 ;
  assign n5430 = n5425 | n5429 ;
  assign n5431 = n2283 | n5430 ;
  assign n5432 = ( n1147 & n5430 ) | ( n1147 & n5431 ) | ( n5430 & n5431 ) ;
  assign n5433 = x26 & n5432 ;
  assign n5434 = x26 & ~n5433 ;
  assign n5435 = ( n5432 & ~n5433 ) | ( n5432 & n5434 ) | ( ~n5433 & n5434 ) ;
  assign n5436 = n5424 & n5435 ;
  assign n5437 = n5424 & ~n5436 ;
  assign n5438 = ~n5424 & n5435 ;
  assign n5439 = n5437 | n5438 ;
  assign n5440 = n5190 | n5439 ;
  assign n5441 = n5190 & n5439 ;
  assign n5442 = n5440 & ~n5441 ;
  assign n5443 = x83 & n1817 ;
  assign n5444 = x82 & n1812 ;
  assign n5445 = x81 & ~n1811 ;
  assign n5446 = n1977 & n5445 ;
  assign n5447 = n5444 | n5446 ;
  assign n5448 = n5443 | n5447 ;
  assign n5449 = n1820 | n5448 ;
  assign n5450 = ( n1510 & n5448 ) | ( n1510 & n5449 ) | ( n5448 & n5449 ) ;
  assign n5451 = x23 & n5450 ;
  assign n5452 = x23 & ~n5451 ;
  assign n5453 = ( n5450 & ~n5451 ) | ( n5450 & n5452 ) | ( ~n5451 & n5452 ) ;
  assign n5454 = n5442 & n5453 ;
  assign n5455 = n5442 & ~n5454 ;
  assign n5456 = ~n5442 & n5453 ;
  assign n5457 = n5455 | n5456 ;
  assign n5458 = n5193 | n5197 ;
  assign n5459 = n5457 | n5458 ;
  assign n5460 = n5457 & n5458 ;
  assign n5461 = n5459 & ~n5460 ;
  assign n5462 = x86 & n1421 ;
  assign n5463 = x85 & n1416 ;
  assign n5464 = x84 & ~n1415 ;
  assign n5465 = n1584 & n5464 ;
  assign n5466 = n5463 | n5465 ;
  assign n5467 = n5462 | n5466 ;
  assign n5468 = n1424 | n5467 ;
  assign n5469 = ( n1921 & n5467 ) | ( n1921 & n5468 ) | ( n5467 & n5468 ) ;
  assign n5470 = x20 & n5469 ;
  assign n5471 = x20 & ~n5470 ;
  assign n5472 = ( n5469 & ~n5470 ) | ( n5469 & n5471 ) | ( ~n5470 & n5471 ) ;
  assign n5473 = n5461 & n5472 ;
  assign n5474 = n5461 & ~n5473 ;
  assign n5475 = ~n5461 & n5472 ;
  assign n5476 = n5474 | n5475 ;
  assign n5477 = n5210 | n5216 ;
  assign n5478 = n5476 | n5477 ;
  assign n5479 = n5476 & n5477 ;
  assign n5480 = n5478 & ~n5479 ;
  assign n5481 = x89 & n1071 ;
  assign n5482 = x88 & n1066 ;
  assign n5483 = x87 & ~n1065 ;
  assign n5484 = n1189 & n5483 ;
  assign n5485 = n5482 | n5484 ;
  assign n5486 = n5481 | n5485 ;
  assign n5487 = n1074 | n5486 ;
  assign n5488 = ( n2244 & n5486 ) | ( n2244 & n5487 ) | ( n5486 & n5487 ) ;
  assign n5489 = x17 & n5488 ;
  assign n5490 = x17 & ~n5489 ;
  assign n5491 = ( n5488 & ~n5489 ) | ( n5488 & n5490 ) | ( ~n5489 & n5490 ) ;
  assign n5492 = n5480 & n5491 ;
  assign n5493 = n5480 & ~n5492 ;
  assign n5494 = ~n5480 & n5491 ;
  assign n5495 = n5493 | n5494 ;
  assign n5496 = n5230 | n5232 ;
  assign n5497 = n5495 & n5496 ;
  assign n5498 = n5495 | n5496 ;
  assign n5499 = ~n5497 & n5498 ;
  assign n5500 = x92 & n771 ;
  assign n5501 = x91 & n766 ;
  assign n5502 = x90 & ~n765 ;
  assign n5503 = n905 & n5502 ;
  assign n5504 = n5501 | n5503 ;
  assign n5505 = n5500 | n5504 ;
  assign n5506 = n774 | n5505 ;
  assign n5507 = ( n2904 & n5505 ) | ( n2904 & n5506 ) | ( n5505 & n5506 ) ;
  assign n5508 = x14 & n5507 ;
  assign n5509 = x14 & ~n5508 ;
  assign n5510 = ( n5507 & ~n5508 ) | ( n5507 & n5509 ) | ( ~n5508 & n5509 ) ;
  assign n5511 = n5499 & n5510 ;
  assign n5512 = n5499 & ~n5511 ;
  assign n5513 = ~n5499 & n5510 ;
  assign n5514 = n5512 | n5513 ;
  assign n5515 = n5330 & n5514 ;
  assign n5516 = n5514 & ~n5515 ;
  assign n5517 = ( n5330 & ~n5515 ) | ( n5330 & n5516 ) | ( ~n5515 & n5516 ) ;
  assign n5518 = n5329 | n5517 ;
  assign n5519 = n5329 & n5517 ;
  assign n5520 = n5518 & ~n5519 ;
  assign n5521 = n5318 & n5520 ;
  assign n5522 = n5318 | n5520 ;
  assign n5523 = ~n5521 & n5522 ;
  assign n5524 = x98 & n337 ;
  assign n5525 = x97 & n332 ;
  assign n5526 = x96 & ~n331 ;
  assign n5527 = n396 & n5526 ;
  assign n5528 = n5525 | n5527 ;
  assign n5529 = n5524 | n5528 ;
  assign n5530 = n340 | n5529 ;
  assign n5531 = ( n4105 & n5529 ) | ( n4105 & n5530 ) | ( n5529 & n5530 ) ;
  assign n5532 = x8 & n5531 ;
  assign n5533 = x8 & ~n5532 ;
  assign n5534 = ( n5531 & ~n5532 ) | ( n5531 & n5533 ) | ( ~n5532 & n5533 ) ;
  assign n5535 = n5523 | n5534 ;
  assign n5536 = n5523 & n5534 ;
  assign n5537 = n5535 & ~n5536 ;
  assign n5538 = ( n5067 & n5068 ) | ( n5067 & n5244 ) | ( n5068 & n5244 ) ;
  assign n5539 = n5537 | n5538 ;
  assign n5540 = n5537 & n5538 ;
  assign n5541 = n5539 & ~n5540 ;
  assign n5542 = n5249 | n5251 ;
  assign n5543 = ( n5317 & n5541 ) | ( n5317 & n5542 ) | ( n5541 & n5542 ) ;
  assign n5544 = ( n5541 & n5542 ) | ( n5541 & ~n5543 ) | ( n5542 & ~n5543 ) ;
  assign n5545 = ( n5317 & ~n5543 ) | ( n5317 & n5544 ) | ( ~n5543 & n5544 ) ;
  assign n5546 = n5306 & n5545 ;
  assign n5547 = n5306 | n5545 ;
  assign n5548 = ~n5546 & n5547 ;
  assign n5549 = n5284 & n5548 ;
  assign n5550 = n5284 | n5548 ;
  assign n5551 = ~n5549 & n5550 ;
  assign n5552 = x102 & n206 ;
  assign n5553 = x101 & n201 ;
  assign n5554 = x100 & ~n200 ;
  assign n5555 = n243 & n5554 ;
  assign n5556 = n5553 | n5555 ;
  assign n5557 = n5552 | n5556 ;
  assign n5558 = n209 | n5557 ;
  assign n5559 = ( n5025 & n5557 ) | ( n5025 & n5558 ) | ( n5557 & n5558 ) ;
  assign n5560 = x5 & n5559 ;
  assign n5561 = x5 & ~n5560 ;
  assign n5562 = ( n5559 & ~n5560 ) | ( n5559 & n5561 ) | ( ~n5560 & n5561 ) ;
  assign n5563 = x99 & n337 ;
  assign n5564 = x98 & n332 ;
  assign n5565 = x97 & ~n331 ;
  assign n5566 = n396 & n5565 ;
  assign n5567 = n5564 | n5566 ;
  assign n5568 = n5563 | n5567 ;
  assign n5569 = n340 | n5568 ;
  assign n5570 = ( n4325 & n5568 ) | ( n4325 & n5569 ) | ( n5568 & n5569 ) ;
  assign n5571 = x8 & n5570 ;
  assign n5572 = x8 & ~n5571 ;
  assign n5573 = ( n5570 & ~n5571 ) | ( n5570 & n5572 ) | ( ~n5571 & n5572 ) ;
  assign n5574 = n5536 | n5540 ;
  assign n5575 = n5436 | n5441 ;
  assign n5576 = n5419 | n5422 ;
  assign n5577 = n5381 | n5387 ;
  assign n5578 = x66 & n5340 ;
  assign n5579 = x65 & n5335 ;
  assign n5580 = ~n5118 & n5339 ;
  assign n5581 = x64 & ~n5334 ;
  assign n5582 = n5580 & n5581 ;
  assign n5583 = n5579 | n5582 ;
  assign n5584 = n5578 | n5583 ;
  assign n5585 = n153 & n5343 ;
  assign n5586 = n5584 | n5585 ;
  assign n5587 = x41 | n5586 ;
  assign n5588 = ~x41 & n5587 ;
  assign n5589 = ( ~n5586 & n5587 ) | ( ~n5586 & n5588 ) | ( n5587 & n5588 ) ;
  assign n5590 = n5350 | n5589 ;
  assign n5591 = n5350 & n5589 ;
  assign n5592 = n5590 & ~n5591 ;
  assign n5593 = n264 & n4575 ;
  assign n5594 = x69 & n4572 ;
  assign n5595 = x68 & n4567 ;
  assign n5596 = x67 & ~n4566 ;
  assign n5597 = n4828 & n5596 ;
  assign n5598 = n5595 | n5597 ;
  assign n5599 = n5594 | n5598 ;
  assign n5600 = n5593 | n5599 ;
  assign n5601 = x38 | n5600 ;
  assign n5602 = ~x38 & n5601 ;
  assign n5603 = ( ~n5600 & n5601 ) | ( ~n5600 & n5602 ) | ( n5601 & n5602 ) ;
  assign n5604 = n5592 & n5603 ;
  assign n5605 = n5592 & ~n5604 ;
  assign n5606 = ~n5592 & n5603 ;
  assign n5607 = n5605 | n5606 ;
  assign n5608 = n5365 | n5368 ;
  assign n5609 = n5607 & n5608 ;
  assign n5610 = n5607 | n5608 ;
  assign n5611 = ~n5609 & n5610 ;
  assign n5612 = x72 & n3913 ;
  assign n5613 = x71 & n3908 ;
  assign n5614 = x70 & ~n3907 ;
  assign n5615 = n4152 & n5614 ;
  assign n5616 = n5613 | n5615 ;
  assign n5617 = n5612 | n5616 ;
  assign n5618 = ( n435 & n3916 ) | ( n435 & n5617 ) | ( n3916 & n5617 ) ;
  assign n5619 = ( x35 & ~n5617 ) | ( x35 & n5618 ) | ( ~n5617 & n5618 ) ;
  assign n5620 = ~n5618 & n5619 ;
  assign n5621 = n5617 | n5619 ;
  assign n5622 = ( ~x35 & n5620 ) | ( ~x35 & n5621 ) | ( n5620 & n5621 ) ;
  assign n5623 = ~n5611 & n5622 ;
  assign n5624 = n5611 & ~n5622 ;
  assign n5625 = n5623 | n5624 ;
  assign n5626 = n5577 & ~n5625 ;
  assign n5627 = ~n5577 & n5625 ;
  assign n5628 = x75 & n3314 ;
  assign n5629 = x74 & n3309 ;
  assign n5630 = x73 & ~n3308 ;
  assign n5631 = n3570 & n5630 ;
  assign n5632 = n5629 | n5631 ;
  assign n5633 = n5628 | n5632 ;
  assign n5634 = n3317 | n5633 ;
  assign n5635 = ( n609 & n5633 ) | ( n609 & n5634 ) | ( n5633 & n5634 ) ;
  assign n5636 = x32 & n5635 ;
  assign n5637 = x32 & ~n5636 ;
  assign n5638 = ( n5635 & ~n5636 ) | ( n5635 & n5637 ) | ( ~n5636 & n5637 ) ;
  assign n5639 = n5627 | n5638 ;
  assign n5640 = n5626 | n5639 ;
  assign n5641 = ( n5626 & n5627 ) | ( n5626 & n5638 ) | ( n5627 & n5638 ) ;
  assign n5642 = n5640 & ~n5641 ;
  assign n5643 = n5401 | n5402 ;
  assign n5644 = n5642 & n5643 ;
  assign n5645 = n5642 | n5643 ;
  assign n5646 = ~n5644 & n5645 ;
  assign n5647 = x78 & n2775 ;
  assign n5648 = x77 & n2770 ;
  assign n5649 = x76 & ~n2769 ;
  assign n5650 = n2978 & n5649 ;
  assign n5651 = n5648 | n5650 ;
  assign n5652 = n5647 | n5651 ;
  assign n5653 = n2778 | n5652 ;
  assign n5654 = ( n868 & n5652 ) | ( n868 & n5653 ) | ( n5652 & n5653 ) ;
  assign n5655 = x29 & n5654 ;
  assign n5656 = x29 & ~n5655 ;
  assign n5657 = ( n5654 & ~n5655 ) | ( n5654 & n5656 ) | ( ~n5655 & n5656 ) ;
  assign n5658 = n5646 | n5657 ;
  assign n5659 = n5646 & n5657 ;
  assign n5660 = n5658 & ~n5659 ;
  assign n5661 = n5576 & n5660 ;
  assign n5662 = n5576 | n5660 ;
  assign n5663 = ~n5661 & n5662 ;
  assign n5664 = x81 & n2280 ;
  assign n5665 = x80 & n2275 ;
  assign n5666 = x79 & ~n2274 ;
  assign n5667 = n2481 & n5666 ;
  assign n5668 = n5665 | n5667 ;
  assign n5669 = n5664 | n5668 ;
  assign n5670 = n2283 | n5669 ;
  assign n5671 = ( n1256 & n5669 ) | ( n1256 & n5670 ) | ( n5669 & n5670 ) ;
  assign n5672 = x26 & n5671 ;
  assign n5673 = x26 & ~n5672 ;
  assign n5674 = ( n5671 & ~n5672 ) | ( n5671 & n5673 ) | ( ~n5672 & n5673 ) ;
  assign n5675 = n5663 | n5674 ;
  assign n5676 = n5663 & n5674 ;
  assign n5677 = n5675 & ~n5676 ;
  assign n5678 = n5575 & n5677 ;
  assign n5679 = n5575 | n5677 ;
  assign n5680 = ~n5678 & n5679 ;
  assign n5681 = x84 & n1817 ;
  assign n5682 = x83 & n1812 ;
  assign n5683 = x82 & ~n1811 ;
  assign n5684 = n1977 & n5683 ;
  assign n5685 = n5682 | n5684 ;
  assign n5686 = n5681 | n5685 ;
  assign n5687 = n1820 | n5686 ;
  assign n5688 = ( n1537 & n5686 ) | ( n1537 & n5687 ) | ( n5686 & n5687 ) ;
  assign n5689 = x23 & n5688 ;
  assign n5690 = x23 & ~n5689 ;
  assign n5691 = ( n5688 & ~n5689 ) | ( n5688 & n5690 ) | ( ~n5689 & n5690 ) ;
  assign n5692 = n5680 & n5691 ;
  assign n5693 = n5680 & ~n5692 ;
  assign n5694 = ~n5680 & n5691 ;
  assign n5695 = n5693 | n5694 ;
  assign n5696 = n5454 | n5460 ;
  assign n5697 = n5695 | n5696 ;
  assign n5698 = n5695 & n5696 ;
  assign n5699 = n5697 & ~n5698 ;
  assign n5700 = x87 & n1421 ;
  assign n5701 = x86 & n1416 ;
  assign n5702 = x85 & ~n1415 ;
  assign n5703 = n1584 & n5702 ;
  assign n5704 = n5701 | n5703 ;
  assign n5705 = n5700 | n5704 ;
  assign n5706 = n1424 | n5705 ;
  assign n5707 = ( n2067 & n5705 ) | ( n2067 & n5706 ) | ( n5705 & n5706 ) ;
  assign n5708 = x20 & n5707 ;
  assign n5709 = x20 & ~n5708 ;
  assign n5710 = ( n5707 & ~n5708 ) | ( n5707 & n5709 ) | ( ~n5708 & n5709 ) ;
  assign n5711 = n5699 | n5710 ;
  assign n5712 = n5473 | n5479 ;
  assign n5713 = ( n5699 & n5710 ) | ( n5699 & n5712 ) | ( n5710 & n5712 ) ;
  assign n5714 = n5711 & ~n5713 ;
  assign n5715 = n5699 & n5710 ;
  assign n5716 = n5711 & ~n5715 ;
  assign n5717 = n5712 & ~n5716 ;
  assign n5718 = n5714 | n5717 ;
  assign n5719 = x90 & n1071 ;
  assign n5720 = x89 & n1066 ;
  assign n5721 = x88 & ~n1065 ;
  assign n5722 = n1189 & n5721 ;
  assign n5723 = n5720 | n5722 ;
  assign n5724 = n5719 | n5723 ;
  assign n5725 = n1074 | n5724 ;
  assign n5726 = ( n2410 & n5724 ) | ( n2410 & n5725 ) | ( n5724 & n5725 ) ;
  assign n5727 = x17 & n5726 ;
  assign n5728 = x17 & ~n5727 ;
  assign n5729 = ( n5726 & ~n5727 ) | ( n5726 & n5728 ) | ( ~n5727 & n5728 ) ;
  assign n5730 = n5718 | n5729 ;
  assign n5731 = n5718 & n5729 ;
  assign n5732 = n5730 & ~n5731 ;
  assign n5733 = n5492 | n5497 ;
  assign n5734 = n5732 & n5733 ;
  assign n5735 = n5732 | n5733 ;
  assign n5736 = ~n5734 & n5735 ;
  assign n5737 = x93 & n771 ;
  assign n5738 = x92 & n766 ;
  assign n5739 = x91 & ~n765 ;
  assign n5740 = n905 & n5739 ;
  assign n5741 = n5738 | n5740 ;
  assign n5742 = n5737 | n5741 ;
  assign n5743 = n774 | n5742 ;
  assign n5744 = ( n2931 & n5742 ) | ( n2931 & n5743 ) | ( n5742 & n5743 ) ;
  assign n5745 = x14 & n5744 ;
  assign n5746 = x14 & ~n5745 ;
  assign n5747 = ( n5744 & ~n5745 ) | ( n5744 & n5746 ) | ( ~n5745 & n5746 ) ;
  assign n5748 = n5736 | n5747 ;
  assign n5749 = n5736 & n5747 ;
  assign n5750 = n5748 & ~n5749 ;
  assign n5751 = n5511 | n5750 ;
  assign n5752 = n5515 | n5751 ;
  assign n5753 = ( n5511 & n5515 ) | ( n5511 & n5750 ) | ( n5515 & n5750 ) ;
  assign n5754 = n5752 & ~n5753 ;
  assign n5755 = x96 & n528 ;
  assign n5756 = x95 & n523 ;
  assign n5757 = x94 & ~n522 ;
  assign n5758 = n635 & n5757 ;
  assign n5759 = n5756 | n5758 ;
  assign n5760 = n5755 | n5759 ;
  assign n5761 = n531 | n5760 ;
  assign n5762 = ( n3509 & n5760 ) | ( n3509 & n5761 ) | ( n5760 & n5761 ) ;
  assign n5763 = x11 & n5762 ;
  assign n5764 = x11 & ~n5763 ;
  assign n5765 = ( n5762 & ~n5763 ) | ( n5762 & n5764 ) | ( ~n5763 & n5764 ) ;
  assign n5766 = n5754 | n5765 ;
  assign n5767 = n5754 & n5765 ;
  assign n5768 = n5766 & ~n5767 ;
  assign n5769 = n5519 | n5521 ;
  assign n5770 = n5768 & n5769 ;
  assign n5771 = n5768 | n5769 ;
  assign n5772 = ~n5770 & n5771 ;
  assign n5773 = ( n5573 & n5574 ) | ( n5573 & ~n5772 ) | ( n5574 & ~n5772 ) ;
  assign n5774 = ( ~n5574 & n5772 ) | ( ~n5574 & n5773 ) | ( n5772 & n5773 ) ;
  assign n5775 = ( ~n5573 & n5773 ) | ( ~n5573 & n5774 ) | ( n5773 & n5774 ) ;
  assign n5776 = n5562 & n5775 ;
  assign n5777 = n5562 | n5775 ;
  assign n5778 = ~n5776 & n5777 ;
  assign n5779 = n5543 | n5778 ;
  assign n5780 = n5543 & n5778 ;
  assign n5781 = n5779 & ~n5780 ;
  assign n5782 = x104 | x105 ;
  assign n5783 = x104 & x105 ;
  assign n5784 = n5782 & ~n5783 ;
  assign n5785 = n5286 | n5292 ;
  assign n5786 = n5784 & n5785 ;
  assign n5787 = n5784 | n5785 ;
  assign n5788 = ~n5786 & n5787 ;
  assign n5789 = x104 & n131 ;
  assign n5790 = x103 & ~n156 ;
  assign n5791 = ( n135 & n5789 ) | ( n135 & n5790 ) | ( n5789 & n5790 ) ;
  assign n5792 = x0 & x105 ;
  assign n5793 = ( ~n135 & n5789 ) | ( ~n135 & n5792 ) | ( n5789 & n5792 ) ;
  assign n5794 = n5791 | n5793 ;
  assign n5795 = n139 | n5794 ;
  assign n5796 = ( n5788 & n5794 ) | ( n5788 & n5795 ) | ( n5794 & n5795 ) ;
  assign n5797 = x2 & n5796 ;
  assign n5798 = x2 & ~n5797 ;
  assign n5799 = ( n5796 & ~n5797 ) | ( n5796 & n5798 ) | ( ~n5797 & n5798 ) ;
  assign n5800 = n5781 | n5799 ;
  assign n5801 = n5781 & n5799 ;
  assign n5802 = n5800 & ~n5801 ;
  assign n5803 = n5546 | n5549 ;
  assign n5804 = n5802 & n5803 ;
  assign n5805 = n5802 | n5803 ;
  assign n5806 = ~n5804 & n5805 ;
  assign n5807 = x105 | x106 ;
  assign n5808 = x105 & x106 ;
  assign n5809 = n5807 & ~n5808 ;
  assign n5810 = n5783 & n5809 ;
  assign n5811 = ( n5786 & n5809 ) | ( n5786 & n5810 ) | ( n5809 & n5810 ) ;
  assign n5812 = n5783 | n5809 ;
  assign n5813 = n5786 | n5812 ;
  assign n5814 = ~n5811 & n5813 ;
  assign n5815 = x105 & n131 ;
  assign n5816 = x104 & ~n156 ;
  assign n5817 = ( n135 & n5815 ) | ( n135 & n5816 ) | ( n5815 & n5816 ) ;
  assign n5818 = x0 & x106 ;
  assign n5819 = ( ~n135 & n5815 ) | ( ~n135 & n5818 ) | ( n5815 & n5818 ) ;
  assign n5820 = n5817 | n5819 ;
  assign n5821 = n139 | n5820 ;
  assign n5822 = ( n5814 & n5820 ) | ( n5814 & n5821 ) | ( n5820 & n5821 ) ;
  assign n5823 = x2 & n5822 ;
  assign n5824 = x2 & ~n5823 ;
  assign n5825 = ( n5822 & ~n5823 ) | ( n5822 & n5824 ) | ( ~n5823 & n5824 ) ;
  assign n5826 = n5776 | n5780 ;
  assign n5827 = x100 & n337 ;
  assign n5828 = x99 & n332 ;
  assign n5829 = x98 & ~n331 ;
  assign n5830 = n396 & n5829 ;
  assign n5831 = n5828 | n5830 ;
  assign n5832 = n5827 | n5831 ;
  assign n5833 = n340 | n5832 ;
  assign n5834 = ( n4532 & n5832 ) | ( n4532 & n5833 ) | ( n5832 & n5833 ) ;
  assign n5835 = x8 & n5834 ;
  assign n5836 = x8 & ~n5835 ;
  assign n5837 = ( n5834 & ~n5835 ) | ( n5834 & n5836 ) | ( ~n5835 & n5836 ) ;
  assign n5838 = x97 & n528 ;
  assign n5839 = x96 & n523 ;
  assign n5840 = x95 & ~n522 ;
  assign n5841 = n635 & n5840 ;
  assign n5842 = n5839 | n5841 ;
  assign n5843 = n5838 | n5842 ;
  assign n5844 = n531 | n5843 ;
  assign n5845 = ( n3707 & n5843 ) | ( n3707 & n5844 ) | ( n5843 & n5844 ) ;
  assign n5846 = x11 & n5845 ;
  assign n5847 = x11 & ~n5846 ;
  assign n5848 = ( n5845 & ~n5846 ) | ( n5845 & n5847 ) | ( ~n5846 & n5847 ) ;
  assign n5849 = n5749 | n5753 ;
  assign n5850 = x94 & n771 ;
  assign n5851 = x93 & n766 ;
  assign n5852 = x92 & ~n765 ;
  assign n5853 = n905 & n5852 ;
  assign n5854 = n5851 | n5853 ;
  assign n5855 = n5850 | n5854 ;
  assign n5856 = n774 | n5855 ;
  assign n5857 = ( n3271 & n5855 ) | ( n3271 & n5856 ) | ( n5855 & n5856 ) ;
  assign n5858 = x14 & n5857 ;
  assign n5859 = x14 & ~n5858 ;
  assign n5860 = ( n5857 & ~n5858 ) | ( n5857 & n5859 ) | ( ~n5858 & n5859 ) ;
  assign n5861 = x91 & n1071 ;
  assign n5862 = x90 & n1066 ;
  assign n5863 = x89 & ~n1065 ;
  assign n5864 = n1189 & n5863 ;
  assign n5865 = n5862 | n5864 ;
  assign n5866 = n5861 | n5865 ;
  assign n5867 = n1074 | n5866 ;
  assign n5868 = ( n2714 & n5866 ) | ( n2714 & n5867 ) | ( n5866 & n5867 ) ;
  assign n5869 = x17 & n5868 ;
  assign n5870 = x17 & ~n5869 ;
  assign n5871 = ( n5868 & ~n5869 ) | ( n5868 & n5870 ) | ( ~n5869 & n5870 ) ;
  assign n5872 = n5731 | n5734 ;
  assign n5873 = n5659 | n5661 ;
  assign n5874 = n5641 | n5644 ;
  assign n5875 = x41 & ~x42 ;
  assign n5876 = ~x41 & x42 ;
  assign n5877 = n5875 | n5876 ;
  assign n5878 = x64 & n5877 ;
  assign n5879 = x67 & n5340 ;
  assign n5880 = x66 & n5335 ;
  assign n5881 = x65 & ~n5334 ;
  assign n5882 = n5580 & n5881 ;
  assign n5883 = n5880 | n5882 ;
  assign n5884 = n5879 | n5883 ;
  assign n5885 = n180 & n5343 ;
  assign n5886 = n5884 | n5885 ;
  assign n5887 = x41 & ~n5886 ;
  assign n5888 = ~x41 & n5886 ;
  assign n5889 = n5887 | n5888 ;
  assign n5890 = ( n5591 & n5878 ) | ( n5591 & n5889 ) | ( n5878 & n5889 ) ;
  assign n5891 = ( n5591 & n5889 ) | ( n5591 & ~n5890 ) | ( n5889 & ~n5890 ) ;
  assign n5892 = ( n5878 & ~n5890 ) | ( n5878 & n5891 ) | ( ~n5890 & n5891 ) ;
  assign n5893 = x70 & n4572 ;
  assign n5894 = x69 & n4567 ;
  assign n5895 = x68 & ~n4566 ;
  assign n5896 = n4828 & n5895 ;
  assign n5897 = n5894 | n5896 ;
  assign n5898 = n5893 | n5897 ;
  assign n5899 = n4575 | n5898 ;
  assign n5900 = ( n310 & n5898 ) | ( n310 & n5899 ) | ( n5898 & n5899 ) ;
  assign n5901 = x38 & ~n5900 ;
  assign n5902 = ~x38 & n5900 ;
  assign n5903 = n5901 | n5902 ;
  assign n5904 = n5892 & n5903 ;
  assign n5905 = n5892 & ~n5904 ;
  assign n5906 = ~n5892 & n5903 ;
  assign n5907 = n5905 | n5906 ;
  assign n5908 = n5604 | n5609 ;
  assign n5909 = n5907 | n5908 ;
  assign n5910 = n5907 & n5908 ;
  assign n5911 = n5909 & ~n5910 ;
  assign n5912 = x73 & n3913 ;
  assign n5913 = x72 & n3908 ;
  assign n5914 = x71 & ~n3907 ;
  assign n5915 = n4152 & n5914 ;
  assign n5916 = n5913 | n5915 ;
  assign n5917 = n5912 | n5916 ;
  assign n5918 = ( n499 & n3916 ) | ( n499 & n5917 ) | ( n3916 & n5917 ) ;
  assign n5919 = ( x35 & ~n5917 ) | ( x35 & n5918 ) | ( ~n5917 & n5918 ) ;
  assign n5920 = ~n5918 & n5919 ;
  assign n5921 = n5917 | n5919 ;
  assign n5922 = ( ~x35 & n5920 ) | ( ~x35 & n5921 ) | ( n5920 & n5921 ) ;
  assign n5923 = n5911 | n5922 ;
  assign n5924 = n5911 & n5922 ;
  assign n5925 = n5923 & ~n5924 ;
  assign n5926 = ( n5577 & n5611 ) | ( n5577 & n5622 ) | ( n5611 & n5622 ) ;
  assign n5927 = n5925 & n5926 ;
  assign n5928 = n5925 | n5926 ;
  assign n5929 = ~n5927 & n5928 ;
  assign n5930 = x76 & n3314 ;
  assign n5931 = x75 & n3309 ;
  assign n5932 = x74 & ~n3308 ;
  assign n5933 = n3570 & n5932 ;
  assign n5934 = n5931 | n5933 ;
  assign n5935 = n5930 | n5934 ;
  assign n5936 = n3317 | n5935 ;
  assign n5937 = ( n740 & n5935 ) | ( n740 & n5936 ) | ( n5935 & n5936 ) ;
  assign n5938 = x32 & n5937 ;
  assign n5939 = x32 & ~n5938 ;
  assign n5940 = ( n5937 & ~n5938 ) | ( n5937 & n5939 ) | ( ~n5938 & n5939 ) ;
  assign n5941 = n5929 & n5940 ;
  assign n5942 = n5929 & ~n5941 ;
  assign n5943 = ~n5929 & n5940 ;
  assign n5944 = n5942 | n5943 ;
  assign n5945 = n5874 & n5944 ;
  assign n5946 = n5874 & ~n5945 ;
  assign n5947 = n5944 & ~n5945 ;
  assign n5948 = n5946 | n5947 ;
  assign n5949 = x79 & n2775 ;
  assign n5950 = x78 & n2770 ;
  assign n5951 = x77 & ~n2769 ;
  assign n5952 = n2978 & n5951 ;
  assign n5953 = n5950 | n5952 ;
  assign n5954 = n5949 | n5953 ;
  assign n5955 = n2778 | n5954 ;
  assign n5956 = ( n961 & n5954 ) | ( n961 & n5955 ) | ( n5954 & n5955 ) ;
  assign n5957 = x29 & n5956 ;
  assign n5958 = x29 & ~n5957 ;
  assign n5959 = ( n5956 & ~n5957 ) | ( n5956 & n5958 ) | ( ~n5957 & n5958 ) ;
  assign n5960 = ( n5873 & n5948 ) | ( n5873 & ~n5959 ) | ( n5948 & ~n5959 ) ;
  assign n5961 = ( ~n5948 & n5959 ) | ( ~n5948 & n5960 ) | ( n5959 & n5960 ) ;
  assign n5962 = ( ~n5873 & n5960 ) | ( ~n5873 & n5961 ) | ( n5960 & n5961 ) ;
  assign n5963 = x82 & n2280 ;
  assign n5964 = x81 & n2275 ;
  assign n5965 = x80 & ~n2274 ;
  assign n5966 = n2481 & n5965 ;
  assign n5967 = n5964 | n5966 ;
  assign n5968 = n5963 | n5967 ;
  assign n5969 = n2283 | n5968 ;
  assign n5970 = ( n1371 & n5968 ) | ( n1371 & n5969 ) | ( n5968 & n5969 ) ;
  assign n5971 = x26 & n5970 ;
  assign n5972 = x26 & ~n5971 ;
  assign n5973 = ( n5970 & ~n5971 ) | ( n5970 & n5972 ) | ( ~n5971 & n5972 ) ;
  assign n5974 = n5962 & n5973 ;
  assign n5975 = n5962 | n5973 ;
  assign n5976 = ~n5974 & n5975 ;
  assign n5977 = n5676 | n5678 ;
  assign n5978 = n5976 & n5977 ;
  assign n5979 = n5976 | n5977 ;
  assign n5980 = ~n5978 & n5979 ;
  assign n5981 = x85 & n1817 ;
  assign n5982 = x84 & n1812 ;
  assign n5983 = x83 & ~n1811 ;
  assign n5984 = n1977 & n5983 ;
  assign n5985 = n5982 | n5984 ;
  assign n5986 = n5981 | n5985 ;
  assign n5987 = n1820 | n5986 ;
  assign n5988 = ( n1765 & n5986 ) | ( n1765 & n5987 ) | ( n5986 & n5987 ) ;
  assign n5989 = x23 & n5988 ;
  assign n5990 = x23 & ~n5989 ;
  assign n5991 = ( n5988 & ~n5989 ) | ( n5988 & n5990 ) | ( ~n5989 & n5990 ) ;
  assign n5992 = n5980 & n5991 ;
  assign n5993 = n5980 & ~n5992 ;
  assign n5994 = ~n5980 & n5991 ;
  assign n5995 = n5993 | n5994 ;
  assign n5996 = n5692 | n5698 ;
  assign n5997 = n5995 | n5996 ;
  assign n5998 = n5995 & n5996 ;
  assign n5999 = n5997 & ~n5998 ;
  assign n6000 = x88 & n1421 ;
  assign n6001 = x87 & n1416 ;
  assign n6002 = x86 & ~n1415 ;
  assign n6003 = n1584 & n6002 ;
  assign n6004 = n6001 | n6003 ;
  assign n6005 = n6000 | n6004 ;
  assign n6006 = n1424 | n6005 ;
  assign n6007 = ( n2095 & n6005 ) | ( n2095 & n6006 ) | ( n6005 & n6006 ) ;
  assign n6008 = x20 & n6007 ;
  assign n6009 = x20 & ~n6008 ;
  assign n6010 = ( n6007 & ~n6008 ) | ( n6007 & n6009 ) | ( ~n6008 & n6009 ) ;
  assign n6011 = n5999 | n6010 ;
  assign n6012 = n5999 & n6010 ;
  assign n6013 = n6011 & ~n6012 ;
  assign n6014 = n5713 | n6013 ;
  assign n6015 = n5713 & n6013 ;
  assign n6016 = n6014 & ~n6015 ;
  assign n6017 = ( n5871 & n5872 ) | ( n5871 & ~n6016 ) | ( n5872 & ~n6016 ) ;
  assign n6018 = ( ~n5872 & n6016 ) | ( ~n5872 & n6017 ) | ( n6016 & n6017 ) ;
  assign n6019 = ( ~n5871 & n6017 ) | ( ~n5871 & n6018 ) | ( n6017 & n6018 ) ;
  assign n6020 = n5860 & n6019 ;
  assign n6021 = n5860 | n6019 ;
  assign n6022 = ~n6020 & n6021 ;
  assign n6023 = n5849 & n6022 ;
  assign n6024 = n5849 | n6022 ;
  assign n6025 = ~n6023 & n6024 ;
  assign n6026 = n5767 | n5770 ;
  assign n6027 = ( n5848 & n6025 ) | ( n5848 & n6026 ) | ( n6025 & n6026 ) ;
  assign n6028 = ( n6025 & n6026 ) | ( n6025 & ~n6027 ) | ( n6026 & ~n6027 ) ;
  assign n6029 = ( n5848 & ~n6027 ) | ( n5848 & n6028 ) | ( ~n6027 & n6028 ) ;
  assign n6030 = n5837 | n6029 ;
  assign n6031 = n5837 & n6029 ;
  assign n6032 = n6030 & ~n6031 ;
  assign n6033 = ( n5573 & n5574 ) | ( n5573 & n5772 ) | ( n5574 & n5772 ) ;
  assign n6034 = n6032 | n6033 ;
  assign n6035 = n6032 & n6033 ;
  assign n6036 = n6034 & ~n6035 ;
  assign n6037 = x103 & n206 ;
  assign n6038 = x102 & n201 ;
  assign n6039 = x101 & ~n200 ;
  assign n6040 = n243 & n6039 ;
  assign n6041 = n6038 | n6040 ;
  assign n6042 = n6037 | n6041 ;
  assign n6043 = n209 | n6042 ;
  assign n6044 = ( n5264 & n6042 ) | ( n5264 & n6043 ) | ( n6042 & n6043 ) ;
  assign n6045 = x5 & n6044 ;
  assign n6046 = x5 & ~n6045 ;
  assign n6047 = ( n6044 & ~n6045 ) | ( n6044 & n6046 ) | ( ~n6045 & n6046 ) ;
  assign n6048 = ( n5826 & n6036 ) | ( n5826 & ~n6047 ) | ( n6036 & ~n6047 ) ;
  assign n6049 = ( ~n6036 & n6047 ) | ( ~n6036 & n6048 ) | ( n6047 & n6048 ) ;
  assign n6050 = ( ~n5826 & n6048 ) | ( ~n5826 & n6049 ) | ( n6048 & n6049 ) ;
  assign n6051 = n5825 & n6050 ;
  assign n6052 = n5825 | n6050 ;
  assign n6053 = ~n6051 & n6052 ;
  assign n6054 = n5801 | n5804 ;
  assign n6055 = n6053 & n6054 ;
  assign n6056 = n6053 | n6054 ;
  assign n6057 = ~n6055 & n6056 ;
  assign n6058 = n5941 | n5945 ;
  assign n6059 = n5924 | n5927 ;
  assign n6060 = ~x42 & x43 ;
  assign n6061 = x42 & ~x43 ;
  assign n6062 = n6060 | n6061 ;
  assign n6063 = ~n5877 & n6062 ;
  assign n6064 = x64 & n6063 ;
  assign n6065 = ~x43 & x44 ;
  assign n6066 = x43 & ~x44 ;
  assign n6067 = n6065 | n6066 ;
  assign n6068 = n5877 & ~n6067 ;
  assign n6069 = x65 & n6068 ;
  assign n6070 = n6064 | n6069 ;
  assign n6071 = n5877 & n6067 ;
  assign n6072 = n142 & n6071 ;
  assign n6073 = n6070 | n6072 ;
  assign n6074 = x44 | n6073 ;
  assign n6075 = ~x44 & n6074 ;
  assign n6076 = ( ~n6073 & n6074 ) | ( ~n6073 & n6075 ) | ( n6074 & n6075 ) ;
  assign n6077 = x44 & ~n5878 ;
  assign n6078 = n6076 & n6077 ;
  assign n6079 = n6076 | n6077 ;
  assign n6080 = ~n6078 & n6079 ;
  assign n6081 = n229 & n5343 ;
  assign n6082 = x68 & n5340 ;
  assign n6083 = x67 & n5335 ;
  assign n6084 = x66 & ~n5334 ;
  assign n6085 = n5580 & n6084 ;
  assign n6086 = n6083 | n6085 ;
  assign n6087 = n6082 | n6086 ;
  assign n6088 = n6081 | n6087 ;
  assign n6089 = x41 | n6088 ;
  assign n6090 = ~x41 & n6089 ;
  assign n6091 = ( ~n6088 & n6089 ) | ( ~n6088 & n6090 ) | ( n6089 & n6090 ) ;
  assign n6092 = n6080 | n6091 ;
  assign n6093 = n6080 & n6091 ;
  assign n6094 = n6092 & ~n6093 ;
  assign n6095 = n5890 | n6094 ;
  assign n6096 = n5890 & n6094 ;
  assign n6097 = n6095 & ~n6096 ;
  assign n6098 = x71 & n4572 ;
  assign n6099 = x70 & n4567 ;
  assign n6100 = x69 & ~n4566 ;
  assign n6101 = n4828 & n6100 ;
  assign n6102 = n6099 | n6101 ;
  assign n6103 = n6098 | n6102 ;
  assign n6104 = n4575 | n6103 ;
  assign n6105 = ( n376 & n6103 ) | ( n376 & n6104 ) | ( n6103 & n6104 ) ;
  assign n6106 = x38 & ~n6105 ;
  assign n6107 = ~x38 & n6105 ;
  assign n6108 = n6106 | n6107 ;
  assign n6109 = n6097 & n6108 ;
  assign n6110 = n6097 & ~n6109 ;
  assign n6111 = ~n6097 & n6108 ;
  assign n6112 = n6110 | n6111 ;
  assign n6113 = n5904 | n5910 ;
  assign n6114 = n6112 | n6113 ;
  assign n6115 = n6112 & n6113 ;
  assign n6116 = n6114 & ~n6115 ;
  assign n6117 = x74 & n3913 ;
  assign n6118 = x73 & n3908 ;
  assign n6119 = x72 & ~n3907 ;
  assign n6120 = n4152 & n6119 ;
  assign n6121 = n6118 | n6120 ;
  assign n6122 = n6117 | n6121 ;
  assign n6123 = n3916 | n6122 ;
  assign n6124 = ( n587 & n6122 ) | ( n587 & n6123 ) | ( n6122 & n6123 ) ;
  assign n6125 = x35 & n6124 ;
  assign n6126 = x35 & ~n6125 ;
  assign n6127 = ( n6124 & ~n6125 ) | ( n6124 & n6126 ) | ( ~n6125 & n6126 ) ;
  assign n6128 = n6116 | n6127 ;
  assign n6129 = n6059 & n6128 ;
  assign n6130 = n6116 & n6127 ;
  assign n6131 = n6128 & ~n6130 ;
  assign n6132 = ~n6129 & n6131 ;
  assign n6133 = x77 & n3314 ;
  assign n6134 = x76 & n3309 ;
  assign n6135 = x75 & ~n3308 ;
  assign n6136 = n3570 & n6135 ;
  assign n6137 = n6134 | n6136 ;
  assign n6138 = n6133 | n6137 ;
  assign n6139 = n3317 | n6138 ;
  assign n6140 = ( n846 & n6138 ) | ( n846 & n6139 ) | ( n6138 & n6139 ) ;
  assign n6141 = x32 & n6140 ;
  assign n6142 = x32 & ~n6141 ;
  assign n6143 = ( n6140 & ~n6141 ) | ( n6140 & n6142 ) | ( ~n6141 & n6142 ) ;
  assign n6144 = n6132 | n6143 ;
  assign n6145 = n6059 & ~n6131 ;
  assign n6146 = n6144 | n6145 ;
  assign n6147 = ( n6132 & n6143 ) | ( n6132 & n6145 ) | ( n6143 & n6145 ) ;
  assign n6148 = n6146 & ~n6147 ;
  assign n6149 = n6058 & n6148 ;
  assign n6150 = n6058 | n6148 ;
  assign n6151 = ~n6149 & n6150 ;
  assign n6152 = x80 & n2775 ;
  assign n6153 = x79 & n2770 ;
  assign n6154 = x78 & ~n2769 ;
  assign n6155 = n2978 & n6154 ;
  assign n6156 = n6153 | n6155 ;
  assign n6157 = n6152 | n6156 ;
  assign n6158 = n2778 | n6157 ;
  assign n6159 = ( n1147 & n6157 ) | ( n1147 & n6158 ) | ( n6157 & n6158 ) ;
  assign n6160 = x29 & n6159 ;
  assign n6161 = x29 & ~n6160 ;
  assign n6162 = ( n6159 & ~n6160 ) | ( n6159 & n6161 ) | ( ~n6160 & n6161 ) ;
  assign n6163 = n6151 & n6162 ;
  assign n6164 = n6151 & ~n6163 ;
  assign n6165 = ~n6151 & n6162 ;
  assign n6166 = n6164 | n6165 ;
  assign n6167 = ( n5873 & n5948 ) | ( n5873 & n5959 ) | ( n5948 & n5959 ) ;
  assign n6168 = n6166 | n6167 ;
  assign n6169 = n6166 & n6167 ;
  assign n6170 = n6168 & ~n6169 ;
  assign n6171 = x83 & n2280 ;
  assign n6172 = x82 & n2275 ;
  assign n6173 = x81 & ~n2274 ;
  assign n6174 = n2481 & n6173 ;
  assign n6175 = n6172 | n6174 ;
  assign n6176 = n6171 | n6175 ;
  assign n6177 = n2283 | n6176 ;
  assign n6178 = ( n1510 & n6176 ) | ( n1510 & n6177 ) | ( n6176 & n6177 ) ;
  assign n6179 = x26 & n6178 ;
  assign n6180 = x26 & ~n6179 ;
  assign n6181 = ( n6178 & ~n6179 ) | ( n6178 & n6180 ) | ( ~n6179 & n6180 ) ;
  assign n6182 = n6170 & n6181 ;
  assign n6183 = n6170 & ~n6182 ;
  assign n6184 = ~n6170 & n6181 ;
  assign n6185 = n6183 | n6184 ;
  assign n6186 = n5974 | n5978 ;
  assign n6187 = n6185 | n6186 ;
  assign n6188 = n6185 & n6186 ;
  assign n6189 = n6187 & ~n6188 ;
  assign n6190 = x86 & n1817 ;
  assign n6191 = x85 & n1812 ;
  assign n6192 = x84 & ~n1811 ;
  assign n6193 = n1977 & n6192 ;
  assign n6194 = n6191 | n6193 ;
  assign n6195 = n6190 | n6194 ;
  assign n6196 = n1820 | n6195 ;
  assign n6197 = ( n1921 & n6195 ) | ( n1921 & n6196 ) | ( n6195 & n6196 ) ;
  assign n6198 = x23 & n6197 ;
  assign n6199 = x23 & ~n6198 ;
  assign n6200 = ( n6197 & ~n6198 ) | ( n6197 & n6199 ) | ( ~n6198 & n6199 ) ;
  assign n6201 = n6189 & n6200 ;
  assign n6202 = n6189 & ~n6201 ;
  assign n6203 = ~n6189 & n6200 ;
  assign n6204 = n6202 | n6203 ;
  assign n6205 = n5992 | n5998 ;
  assign n6206 = n6204 | n6205 ;
  assign n6207 = n6204 & n6205 ;
  assign n6208 = n6206 & ~n6207 ;
  assign n6209 = x89 & n1421 ;
  assign n6210 = x88 & n1416 ;
  assign n6211 = x87 & ~n1415 ;
  assign n6212 = n1584 & n6211 ;
  assign n6213 = n6210 | n6212 ;
  assign n6214 = n6209 | n6213 ;
  assign n6215 = n1424 | n6214 ;
  assign n6216 = ( n2244 & n6214 ) | ( n2244 & n6215 ) | ( n6214 & n6215 ) ;
  assign n6217 = x20 & n6216 ;
  assign n6218 = x20 & ~n6217 ;
  assign n6219 = ( n6216 & ~n6217 ) | ( n6216 & n6218 ) | ( ~n6217 & n6218 ) ;
  assign n6220 = n6208 & n6219 ;
  assign n6221 = n6208 & ~n6220 ;
  assign n6222 = ~n6208 & n6219 ;
  assign n6223 = n6221 | n6222 ;
  assign n6224 = n6012 | n6015 ;
  assign n6225 = n6223 & n6224 ;
  assign n6226 = n6223 | n6224 ;
  assign n6227 = ~n6225 & n6226 ;
  assign n6228 = x92 & n1071 ;
  assign n6229 = x91 & n1066 ;
  assign n6230 = x90 & ~n1065 ;
  assign n6231 = n1189 & n6230 ;
  assign n6232 = n6229 | n6231 ;
  assign n6233 = n6228 | n6232 ;
  assign n6234 = n1074 | n6233 ;
  assign n6235 = ( n2904 & n6233 ) | ( n2904 & n6234 ) | ( n6233 & n6234 ) ;
  assign n6236 = x17 & n6235 ;
  assign n6237 = x17 & ~n6236 ;
  assign n6238 = ( n6235 & ~n6236 ) | ( n6235 & n6237 ) | ( ~n6236 & n6237 ) ;
  assign n6239 = ~n6227 & n6238 ;
  assign n6240 = n6227 & ~n6238 ;
  assign n6241 = n6239 | n6240 ;
  assign n6242 = ( n5871 & n5872 ) | ( n5871 & n6016 ) | ( n5872 & n6016 ) ;
  assign n6243 = n6241 & ~n6242 ;
  assign n6244 = ~n6241 & n6242 ;
  assign n6245 = x95 & n771 ;
  assign n6246 = x94 & n766 ;
  assign n6247 = x93 & ~n765 ;
  assign n6248 = n905 & n6247 ;
  assign n6249 = n6246 | n6248 ;
  assign n6250 = n6245 | n6249 ;
  assign n6251 = n774 | n6250 ;
  assign n6252 = ( n3479 & n6250 ) | ( n3479 & n6251 ) | ( n6250 & n6251 ) ;
  assign n6253 = x14 & n6252 ;
  assign n6254 = x14 & ~n6253 ;
  assign n6255 = ( n6252 & ~n6253 ) | ( n6252 & n6254 ) | ( ~n6253 & n6254 ) ;
  assign n6256 = n6244 | n6255 ;
  assign n6257 = n6243 | n6256 ;
  assign n6258 = ( n6243 & n6244 ) | ( n6243 & n6255 ) | ( n6244 & n6255 ) ;
  assign n6259 = n6257 & ~n6258 ;
  assign n6260 = n6020 | n6023 ;
  assign n6261 = n6259 & n6260 ;
  assign n6262 = n6259 | n6260 ;
  assign n6263 = ~n6261 & n6262 ;
  assign n6264 = x98 & n528 ;
  assign n6265 = x97 & n523 ;
  assign n6266 = x96 & ~n522 ;
  assign n6267 = n635 & n6266 ;
  assign n6268 = n6265 | n6267 ;
  assign n6269 = n6264 | n6268 ;
  assign n6270 = n531 | n6269 ;
  assign n6271 = ( n4105 & n6269 ) | ( n4105 & n6270 ) | ( n6269 & n6270 ) ;
  assign n6272 = x11 & n6271 ;
  assign n6273 = x11 & ~n6272 ;
  assign n6274 = ( n6271 & ~n6272 ) | ( n6271 & n6273 ) | ( ~n6272 & n6273 ) ;
  assign n6275 = n6263 & n6274 ;
  assign n6276 = n6263 & ~n6275 ;
  assign n6277 = ~n6263 & n6274 ;
  assign n6278 = n6276 | n6277 ;
  assign n6279 = n6027 | n6278 ;
  assign n6280 = n6027 & n6278 ;
  assign n6281 = n6279 & ~n6280 ;
  assign n6282 = x101 & n337 ;
  assign n6283 = x100 & n332 ;
  assign n6284 = x99 & ~n331 ;
  assign n6285 = n396 & n6284 ;
  assign n6286 = n6283 | n6285 ;
  assign n6287 = n6282 | n6286 ;
  assign n6288 = n340 | n6287 ;
  assign n6289 = ( n4783 & n6287 ) | ( n4783 & n6288 ) | ( n6287 & n6288 ) ;
  assign n6290 = x8 & n6289 ;
  assign n6291 = x8 & ~n6290 ;
  assign n6292 = ( n6289 & ~n6290 ) | ( n6289 & n6291 ) | ( ~n6290 & n6291 ) ;
  assign n6293 = n6281 | n6292 ;
  assign n6294 = n6031 | n6035 ;
  assign n6295 = ( n6281 & n6292 ) | ( n6281 & n6294 ) | ( n6292 & n6294 ) ;
  assign n6296 = n6293 & ~n6295 ;
  assign n6297 = n6281 & n6292 ;
  assign n6298 = n6293 & ~n6297 ;
  assign n6299 = n6294 & ~n6298 ;
  assign n6300 = n6296 | n6299 ;
  assign n6301 = x104 & n206 ;
  assign n6302 = x103 & n201 ;
  assign n6303 = x102 & ~n200 ;
  assign n6304 = n243 & n6303 ;
  assign n6305 = n6302 | n6304 ;
  assign n6306 = n6301 | n6305 ;
  assign n6307 = n209 | n6306 ;
  assign n6308 = ( n5295 & n6306 ) | ( n5295 & n6307 ) | ( n6306 & n6307 ) ;
  assign n6309 = x5 & n6308 ;
  assign n6310 = x5 & ~n6309 ;
  assign n6311 = ( n6308 & ~n6309 ) | ( n6308 & n6310 ) | ( ~n6309 & n6310 ) ;
  assign n6312 = n6300 | n6311 ;
  assign n6313 = n6300 & n6311 ;
  assign n6314 = n6312 & ~n6313 ;
  assign n6315 = ( n5826 & n6036 ) | ( n5826 & n6047 ) | ( n6036 & n6047 ) ;
  assign n6316 = n6314 & n6315 ;
  assign n6317 = n6314 | n6315 ;
  assign n6318 = ~n6316 & n6317 ;
  assign n6319 = x106 | x107 ;
  assign n6320 = x106 & x107 ;
  assign n6321 = n6319 & ~n6320 ;
  assign n6322 = n5808 | n5810 ;
  assign n6323 = n6321 & n6322 ;
  assign n6324 = n5807 & n6321 ;
  assign n6325 = ( n5786 & n6323 ) | ( n5786 & n6324 ) | ( n6323 & n6324 ) ;
  assign n6326 = ( n5786 & n5807 ) | ( n5786 & n6322 ) | ( n5807 & n6322 ) ;
  assign n6327 = n6321 | n6326 ;
  assign n6328 = ~n6325 & n6327 ;
  assign n6329 = x106 & n131 ;
  assign n6330 = x105 & ~n156 ;
  assign n6331 = ( n135 & n6329 ) | ( n135 & n6330 ) | ( n6329 & n6330 ) ;
  assign n6332 = x0 & x107 ;
  assign n6333 = ( ~n135 & n6329 ) | ( ~n135 & n6332 ) | ( n6329 & n6332 ) ;
  assign n6334 = n6331 | n6333 ;
  assign n6335 = n139 | n6334 ;
  assign n6336 = ( n6328 & n6334 ) | ( n6328 & n6335 ) | ( n6334 & n6335 ) ;
  assign n6337 = x2 & n6336 ;
  assign n6338 = x2 & ~n6337 ;
  assign n6339 = ( n6336 & ~n6337 ) | ( n6336 & n6338 ) | ( ~n6337 & n6338 ) ;
  assign n6340 = n6318 & n6339 ;
  assign n6341 = n6318 & ~n6340 ;
  assign n6342 = ~n6318 & n6339 ;
  assign n6343 = n6341 | n6342 ;
  assign n6344 = n6051 | n6055 ;
  assign n6345 = n6343 & n6344 ;
  assign n6346 = n6343 | n6344 ;
  assign n6347 = ~n6345 & n6346 ;
  assign n6348 = x107 | x108 ;
  assign n6349 = x107 & x108 ;
  assign n6350 = n6348 & ~n6349 ;
  assign n6351 = n6320 | n6323 ;
  assign n6352 = n6350 & n6351 ;
  assign n6353 = n6320 | n6324 ;
  assign n6354 = n6350 & n6353 ;
  assign n6355 = ( n5786 & n6352 ) | ( n5786 & n6354 ) | ( n6352 & n6354 ) ;
  assign n6356 = ( n5786 & n6351 ) | ( n5786 & n6353 ) | ( n6351 & n6353 ) ;
  assign n6357 = n6350 | n6356 ;
  assign n6358 = ~n6355 & n6357 ;
  assign n6359 = x107 & n131 ;
  assign n6360 = x106 & ~n156 ;
  assign n6361 = ( n135 & n6359 ) | ( n135 & n6360 ) | ( n6359 & n6360 ) ;
  assign n6362 = x0 & x108 ;
  assign n6363 = ( ~n135 & n6359 ) | ( ~n135 & n6362 ) | ( n6359 & n6362 ) ;
  assign n6364 = n6361 | n6363 ;
  assign n6365 = n139 | n6364 ;
  assign n6366 = ( n6358 & n6364 ) | ( n6358 & n6365 ) | ( n6364 & n6365 ) ;
  assign n6367 = x2 & n6366 ;
  assign n6368 = x2 & ~n6367 ;
  assign n6369 = ( n6366 & ~n6367 ) | ( n6366 & n6368 ) | ( ~n6367 & n6368 ) ;
  assign n6370 = n6340 | n6345 ;
  assign n6371 = n6313 | n6316 ;
  assign n6372 = n6258 | n6261 ;
  assign n6373 = x90 & n1421 ;
  assign n6374 = x89 & n1416 ;
  assign n6375 = x88 & ~n1415 ;
  assign n6376 = n1584 & n6375 ;
  assign n6377 = n6374 | n6376 ;
  assign n6378 = n6373 | n6377 ;
  assign n6379 = n1424 | n6378 ;
  assign n6380 = ( n2410 & n6378 ) | ( n2410 & n6379 ) | ( n6378 & n6379 ) ;
  assign n6381 = x20 & n6380 ;
  assign n6382 = x20 & ~n6381 ;
  assign n6383 = ( n6380 & ~n6381 ) | ( n6380 & n6382 ) | ( ~n6381 & n6382 ) ;
  assign n6384 = x87 & n1817 ;
  assign n6385 = x86 & n1812 ;
  assign n6386 = x85 & ~n1811 ;
  assign n6387 = n1977 & n6386 ;
  assign n6388 = n6385 | n6387 ;
  assign n6389 = n6384 | n6388 ;
  assign n6390 = n1820 | n6389 ;
  assign n6391 = ( n2067 & n6389 ) | ( n2067 & n6390 ) | ( n6389 & n6390 ) ;
  assign n6392 = x23 & n6391 ;
  assign n6393 = x23 & ~n6392 ;
  assign n6394 = ( n6391 & ~n6392 ) | ( n6391 & n6393 ) | ( ~n6392 & n6393 ) ;
  assign n6395 = n6109 | n6115 ;
  assign n6396 = x66 & n6068 ;
  assign n6397 = x65 & n6063 ;
  assign n6398 = ~n5877 & n6067 ;
  assign n6399 = x64 & ~n6062 ;
  assign n6400 = n6398 & n6399 ;
  assign n6401 = n6397 | n6400 ;
  assign n6402 = n6396 | n6401 ;
  assign n6403 = n153 & n6071 ;
  assign n6404 = n6402 | n6403 ;
  assign n6405 = x44 | n6404 ;
  assign n6406 = ~x44 & n6405 ;
  assign n6407 = ( ~n6404 & n6405 ) | ( ~n6404 & n6406 ) | ( n6405 & n6406 ) ;
  assign n6408 = n6078 | n6407 ;
  assign n6409 = n6078 & n6407 ;
  assign n6410 = n6408 & ~n6409 ;
  assign n6411 = n264 & n5343 ;
  assign n6412 = x69 & n5340 ;
  assign n6413 = x68 & n5335 ;
  assign n6414 = x67 & ~n5334 ;
  assign n6415 = n5580 & n6414 ;
  assign n6416 = n6413 | n6415 ;
  assign n6417 = n6412 | n6416 ;
  assign n6418 = n6411 | n6417 ;
  assign n6419 = x41 | n6418 ;
  assign n6420 = ~x41 & n6419 ;
  assign n6421 = ( ~n6418 & n6419 ) | ( ~n6418 & n6420 ) | ( n6419 & n6420 ) ;
  assign n6422 = n6410 & n6421 ;
  assign n6423 = n6410 & ~n6422 ;
  assign n6424 = ~n6410 & n6421 ;
  assign n6425 = n6423 | n6424 ;
  assign n6426 = n6093 | n6096 ;
  assign n6427 = n6425 & n6426 ;
  assign n6428 = n6425 | n6426 ;
  assign n6429 = ~n6427 & n6428 ;
  assign n6430 = x72 & n4572 ;
  assign n6431 = x71 & n4567 ;
  assign n6432 = x70 & ~n4566 ;
  assign n6433 = n4828 & n6432 ;
  assign n6434 = n6431 | n6433 ;
  assign n6435 = n6430 | n6434 ;
  assign n6436 = ( n435 & n4575 ) | ( n435 & n6435 ) | ( n4575 & n6435 ) ;
  assign n6437 = ( x38 & ~n6435 ) | ( x38 & n6436 ) | ( ~n6435 & n6436 ) ;
  assign n6438 = ~n6436 & n6437 ;
  assign n6439 = n6435 | n6437 ;
  assign n6440 = ( ~x38 & n6438 ) | ( ~x38 & n6439 ) | ( n6438 & n6439 ) ;
  assign n6441 = ~n6429 & n6440 ;
  assign n6442 = n6429 & ~n6440 ;
  assign n6443 = n6441 | n6442 ;
  assign n6444 = n6395 & ~n6443 ;
  assign n6445 = ~n6395 & n6443 ;
  assign n6446 = x75 & n3913 ;
  assign n6447 = x74 & n3908 ;
  assign n6448 = x73 & ~n3907 ;
  assign n6449 = n4152 & n6448 ;
  assign n6450 = n6447 | n6449 ;
  assign n6451 = n6446 | n6450 ;
  assign n6452 = n3916 | n6451 ;
  assign n6453 = ( n609 & n6451 ) | ( n609 & n6452 ) | ( n6451 & n6452 ) ;
  assign n6454 = x35 & n6453 ;
  assign n6455 = x35 & ~n6454 ;
  assign n6456 = ( n6453 & ~n6454 ) | ( n6453 & n6455 ) | ( ~n6454 & n6455 ) ;
  assign n6457 = n6445 | n6456 ;
  assign n6458 = n6444 | n6457 ;
  assign n6459 = ( n6444 & n6445 ) | ( n6444 & n6456 ) | ( n6445 & n6456 ) ;
  assign n6460 = n6458 & ~n6459 ;
  assign n6461 = n6129 | n6130 ;
  assign n6462 = n6460 & n6461 ;
  assign n6463 = n6460 | n6461 ;
  assign n6464 = ~n6462 & n6463 ;
  assign n6465 = x78 & n3314 ;
  assign n6466 = x77 & n3309 ;
  assign n6467 = x76 & ~n3308 ;
  assign n6468 = n3570 & n6467 ;
  assign n6469 = n6466 | n6468 ;
  assign n6470 = n6465 | n6469 ;
  assign n6471 = n3317 | n6470 ;
  assign n6472 = ( n868 & n6470 ) | ( n868 & n6471 ) | ( n6470 & n6471 ) ;
  assign n6473 = x32 & n6472 ;
  assign n6474 = x32 & ~n6473 ;
  assign n6475 = ( n6472 & ~n6473 ) | ( n6472 & n6474 ) | ( ~n6473 & n6474 ) ;
  assign n6476 = n6464 | n6475 ;
  assign n6477 = n6464 & n6475 ;
  assign n6478 = n6476 & ~n6477 ;
  assign n6479 = n6147 | n6149 ;
  assign n6480 = n6478 & n6479 ;
  assign n6481 = n6478 | n6479 ;
  assign n6482 = ~n6480 & n6481 ;
  assign n6483 = x81 & n2775 ;
  assign n6484 = x80 & n2770 ;
  assign n6485 = x79 & ~n2769 ;
  assign n6486 = n2978 & n6485 ;
  assign n6487 = n6484 | n6486 ;
  assign n6488 = n6483 | n6487 ;
  assign n6489 = n2778 | n6488 ;
  assign n6490 = ( n1256 & n6488 ) | ( n1256 & n6489 ) | ( n6488 & n6489 ) ;
  assign n6491 = x29 & n6490 ;
  assign n6492 = x29 & ~n6491 ;
  assign n6493 = ( n6490 & ~n6491 ) | ( n6490 & n6492 ) | ( ~n6491 & n6492 ) ;
  assign n6494 = n6482 | n6493 ;
  assign n6495 = n6482 & n6493 ;
  assign n6496 = n6494 & ~n6495 ;
  assign n6497 = n6163 & n6496 ;
  assign n6498 = ( n6169 & n6496 ) | ( n6169 & n6497 ) | ( n6496 & n6497 ) ;
  assign n6499 = n6163 | n6496 ;
  assign n6500 = n6169 | n6499 ;
  assign n6501 = ~n6498 & n6500 ;
  assign n6502 = x84 & n2280 ;
  assign n6503 = x83 & n2275 ;
  assign n6504 = x82 & ~n2274 ;
  assign n6505 = n2481 & n6504 ;
  assign n6506 = n6503 | n6505 ;
  assign n6507 = n6502 | n6506 ;
  assign n6508 = n2283 | n6507 ;
  assign n6509 = ( n1537 & n6507 ) | ( n1537 & n6508 ) | ( n6507 & n6508 ) ;
  assign n6510 = x26 & n6509 ;
  assign n6511 = x26 & ~n6510 ;
  assign n6512 = ( n6509 & ~n6510 ) | ( n6509 & n6511 ) | ( ~n6510 & n6511 ) ;
  assign n6513 = n6501 & n6512 ;
  assign n6514 = n6501 & ~n6513 ;
  assign n6515 = ~n6501 & n6512 ;
  assign n6516 = n6514 | n6515 ;
  assign n6517 = n6182 | n6188 ;
  assign n6518 = n6516 | n6517 ;
  assign n6519 = n6516 & n6517 ;
  assign n6520 = n6518 & ~n6519 ;
  assign n6521 = n6201 | n6207 ;
  assign n6522 = ( n6394 & n6520 ) | ( n6394 & n6521 ) | ( n6520 & n6521 ) ;
  assign n6523 = ( n6520 & n6521 ) | ( n6520 & ~n6522 ) | ( n6521 & ~n6522 ) ;
  assign n6524 = ( n6394 & ~n6522 ) | ( n6394 & n6523 ) | ( ~n6522 & n6523 ) ;
  assign n6525 = n6383 | n6524 ;
  assign n6526 = n6383 & n6524 ;
  assign n6527 = n6525 & ~n6526 ;
  assign n6528 = n6220 | n6225 ;
  assign n6529 = n6527 & n6528 ;
  assign n6530 = n6527 | n6528 ;
  assign n6531 = ~n6529 & n6530 ;
  assign n6532 = x93 & n1071 ;
  assign n6533 = x92 & n1066 ;
  assign n6534 = x91 & ~n1065 ;
  assign n6535 = n1189 & n6534 ;
  assign n6536 = n6533 | n6535 ;
  assign n6537 = n6532 | n6536 ;
  assign n6538 = n1074 | n6537 ;
  assign n6539 = ( n2931 & n6537 ) | ( n2931 & n6538 ) | ( n6537 & n6538 ) ;
  assign n6540 = x17 & n6539 ;
  assign n6541 = x17 & ~n6540 ;
  assign n6542 = ( n6539 & ~n6540 ) | ( n6539 & n6541 ) | ( ~n6540 & n6541 ) ;
  assign n6543 = n6531 | n6542 ;
  assign n6544 = n6531 & n6542 ;
  assign n6545 = n6543 & ~n6544 ;
  assign n6546 = ( n6227 & n6238 ) | ( n6227 & n6242 ) | ( n6238 & n6242 ) ;
  assign n6547 = n6545 & n6546 ;
  assign n6548 = n6545 | n6546 ;
  assign n6549 = ~n6547 & n6548 ;
  assign n6550 = x96 & n771 ;
  assign n6551 = x95 & n766 ;
  assign n6552 = x94 & ~n765 ;
  assign n6553 = n905 & n6552 ;
  assign n6554 = n6551 | n6553 ;
  assign n6555 = n6550 | n6554 ;
  assign n6556 = n774 | n6555 ;
  assign n6557 = ( n3509 & n6555 ) | ( n3509 & n6556 ) | ( n6555 & n6556 ) ;
  assign n6558 = x14 & n6557 ;
  assign n6559 = x14 & ~n6558 ;
  assign n6560 = ( n6557 & ~n6558 ) | ( n6557 & n6559 ) | ( ~n6558 & n6559 ) ;
  assign n6561 = n6549 | n6560 ;
  assign n6562 = n6549 & n6560 ;
  assign n6563 = n6561 & ~n6562 ;
  assign n6564 = n6372 & n6563 ;
  assign n6565 = n6372 | n6563 ;
  assign n6566 = ~n6564 & n6565 ;
  assign n6567 = x99 & n528 ;
  assign n6568 = x98 & n523 ;
  assign n6569 = x97 & ~n522 ;
  assign n6570 = n635 & n6569 ;
  assign n6571 = n6568 | n6570 ;
  assign n6572 = n6567 | n6571 ;
  assign n6573 = n531 | n6572 ;
  assign n6574 = ( n4325 & n6572 ) | ( n4325 & n6573 ) | ( n6572 & n6573 ) ;
  assign n6575 = x11 & n6574 ;
  assign n6576 = x11 & ~n6575 ;
  assign n6577 = ( n6574 & ~n6575 ) | ( n6574 & n6576 ) | ( ~n6575 & n6576 ) ;
  assign n6578 = n6566 & n6577 ;
  assign n6579 = n6566 & ~n6578 ;
  assign n6580 = ~n6566 & n6577 ;
  assign n6581 = n6579 | n6580 ;
  assign n6582 = n6275 | n6280 ;
  assign n6583 = n6581 | n6582 ;
  assign n6584 = n6581 & n6582 ;
  assign n6585 = n6583 & ~n6584 ;
  assign n6586 = x102 & n337 ;
  assign n6587 = x101 & n332 ;
  assign n6588 = x100 & ~n331 ;
  assign n6589 = n396 & n6588 ;
  assign n6590 = n6587 | n6589 ;
  assign n6591 = n6586 | n6590 ;
  assign n6592 = n340 | n6591 ;
  assign n6593 = ( n5025 & n6591 ) | ( n5025 & n6592 ) | ( n6591 & n6592 ) ;
  assign n6594 = x8 & n6593 ;
  assign n6595 = x8 & ~n6594 ;
  assign n6596 = ( n6593 & ~n6594 ) | ( n6593 & n6595 ) | ( ~n6594 & n6595 ) ;
  assign n6597 = n6585 & n6596 ;
  assign n6598 = n6585 & ~n6597 ;
  assign n6599 = ~n6585 & n6596 ;
  assign n6600 = n6598 | n6599 ;
  assign n6601 = n6295 | n6600 ;
  assign n6602 = n6295 & n6600 ;
  assign n6603 = n6601 & ~n6602 ;
  assign n6604 = x105 & n206 ;
  assign n6605 = x104 & n201 ;
  assign n6606 = x103 & ~n200 ;
  assign n6607 = n243 & n6606 ;
  assign n6608 = n6605 | n6607 ;
  assign n6609 = n6604 | n6608 ;
  assign n6610 = n209 | n6609 ;
  assign n6611 = ( n5788 & n6609 ) | ( n5788 & n6610 ) | ( n6609 & n6610 ) ;
  assign n6612 = x5 & n6611 ;
  assign n6613 = x5 & ~n6612 ;
  assign n6614 = ( n6611 & ~n6612 ) | ( n6611 & n6613 ) | ( ~n6612 & n6613 ) ;
  assign n6615 = n6603 & n6614 ;
  assign n6616 = n6603 & ~n6615 ;
  assign n6617 = ~n6603 & n6614 ;
  assign n6618 = n6616 | n6617 ;
  assign n6619 = n6371 & n6618 ;
  assign n6620 = n6371 & ~n6619 ;
  assign n6621 = n6618 & ~n6619 ;
  assign n6622 = n6620 | n6621 ;
  assign n6623 = ( n6369 & n6370 ) | ( n6369 & ~n6622 ) | ( n6370 & ~n6622 ) ;
  assign n6624 = ( ~n6370 & n6622 ) | ( ~n6370 & n6623 ) | ( n6622 & n6623 ) ;
  assign n6625 = ( ~n6369 & n6623 ) | ( ~n6369 & n6624 ) | ( n6623 & n6624 ) ;
  assign n6626 = x100 & n528 ;
  assign n6627 = x99 & n523 ;
  assign n6628 = x98 & ~n522 ;
  assign n6629 = n635 & n6628 ;
  assign n6630 = n6627 | n6629 ;
  assign n6631 = n6626 | n6630 ;
  assign n6632 = n531 | n6631 ;
  assign n6633 = ( n4532 & n6631 ) | ( n4532 & n6632 ) | ( n6631 & n6632 ) ;
  assign n6634 = x11 & n6633 ;
  assign n6635 = x11 & ~n6634 ;
  assign n6636 = ( n6633 & ~n6634 ) | ( n6633 & n6635 ) | ( ~n6634 & n6635 ) ;
  assign n6637 = x97 & n771 ;
  assign n6638 = x96 & n766 ;
  assign n6639 = x95 & ~n765 ;
  assign n6640 = n905 & n6639 ;
  assign n6641 = n6638 | n6640 ;
  assign n6642 = n6637 | n6641 ;
  assign n6643 = n774 | n6642 ;
  assign n6644 = ( n3707 & n6642 ) | ( n3707 & n6643 ) | ( n6642 & n6643 ) ;
  assign n6645 = x14 & n6644 ;
  assign n6646 = x14 & ~n6645 ;
  assign n6647 = ( n6644 & ~n6645 ) | ( n6644 & n6646 ) | ( ~n6645 & n6646 ) ;
  assign n6648 = x94 & n1071 ;
  assign n6649 = x93 & n1066 ;
  assign n6650 = x92 & ~n1065 ;
  assign n6651 = n1189 & n6650 ;
  assign n6652 = n6649 | n6651 ;
  assign n6653 = n6648 | n6652 ;
  assign n6654 = n1074 | n6653 ;
  assign n6655 = ( n3271 & n6653 ) | ( n3271 & n6654 ) | ( n6653 & n6654 ) ;
  assign n6656 = x17 & n6655 ;
  assign n6657 = x17 & ~n6656 ;
  assign n6658 = ( n6655 & ~n6656 ) | ( n6655 & n6657 ) | ( ~n6656 & n6657 ) ;
  assign n6659 = x91 & n1421 ;
  assign n6660 = x90 & n1416 ;
  assign n6661 = x89 & ~n1415 ;
  assign n6662 = n1584 & n6661 ;
  assign n6663 = n6660 | n6662 ;
  assign n6664 = n6659 | n6663 ;
  assign n6665 = n1424 | n6664 ;
  assign n6666 = ( n2714 & n6664 ) | ( n2714 & n6665 ) | ( n6664 & n6665 ) ;
  assign n6667 = x20 & n6666 ;
  assign n6668 = x20 & ~n6667 ;
  assign n6669 = ( n6666 & ~n6667 ) | ( n6666 & n6668 ) | ( ~n6667 & n6668 ) ;
  assign n6670 = n6526 | n6529 ;
  assign n6671 = n6495 | n6498 ;
  assign n6672 = n6477 | n6480 ;
  assign n6673 = n6459 | n6462 ;
  assign n6674 = x44 & ~x45 ;
  assign n6675 = ~x44 & x45 ;
  assign n6676 = n6674 | n6675 ;
  assign n6677 = x64 & n6676 ;
  assign n6678 = x67 & n6068 ;
  assign n6679 = x66 & n6063 ;
  assign n6680 = x65 & ~n6062 ;
  assign n6681 = n6398 & n6680 ;
  assign n6682 = n6679 | n6681 ;
  assign n6683 = n6678 | n6682 ;
  assign n6684 = n180 & n6071 ;
  assign n6685 = n6683 | n6684 ;
  assign n6686 = x44 & ~n6685 ;
  assign n6687 = ~x44 & n6685 ;
  assign n6688 = n6686 | n6687 ;
  assign n6689 = ( n6409 & n6677 ) | ( n6409 & n6688 ) | ( n6677 & n6688 ) ;
  assign n6690 = ( n6409 & n6688 ) | ( n6409 & ~n6689 ) | ( n6688 & ~n6689 ) ;
  assign n6691 = ( n6677 & ~n6689 ) | ( n6677 & n6690 ) | ( ~n6689 & n6690 ) ;
  assign n6692 = x70 & n5340 ;
  assign n6693 = x69 & n5335 ;
  assign n6694 = x68 & ~n5334 ;
  assign n6695 = n5580 & n6694 ;
  assign n6696 = n6693 | n6695 ;
  assign n6697 = n6692 | n6696 ;
  assign n6698 = n5343 | n6697 ;
  assign n6699 = ( n310 & n6697 ) | ( n310 & n6698 ) | ( n6697 & n6698 ) ;
  assign n6700 = x41 & ~n6699 ;
  assign n6701 = ~x41 & n6699 ;
  assign n6702 = n6700 | n6701 ;
  assign n6703 = n6691 & n6702 ;
  assign n6704 = n6691 & ~n6703 ;
  assign n6705 = ~n6691 & n6702 ;
  assign n6706 = n6704 | n6705 ;
  assign n6707 = n6422 | n6427 ;
  assign n6708 = n6706 | n6707 ;
  assign n6709 = n6706 & n6707 ;
  assign n6710 = n6708 & ~n6709 ;
  assign n6711 = x73 & n4572 ;
  assign n6712 = x72 & n4567 ;
  assign n6713 = x71 & ~n4566 ;
  assign n6714 = n4828 & n6713 ;
  assign n6715 = n6712 | n6714 ;
  assign n6716 = n6711 | n6715 ;
  assign n6717 = ( n499 & n4575 ) | ( n499 & n6716 ) | ( n4575 & n6716 ) ;
  assign n6718 = ( x38 & ~n6716 ) | ( x38 & n6717 ) | ( ~n6716 & n6717 ) ;
  assign n6719 = ~n6717 & n6718 ;
  assign n6720 = n6716 | n6718 ;
  assign n6721 = ( ~x38 & n6719 ) | ( ~x38 & n6720 ) | ( n6719 & n6720 ) ;
  assign n6722 = n6710 | n6721 ;
  assign n6723 = n6710 & n6721 ;
  assign n6724 = n6722 & ~n6723 ;
  assign n6725 = ( n6395 & n6429 ) | ( n6395 & n6440 ) | ( n6429 & n6440 ) ;
  assign n6726 = n6724 & n6725 ;
  assign n6727 = n6724 | n6725 ;
  assign n6728 = ~n6726 & n6727 ;
  assign n6729 = x76 & n3913 ;
  assign n6730 = x75 & n3908 ;
  assign n6731 = x74 & ~n3907 ;
  assign n6732 = n4152 & n6731 ;
  assign n6733 = n6730 | n6732 ;
  assign n6734 = n6729 | n6733 ;
  assign n6735 = n3916 | n6734 ;
  assign n6736 = ( n740 & n6734 ) | ( n740 & n6735 ) | ( n6734 & n6735 ) ;
  assign n6737 = x35 & n6736 ;
  assign n6738 = x35 & ~n6737 ;
  assign n6739 = ( n6736 & ~n6737 ) | ( n6736 & n6738 ) | ( ~n6737 & n6738 ) ;
  assign n6740 = n6728 & n6739 ;
  assign n6741 = n6728 & ~n6740 ;
  assign n6742 = ~n6728 & n6739 ;
  assign n6743 = n6741 | n6742 ;
  assign n6744 = n6673 & n6743 ;
  assign n6745 = n6673 & ~n6744 ;
  assign n6746 = n6743 & ~n6744 ;
  assign n6747 = n6745 | n6746 ;
  assign n6748 = x79 & n3314 ;
  assign n6749 = x78 & n3309 ;
  assign n6750 = x77 & ~n3308 ;
  assign n6751 = n3570 & n6750 ;
  assign n6752 = n6749 | n6751 ;
  assign n6753 = n6748 | n6752 ;
  assign n6754 = n3317 | n6753 ;
  assign n6755 = ( n961 & n6753 ) | ( n961 & n6754 ) | ( n6753 & n6754 ) ;
  assign n6756 = x32 & n6755 ;
  assign n6757 = x32 & ~n6756 ;
  assign n6758 = ( n6755 & ~n6756 ) | ( n6755 & n6757 ) | ( ~n6756 & n6757 ) ;
  assign n6759 = ( n6672 & n6747 ) | ( n6672 & ~n6758 ) | ( n6747 & ~n6758 ) ;
  assign n6760 = ( ~n6747 & n6758 ) | ( ~n6747 & n6759 ) | ( n6758 & n6759 ) ;
  assign n6761 = ( ~n6672 & n6759 ) | ( ~n6672 & n6760 ) | ( n6759 & n6760 ) ;
  assign n6762 = x82 & n2775 ;
  assign n6763 = x81 & n2770 ;
  assign n6764 = x80 & ~n2769 ;
  assign n6765 = n2978 & n6764 ;
  assign n6766 = n6763 | n6765 ;
  assign n6767 = n6762 | n6766 ;
  assign n6768 = n2778 | n6767 ;
  assign n6769 = ( n1371 & n6767 ) | ( n1371 & n6768 ) | ( n6767 & n6768 ) ;
  assign n6770 = x29 & n6769 ;
  assign n6771 = x29 & ~n6770 ;
  assign n6772 = ( n6769 & ~n6770 ) | ( n6769 & n6771 ) | ( ~n6770 & n6771 ) ;
  assign n6773 = n6761 & n6772 ;
  assign n6774 = n6761 | n6772 ;
  assign n6775 = ~n6773 & n6774 ;
  assign n6776 = n6671 & n6775 ;
  assign n6777 = n6671 | n6775 ;
  assign n6778 = ~n6776 & n6777 ;
  assign n6779 = x85 & n2280 ;
  assign n6780 = x84 & n2275 ;
  assign n6781 = x83 & ~n2274 ;
  assign n6782 = n2481 & n6781 ;
  assign n6783 = n6780 | n6782 ;
  assign n6784 = n6779 | n6783 ;
  assign n6785 = n2283 | n6784 ;
  assign n6786 = ( n1765 & n6784 ) | ( n1765 & n6785 ) | ( n6784 & n6785 ) ;
  assign n6787 = x26 & n6786 ;
  assign n6788 = x26 & ~n6787 ;
  assign n6789 = ( n6786 & ~n6787 ) | ( n6786 & n6788 ) | ( ~n6787 & n6788 ) ;
  assign n6790 = n6778 & n6789 ;
  assign n6791 = n6778 & ~n6790 ;
  assign n6792 = ~n6778 & n6789 ;
  assign n6793 = n6791 | n6792 ;
  assign n6794 = n6513 | n6519 ;
  assign n6795 = n6793 | n6794 ;
  assign n6796 = n6793 & n6794 ;
  assign n6797 = n6795 & ~n6796 ;
  assign n6798 = x88 & n1817 ;
  assign n6799 = x87 & n1812 ;
  assign n6800 = x86 & ~n1811 ;
  assign n6801 = n1977 & n6800 ;
  assign n6802 = n6799 | n6801 ;
  assign n6803 = n6798 | n6802 ;
  assign n6804 = n1820 | n6803 ;
  assign n6805 = ( n2095 & n6803 ) | ( n2095 & n6804 ) | ( n6803 & n6804 ) ;
  assign n6806 = x23 & n6805 ;
  assign n6807 = x23 & ~n6806 ;
  assign n6808 = ( n6805 & ~n6806 ) | ( n6805 & n6807 ) | ( ~n6806 & n6807 ) ;
  assign n6809 = n6797 | n6808 ;
  assign n6810 = n6797 & n6808 ;
  assign n6811 = n6809 & ~n6810 ;
  assign n6812 = n6522 & n6811 ;
  assign n6813 = n6522 | n6811 ;
  assign n6814 = ~n6812 & n6813 ;
  assign n6815 = ( n6669 & n6670 ) | ( n6669 & ~n6814 ) | ( n6670 & ~n6814 ) ;
  assign n6816 = ( ~n6670 & n6814 ) | ( ~n6670 & n6815 ) | ( n6814 & n6815 ) ;
  assign n6817 = ( ~n6669 & n6815 ) | ( ~n6669 & n6816 ) | ( n6815 & n6816 ) ;
  assign n6818 = n6658 & n6817 ;
  assign n6819 = n6658 | n6817 ;
  assign n6820 = ~n6818 & n6819 ;
  assign n6821 = n6544 | n6547 ;
  assign n6822 = n6820 & n6821 ;
  assign n6823 = n6820 | n6821 ;
  assign n6824 = ~n6822 & n6823 ;
  assign n6825 = n6562 | n6564 ;
  assign n6826 = ( n6647 & n6824 ) | ( n6647 & n6825 ) | ( n6824 & n6825 ) ;
  assign n6827 = ( n6824 & n6825 ) | ( n6824 & ~n6826 ) | ( n6825 & ~n6826 ) ;
  assign n6828 = ( n6647 & ~n6826 ) | ( n6647 & n6827 ) | ( ~n6826 & n6827 ) ;
  assign n6829 = n6636 & n6828 ;
  assign n6830 = n6636 | n6828 ;
  assign n6831 = ~n6829 & n6830 ;
  assign n6832 = n6578 | n6831 ;
  assign n6833 = n6584 | n6832 ;
  assign n6834 = ( n6578 & n6584 ) | ( n6578 & n6831 ) | ( n6584 & n6831 ) ;
  assign n6835 = n6833 & ~n6834 ;
  assign n6836 = x103 & n337 ;
  assign n6837 = x102 & n332 ;
  assign n6838 = x101 & ~n331 ;
  assign n6839 = n396 & n6838 ;
  assign n6840 = n6837 | n6839 ;
  assign n6841 = n6836 | n6840 ;
  assign n6842 = n340 | n6841 ;
  assign n6843 = ( n5264 & n6841 ) | ( n5264 & n6842 ) | ( n6841 & n6842 ) ;
  assign n6844 = x8 & n6843 ;
  assign n6845 = x8 & ~n6844 ;
  assign n6846 = ( n6843 & ~n6844 ) | ( n6843 & n6845 ) | ( ~n6844 & n6845 ) ;
  assign n6847 = n6835 & n6846 ;
  assign n6848 = n6835 & ~n6847 ;
  assign n6849 = ~n6835 & n6846 ;
  assign n6850 = n6848 | n6849 ;
  assign n6851 = n6597 | n6602 ;
  assign n6852 = n6850 | n6851 ;
  assign n6853 = n6850 & n6851 ;
  assign n6854 = n6852 & ~n6853 ;
  assign n6855 = x106 & n206 ;
  assign n6856 = x105 & n201 ;
  assign n6857 = x104 & ~n200 ;
  assign n6858 = n243 & n6857 ;
  assign n6859 = n6856 | n6858 ;
  assign n6860 = n6855 | n6859 ;
  assign n6861 = n209 | n6860 ;
  assign n6862 = ( n5814 & n6860 ) | ( n5814 & n6861 ) | ( n6860 & n6861 ) ;
  assign n6863 = x5 & n6862 ;
  assign n6864 = x5 & ~n6863 ;
  assign n6865 = ( n6862 & ~n6863 ) | ( n6862 & n6864 ) | ( ~n6863 & n6864 ) ;
  assign n6866 = n6854 & n6865 ;
  assign n6867 = n6854 & ~n6866 ;
  assign n6868 = ~n6854 & n6865 ;
  assign n6869 = n6867 | n6868 ;
  assign n6870 = n6615 | n6619 ;
  assign n6871 = n6869 | n6870 ;
  assign n6872 = n6869 & n6870 ;
  assign n6873 = n6871 & ~n6872 ;
  assign n6874 = x108 | x109 ;
  assign n6875 = x108 & x109 ;
  assign n6876 = n6874 & ~n6875 ;
  assign n6877 = n6349 | n6352 ;
  assign n6878 = n6876 & n6877 ;
  assign n6879 = n6349 | n6354 ;
  assign n6880 = n6876 & n6879 ;
  assign n6881 = ( n5786 & n6878 ) | ( n5786 & n6880 ) | ( n6878 & n6880 ) ;
  assign n6882 = ( n5786 & n6877 ) | ( n5786 & n6879 ) | ( n6877 & n6879 ) ;
  assign n6883 = n6876 | n6882 ;
  assign n6884 = ~n6881 & n6883 ;
  assign n6885 = x108 & n131 ;
  assign n6886 = x107 & ~n156 ;
  assign n6887 = ( n135 & n6885 ) | ( n135 & n6886 ) | ( n6885 & n6886 ) ;
  assign n6888 = x0 & x109 ;
  assign n6889 = ( ~n135 & n6885 ) | ( ~n135 & n6888 ) | ( n6885 & n6888 ) ;
  assign n6890 = n6887 | n6889 ;
  assign n6891 = n139 | n6890 ;
  assign n6892 = ( n6884 & n6890 ) | ( n6884 & n6891 ) | ( n6890 & n6891 ) ;
  assign n6893 = x2 & n6892 ;
  assign n6894 = x2 & ~n6893 ;
  assign n6895 = ( n6892 & ~n6893 ) | ( n6892 & n6894 ) | ( ~n6893 & n6894 ) ;
  assign n6896 = n6873 | n6895 ;
  assign n6897 = n6873 & n6895 ;
  assign n6898 = n6896 & ~n6897 ;
  assign n6899 = ( n6369 & n6370 ) | ( n6369 & n6622 ) | ( n6370 & n6622 ) ;
  assign n6900 = n6898 | n6899 ;
  assign n6901 = n6898 & n6899 ;
  assign n6902 = n6900 & ~n6901 ;
  assign n6903 = x107 & n206 ;
  assign n6904 = x106 & n201 ;
  assign n6905 = x105 & ~n200 ;
  assign n6906 = n243 & n6905 ;
  assign n6907 = n6904 | n6906 ;
  assign n6908 = n6903 | n6907 ;
  assign n6909 = n209 | n6908 ;
  assign n6910 = ( n6328 & n6908 ) | ( n6328 & n6909 ) | ( n6908 & n6909 ) ;
  assign n6911 = x5 & n6910 ;
  assign n6912 = x5 & ~n6911 ;
  assign n6913 = ( n6910 & ~n6911 ) | ( n6910 & n6912 ) | ( ~n6911 & n6912 ) ;
  assign n6914 = x104 & n337 ;
  assign n6915 = x103 & n332 ;
  assign n6916 = x102 & ~n331 ;
  assign n6917 = n396 & n6916 ;
  assign n6918 = n6915 | n6917 ;
  assign n6919 = n6914 | n6918 ;
  assign n6920 = n340 | n6919 ;
  assign n6921 = ( n5295 & n6919 ) | ( n5295 & n6920 ) | ( n6919 & n6920 ) ;
  assign n6922 = x8 & n6921 ;
  assign n6923 = x8 & ~n6922 ;
  assign n6924 = ( n6921 & ~n6922 ) | ( n6921 & n6923 ) | ( ~n6922 & n6923 ) ;
  assign n6925 = n6847 | n6853 ;
  assign n6926 = n6818 | n6822 ;
  assign n6927 = n6740 | n6744 ;
  assign n6928 = n6723 | n6726 ;
  assign n6929 = ~x45 & x46 ;
  assign n6930 = x45 & ~x46 ;
  assign n6931 = n6929 | n6930 ;
  assign n6932 = ~n6676 & n6931 ;
  assign n6933 = x64 & n6932 ;
  assign n6934 = ~x46 & x47 ;
  assign n6935 = x46 & ~x47 ;
  assign n6936 = n6934 | n6935 ;
  assign n6937 = n6676 & ~n6936 ;
  assign n6938 = x65 & n6937 ;
  assign n6939 = n6933 | n6938 ;
  assign n6940 = n6676 & n6936 ;
  assign n6941 = n142 & n6940 ;
  assign n6942 = n6939 | n6941 ;
  assign n6943 = x47 | n6942 ;
  assign n6944 = ~x47 & n6943 ;
  assign n6945 = ( ~n6942 & n6943 ) | ( ~n6942 & n6944 ) | ( n6943 & n6944 ) ;
  assign n6946 = x47 & ~n6677 ;
  assign n6947 = n6945 & n6946 ;
  assign n6948 = n6945 | n6946 ;
  assign n6949 = ~n6947 & n6948 ;
  assign n6950 = n229 & n6071 ;
  assign n6951 = x68 & n6068 ;
  assign n6952 = x67 & n6063 ;
  assign n6953 = x66 & ~n6062 ;
  assign n6954 = n6398 & n6953 ;
  assign n6955 = n6952 | n6954 ;
  assign n6956 = n6951 | n6955 ;
  assign n6957 = n6950 | n6956 ;
  assign n6958 = x44 | n6957 ;
  assign n6959 = ~x44 & n6958 ;
  assign n6960 = ( ~n6957 & n6958 ) | ( ~n6957 & n6959 ) | ( n6958 & n6959 ) ;
  assign n6961 = n6949 | n6960 ;
  assign n6962 = n6949 & n6960 ;
  assign n6963 = n6961 & ~n6962 ;
  assign n6964 = n6689 | n6963 ;
  assign n6965 = n6689 & n6963 ;
  assign n6966 = n6964 & ~n6965 ;
  assign n6967 = x71 & n5340 ;
  assign n6968 = x70 & n5335 ;
  assign n6969 = x69 & ~n5334 ;
  assign n6970 = n5580 & n6969 ;
  assign n6971 = n6968 | n6970 ;
  assign n6972 = n6967 | n6971 ;
  assign n6973 = n5343 | n6972 ;
  assign n6974 = ( n376 & n6972 ) | ( n376 & n6973 ) | ( n6972 & n6973 ) ;
  assign n6975 = x41 & ~n6974 ;
  assign n6976 = ~x41 & n6974 ;
  assign n6977 = n6975 | n6976 ;
  assign n6978 = n6966 & n6977 ;
  assign n6979 = n6966 & ~n6978 ;
  assign n6980 = ~n6966 & n6977 ;
  assign n6981 = n6979 | n6980 ;
  assign n6982 = n6703 | n6709 ;
  assign n6983 = n6981 | n6982 ;
  assign n6984 = n6981 & n6982 ;
  assign n6985 = n6983 & ~n6984 ;
  assign n6986 = x74 & n4572 ;
  assign n6987 = x73 & n4567 ;
  assign n6988 = x72 & ~n4566 ;
  assign n6989 = n4828 & n6988 ;
  assign n6990 = n6987 | n6989 ;
  assign n6991 = n6986 | n6990 ;
  assign n6992 = n4575 | n6991 ;
  assign n6993 = ( n587 & n6991 ) | ( n587 & n6992 ) | ( n6991 & n6992 ) ;
  assign n6994 = x38 & n6993 ;
  assign n6995 = x38 & ~n6994 ;
  assign n6996 = ( n6993 & ~n6994 ) | ( n6993 & n6995 ) | ( ~n6994 & n6995 ) ;
  assign n6997 = n6985 | n6996 ;
  assign n6998 = n6928 & n6997 ;
  assign n6999 = n6985 & n6996 ;
  assign n7000 = n6997 & ~n6999 ;
  assign n7001 = ~n6998 & n7000 ;
  assign n7002 = x77 & n3913 ;
  assign n7003 = x76 & n3908 ;
  assign n7004 = x75 & ~n3907 ;
  assign n7005 = n4152 & n7004 ;
  assign n7006 = n7003 | n7005 ;
  assign n7007 = n7002 | n7006 ;
  assign n7008 = n3916 | n7007 ;
  assign n7009 = ( n846 & n7007 ) | ( n846 & n7008 ) | ( n7007 & n7008 ) ;
  assign n7010 = x35 & n7009 ;
  assign n7011 = x35 & ~n7010 ;
  assign n7012 = ( n7009 & ~n7010 ) | ( n7009 & n7011 ) | ( ~n7010 & n7011 ) ;
  assign n7013 = n7001 | n7012 ;
  assign n7014 = n6928 & ~n7000 ;
  assign n7015 = n7013 | n7014 ;
  assign n7016 = ( n7001 & n7012 ) | ( n7001 & n7014 ) | ( n7012 & n7014 ) ;
  assign n7017 = n7015 & ~n7016 ;
  assign n7018 = n6927 & n7017 ;
  assign n7019 = n6927 | n7017 ;
  assign n7020 = ~n7018 & n7019 ;
  assign n7021 = x80 & n3314 ;
  assign n7022 = x79 & n3309 ;
  assign n7023 = x78 & ~n3308 ;
  assign n7024 = n3570 & n7023 ;
  assign n7025 = n7022 | n7024 ;
  assign n7026 = n7021 | n7025 ;
  assign n7027 = n3317 | n7026 ;
  assign n7028 = ( n1147 & n7026 ) | ( n1147 & n7027 ) | ( n7026 & n7027 ) ;
  assign n7029 = x32 & n7028 ;
  assign n7030 = x32 & ~n7029 ;
  assign n7031 = ( n7028 & ~n7029 ) | ( n7028 & n7030 ) | ( ~n7029 & n7030 ) ;
  assign n7032 = n7020 & n7031 ;
  assign n7033 = n7020 & ~n7032 ;
  assign n7034 = ~n7020 & n7031 ;
  assign n7035 = n7033 | n7034 ;
  assign n7036 = ( n6672 & n6747 ) | ( n6672 & n6758 ) | ( n6747 & n6758 ) ;
  assign n7037 = n7035 | n7036 ;
  assign n7038 = n7035 & n7036 ;
  assign n7039 = n7037 & ~n7038 ;
  assign n7040 = x83 & n2775 ;
  assign n7041 = x82 & n2770 ;
  assign n7042 = x81 & ~n2769 ;
  assign n7043 = n2978 & n7042 ;
  assign n7044 = n7041 | n7043 ;
  assign n7045 = n7040 | n7044 ;
  assign n7046 = n2778 | n7045 ;
  assign n7047 = ( n1510 & n7045 ) | ( n1510 & n7046 ) | ( n7045 & n7046 ) ;
  assign n7048 = x29 & n7047 ;
  assign n7049 = x29 & ~n7048 ;
  assign n7050 = ( n7047 & ~n7048 ) | ( n7047 & n7049 ) | ( ~n7048 & n7049 ) ;
  assign n7051 = n7039 & n7050 ;
  assign n7052 = n7039 & ~n7051 ;
  assign n7053 = ~n7039 & n7050 ;
  assign n7054 = n7052 | n7053 ;
  assign n7055 = n6773 | n6776 ;
  assign n7056 = n7054 | n7055 ;
  assign n7057 = n7054 & n7055 ;
  assign n7058 = n7056 & ~n7057 ;
  assign n7059 = x86 & n2280 ;
  assign n7060 = x85 & n2275 ;
  assign n7061 = x84 & ~n2274 ;
  assign n7062 = n2481 & n7061 ;
  assign n7063 = n7060 | n7062 ;
  assign n7064 = n7059 | n7063 ;
  assign n7065 = n2283 | n7064 ;
  assign n7066 = ( n1921 & n7064 ) | ( n1921 & n7065 ) | ( n7064 & n7065 ) ;
  assign n7067 = x26 & n7066 ;
  assign n7068 = x26 & ~n7067 ;
  assign n7069 = ( n7066 & ~n7067 ) | ( n7066 & n7068 ) | ( ~n7067 & n7068 ) ;
  assign n7070 = n7058 & n7069 ;
  assign n7071 = n7058 & ~n7070 ;
  assign n7072 = ~n7058 & n7069 ;
  assign n7073 = n7071 | n7072 ;
  assign n7074 = n6790 | n6796 ;
  assign n7075 = n7073 | n7074 ;
  assign n7076 = n7073 & n7074 ;
  assign n7077 = n7075 & ~n7076 ;
  assign n7078 = x89 & n1817 ;
  assign n7079 = x88 & n1812 ;
  assign n7080 = x87 & ~n1811 ;
  assign n7081 = n1977 & n7080 ;
  assign n7082 = n7079 | n7081 ;
  assign n7083 = n7078 | n7082 ;
  assign n7084 = n1820 | n7083 ;
  assign n7085 = ( n2244 & n7083 ) | ( n2244 & n7084 ) | ( n7083 & n7084 ) ;
  assign n7086 = x23 & n7085 ;
  assign n7087 = x23 & ~n7086 ;
  assign n7088 = ( n7085 & ~n7086 ) | ( n7085 & n7087 ) | ( ~n7086 & n7087 ) ;
  assign n7089 = n7077 & n7088 ;
  assign n7090 = n7077 & ~n7089 ;
  assign n7091 = ~n7077 & n7088 ;
  assign n7092 = n7090 | n7091 ;
  assign n7093 = n6810 | n6812 ;
  assign n7094 = n7092 & n7093 ;
  assign n7095 = n7092 | n7093 ;
  assign n7096 = ~n7094 & n7095 ;
  assign n7097 = x92 & n1421 ;
  assign n7098 = x91 & n1416 ;
  assign n7099 = x90 & ~n1415 ;
  assign n7100 = n1584 & n7099 ;
  assign n7101 = n7098 | n7100 ;
  assign n7102 = n7097 | n7101 ;
  assign n7103 = n1424 | n7102 ;
  assign n7104 = ( n2904 & n7102 ) | ( n2904 & n7103 ) | ( n7102 & n7103 ) ;
  assign n7105 = x20 & n7104 ;
  assign n7106 = x20 & ~n7105 ;
  assign n7107 = ( n7104 & ~n7105 ) | ( n7104 & n7106 ) | ( ~n7105 & n7106 ) ;
  assign n7108 = ~n7096 & n7107 ;
  assign n7109 = n7096 & ~n7107 ;
  assign n7110 = n7108 | n7109 ;
  assign n7111 = ( n6669 & n6670 ) | ( n6669 & n6814 ) | ( n6670 & n6814 ) ;
  assign n7112 = n7110 & ~n7111 ;
  assign n7113 = ~n7110 & n7111 ;
  assign n7114 = x95 & n1071 ;
  assign n7115 = x94 & n1066 ;
  assign n7116 = x93 & ~n1065 ;
  assign n7117 = n1189 & n7116 ;
  assign n7118 = n7115 | n7117 ;
  assign n7119 = n7114 | n7118 ;
  assign n7120 = n1074 | n7119 ;
  assign n7121 = ( n3479 & n7119 ) | ( n3479 & n7120 ) | ( n7119 & n7120 ) ;
  assign n7122 = x17 & n7121 ;
  assign n7123 = x17 & ~n7122 ;
  assign n7124 = ( n7121 & ~n7122 ) | ( n7121 & n7123 ) | ( ~n7122 & n7123 ) ;
  assign n7125 = n7113 | n7124 ;
  assign n7126 = n7112 | n7125 ;
  assign n7127 = ( n7112 & n7113 ) | ( n7112 & n7124 ) | ( n7113 & n7124 ) ;
  assign n7128 = n7126 & ~n7127 ;
  assign n7129 = n6926 & n7128 ;
  assign n7130 = n6926 | n7128 ;
  assign n7131 = ~n7129 & n7130 ;
  assign n7132 = x98 & n771 ;
  assign n7133 = x97 & n766 ;
  assign n7134 = x96 & ~n765 ;
  assign n7135 = n905 & n7134 ;
  assign n7136 = n7133 | n7135 ;
  assign n7137 = n7132 | n7136 ;
  assign n7138 = n774 | n7137 ;
  assign n7139 = ( n4105 & n7137 ) | ( n4105 & n7138 ) | ( n7137 & n7138 ) ;
  assign n7140 = x14 & n7139 ;
  assign n7141 = x14 & ~n7140 ;
  assign n7142 = ( n7139 & ~n7140 ) | ( n7139 & n7141 ) | ( ~n7140 & n7141 ) ;
  assign n7143 = n7131 & n7142 ;
  assign n7144 = n7131 & ~n7143 ;
  assign n7145 = ~n7131 & n7142 ;
  assign n7146 = n7144 | n7145 ;
  assign n7147 = n6826 | n7146 ;
  assign n7148 = n6826 & n7146 ;
  assign n7149 = n7147 & ~n7148 ;
  assign n7150 = x101 & n528 ;
  assign n7151 = x100 & n523 ;
  assign n7152 = x99 & ~n522 ;
  assign n7153 = n635 & n7152 ;
  assign n7154 = n7151 | n7153 ;
  assign n7155 = n7150 | n7154 ;
  assign n7156 = n531 | n7155 ;
  assign n7157 = ( n4783 & n7155 ) | ( n4783 & n7156 ) | ( n7155 & n7156 ) ;
  assign n7158 = x11 & n7157 ;
  assign n7159 = x11 & ~n7158 ;
  assign n7160 = ( n7157 & ~n7158 ) | ( n7157 & n7159 ) | ( ~n7158 & n7159 ) ;
  assign n7161 = n7149 & n7160 ;
  assign n7162 = n7149 & ~n7161 ;
  assign n7163 = ~n7149 & n7160 ;
  assign n7164 = n7162 | n7163 ;
  assign n7165 = n6829 | n6834 ;
  assign n7166 = n7164 | n7165 ;
  assign n7167 = n7164 & n7165 ;
  assign n7168 = n7166 & ~n7167 ;
  assign n7169 = ( n6924 & n6925 ) | ( n6924 & ~n7168 ) | ( n6925 & ~n7168 ) ;
  assign n7170 = ( ~n6925 & n7168 ) | ( ~n6925 & n7169 ) | ( n7168 & n7169 ) ;
  assign n7171 = ( ~n6924 & n7169 ) | ( ~n6924 & n7170 ) | ( n7169 & n7170 ) ;
  assign n7172 = n6913 & n7171 ;
  assign n7173 = n6913 | n7171 ;
  assign n7174 = ~n7172 & n7173 ;
  assign n7175 = n6866 | n6872 ;
  assign n7176 = n7174 | n7175 ;
  assign n7177 = n7174 & n7175 ;
  assign n7178 = n7176 & ~n7177 ;
  assign n7179 = x109 | x110 ;
  assign n7180 = x109 & x110 ;
  assign n7181 = n7179 & ~n7180 ;
  assign n7182 = n6875 | n6878 ;
  assign n7183 = n7181 & n7182 ;
  assign n7184 = n6875 | n6880 ;
  assign n7185 = n7181 & n7184 ;
  assign n7186 = ( n5786 & n7183 ) | ( n5786 & n7185 ) | ( n7183 & n7185 ) ;
  assign n7187 = ( n5786 & n7182 ) | ( n5786 & n7184 ) | ( n7182 & n7184 ) ;
  assign n7188 = n7181 | n7187 ;
  assign n7189 = ~n7186 & n7188 ;
  assign n7190 = x109 & n131 ;
  assign n7191 = x108 & ~n156 ;
  assign n7192 = ( n135 & n7190 ) | ( n135 & n7191 ) | ( n7190 & n7191 ) ;
  assign n7193 = x0 & x110 ;
  assign n7194 = ( ~n135 & n7190 ) | ( ~n135 & n7193 ) | ( n7190 & n7193 ) ;
  assign n7195 = n7192 | n7194 ;
  assign n7196 = n139 | n7195 ;
  assign n7197 = ( n7189 & n7195 ) | ( n7189 & n7196 ) | ( n7195 & n7196 ) ;
  assign n7198 = x2 & n7197 ;
  assign n7199 = x2 & ~n7198 ;
  assign n7200 = ( n7197 & ~n7198 ) | ( n7197 & n7199 ) | ( ~n7198 & n7199 ) ;
  assign n7201 = n7178 & n7200 ;
  assign n7202 = n7178 & ~n7201 ;
  assign n7203 = ~n7178 & n7200 ;
  assign n7204 = n7202 | n7203 ;
  assign n7205 = n6897 | n6901 ;
  assign n7206 = n7204 & n7205 ;
  assign n7207 = n7204 | n7205 ;
  assign n7208 = ~n7206 & n7207 ;
  assign n7209 = n7172 | n7177 ;
  assign n7210 = n7127 | n7129 ;
  assign n7211 = n7070 | n7076 ;
  assign n7212 = n7032 | n7038 ;
  assign n7213 = n6978 | n6984 ;
  assign n7214 = x66 & n6937 ;
  assign n7215 = x65 & n6932 ;
  assign n7216 = ~n6676 & n6936 ;
  assign n7217 = x64 & ~n6931 ;
  assign n7218 = n7216 & n7217 ;
  assign n7219 = n7215 | n7218 ;
  assign n7220 = n7214 | n7219 ;
  assign n7221 = n153 & n6940 ;
  assign n7222 = n7220 | n7221 ;
  assign n7223 = x47 | n7222 ;
  assign n7224 = ~x47 & n7223 ;
  assign n7225 = ( ~n7222 & n7223 ) | ( ~n7222 & n7224 ) | ( n7223 & n7224 ) ;
  assign n7226 = n6947 | n7225 ;
  assign n7227 = n6947 & n7225 ;
  assign n7228 = n7226 & ~n7227 ;
  assign n7229 = n264 & n6071 ;
  assign n7230 = x69 & n6068 ;
  assign n7231 = x68 & n6063 ;
  assign n7232 = x67 & ~n6062 ;
  assign n7233 = n6398 & n7232 ;
  assign n7234 = n7231 | n7233 ;
  assign n7235 = n7230 | n7234 ;
  assign n7236 = n7229 | n7235 ;
  assign n7237 = x44 | n7236 ;
  assign n7238 = ~x44 & n7237 ;
  assign n7239 = ( ~n7236 & n7237 ) | ( ~n7236 & n7238 ) | ( n7237 & n7238 ) ;
  assign n7240 = n7228 & n7239 ;
  assign n7241 = n7228 & ~n7240 ;
  assign n7242 = ~n7228 & n7239 ;
  assign n7243 = n7241 | n7242 ;
  assign n7244 = n6962 | n6965 ;
  assign n7245 = n7243 & n7244 ;
  assign n7246 = n7243 | n7244 ;
  assign n7247 = ~n7245 & n7246 ;
  assign n7248 = x72 & n5340 ;
  assign n7249 = x71 & n5335 ;
  assign n7250 = x70 & ~n5334 ;
  assign n7251 = n5580 & n7250 ;
  assign n7252 = n7249 | n7251 ;
  assign n7253 = n7248 | n7252 ;
  assign n7254 = ( n435 & n5343 ) | ( n435 & n7253 ) | ( n5343 & n7253 ) ;
  assign n7255 = ( x41 & ~n7253 ) | ( x41 & n7254 ) | ( ~n7253 & n7254 ) ;
  assign n7256 = ~n7254 & n7255 ;
  assign n7257 = n7253 | n7255 ;
  assign n7258 = ( ~x41 & n7256 ) | ( ~x41 & n7257 ) | ( n7256 & n7257 ) ;
  assign n7259 = ~n7247 & n7258 ;
  assign n7260 = n7247 & ~n7258 ;
  assign n7261 = n7259 | n7260 ;
  assign n7262 = n7213 & ~n7261 ;
  assign n7263 = ~n7213 & n7261 ;
  assign n7264 = x75 & n4572 ;
  assign n7265 = x74 & n4567 ;
  assign n7266 = x73 & ~n4566 ;
  assign n7267 = n4828 & n7266 ;
  assign n7268 = n7265 | n7267 ;
  assign n7269 = n7264 | n7268 ;
  assign n7270 = n4575 | n7269 ;
  assign n7271 = ( n609 & n7269 ) | ( n609 & n7270 ) | ( n7269 & n7270 ) ;
  assign n7272 = x38 & n7271 ;
  assign n7273 = x38 & ~n7272 ;
  assign n7274 = ( n7271 & ~n7272 ) | ( n7271 & n7273 ) | ( ~n7272 & n7273 ) ;
  assign n7275 = n7263 | n7274 ;
  assign n7276 = n7262 | n7275 ;
  assign n7277 = ( n7262 & n7263 ) | ( n7262 & n7274 ) | ( n7263 & n7274 ) ;
  assign n7278 = n7276 & ~n7277 ;
  assign n7279 = n6998 | n6999 ;
  assign n7280 = n7278 & n7279 ;
  assign n7281 = n7278 | n7279 ;
  assign n7282 = ~n7280 & n7281 ;
  assign n7283 = x78 & n3913 ;
  assign n7284 = x77 & n3908 ;
  assign n7285 = x76 & ~n3907 ;
  assign n7286 = n4152 & n7285 ;
  assign n7287 = n7284 | n7286 ;
  assign n7288 = n7283 | n7287 ;
  assign n7289 = n3916 | n7288 ;
  assign n7290 = ( n868 & n7288 ) | ( n868 & n7289 ) | ( n7288 & n7289 ) ;
  assign n7291 = x35 & n7290 ;
  assign n7292 = x35 & ~n7291 ;
  assign n7293 = ( n7290 & ~n7291 ) | ( n7290 & n7292 ) | ( ~n7291 & n7292 ) ;
  assign n7294 = n7282 & n7293 ;
  assign n7295 = n7282 & ~n7294 ;
  assign n7296 = ~n7282 & n7293 ;
  assign n7297 = n7295 | n7296 ;
  assign n7298 = n7016 | n7018 ;
  assign n7299 = n7297 & n7298 ;
  assign n7300 = n7297 | n7298 ;
  assign n7301 = ~n7299 & n7300 ;
  assign n7302 = x81 & n3314 ;
  assign n7303 = x80 & n3309 ;
  assign n7304 = x79 & ~n3308 ;
  assign n7305 = n3570 & n7304 ;
  assign n7306 = n7303 | n7305 ;
  assign n7307 = n7302 | n7306 ;
  assign n7308 = n3317 | n7307 ;
  assign n7309 = ( n1256 & n7307 ) | ( n1256 & n7308 ) | ( n7307 & n7308 ) ;
  assign n7310 = x32 & n7309 ;
  assign n7311 = x32 & ~n7310 ;
  assign n7312 = ( n7309 & ~n7310 ) | ( n7309 & n7311 ) | ( ~n7310 & n7311 ) ;
  assign n7313 = ~n7301 & n7312 ;
  assign n7314 = n7301 & ~n7312 ;
  assign n7315 = n7313 | n7314 ;
  assign n7316 = ~n7212 & n7315 ;
  assign n7317 = n7212 & ~n7315 ;
  assign n7318 = n7316 | n7317 ;
  assign n7319 = x84 & n2775 ;
  assign n7320 = x83 & n2770 ;
  assign n7321 = x82 & ~n2769 ;
  assign n7322 = n2978 & n7321 ;
  assign n7323 = n7320 | n7322 ;
  assign n7324 = n7319 | n7323 ;
  assign n7325 = n2778 | n7324 ;
  assign n7326 = ( n1537 & n7324 ) | ( n1537 & n7325 ) | ( n7324 & n7325 ) ;
  assign n7327 = x29 & n7326 ;
  assign n7328 = x29 & ~n7327 ;
  assign n7329 = ( n7326 & ~n7327 ) | ( n7326 & n7328 ) | ( ~n7327 & n7328 ) ;
  assign n7330 = n7318 & n7329 ;
  assign n7331 = n7318 | n7329 ;
  assign n7332 = ~n7330 & n7331 ;
  assign n7333 = n7051 | n7057 ;
  assign n7334 = n7332 | n7333 ;
  assign n7335 = n7332 & n7333 ;
  assign n7336 = n7334 & ~n7335 ;
  assign n7337 = x87 & n2280 ;
  assign n7338 = x86 & n2275 ;
  assign n7339 = x85 & ~n2274 ;
  assign n7340 = n2481 & n7339 ;
  assign n7341 = n7338 | n7340 ;
  assign n7342 = n7337 | n7341 ;
  assign n7343 = n2283 | n7342 ;
  assign n7344 = ( n2067 & n7342 ) | ( n2067 & n7343 ) | ( n7342 & n7343 ) ;
  assign n7345 = x26 & n7344 ;
  assign n7346 = x26 & ~n7345 ;
  assign n7347 = ( n7344 & ~n7345 ) | ( n7344 & n7346 ) | ( ~n7345 & n7346 ) ;
  assign n7348 = n7336 | n7347 ;
  assign n7349 = n7211 & n7348 ;
  assign n7350 = n7336 & n7347 ;
  assign n7351 = n7348 & ~n7350 ;
  assign n7352 = ~n7349 & n7351 ;
  assign n7353 = x90 & n1817 ;
  assign n7354 = x89 & n1812 ;
  assign n7355 = x88 & ~n1811 ;
  assign n7356 = n1977 & n7355 ;
  assign n7357 = n7354 | n7356 ;
  assign n7358 = n7353 | n7357 ;
  assign n7359 = n1820 | n7358 ;
  assign n7360 = ( n2410 & n7358 ) | ( n2410 & n7359 ) | ( n7358 & n7359 ) ;
  assign n7361 = x23 & n7360 ;
  assign n7362 = x23 & ~n7361 ;
  assign n7363 = ( n7360 & ~n7361 ) | ( n7360 & n7362 ) | ( ~n7361 & n7362 ) ;
  assign n7364 = n7352 | n7363 ;
  assign n7365 = n7211 & ~n7351 ;
  assign n7366 = n7364 | n7365 ;
  assign n7367 = ( n7352 & n7363 ) | ( n7352 & n7365 ) | ( n7363 & n7365 ) ;
  assign n7368 = n7366 & ~n7367 ;
  assign n7369 = n7089 | n7094 ;
  assign n7370 = n7368 & n7369 ;
  assign n7371 = n7368 | n7369 ;
  assign n7372 = ~n7370 & n7371 ;
  assign n7373 = x93 & n1421 ;
  assign n7374 = x92 & n1416 ;
  assign n7375 = x91 & ~n1415 ;
  assign n7376 = n1584 & n7375 ;
  assign n7377 = n7374 | n7376 ;
  assign n7378 = n7373 | n7377 ;
  assign n7379 = n1424 | n7378 ;
  assign n7380 = ( n2931 & n7378 ) | ( n2931 & n7379 ) | ( n7378 & n7379 ) ;
  assign n7381 = x20 & n7380 ;
  assign n7382 = x20 & ~n7381 ;
  assign n7383 = ( n7380 & ~n7381 ) | ( n7380 & n7382 ) | ( ~n7381 & n7382 ) ;
  assign n7384 = n7372 | n7383 ;
  assign n7385 = n7372 & n7383 ;
  assign n7386 = n7384 & ~n7385 ;
  assign n7387 = ( n7096 & n7107 ) | ( n7096 & n7111 ) | ( n7107 & n7111 ) ;
  assign n7388 = n7386 & n7387 ;
  assign n7389 = n7386 | n7387 ;
  assign n7390 = ~n7388 & n7389 ;
  assign n7391 = x96 & n1071 ;
  assign n7392 = x95 & n1066 ;
  assign n7393 = x94 & ~n1065 ;
  assign n7394 = n1189 & n7393 ;
  assign n7395 = n7392 | n7394 ;
  assign n7396 = n7391 | n7395 ;
  assign n7397 = n1074 | n7396 ;
  assign n7398 = ( n3509 & n7396 ) | ( n3509 & n7397 ) | ( n7396 & n7397 ) ;
  assign n7399 = x17 & n7398 ;
  assign n7400 = x17 & ~n7399 ;
  assign n7401 = ( n7398 & ~n7399 ) | ( n7398 & n7400 ) | ( ~n7399 & n7400 ) ;
  assign n7402 = n7390 | n7401 ;
  assign n7403 = n7390 & n7401 ;
  assign n7404 = n7402 & ~n7403 ;
  assign n7405 = n7210 & n7404 ;
  assign n7406 = n7210 | n7404 ;
  assign n7407 = ~n7405 & n7406 ;
  assign n7408 = x99 & n771 ;
  assign n7409 = x98 & n766 ;
  assign n7410 = x97 & ~n765 ;
  assign n7411 = n905 & n7410 ;
  assign n7412 = n7409 | n7411 ;
  assign n7413 = n7408 | n7412 ;
  assign n7414 = n774 | n7413 ;
  assign n7415 = ( n4325 & n7413 ) | ( n4325 & n7414 ) | ( n7413 & n7414 ) ;
  assign n7416 = x14 & n7415 ;
  assign n7417 = x14 & ~n7416 ;
  assign n7418 = ( n7415 & ~n7416 ) | ( n7415 & n7417 ) | ( ~n7416 & n7417 ) ;
  assign n7419 = n7407 & n7418 ;
  assign n7420 = n7407 & ~n7419 ;
  assign n7421 = ~n7407 & n7418 ;
  assign n7422 = n7420 | n7421 ;
  assign n7423 = n7143 | n7148 ;
  assign n7424 = n7422 | n7423 ;
  assign n7425 = n7422 & n7423 ;
  assign n7426 = n7424 & ~n7425 ;
  assign n7427 = x102 & n528 ;
  assign n7428 = x101 & n523 ;
  assign n7429 = x100 & ~n522 ;
  assign n7430 = n635 & n7429 ;
  assign n7431 = n7428 | n7430 ;
  assign n7432 = n7427 | n7431 ;
  assign n7433 = n531 | n7432 ;
  assign n7434 = ( n5025 & n7432 ) | ( n5025 & n7433 ) | ( n7432 & n7433 ) ;
  assign n7435 = x11 & n7434 ;
  assign n7436 = x11 & ~n7435 ;
  assign n7437 = ( n7434 & ~n7435 ) | ( n7434 & n7436 ) | ( ~n7435 & n7436 ) ;
  assign n7438 = n7426 & n7437 ;
  assign n7439 = n7426 & ~n7438 ;
  assign n7440 = ~n7426 & n7437 ;
  assign n7441 = n7439 | n7440 ;
  assign n7442 = n7161 | n7167 ;
  assign n7443 = n7441 | n7442 ;
  assign n7444 = n7441 & n7442 ;
  assign n7445 = n7443 & ~n7444 ;
  assign n7446 = x105 & n337 ;
  assign n7447 = x104 & n332 ;
  assign n7448 = x103 & ~n331 ;
  assign n7449 = n396 & n7448 ;
  assign n7450 = n7447 | n7449 ;
  assign n7451 = n7446 | n7450 ;
  assign n7452 = n340 | n7451 ;
  assign n7453 = ( n5788 & n7451 ) | ( n5788 & n7452 ) | ( n7451 & n7452 ) ;
  assign n7454 = x8 & n7453 ;
  assign n7455 = x8 & ~n7454 ;
  assign n7456 = ( n7453 & ~n7454 ) | ( n7453 & n7455 ) | ( ~n7454 & n7455 ) ;
  assign n7457 = n7445 & n7456 ;
  assign n7458 = n7445 | n7456 ;
  assign n7459 = ~n7457 & n7458 ;
  assign n7460 = n6924 | n7168 ;
  assign n7461 = n6925 & n7460 ;
  assign n7462 = n6924 & n7168 ;
  assign n7463 = n7461 | n7462 ;
  assign n7464 = n7459 & n7463 ;
  assign n7465 = n7463 & ~n7464 ;
  assign n7466 = ( n7459 & ~n7464 ) | ( n7459 & n7465 ) | ( ~n7464 & n7465 ) ;
  assign n7467 = x108 & n206 ;
  assign n7468 = x107 & n201 ;
  assign n7469 = x106 & ~n200 ;
  assign n7470 = n243 & n7469 ;
  assign n7471 = n7468 | n7470 ;
  assign n7472 = n7467 | n7471 ;
  assign n7473 = n209 | n7472 ;
  assign n7474 = ( n6358 & n7472 ) | ( n6358 & n7473 ) | ( n7472 & n7473 ) ;
  assign n7475 = x5 & n7474 ;
  assign n7476 = x5 & ~n7475 ;
  assign n7477 = ( n7474 & ~n7475 ) | ( n7474 & n7476 ) | ( ~n7475 & n7476 ) ;
  assign n7478 = n7466 | n7477 ;
  assign n7479 = n7466 & n7477 ;
  assign n7480 = n7478 & ~n7479 ;
  assign n7481 = n7209 & n7480 ;
  assign n7482 = n7209 | n7480 ;
  assign n7483 = ~n7481 & n7482 ;
  assign n7484 = x110 | x111 ;
  assign n7485 = x110 & x111 ;
  assign n7486 = n7484 & ~n7485 ;
  assign n7487 = n7180 | n7183 ;
  assign n7488 = n7180 | n7185 ;
  assign n7489 = ( n5786 & n7487 ) | ( n5786 & n7488 ) | ( n7487 & n7488 ) ;
  assign n7490 = n7486 | n7489 ;
  assign n7491 = n7486 & n7489 ;
  assign n7492 = n7490 & ~n7491 ;
  assign n7493 = x110 & n131 ;
  assign n7494 = x109 & ~n156 ;
  assign n7495 = ( n135 & n7493 ) | ( n135 & n7494 ) | ( n7493 & n7494 ) ;
  assign n7496 = x0 & x111 ;
  assign n7497 = ( ~n135 & n7493 ) | ( ~n135 & n7496 ) | ( n7493 & n7496 ) ;
  assign n7498 = n7495 | n7497 ;
  assign n7499 = n139 | n7498 ;
  assign n7500 = ( n7492 & n7498 ) | ( n7492 & n7499 ) | ( n7498 & n7499 ) ;
  assign n7501 = x2 & n7500 ;
  assign n7502 = x2 & ~n7501 ;
  assign n7503 = ( n7500 & ~n7501 ) | ( n7500 & n7502 ) | ( ~n7501 & n7502 ) ;
  assign n7504 = n7483 & n7503 ;
  assign n7505 = n7483 & ~n7504 ;
  assign n7506 = ~n7483 & n7503 ;
  assign n7507 = n7505 | n7506 ;
  assign n7508 = n7201 | n7206 ;
  assign n7509 = n7507 & n7508 ;
  assign n7510 = n7507 | n7508 ;
  assign n7511 = ~n7509 & n7510 ;
  assign n7512 = n7504 | n7509 ;
  assign n7513 = x109 & n206 ;
  assign n7514 = x108 & n201 ;
  assign n7515 = x107 & ~n200 ;
  assign n7516 = n243 & n7515 ;
  assign n7517 = n7514 | n7516 ;
  assign n7518 = n7513 | n7517 ;
  assign n7519 = n209 | n7518 ;
  assign n7520 = ( n6884 & n7518 ) | ( n6884 & n7519 ) | ( n7518 & n7519 ) ;
  assign n7521 = x5 & n7520 ;
  assign n7522 = x5 & ~n7521 ;
  assign n7523 = ( n7520 & ~n7521 ) | ( n7520 & n7522 ) | ( ~n7521 & n7522 ) ;
  assign n7524 = x106 & n337 ;
  assign n7525 = x105 & n332 ;
  assign n7526 = x104 & ~n331 ;
  assign n7527 = n396 & n7526 ;
  assign n7528 = n7525 | n7527 ;
  assign n7529 = n7524 | n7528 ;
  assign n7530 = n340 | n7529 ;
  assign n7531 = ( n5814 & n7529 ) | ( n5814 & n7530 ) | ( n7529 & n7530 ) ;
  assign n7532 = x8 & n7531 ;
  assign n7533 = x8 & ~n7532 ;
  assign n7534 = ( n7531 & ~n7532 ) | ( n7531 & n7533 ) | ( ~n7532 & n7533 ) ;
  assign n7535 = n7457 | n7464 ;
  assign n7536 = x100 & n771 ;
  assign n7537 = x99 & n766 ;
  assign n7538 = x98 & ~n765 ;
  assign n7539 = n905 & n7538 ;
  assign n7540 = n7537 | n7539 ;
  assign n7541 = n7536 | n7540 ;
  assign n7542 = n774 | n7541 ;
  assign n7543 = ( n4532 & n7541 ) | ( n4532 & n7542 ) | ( n7541 & n7542 ) ;
  assign n7544 = x14 & n7543 ;
  assign n7545 = x14 & ~n7544 ;
  assign n7546 = ( n7543 & ~n7544 ) | ( n7543 & n7545 ) | ( ~n7544 & n7545 ) ;
  assign n7547 = x97 & n1071 ;
  assign n7548 = x96 & n1066 ;
  assign n7549 = x95 & ~n1065 ;
  assign n7550 = n1189 & n7549 ;
  assign n7551 = n7548 | n7550 ;
  assign n7552 = n7547 | n7551 ;
  assign n7553 = n1074 | n7552 ;
  assign n7554 = ( n3707 & n7552 ) | ( n3707 & n7553 ) | ( n7552 & n7553 ) ;
  assign n7555 = x17 & n7554 ;
  assign n7556 = x17 & ~n7555 ;
  assign n7557 = ( n7554 & ~n7555 ) | ( n7554 & n7556 ) | ( ~n7555 & n7556 ) ;
  assign n7558 = x94 & n1421 ;
  assign n7559 = x93 & n1416 ;
  assign n7560 = x92 & ~n1415 ;
  assign n7561 = n1584 & n7560 ;
  assign n7562 = n7559 | n7561 ;
  assign n7563 = n7558 | n7562 ;
  assign n7564 = n1424 | n7563 ;
  assign n7565 = ( n3271 & n7563 ) | ( n3271 & n7564 ) | ( n7563 & n7564 ) ;
  assign n7566 = x20 & n7565 ;
  assign n7567 = x20 & ~n7566 ;
  assign n7568 = ( n7565 & ~n7566 ) | ( n7565 & n7567 ) | ( ~n7566 & n7567 ) ;
  assign n7569 = x91 & n1817 ;
  assign n7570 = x90 & n1812 ;
  assign n7571 = x89 & ~n1811 ;
  assign n7572 = n1977 & n7571 ;
  assign n7573 = n7570 | n7572 ;
  assign n7574 = n7569 | n7573 ;
  assign n7575 = n1820 | n7574 ;
  assign n7576 = ( n2714 & n7574 ) | ( n2714 & n7575 ) | ( n7574 & n7575 ) ;
  assign n7577 = x23 & n7576 ;
  assign n7578 = x23 & ~n7577 ;
  assign n7579 = ( n7576 & ~n7577 ) | ( n7576 & n7578 ) | ( ~n7577 & n7578 ) ;
  assign n7580 = n7367 | n7370 ;
  assign n7581 = n7294 | n7299 ;
  assign n7582 = n7277 | n7280 ;
  assign n7583 = x47 & ~x48 ;
  assign n7584 = ~x47 & x48 ;
  assign n7585 = n7583 | n7584 ;
  assign n7586 = x64 & n7585 ;
  assign n7587 = x67 & n6937 ;
  assign n7588 = x66 & n6932 ;
  assign n7589 = x65 & ~n6931 ;
  assign n7590 = n7216 & n7589 ;
  assign n7591 = n7588 | n7590 ;
  assign n7592 = n7587 | n7591 ;
  assign n7593 = n180 & n6940 ;
  assign n7594 = n7592 | n7593 ;
  assign n7595 = x47 & ~n7594 ;
  assign n7596 = ~x47 & n7594 ;
  assign n7597 = n7595 | n7596 ;
  assign n7598 = ( n7227 & n7586 ) | ( n7227 & n7597 ) | ( n7586 & n7597 ) ;
  assign n7599 = ( n7227 & n7597 ) | ( n7227 & ~n7598 ) | ( n7597 & ~n7598 ) ;
  assign n7600 = ( n7586 & ~n7598 ) | ( n7586 & n7599 ) | ( ~n7598 & n7599 ) ;
  assign n7601 = x70 & n6068 ;
  assign n7602 = x69 & n6063 ;
  assign n7603 = x68 & ~n6062 ;
  assign n7604 = n6398 & n7603 ;
  assign n7605 = n7602 | n7604 ;
  assign n7606 = n7601 | n7605 ;
  assign n7607 = n6071 | n7606 ;
  assign n7608 = ( n310 & n7606 ) | ( n310 & n7607 ) | ( n7606 & n7607 ) ;
  assign n7609 = x44 & ~n7608 ;
  assign n7610 = ~x44 & n7608 ;
  assign n7611 = n7609 | n7610 ;
  assign n7612 = n7600 & n7611 ;
  assign n7613 = n7600 & ~n7612 ;
  assign n7614 = ~n7600 & n7611 ;
  assign n7615 = n7613 | n7614 ;
  assign n7616 = n7240 | n7245 ;
  assign n7617 = n7615 | n7616 ;
  assign n7618 = n7615 & n7616 ;
  assign n7619 = n7617 & ~n7618 ;
  assign n7620 = x73 & n5340 ;
  assign n7621 = x72 & n5335 ;
  assign n7622 = x71 & ~n5334 ;
  assign n7623 = n5580 & n7622 ;
  assign n7624 = n7621 | n7623 ;
  assign n7625 = n7620 | n7624 ;
  assign n7626 = ( n499 & n5343 ) | ( n499 & n7625 ) | ( n5343 & n7625 ) ;
  assign n7627 = ( x41 & ~n7625 ) | ( x41 & n7626 ) | ( ~n7625 & n7626 ) ;
  assign n7628 = ~n7626 & n7627 ;
  assign n7629 = n7625 | n7627 ;
  assign n7630 = ( ~x41 & n7628 ) | ( ~x41 & n7629 ) | ( n7628 & n7629 ) ;
  assign n7631 = n7619 | n7630 ;
  assign n7632 = n7619 & n7630 ;
  assign n7633 = n7631 & ~n7632 ;
  assign n7634 = ( n7213 & n7247 ) | ( n7213 & n7258 ) | ( n7247 & n7258 ) ;
  assign n7635 = n7633 & n7634 ;
  assign n7636 = n7633 | n7634 ;
  assign n7637 = ~n7635 & n7636 ;
  assign n7638 = x76 & n4572 ;
  assign n7639 = x75 & n4567 ;
  assign n7640 = x74 & ~n4566 ;
  assign n7641 = n4828 & n7640 ;
  assign n7642 = n7639 | n7641 ;
  assign n7643 = n7638 | n7642 ;
  assign n7644 = n4575 | n7643 ;
  assign n7645 = ( n740 & n7643 ) | ( n740 & n7644 ) | ( n7643 & n7644 ) ;
  assign n7646 = x38 & n7645 ;
  assign n7647 = x38 & ~n7646 ;
  assign n7648 = ( n7645 & ~n7646 ) | ( n7645 & n7647 ) | ( ~n7646 & n7647 ) ;
  assign n7649 = n7637 & n7648 ;
  assign n7650 = n7637 & ~n7649 ;
  assign n7651 = ~n7637 & n7648 ;
  assign n7652 = n7650 | n7651 ;
  assign n7653 = n7582 & n7652 ;
  assign n7654 = n7582 | n7652 ;
  assign n7655 = ~n7653 & n7654 ;
  assign n7656 = x79 & n3913 ;
  assign n7657 = x78 & n3908 ;
  assign n7658 = x77 & ~n3907 ;
  assign n7659 = n4152 & n7658 ;
  assign n7660 = n7657 | n7659 ;
  assign n7661 = n7656 | n7660 ;
  assign n7662 = n3916 | n7661 ;
  assign n7663 = ( n961 & n7661 ) | ( n961 & n7662 ) | ( n7661 & n7662 ) ;
  assign n7664 = x35 & n7663 ;
  assign n7665 = x35 & ~n7664 ;
  assign n7666 = ( n7663 & ~n7664 ) | ( n7663 & n7665 ) | ( ~n7664 & n7665 ) ;
  assign n7667 = n7655 & n7666 ;
  assign n7668 = n7655 | n7666 ;
  assign n7669 = ~n7667 & n7668 ;
  assign n7670 = n7581 & n7669 ;
  assign n7671 = n7581 | n7669 ;
  assign n7672 = ~n7670 & n7671 ;
  assign n7673 = x82 & n3314 ;
  assign n7674 = x81 & n3309 ;
  assign n7675 = x80 & ~n3308 ;
  assign n7676 = n3570 & n7675 ;
  assign n7677 = n7674 | n7676 ;
  assign n7678 = n7673 | n7677 ;
  assign n7679 = n3317 | n7678 ;
  assign n7680 = ( n1371 & n7678 ) | ( n1371 & n7679 ) | ( n7678 & n7679 ) ;
  assign n7681 = x32 & n7680 ;
  assign n7682 = x32 & ~n7681 ;
  assign n7683 = ( n7680 & ~n7681 ) | ( n7680 & n7682 ) | ( ~n7681 & n7682 ) ;
  assign n7684 = n7672 & n7683 ;
  assign n7685 = n7672 & ~n7684 ;
  assign n7686 = ~n7672 & n7683 ;
  assign n7687 = n7685 | n7686 ;
  assign n7688 = ( n7212 & n7301 ) | ( n7212 & n7312 ) | ( n7301 & n7312 ) ;
  assign n7689 = n7687 | n7688 ;
  assign n7690 = n7687 & n7688 ;
  assign n7691 = n7689 & ~n7690 ;
  assign n7692 = x85 & n2775 ;
  assign n7693 = x84 & n2770 ;
  assign n7694 = x83 & ~n2769 ;
  assign n7695 = n2978 & n7694 ;
  assign n7696 = n7693 | n7695 ;
  assign n7697 = n7692 | n7696 ;
  assign n7698 = n2778 | n7697 ;
  assign n7699 = ( n1765 & n7697 ) | ( n1765 & n7698 ) | ( n7697 & n7698 ) ;
  assign n7700 = x29 & n7699 ;
  assign n7701 = x29 & ~n7700 ;
  assign n7702 = ( n7699 & ~n7700 ) | ( n7699 & n7701 ) | ( ~n7700 & n7701 ) ;
  assign n7703 = n7691 & n7702 ;
  assign n7704 = n7691 & ~n7703 ;
  assign n7705 = ~n7691 & n7702 ;
  assign n7706 = n7704 | n7705 ;
  assign n7707 = n7330 | n7335 ;
  assign n7708 = n7706 | n7707 ;
  assign n7709 = n7706 & n7707 ;
  assign n7710 = n7708 & ~n7709 ;
  assign n7711 = x88 & n2280 ;
  assign n7712 = x87 & n2275 ;
  assign n7713 = x86 & ~n2274 ;
  assign n7714 = n2481 & n7713 ;
  assign n7715 = n7712 | n7714 ;
  assign n7716 = n7711 | n7715 ;
  assign n7717 = n2283 | n7716 ;
  assign n7718 = ( n2095 & n7716 ) | ( n2095 & n7717 ) | ( n7716 & n7717 ) ;
  assign n7719 = x26 & n7718 ;
  assign n7720 = x26 & ~n7719 ;
  assign n7721 = ( n7718 & ~n7719 ) | ( n7718 & n7720 ) | ( ~n7719 & n7720 ) ;
  assign n7722 = n7710 | n7721 ;
  assign n7723 = n7710 & n7721 ;
  assign n7724 = n7722 & ~n7723 ;
  assign n7725 = n7349 | n7350 ;
  assign n7726 = n7724 & n7725 ;
  assign n7727 = n7724 | n7725 ;
  assign n7728 = ~n7726 & n7727 ;
  assign n7729 = ( n7579 & n7580 ) | ( n7579 & ~n7728 ) | ( n7580 & ~n7728 ) ;
  assign n7730 = ( ~n7580 & n7728 ) | ( ~n7580 & n7729 ) | ( n7728 & n7729 ) ;
  assign n7731 = ( ~n7579 & n7729 ) | ( ~n7579 & n7730 ) | ( n7729 & n7730 ) ;
  assign n7732 = n7568 & n7731 ;
  assign n7733 = n7568 | n7731 ;
  assign n7734 = ~n7732 & n7733 ;
  assign n7735 = n7385 | n7388 ;
  assign n7736 = n7734 & n7735 ;
  assign n7737 = n7734 | n7735 ;
  assign n7738 = ~n7736 & n7737 ;
  assign n7739 = n7403 | n7405 ;
  assign n7740 = ( n7557 & n7738 ) | ( n7557 & n7739 ) | ( n7738 & n7739 ) ;
  assign n7741 = ( n7738 & n7739 ) | ( n7738 & ~n7740 ) | ( n7739 & ~n7740 ) ;
  assign n7742 = ( n7557 & ~n7740 ) | ( n7557 & n7741 ) | ( ~n7740 & n7741 ) ;
  assign n7743 = n7546 & n7742 ;
  assign n7744 = n7546 | n7742 ;
  assign n7745 = ~n7743 & n7744 ;
  assign n7746 = n7419 | n7745 ;
  assign n7747 = n7425 | n7746 ;
  assign n7748 = ( n7419 & n7425 ) | ( n7419 & n7745 ) | ( n7425 & n7745 ) ;
  assign n7749 = n7747 & ~n7748 ;
  assign n7750 = x103 & n528 ;
  assign n7751 = x102 & n523 ;
  assign n7752 = x101 & ~n522 ;
  assign n7753 = n635 & n7752 ;
  assign n7754 = n7751 | n7753 ;
  assign n7755 = n7750 | n7754 ;
  assign n7756 = n531 | n7755 ;
  assign n7757 = ( n5264 & n7755 ) | ( n5264 & n7756 ) | ( n7755 & n7756 ) ;
  assign n7758 = x11 & n7757 ;
  assign n7759 = x11 & ~n7758 ;
  assign n7760 = ( n7757 & ~n7758 ) | ( n7757 & n7759 ) | ( ~n7758 & n7759 ) ;
  assign n7761 = n7749 & n7760 ;
  assign n7762 = n7749 & ~n7761 ;
  assign n7763 = ~n7749 & n7760 ;
  assign n7764 = n7762 | n7763 ;
  assign n7765 = n7438 | n7444 ;
  assign n7766 = n7764 | n7765 ;
  assign n7767 = n7764 & n7765 ;
  assign n7768 = n7766 & ~n7767 ;
  assign n7769 = ( n7534 & n7535 ) | ( n7534 & ~n7768 ) | ( n7535 & ~n7768 ) ;
  assign n7770 = ( ~n7535 & n7768 ) | ( ~n7535 & n7769 ) | ( n7768 & n7769 ) ;
  assign n7771 = ( ~n7534 & n7769 ) | ( ~n7534 & n7770 ) | ( n7769 & n7770 ) ;
  assign n7772 = n7523 & n7771 ;
  assign n7773 = n7523 | n7771 ;
  assign n7774 = ~n7772 & n7773 ;
  assign n7775 = n7479 | n7481 ;
  assign n7776 = n7774 & n7775 ;
  assign n7777 = n7774 | n7775 ;
  assign n7778 = ~n7776 & n7777 ;
  assign n7779 = x111 & n131 ;
  assign n7780 = x110 & ~n156 ;
  assign n7781 = ( n135 & n7779 ) | ( n135 & n7780 ) | ( n7779 & n7780 ) ;
  assign n7782 = x0 & x112 ;
  assign n7783 = ( ~n135 & n7779 ) | ( ~n135 & n7782 ) | ( n7779 & n7782 ) ;
  assign n7784 = n7781 | n7783 ;
  assign n7785 = n139 | n7784 ;
  assign n7786 = n7485 | n7491 ;
  assign n7787 = ( x111 & ~x112 ) | ( x111 & n7786 ) | ( ~x112 & n7786 ) ;
  assign n7788 = ( ~x111 & x112 ) | ( ~x111 & n7787 ) | ( x112 & n7787 ) ;
  assign n7789 = ( ~n7786 & n7787 ) | ( ~n7786 & n7788 ) | ( n7787 & n7788 ) ;
  assign n7790 = ( n7784 & n7785 ) | ( n7784 & n7789 ) | ( n7785 & n7789 ) ;
  assign n7791 = x2 & n7790 ;
  assign n7792 = x2 & ~n7791 ;
  assign n7793 = ( n7790 & ~n7791 ) | ( n7790 & n7792 ) | ( ~n7791 & n7792 ) ;
  assign n7794 = n7778 | n7793 ;
  assign n7795 = n7778 & n7793 ;
  assign n7796 = n7794 & ~n7795 ;
  assign n7797 = n7512 | n7796 ;
  assign n7798 = n7512 & n7796 ;
  assign n7799 = n7797 & ~n7798 ;
  assign n7800 = n7795 | n7798 ;
  assign n7801 = ( n7579 & n7580 ) | ( n7579 & n7728 ) | ( n7580 & n7728 ) ;
  assign n7802 = n7649 | n7653 ;
  assign n7803 = n7632 | n7635 ;
  assign n7804 = ~x48 & x49 ;
  assign n7805 = x48 & ~x49 ;
  assign n7806 = n7804 | n7805 ;
  assign n7807 = ~n7585 & n7806 ;
  assign n7808 = x64 & n7807 ;
  assign n7809 = ~x49 & x50 ;
  assign n7810 = x49 & ~x50 ;
  assign n7811 = n7809 | n7810 ;
  assign n7812 = n7585 & ~n7811 ;
  assign n7813 = x65 & n7812 ;
  assign n7814 = n7808 | n7813 ;
  assign n7815 = n7585 & n7811 ;
  assign n7816 = n142 & n7815 ;
  assign n7817 = n7814 | n7816 ;
  assign n7818 = x50 | n7817 ;
  assign n7819 = ~x50 & n7818 ;
  assign n7820 = ( ~n7817 & n7818 ) | ( ~n7817 & n7819 ) | ( n7818 & n7819 ) ;
  assign n7821 = x50 & ~n7586 ;
  assign n7822 = n7820 & n7821 ;
  assign n7823 = n7820 | n7821 ;
  assign n7824 = ~n7822 & n7823 ;
  assign n7825 = n229 & n6940 ;
  assign n7826 = x68 & n6937 ;
  assign n7827 = x67 & n6932 ;
  assign n7828 = x66 & ~n6931 ;
  assign n7829 = n7216 & n7828 ;
  assign n7830 = n7827 | n7829 ;
  assign n7831 = n7826 | n7830 ;
  assign n7832 = n7825 | n7831 ;
  assign n7833 = x47 | n7832 ;
  assign n7834 = ~x47 & n7833 ;
  assign n7835 = ( ~n7832 & n7833 ) | ( ~n7832 & n7834 ) | ( n7833 & n7834 ) ;
  assign n7836 = n7824 | n7835 ;
  assign n7837 = n7824 & n7835 ;
  assign n7838 = n7836 & ~n7837 ;
  assign n7839 = n7598 | n7838 ;
  assign n7840 = n7598 & n7838 ;
  assign n7841 = n7839 & ~n7840 ;
  assign n7842 = x71 & n6068 ;
  assign n7843 = x70 & n6063 ;
  assign n7844 = x69 & ~n6062 ;
  assign n7845 = n6398 & n7844 ;
  assign n7846 = n7843 | n7845 ;
  assign n7847 = n7842 | n7846 ;
  assign n7848 = n6071 | n7847 ;
  assign n7849 = ( n376 & n7847 ) | ( n376 & n7848 ) | ( n7847 & n7848 ) ;
  assign n7850 = x44 & ~n7849 ;
  assign n7851 = ~x44 & n7849 ;
  assign n7852 = n7850 | n7851 ;
  assign n7853 = n7841 & n7852 ;
  assign n7854 = n7841 & ~n7853 ;
  assign n7855 = ~n7841 & n7852 ;
  assign n7856 = n7854 | n7855 ;
  assign n7857 = n7612 | n7618 ;
  assign n7858 = n7856 | n7857 ;
  assign n7859 = n7856 & n7857 ;
  assign n7860 = n7858 & ~n7859 ;
  assign n7861 = x74 & n5340 ;
  assign n7862 = x73 & n5335 ;
  assign n7863 = x72 & ~n5334 ;
  assign n7864 = n5580 & n7863 ;
  assign n7865 = n7862 | n7864 ;
  assign n7866 = n7861 | n7865 ;
  assign n7867 = n5343 | n7866 ;
  assign n7868 = ( n587 & n7866 ) | ( n587 & n7867 ) | ( n7866 & n7867 ) ;
  assign n7869 = x41 & n7868 ;
  assign n7870 = x41 & ~n7869 ;
  assign n7871 = ( n7868 & ~n7869 ) | ( n7868 & n7870 ) | ( ~n7869 & n7870 ) ;
  assign n7872 = n7860 | n7871 ;
  assign n7873 = n7803 & n7872 ;
  assign n7874 = n7860 & n7871 ;
  assign n7875 = n7872 & ~n7874 ;
  assign n7876 = ~n7873 & n7875 ;
  assign n7877 = x77 & n4572 ;
  assign n7878 = x76 & n4567 ;
  assign n7879 = x75 & ~n4566 ;
  assign n7880 = n4828 & n7879 ;
  assign n7881 = n7878 | n7880 ;
  assign n7882 = n7877 | n7881 ;
  assign n7883 = n4575 | n7882 ;
  assign n7884 = ( n846 & n7882 ) | ( n846 & n7883 ) | ( n7882 & n7883 ) ;
  assign n7885 = x38 & n7884 ;
  assign n7886 = x38 & ~n7885 ;
  assign n7887 = ( n7884 & ~n7885 ) | ( n7884 & n7886 ) | ( ~n7885 & n7886 ) ;
  assign n7888 = n7876 | n7887 ;
  assign n7889 = n7803 & ~n7875 ;
  assign n7890 = n7888 | n7889 ;
  assign n7891 = ( n7876 & n7887 ) | ( n7876 & n7889 ) | ( n7887 & n7889 ) ;
  assign n7892 = n7890 & ~n7891 ;
  assign n7893 = n7802 & n7892 ;
  assign n7894 = n7802 | n7892 ;
  assign n7895 = ~n7893 & n7894 ;
  assign n7896 = x80 & n3913 ;
  assign n7897 = x79 & n3908 ;
  assign n7898 = x78 & ~n3907 ;
  assign n7899 = n4152 & n7898 ;
  assign n7900 = n7897 | n7899 ;
  assign n7901 = n7896 | n7900 ;
  assign n7902 = n3916 | n7901 ;
  assign n7903 = ( n1147 & n7901 ) | ( n1147 & n7902 ) | ( n7901 & n7902 ) ;
  assign n7904 = x35 & n7903 ;
  assign n7905 = x35 & ~n7904 ;
  assign n7906 = ( n7903 & ~n7904 ) | ( n7903 & n7905 ) | ( ~n7904 & n7905 ) ;
  assign n7907 = n7895 & n7906 ;
  assign n7908 = n7895 & ~n7907 ;
  assign n7909 = ~n7895 & n7906 ;
  assign n7910 = n7908 | n7909 ;
  assign n7911 = n7667 | n7670 ;
  assign n7912 = n7910 | n7911 ;
  assign n7913 = n7910 & n7911 ;
  assign n7914 = n7912 & ~n7913 ;
  assign n7915 = x83 & n3314 ;
  assign n7916 = x82 & n3309 ;
  assign n7917 = x81 & ~n3308 ;
  assign n7918 = n3570 & n7917 ;
  assign n7919 = n7916 | n7918 ;
  assign n7920 = n7915 | n7919 ;
  assign n7921 = n3317 | n7920 ;
  assign n7922 = ( n1510 & n7920 ) | ( n1510 & n7921 ) | ( n7920 & n7921 ) ;
  assign n7923 = x32 & n7922 ;
  assign n7924 = x32 & ~n7923 ;
  assign n7925 = ( n7922 & ~n7923 ) | ( n7922 & n7924 ) | ( ~n7923 & n7924 ) ;
  assign n7926 = n7914 & n7925 ;
  assign n7927 = n7914 & ~n7926 ;
  assign n7928 = ~n7914 & n7925 ;
  assign n7929 = n7927 | n7928 ;
  assign n7930 = n7684 | n7690 ;
  assign n7931 = n7929 | n7930 ;
  assign n7932 = n7929 & n7930 ;
  assign n7933 = n7931 & ~n7932 ;
  assign n7934 = x86 & n2775 ;
  assign n7935 = x85 & n2770 ;
  assign n7936 = x84 & ~n2769 ;
  assign n7937 = n2978 & n7936 ;
  assign n7938 = n7935 | n7937 ;
  assign n7939 = n7934 | n7938 ;
  assign n7940 = n2778 | n7939 ;
  assign n7941 = ( n1921 & n7939 ) | ( n1921 & n7940 ) | ( n7939 & n7940 ) ;
  assign n7942 = x29 & n7941 ;
  assign n7943 = x29 & ~n7942 ;
  assign n7944 = ( n7941 & ~n7942 ) | ( n7941 & n7943 ) | ( ~n7942 & n7943 ) ;
  assign n7945 = n7933 & n7944 ;
  assign n7946 = n7933 & ~n7945 ;
  assign n7947 = ~n7933 & n7944 ;
  assign n7948 = n7946 | n7947 ;
  assign n7949 = n7703 | n7709 ;
  assign n7950 = n7948 | n7949 ;
  assign n7951 = n7948 & n7949 ;
  assign n7952 = n7950 & ~n7951 ;
  assign n7953 = x89 & n2280 ;
  assign n7954 = x88 & n2275 ;
  assign n7955 = x87 & ~n2274 ;
  assign n7956 = n2481 & n7955 ;
  assign n7957 = n7954 | n7956 ;
  assign n7958 = n7953 | n7957 ;
  assign n7959 = n2283 | n7958 ;
  assign n7960 = ( n2244 & n7958 ) | ( n2244 & n7959 ) | ( n7958 & n7959 ) ;
  assign n7961 = x26 & n7960 ;
  assign n7962 = x26 & ~n7961 ;
  assign n7963 = ( n7960 & ~n7961 ) | ( n7960 & n7962 ) | ( ~n7961 & n7962 ) ;
  assign n7964 = n7952 & n7963 ;
  assign n7965 = n7952 & ~n7964 ;
  assign n7966 = ~n7952 & n7963 ;
  assign n7967 = n7965 | n7966 ;
  assign n7968 = n7723 | n7726 ;
  assign n7969 = n7967 & n7968 ;
  assign n7970 = n7967 | n7968 ;
  assign n7971 = ~n7969 & n7970 ;
  assign n7972 = x92 & n1817 ;
  assign n7973 = x91 & n1812 ;
  assign n7974 = x90 & ~n1811 ;
  assign n7975 = n1977 & n7974 ;
  assign n7976 = n7973 | n7975 ;
  assign n7977 = n7972 | n7976 ;
  assign n7978 = n1820 | n7977 ;
  assign n7979 = ( n2904 & n7977 ) | ( n2904 & n7978 ) | ( n7977 & n7978 ) ;
  assign n7980 = x23 & n7979 ;
  assign n7981 = x23 & ~n7980 ;
  assign n7982 = ( n7979 & ~n7980 ) | ( n7979 & n7981 ) | ( ~n7980 & n7981 ) ;
  assign n7983 = n7971 & n7982 ;
  assign n7984 = n7971 & ~n7983 ;
  assign n7985 = ~n7971 & n7982 ;
  assign n7986 = n7984 | n7985 ;
  assign n7987 = n7801 & n7986 ;
  assign n7988 = n7986 & ~n7987 ;
  assign n7989 = ( n7801 & ~n7987 ) | ( n7801 & n7988 ) | ( ~n7987 & n7988 ) ;
  assign n7990 = x95 & n1421 ;
  assign n7991 = x94 & n1416 ;
  assign n7992 = x93 & ~n1415 ;
  assign n7993 = n1584 & n7992 ;
  assign n7994 = n7991 | n7993 ;
  assign n7995 = n7990 | n7994 ;
  assign n7996 = n1424 | n7995 ;
  assign n7997 = ( n3479 & n7995 ) | ( n3479 & n7996 ) | ( n7995 & n7996 ) ;
  assign n7998 = x20 & n7997 ;
  assign n7999 = x20 & ~n7998 ;
  assign n8000 = ( n7997 & ~n7998 ) | ( n7997 & n7999 ) | ( ~n7998 & n7999 ) ;
  assign n8001 = n7989 & n8000 ;
  assign n8002 = n7989 & ~n8001 ;
  assign n8003 = n7732 | n7736 ;
  assign n8004 = ~n7989 & n8000 ;
  assign n8005 = n8003 | n8004 ;
  assign n8006 = n8002 | n8005 ;
  assign n8007 = ( n8002 & n8003 ) | ( n8002 & n8004 ) | ( n8003 & n8004 ) ;
  assign n8008 = n8006 & ~n8007 ;
  assign n8009 = x98 & n1071 ;
  assign n8010 = x97 & n1066 ;
  assign n8011 = x96 & ~n1065 ;
  assign n8012 = n1189 & n8011 ;
  assign n8013 = n8010 | n8012 ;
  assign n8014 = n8009 | n8013 ;
  assign n8015 = n1074 | n8014 ;
  assign n8016 = ( n4105 & n8014 ) | ( n4105 & n8015 ) | ( n8014 & n8015 ) ;
  assign n8017 = x17 & n8016 ;
  assign n8018 = x17 & ~n8017 ;
  assign n8019 = ( n8016 & ~n8017 ) | ( n8016 & n8018 ) | ( ~n8017 & n8018 ) ;
  assign n8020 = n8008 & n8019 ;
  assign n8021 = n8008 & ~n8020 ;
  assign n8022 = ~n8008 & n8019 ;
  assign n8023 = n8021 | n8022 ;
  assign n8024 = n7740 | n8023 ;
  assign n8025 = n7740 & n8023 ;
  assign n8026 = n8024 & ~n8025 ;
  assign n8027 = x101 & n771 ;
  assign n8028 = x100 & n766 ;
  assign n8029 = x99 & ~n765 ;
  assign n8030 = n905 & n8029 ;
  assign n8031 = n8028 | n8030 ;
  assign n8032 = n8027 | n8031 ;
  assign n8033 = n774 | n8032 ;
  assign n8034 = ( n4783 & n8032 ) | ( n4783 & n8033 ) | ( n8032 & n8033 ) ;
  assign n8035 = x14 & n8034 ;
  assign n8036 = x14 & ~n8035 ;
  assign n8037 = ( n8034 & ~n8035 ) | ( n8034 & n8036 ) | ( ~n8035 & n8036 ) ;
  assign n8038 = n8026 & n8037 ;
  assign n8039 = n8026 & ~n8038 ;
  assign n8040 = ~n8026 & n8037 ;
  assign n8041 = n8039 | n8040 ;
  assign n8042 = n7743 | n7748 ;
  assign n8043 = n8041 | n8042 ;
  assign n8044 = n8041 & n8042 ;
  assign n8045 = n8043 & ~n8044 ;
  assign n8046 = x104 & n528 ;
  assign n8047 = x103 & n523 ;
  assign n8048 = x102 & ~n522 ;
  assign n8049 = n635 & n8048 ;
  assign n8050 = n8047 | n8049 ;
  assign n8051 = n8046 | n8050 ;
  assign n8052 = n531 | n8051 ;
  assign n8053 = ( n5295 & n8051 ) | ( n5295 & n8052 ) | ( n8051 & n8052 ) ;
  assign n8054 = x11 & n8053 ;
  assign n8055 = x11 & ~n8054 ;
  assign n8056 = ( n8053 & ~n8054 ) | ( n8053 & n8055 ) | ( ~n8054 & n8055 ) ;
  assign n8057 = n8045 & n8056 ;
  assign n8058 = n8045 & ~n8057 ;
  assign n8059 = ~n8045 & n8056 ;
  assign n8060 = n8058 | n8059 ;
  assign n8061 = n7761 | n7767 ;
  assign n8062 = n8060 | n8061 ;
  assign n8063 = n8060 & n8061 ;
  assign n8064 = n8062 & ~n8063 ;
  assign n8065 = x107 & n337 ;
  assign n8066 = x106 & n332 ;
  assign n8067 = x105 & ~n331 ;
  assign n8068 = n396 & n8067 ;
  assign n8069 = n8066 | n8068 ;
  assign n8070 = n8065 | n8069 ;
  assign n8071 = n340 | n8070 ;
  assign n8072 = ( n6328 & n8070 ) | ( n6328 & n8071 ) | ( n8070 & n8071 ) ;
  assign n8073 = x8 & n8072 ;
  assign n8074 = x8 & ~n8073 ;
  assign n8075 = ( n8072 & ~n8073 ) | ( n8072 & n8074 ) | ( ~n8073 & n8074 ) ;
  assign n8076 = n8064 & n8075 ;
  assign n8077 = n8064 & ~n8076 ;
  assign n8078 = ~n8064 & n8075 ;
  assign n8079 = n8077 | n8078 ;
  assign n8080 = ( n7534 & n7535 ) | ( n7534 & n7768 ) | ( n7535 & n7768 ) ;
  assign n8081 = n8079 | n8080 ;
  assign n8082 = n8079 & n8080 ;
  assign n8083 = n8081 & ~n8082 ;
  assign n8084 = x110 & n206 ;
  assign n8085 = x109 & n201 ;
  assign n8086 = x108 & ~n200 ;
  assign n8087 = n243 & n8086 ;
  assign n8088 = n8085 | n8087 ;
  assign n8089 = n8084 | n8088 ;
  assign n8090 = n209 | n8089 ;
  assign n8091 = ( n7189 & n8089 ) | ( n7189 & n8090 ) | ( n8089 & n8090 ) ;
  assign n8092 = x5 & n8091 ;
  assign n8093 = x5 & ~n8092 ;
  assign n8094 = ( n8091 & ~n8092 ) | ( n8091 & n8093 ) | ( ~n8092 & n8093 ) ;
  assign n8095 = n8083 & n8094 ;
  assign n8096 = n8083 & ~n8095 ;
  assign n8097 = ~n8083 & n8094 ;
  assign n8098 = n8096 | n8097 ;
  assign n8099 = n7772 | n7776 ;
  assign n8100 = n8098 | n8099 ;
  assign n8101 = n8098 & n8099 ;
  assign n8102 = n8100 & ~n8101 ;
  assign n8103 = x111 | x112 ;
  assign n8104 = x112 | x113 ;
  assign n8105 = x112 & x113 ;
  assign n8106 = n8104 & ~n8105 ;
  assign n8107 = n8103 & n8106 ;
  assign n8108 = x111 & x112 ;
  assign n8109 = n8106 & n8108 ;
  assign n8110 = ( n7786 & n8107 ) | ( n7786 & n8109 ) | ( n8107 & n8109 ) ;
  assign n8111 = ( n7786 & n8103 ) | ( n7786 & n8108 ) | ( n8103 & n8108 ) ;
  assign n8112 = n8106 | n8111 ;
  assign n8113 = ~n8110 & n8112 ;
  assign n8114 = x112 & n131 ;
  assign n8115 = x111 & ~n156 ;
  assign n8116 = ( n135 & n8114 ) | ( n135 & n8115 ) | ( n8114 & n8115 ) ;
  assign n8117 = x0 & x113 ;
  assign n8118 = ( ~n135 & n8114 ) | ( ~n135 & n8117 ) | ( n8114 & n8117 ) ;
  assign n8119 = n8116 | n8118 ;
  assign n8120 = n139 | n8119 ;
  assign n8121 = ( n8113 & n8119 ) | ( n8113 & n8120 ) | ( n8119 & n8120 ) ;
  assign n8122 = x2 & n8121 ;
  assign n8123 = x2 & ~n8122 ;
  assign n8124 = ( n8121 & ~n8122 ) | ( n8121 & n8123 ) | ( ~n8122 & n8123 ) ;
  assign n8125 = n8102 | n8124 ;
  assign n8126 = n8102 & n8124 ;
  assign n8127 = n8125 & ~n8126 ;
  assign n8128 = n7800 & n8127 ;
  assign n8129 = n7800 | n8127 ;
  assign n8130 = ~n8128 & n8129 ;
  assign n8131 = n7945 | n7951 ;
  assign n8132 = n7907 | n7913 ;
  assign n8133 = n7853 | n7859 ;
  assign n8134 = x66 & n7812 ;
  assign n8135 = x65 & n7807 ;
  assign n8136 = ~n7585 & n7811 ;
  assign n8137 = x64 & ~n7806 ;
  assign n8138 = n8136 & n8137 ;
  assign n8139 = n8135 | n8138 ;
  assign n8140 = n8134 | n8139 ;
  assign n8141 = n153 & n7815 ;
  assign n8142 = n8140 | n8141 ;
  assign n8143 = x50 | n8142 ;
  assign n8144 = ~x50 & n8143 ;
  assign n8145 = ( ~n8142 & n8143 ) | ( ~n8142 & n8144 ) | ( n8143 & n8144 ) ;
  assign n8146 = n7822 | n8145 ;
  assign n8147 = n7822 & n8145 ;
  assign n8148 = n8146 & ~n8147 ;
  assign n8149 = n264 & n6940 ;
  assign n8150 = x69 & n6937 ;
  assign n8151 = x68 & n6932 ;
  assign n8152 = x67 & ~n6931 ;
  assign n8153 = n7216 & n8152 ;
  assign n8154 = n8151 | n8153 ;
  assign n8155 = n8150 | n8154 ;
  assign n8156 = n8149 | n8155 ;
  assign n8157 = x47 | n8156 ;
  assign n8158 = ~x47 & n8157 ;
  assign n8159 = ( ~n8156 & n8157 ) | ( ~n8156 & n8158 ) | ( n8157 & n8158 ) ;
  assign n8160 = n8148 & n8159 ;
  assign n8161 = n8148 & ~n8160 ;
  assign n8162 = ~n8148 & n8159 ;
  assign n8163 = n8161 | n8162 ;
  assign n8164 = n7837 | n7840 ;
  assign n8165 = n8163 & n8164 ;
  assign n8166 = n8163 | n8164 ;
  assign n8167 = ~n8165 & n8166 ;
  assign n8168 = x72 & n6068 ;
  assign n8169 = x71 & n6063 ;
  assign n8170 = x70 & ~n6062 ;
  assign n8171 = n6398 & n8170 ;
  assign n8172 = n8169 | n8171 ;
  assign n8173 = n8168 | n8172 ;
  assign n8174 = ( n435 & n6071 ) | ( n435 & n8173 ) | ( n6071 & n8173 ) ;
  assign n8175 = ( x44 & ~n8173 ) | ( x44 & n8174 ) | ( ~n8173 & n8174 ) ;
  assign n8176 = ~n8174 & n8175 ;
  assign n8177 = n8173 | n8175 ;
  assign n8178 = ( ~x44 & n8176 ) | ( ~x44 & n8177 ) | ( n8176 & n8177 ) ;
  assign n8179 = ~n8167 & n8178 ;
  assign n8180 = n8167 & ~n8178 ;
  assign n8181 = n8179 | n8180 ;
  assign n8182 = n8133 & ~n8181 ;
  assign n8183 = ~n8133 & n8181 ;
  assign n8184 = x75 & n5340 ;
  assign n8185 = x74 & n5335 ;
  assign n8186 = x73 & ~n5334 ;
  assign n8187 = n5580 & n8186 ;
  assign n8188 = n8185 | n8187 ;
  assign n8189 = n8184 | n8188 ;
  assign n8190 = n5343 | n8189 ;
  assign n8191 = ( n609 & n8189 ) | ( n609 & n8190 ) | ( n8189 & n8190 ) ;
  assign n8192 = x41 & n8191 ;
  assign n8193 = x41 & ~n8192 ;
  assign n8194 = ( n8191 & ~n8192 ) | ( n8191 & n8193 ) | ( ~n8192 & n8193 ) ;
  assign n8195 = n8183 | n8194 ;
  assign n8196 = n8182 | n8195 ;
  assign n8197 = ( n8182 & n8183 ) | ( n8182 & n8194 ) | ( n8183 & n8194 ) ;
  assign n8198 = n8196 & ~n8197 ;
  assign n8199 = n7873 | n7874 ;
  assign n8200 = n8198 & n8199 ;
  assign n8201 = n8198 | n8199 ;
  assign n8202 = ~n8200 & n8201 ;
  assign n8203 = x78 & n4572 ;
  assign n8204 = x77 & n4567 ;
  assign n8205 = x76 & ~n4566 ;
  assign n8206 = n4828 & n8205 ;
  assign n8207 = n8204 | n8206 ;
  assign n8208 = n8203 | n8207 ;
  assign n8209 = n4575 | n8208 ;
  assign n8210 = ( n868 & n8208 ) | ( n868 & n8209 ) | ( n8208 & n8209 ) ;
  assign n8211 = x38 & n8210 ;
  assign n8212 = x38 & ~n8211 ;
  assign n8213 = ( n8210 & ~n8211 ) | ( n8210 & n8212 ) | ( ~n8211 & n8212 ) ;
  assign n8214 = n8202 & n8213 ;
  assign n8215 = n8202 & ~n8214 ;
  assign n8216 = ~n8202 & n8213 ;
  assign n8217 = n8215 | n8216 ;
  assign n8218 = n7891 | n7893 ;
  assign n8219 = n8217 & n8218 ;
  assign n8220 = n8217 | n8218 ;
  assign n8221 = ~n8219 & n8220 ;
  assign n8222 = x81 & n3913 ;
  assign n8223 = x80 & n3908 ;
  assign n8224 = x79 & ~n3907 ;
  assign n8225 = n4152 & n8224 ;
  assign n8226 = n8223 | n8225 ;
  assign n8227 = n8222 | n8226 ;
  assign n8228 = n3916 | n8227 ;
  assign n8229 = ( n1256 & n8227 ) | ( n1256 & n8228 ) | ( n8227 & n8228 ) ;
  assign n8230 = x35 & n8229 ;
  assign n8231 = x35 & ~n8230 ;
  assign n8232 = ( n8229 & ~n8230 ) | ( n8229 & n8231 ) | ( ~n8230 & n8231 ) ;
  assign n8233 = n8221 & n8232 ;
  assign n8234 = n8221 & ~n8233 ;
  assign n8235 = ~n8221 & n8232 ;
  assign n8236 = n8234 | n8235 ;
  assign n8237 = n8132 & n8236 ;
  assign n8238 = n8132 & ~n8237 ;
  assign n8239 = n8236 & ~n8237 ;
  assign n8240 = n8238 | n8239 ;
  assign n8241 = x84 & n3314 ;
  assign n8242 = x83 & n3309 ;
  assign n8243 = x82 & ~n3308 ;
  assign n8244 = n3570 & n8243 ;
  assign n8245 = n8242 | n8244 ;
  assign n8246 = n8241 | n8245 ;
  assign n8247 = n3317 | n8246 ;
  assign n8248 = ( n1537 & n8246 ) | ( n1537 & n8247 ) | ( n8246 & n8247 ) ;
  assign n8249 = x32 & n8248 ;
  assign n8250 = x32 & ~n8249 ;
  assign n8251 = ( n8248 & ~n8249 ) | ( n8248 & n8250 ) | ( ~n8249 & n8250 ) ;
  assign n8252 = n8240 & n8251 ;
  assign n8253 = n8240 & ~n8252 ;
  assign n8254 = ~n8240 & n8251 ;
  assign n8255 = n8253 | n8254 ;
  assign n8256 = n7926 | n7932 ;
  assign n8257 = n8255 | n8256 ;
  assign n8258 = n8255 & n8256 ;
  assign n8259 = n8257 & ~n8258 ;
  assign n8260 = x87 & n2775 ;
  assign n8261 = x86 & n2770 ;
  assign n8262 = x85 & ~n2769 ;
  assign n8263 = n2978 & n8262 ;
  assign n8264 = n8261 | n8263 ;
  assign n8265 = n8260 | n8264 ;
  assign n8266 = n2778 | n8265 ;
  assign n8267 = ( n2067 & n8265 ) | ( n2067 & n8266 ) | ( n8265 & n8266 ) ;
  assign n8268 = x29 & n8267 ;
  assign n8269 = x29 & ~n8268 ;
  assign n8270 = ( n8267 & ~n8268 ) | ( n8267 & n8269 ) | ( ~n8268 & n8269 ) ;
  assign n8271 = n8259 | n8270 ;
  assign n8272 = n8131 & n8271 ;
  assign n8273 = n8259 & n8270 ;
  assign n8274 = n8271 & ~n8273 ;
  assign n8275 = ~n8272 & n8274 ;
  assign n8276 = x90 & n2280 ;
  assign n8277 = x89 & n2275 ;
  assign n8278 = x88 & ~n2274 ;
  assign n8279 = n2481 & n8278 ;
  assign n8280 = n8277 | n8279 ;
  assign n8281 = n8276 | n8280 ;
  assign n8282 = n2283 | n8281 ;
  assign n8283 = ( n2410 & n8281 ) | ( n2410 & n8282 ) | ( n8281 & n8282 ) ;
  assign n8284 = x26 & n8283 ;
  assign n8285 = x26 & ~n8284 ;
  assign n8286 = ( n8283 & ~n8284 ) | ( n8283 & n8285 ) | ( ~n8284 & n8285 ) ;
  assign n8287 = n8275 | n8286 ;
  assign n8288 = n8131 & ~n8274 ;
  assign n8289 = n8287 | n8288 ;
  assign n8290 = ( n8275 & n8286 ) | ( n8275 & n8288 ) | ( n8286 & n8288 ) ;
  assign n8291 = n8289 & ~n8290 ;
  assign n8292 = n7964 | n7969 ;
  assign n8293 = n8291 & n8292 ;
  assign n8294 = n8291 | n8292 ;
  assign n8295 = ~n8293 & n8294 ;
  assign n8296 = x93 & n1817 ;
  assign n8297 = x92 & n1812 ;
  assign n8298 = x91 & ~n1811 ;
  assign n8299 = n1977 & n8298 ;
  assign n8300 = n8297 | n8299 ;
  assign n8301 = n8296 | n8300 ;
  assign n8302 = n1820 | n8301 ;
  assign n8303 = ( n2931 & n8301 ) | ( n2931 & n8302 ) | ( n8301 & n8302 ) ;
  assign n8304 = x23 & n8303 ;
  assign n8305 = x23 & ~n8304 ;
  assign n8306 = ( n8303 & ~n8304 ) | ( n8303 & n8305 ) | ( ~n8304 & n8305 ) ;
  assign n8307 = n8295 | n8306 ;
  assign n8308 = n8295 & n8306 ;
  assign n8309 = n8307 & ~n8308 ;
  assign n8310 = n7983 | n8309 ;
  assign n8311 = n7987 | n8310 ;
  assign n8312 = ( n7983 & n7987 ) | ( n7983 & n8309 ) | ( n7987 & n8309 ) ;
  assign n8313 = n8311 & ~n8312 ;
  assign n8314 = x96 & n1421 ;
  assign n8315 = x95 & n1416 ;
  assign n8316 = x94 & ~n1415 ;
  assign n8317 = n1584 & n8316 ;
  assign n8318 = n8315 | n8317 ;
  assign n8319 = n8314 | n8318 ;
  assign n8320 = n1424 | n8319 ;
  assign n8321 = ( n3509 & n8319 ) | ( n3509 & n8320 ) | ( n8319 & n8320 ) ;
  assign n8322 = x20 & n8321 ;
  assign n8323 = x20 & ~n8322 ;
  assign n8324 = ( n8321 & ~n8322 ) | ( n8321 & n8323 ) | ( ~n8322 & n8323 ) ;
  assign n8325 = n8313 | n8324 ;
  assign n8326 = n8313 & n8324 ;
  assign n8327 = n8325 & ~n8326 ;
  assign n8328 = n8001 | n8327 ;
  assign n8329 = n8007 | n8328 ;
  assign n8330 = ( n8001 & n8007 ) | ( n8001 & n8327 ) | ( n8007 & n8327 ) ;
  assign n8331 = n8329 & ~n8330 ;
  assign n8332 = x99 & n1071 ;
  assign n8333 = x98 & n1066 ;
  assign n8334 = x97 & ~n1065 ;
  assign n8335 = n1189 & n8334 ;
  assign n8336 = n8333 | n8335 ;
  assign n8337 = n8332 | n8336 ;
  assign n8338 = n1074 | n8337 ;
  assign n8339 = ( n4325 & n8337 ) | ( n4325 & n8338 ) | ( n8337 & n8338 ) ;
  assign n8340 = x17 & n8339 ;
  assign n8341 = x17 & ~n8340 ;
  assign n8342 = ( n8339 & ~n8340 ) | ( n8339 & n8341 ) | ( ~n8340 & n8341 ) ;
  assign n8343 = n8331 & n8342 ;
  assign n8344 = n8331 & ~n8343 ;
  assign n8345 = ~n8331 & n8342 ;
  assign n8346 = n8344 | n8345 ;
  assign n8347 = n8020 | n8025 ;
  assign n8348 = n8346 | n8347 ;
  assign n8349 = n8346 & n8347 ;
  assign n8350 = n8348 & ~n8349 ;
  assign n8351 = x102 & n771 ;
  assign n8352 = x101 & n766 ;
  assign n8353 = x100 & ~n765 ;
  assign n8354 = n905 & n8353 ;
  assign n8355 = n8352 | n8354 ;
  assign n8356 = n8351 | n8355 ;
  assign n8357 = n774 | n8356 ;
  assign n8358 = ( n5025 & n8356 ) | ( n5025 & n8357 ) | ( n8356 & n8357 ) ;
  assign n8359 = x14 & n8358 ;
  assign n8360 = x14 & ~n8359 ;
  assign n8361 = ( n8358 & ~n8359 ) | ( n8358 & n8360 ) | ( ~n8359 & n8360 ) ;
  assign n8362 = n8350 & n8361 ;
  assign n8363 = n8350 & ~n8362 ;
  assign n8364 = ~n8350 & n8361 ;
  assign n8365 = n8363 | n8364 ;
  assign n8366 = n8038 | n8044 ;
  assign n8367 = n8365 | n8366 ;
  assign n8368 = n8365 & n8366 ;
  assign n8369 = n8367 & ~n8368 ;
  assign n8370 = x105 & n528 ;
  assign n8371 = x104 & n523 ;
  assign n8372 = x103 & ~n522 ;
  assign n8373 = n635 & n8372 ;
  assign n8374 = n8371 | n8373 ;
  assign n8375 = n8370 | n8374 ;
  assign n8376 = n531 | n8375 ;
  assign n8377 = ( n5788 & n8375 ) | ( n5788 & n8376 ) | ( n8375 & n8376 ) ;
  assign n8378 = x11 & n8377 ;
  assign n8379 = x11 & ~n8378 ;
  assign n8380 = ( n8377 & ~n8378 ) | ( n8377 & n8379 ) | ( ~n8378 & n8379 ) ;
  assign n8381 = n8369 & n8380 ;
  assign n8382 = n8369 & ~n8381 ;
  assign n8383 = ~n8369 & n8380 ;
  assign n8384 = n8382 | n8383 ;
  assign n8385 = n8057 | n8063 ;
  assign n8386 = n8384 | n8385 ;
  assign n8387 = n8384 & n8385 ;
  assign n8388 = n8386 & ~n8387 ;
  assign n8389 = x108 & n337 ;
  assign n8390 = x107 & n332 ;
  assign n8391 = x106 & ~n331 ;
  assign n8392 = n396 & n8391 ;
  assign n8393 = n8390 | n8392 ;
  assign n8394 = n8389 | n8393 ;
  assign n8395 = n340 | n8394 ;
  assign n8396 = ( n6358 & n8394 ) | ( n6358 & n8395 ) | ( n8394 & n8395 ) ;
  assign n8397 = x8 & n8396 ;
  assign n8398 = x8 & ~n8397 ;
  assign n8399 = ( n8396 & ~n8397 ) | ( n8396 & n8398 ) | ( ~n8397 & n8398 ) ;
  assign n8400 = n8388 | n8399 ;
  assign n8401 = n8076 | n8082 ;
  assign n8402 = ( n8388 & n8399 ) | ( n8388 & n8401 ) | ( n8399 & n8401 ) ;
  assign n8403 = n8400 & ~n8402 ;
  assign n8404 = n8388 & n8399 ;
  assign n8405 = n8400 & ~n8404 ;
  assign n8406 = n8401 & ~n8405 ;
  assign n8407 = n8403 | n8406 ;
  assign n8408 = x111 & n206 ;
  assign n8409 = x110 & n201 ;
  assign n8410 = x109 & ~n200 ;
  assign n8411 = n243 & n8410 ;
  assign n8412 = n8409 | n8411 ;
  assign n8413 = n8408 | n8412 ;
  assign n8414 = n209 | n8413 ;
  assign n8415 = ( n7492 & n8413 ) | ( n7492 & n8414 ) | ( n8413 & n8414 ) ;
  assign n8416 = x5 & n8415 ;
  assign n8417 = x5 & ~n8416 ;
  assign n8418 = ( n8415 & ~n8416 ) | ( n8415 & n8417 ) | ( ~n8416 & n8417 ) ;
  assign n8419 = n8407 & n8418 ;
  assign n8420 = n8407 & ~n8419 ;
  assign n8421 = ~n8407 & n8418 ;
  assign n8422 = n8420 | n8421 ;
  assign n8423 = n8095 | n8101 ;
  assign n8424 = n8422 | n8423 ;
  assign n8425 = n8422 & n8423 ;
  assign n8426 = n8424 & ~n8425 ;
  assign n8427 = x113 | x114 ;
  assign n8428 = x113 & x114 ;
  assign n8429 = n8427 & ~n8428 ;
  assign n8430 = n8105 | n8107 ;
  assign n8431 = n8429 & n8430 ;
  assign n8432 = n8105 | n8109 ;
  assign n8433 = n8429 & n8432 ;
  assign n8434 = ( n7786 & n8431 ) | ( n7786 & n8433 ) | ( n8431 & n8433 ) ;
  assign n8435 = ( n7786 & n8430 ) | ( n7786 & n8432 ) | ( n8430 & n8432 ) ;
  assign n8436 = n8429 | n8435 ;
  assign n8437 = ~n8434 & n8436 ;
  assign n8438 = x113 & n131 ;
  assign n8439 = x112 & ~n156 ;
  assign n8440 = ( n135 & n8438 ) | ( n135 & n8439 ) | ( n8438 & n8439 ) ;
  assign n8441 = x0 & x114 ;
  assign n8442 = ( ~n135 & n8438 ) | ( ~n135 & n8441 ) | ( n8438 & n8441 ) ;
  assign n8443 = n8440 | n8442 ;
  assign n8444 = n139 | n8443 ;
  assign n8445 = ( n8437 & n8443 ) | ( n8437 & n8444 ) | ( n8443 & n8444 ) ;
  assign n8446 = x2 & n8445 ;
  assign n8447 = x2 & ~n8446 ;
  assign n8448 = ( n8445 & ~n8446 ) | ( n8445 & n8447 ) | ( ~n8446 & n8447 ) ;
  assign n8449 = n8426 & n8448 ;
  assign n8450 = n8426 & ~n8449 ;
  assign n8451 = ~n8426 & n8448 ;
  assign n8452 = n8450 | n8451 ;
  assign n8453 = n8126 | n8128 ;
  assign n8454 = n8452 & n8453 ;
  assign n8455 = n8452 | n8453 ;
  assign n8456 = ~n8454 & n8455 ;
  assign n8457 = x112 & n206 ;
  assign n8458 = x111 & n201 ;
  assign n8459 = x110 & ~n200 ;
  assign n8460 = n243 & n8459 ;
  assign n8461 = n8458 | n8460 ;
  assign n8462 = n8457 | n8461 ;
  assign n8463 = n209 | n8462 ;
  assign n8464 = ( n7789 & n8462 ) | ( n7789 & n8463 ) | ( n8462 & n8463 ) ;
  assign n8465 = x5 & n8464 ;
  assign n8466 = x5 & ~n8465 ;
  assign n8467 = ( n8464 & ~n8465 ) | ( n8464 & n8466 ) | ( ~n8465 & n8466 ) ;
  assign n8468 = x109 & n337 ;
  assign n8469 = x108 & n332 ;
  assign n8470 = x107 & ~n331 ;
  assign n8471 = n396 & n8470 ;
  assign n8472 = n8469 | n8471 ;
  assign n8473 = n8468 | n8472 ;
  assign n8474 = n340 | n8473 ;
  assign n8475 = ( n6884 & n8473 ) | ( n6884 & n8474 ) | ( n8473 & n8474 ) ;
  assign n8476 = x8 & n8475 ;
  assign n8477 = x8 & ~n8476 ;
  assign n8478 = ( n8475 & ~n8476 ) | ( n8475 & n8477 ) | ( ~n8476 & n8477 ) ;
  assign n8479 = n8343 | n8349 ;
  assign n8480 = x100 & n1071 ;
  assign n8481 = x99 & n1066 ;
  assign n8482 = x98 & ~n1065 ;
  assign n8483 = n1189 & n8482 ;
  assign n8484 = n8481 | n8483 ;
  assign n8485 = n8480 | n8484 ;
  assign n8486 = n1074 | n8485 ;
  assign n8487 = ( n4532 & n8485 ) | ( n4532 & n8486 ) | ( n8485 & n8486 ) ;
  assign n8488 = x17 & n8487 ;
  assign n8489 = x17 & ~n8488 ;
  assign n8490 = ( n8487 & ~n8488 ) | ( n8487 & n8489 ) | ( ~n8488 & n8489 ) ;
  assign n8491 = x97 & n1421 ;
  assign n8492 = x96 & n1416 ;
  assign n8493 = x95 & ~n1415 ;
  assign n8494 = n1584 & n8493 ;
  assign n8495 = n8492 | n8494 ;
  assign n8496 = n8491 | n8495 ;
  assign n8497 = n1424 | n8496 ;
  assign n8498 = ( n3707 & n8496 ) | ( n3707 & n8497 ) | ( n8496 & n8497 ) ;
  assign n8499 = x20 & n8498 ;
  assign n8500 = x20 & ~n8499 ;
  assign n8501 = ( n8498 & ~n8499 ) | ( n8498 & n8500 ) | ( ~n8499 & n8500 ) ;
  assign n8502 = n8326 | n8330 ;
  assign n8503 = n8308 | n8312 ;
  assign n8504 = x94 & n1817 ;
  assign n8505 = x93 & n1812 ;
  assign n8506 = x92 & ~n1811 ;
  assign n8507 = n1977 & n8506 ;
  assign n8508 = n8505 | n8507 ;
  assign n8509 = n8504 | n8508 ;
  assign n8510 = n1820 | n8509 ;
  assign n8511 = ( n3271 & n8509 ) | ( n3271 & n8510 ) | ( n8509 & n8510 ) ;
  assign n8512 = x23 & n8511 ;
  assign n8513 = x23 & ~n8512 ;
  assign n8514 = ( n8511 & ~n8512 ) | ( n8511 & n8513 ) | ( ~n8512 & n8513 ) ;
  assign n8515 = x91 & n2280 ;
  assign n8516 = x90 & n2275 ;
  assign n8517 = x89 & ~n2274 ;
  assign n8518 = n2481 & n8517 ;
  assign n8519 = n8516 | n8518 ;
  assign n8520 = n8515 | n8519 ;
  assign n8521 = n2283 | n8520 ;
  assign n8522 = ( n2714 & n8520 ) | ( n2714 & n8521 ) | ( n8520 & n8521 ) ;
  assign n8523 = x26 & n8522 ;
  assign n8524 = x26 & ~n8523 ;
  assign n8525 = ( n8522 & ~n8523 ) | ( n8522 & n8524 ) | ( ~n8523 & n8524 ) ;
  assign n8526 = n8290 | n8293 ;
  assign n8527 = n8233 | n8237 ;
  assign n8528 = n8214 | n8219 ;
  assign n8529 = n8197 | n8200 ;
  assign n8530 = x50 & ~x51 ;
  assign n8531 = ~x50 & x51 ;
  assign n8532 = n8530 | n8531 ;
  assign n8533 = x64 & n8532 ;
  assign n8534 = x67 & n7812 ;
  assign n8535 = x66 & n7807 ;
  assign n8536 = x65 & ~n7806 ;
  assign n8537 = n8136 & n8536 ;
  assign n8538 = n8535 | n8537 ;
  assign n8539 = n8534 | n8538 ;
  assign n8540 = n180 & n7815 ;
  assign n8541 = n8539 | n8540 ;
  assign n8542 = x50 & ~n8541 ;
  assign n8543 = ~x50 & n8541 ;
  assign n8544 = n8542 | n8543 ;
  assign n8545 = ( n8147 & n8533 ) | ( n8147 & n8544 ) | ( n8533 & n8544 ) ;
  assign n8546 = ( n8147 & n8544 ) | ( n8147 & ~n8545 ) | ( n8544 & ~n8545 ) ;
  assign n8547 = ( n8533 & ~n8545 ) | ( n8533 & n8546 ) | ( ~n8545 & n8546 ) ;
  assign n8548 = x70 & n6937 ;
  assign n8549 = x69 & n6932 ;
  assign n8550 = x68 & ~n6931 ;
  assign n8551 = n7216 & n8550 ;
  assign n8552 = n8549 | n8551 ;
  assign n8553 = n8548 | n8552 ;
  assign n8554 = n6940 | n8553 ;
  assign n8555 = ( n310 & n8553 ) | ( n310 & n8554 ) | ( n8553 & n8554 ) ;
  assign n8556 = x47 & ~n8555 ;
  assign n8557 = ~x47 & n8555 ;
  assign n8558 = n8556 | n8557 ;
  assign n8559 = n8547 & n8558 ;
  assign n8560 = n8547 & ~n8559 ;
  assign n8561 = ~n8547 & n8558 ;
  assign n8562 = n8560 | n8561 ;
  assign n8563 = n8160 | n8165 ;
  assign n8564 = n8562 | n8563 ;
  assign n8565 = n8562 & n8563 ;
  assign n8566 = n8564 & ~n8565 ;
  assign n8567 = x73 & n6068 ;
  assign n8568 = x72 & n6063 ;
  assign n8569 = x71 & ~n6062 ;
  assign n8570 = n6398 & n8569 ;
  assign n8571 = n8568 | n8570 ;
  assign n8572 = n8567 | n8571 ;
  assign n8573 = ( n499 & n6071 ) | ( n499 & n8572 ) | ( n6071 & n8572 ) ;
  assign n8574 = ( x44 & ~n8572 ) | ( x44 & n8573 ) | ( ~n8572 & n8573 ) ;
  assign n8575 = ~n8573 & n8574 ;
  assign n8576 = n8572 | n8574 ;
  assign n8577 = ( ~x44 & n8575 ) | ( ~x44 & n8576 ) | ( n8575 & n8576 ) ;
  assign n8578 = n8566 | n8577 ;
  assign n8579 = n8566 & n8577 ;
  assign n8580 = n8578 & ~n8579 ;
  assign n8581 = ( n8133 & n8167 ) | ( n8133 & n8178 ) | ( n8167 & n8178 ) ;
  assign n8582 = n8580 & n8581 ;
  assign n8583 = n8580 | n8581 ;
  assign n8584 = ~n8582 & n8583 ;
  assign n8585 = x76 & n5340 ;
  assign n8586 = x75 & n5335 ;
  assign n8587 = x74 & ~n5334 ;
  assign n8588 = n5580 & n8587 ;
  assign n8589 = n8586 | n8588 ;
  assign n8590 = n8585 | n8589 ;
  assign n8591 = n5343 | n8590 ;
  assign n8592 = ( n740 & n8590 ) | ( n740 & n8591 ) | ( n8590 & n8591 ) ;
  assign n8593 = x41 & n8592 ;
  assign n8594 = x41 & ~n8593 ;
  assign n8595 = ( n8592 & ~n8593 ) | ( n8592 & n8594 ) | ( ~n8593 & n8594 ) ;
  assign n8596 = n8584 & n8595 ;
  assign n8597 = n8584 & ~n8596 ;
  assign n8598 = ~n8584 & n8595 ;
  assign n8599 = n8597 | n8598 ;
  assign n8600 = n8529 & n8599 ;
  assign n8601 = n8529 | n8599 ;
  assign n8602 = ~n8600 & n8601 ;
  assign n8603 = x79 & n4572 ;
  assign n8604 = x78 & n4567 ;
  assign n8605 = x77 & ~n4566 ;
  assign n8606 = n4828 & n8605 ;
  assign n8607 = n8604 | n8606 ;
  assign n8608 = n8603 | n8607 ;
  assign n8609 = n4575 | n8608 ;
  assign n8610 = ( n961 & n8608 ) | ( n961 & n8609 ) | ( n8608 & n8609 ) ;
  assign n8611 = x38 & n8610 ;
  assign n8612 = x38 & ~n8611 ;
  assign n8613 = ( n8610 & ~n8611 ) | ( n8610 & n8612 ) | ( ~n8611 & n8612 ) ;
  assign n8614 = n8602 & n8613 ;
  assign n8615 = n8602 | n8613 ;
  assign n8616 = ~n8614 & n8615 ;
  assign n8617 = n8528 & n8616 ;
  assign n8618 = n8528 | n8616 ;
  assign n8619 = ~n8617 & n8618 ;
  assign n8620 = x82 & n3913 ;
  assign n8621 = x81 & n3908 ;
  assign n8622 = x80 & ~n3907 ;
  assign n8623 = n4152 & n8622 ;
  assign n8624 = n8621 | n8623 ;
  assign n8625 = n8620 | n8624 ;
  assign n8626 = n3916 | n8625 ;
  assign n8627 = ( n1371 & n8625 ) | ( n1371 & n8626 ) | ( n8625 & n8626 ) ;
  assign n8628 = x35 & n8627 ;
  assign n8629 = x35 & ~n8628 ;
  assign n8630 = ( n8627 & ~n8628 ) | ( n8627 & n8629 ) | ( ~n8628 & n8629 ) ;
  assign n8631 = n8619 & n8630 ;
  assign n8632 = n8619 | n8630 ;
  assign n8633 = ~n8631 & n8632 ;
  assign n8634 = n8527 & n8633 ;
  assign n8635 = n8527 | n8633 ;
  assign n8636 = ~n8634 & n8635 ;
  assign n8637 = x85 & n3314 ;
  assign n8638 = x84 & n3309 ;
  assign n8639 = x83 & ~n3308 ;
  assign n8640 = n3570 & n8639 ;
  assign n8641 = n8638 | n8640 ;
  assign n8642 = n8637 | n8641 ;
  assign n8643 = n3317 | n8642 ;
  assign n8644 = ( n1765 & n8642 ) | ( n1765 & n8643 ) | ( n8642 & n8643 ) ;
  assign n8645 = x32 & n8644 ;
  assign n8646 = x32 & ~n8645 ;
  assign n8647 = ( n8644 & ~n8645 ) | ( n8644 & n8646 ) | ( ~n8645 & n8646 ) ;
  assign n8648 = n8636 & n8647 ;
  assign n8649 = n8636 & ~n8648 ;
  assign n8650 = ~n8636 & n8647 ;
  assign n8651 = n8649 | n8650 ;
  assign n8652 = n8252 | n8258 ;
  assign n8653 = n8651 | n8652 ;
  assign n8654 = n8651 & n8652 ;
  assign n8655 = n8653 & ~n8654 ;
  assign n8656 = x88 & n2775 ;
  assign n8657 = x87 & n2770 ;
  assign n8658 = x86 & ~n2769 ;
  assign n8659 = n2978 & n8658 ;
  assign n8660 = n8657 | n8659 ;
  assign n8661 = n8656 | n8660 ;
  assign n8662 = n2778 | n8661 ;
  assign n8663 = ( n2095 & n8661 ) | ( n2095 & n8662 ) | ( n8661 & n8662 ) ;
  assign n8664 = x29 & n8663 ;
  assign n8665 = x29 & ~n8664 ;
  assign n8666 = ( n8663 & ~n8664 ) | ( n8663 & n8665 ) | ( ~n8664 & n8665 ) ;
  assign n8667 = n8655 | n8666 ;
  assign n8668 = n8655 & n8666 ;
  assign n8669 = n8667 & ~n8668 ;
  assign n8670 = n8272 | n8273 ;
  assign n8671 = n8669 & n8670 ;
  assign n8672 = n8669 | n8670 ;
  assign n8673 = ~n8671 & n8672 ;
  assign n8674 = ( n8525 & n8526 ) | ( n8525 & ~n8673 ) | ( n8526 & ~n8673 ) ;
  assign n8675 = ( ~n8526 & n8673 ) | ( ~n8526 & n8674 ) | ( n8673 & n8674 ) ;
  assign n8676 = ( ~n8525 & n8674 ) | ( ~n8525 & n8675 ) | ( n8674 & n8675 ) ;
  assign n8677 = n8514 & n8676 ;
  assign n8678 = n8514 | n8676 ;
  assign n8679 = ~n8677 & n8678 ;
  assign n8680 = n8503 & n8679 ;
  assign n8681 = n8503 | n8679 ;
  assign n8682 = ~n8680 & n8681 ;
  assign n8683 = ( n8501 & n8502 ) | ( n8501 & ~n8682 ) | ( n8502 & ~n8682 ) ;
  assign n8684 = ( ~n8502 & n8682 ) | ( ~n8502 & n8683 ) | ( n8682 & n8683 ) ;
  assign n8685 = ( ~n8501 & n8683 ) | ( ~n8501 & n8684 ) | ( n8683 & n8684 ) ;
  assign n8686 = n8490 & n8685 ;
  assign n8687 = n8490 | n8685 ;
  assign n8688 = ~n8686 & n8687 ;
  assign n8689 = n8479 | n8688 ;
  assign n8690 = n8479 & n8688 ;
  assign n8691 = n8689 & ~n8690 ;
  assign n8692 = x103 & n771 ;
  assign n8693 = x102 & n766 ;
  assign n8694 = x101 & ~n765 ;
  assign n8695 = n905 & n8694 ;
  assign n8696 = n8693 | n8695 ;
  assign n8697 = n8692 | n8696 ;
  assign n8698 = n774 | n8697 ;
  assign n8699 = ( n5264 & n8697 ) | ( n5264 & n8698 ) | ( n8697 & n8698 ) ;
  assign n8700 = x14 & n8699 ;
  assign n8701 = x14 & ~n8700 ;
  assign n8702 = ( n8699 & ~n8700 ) | ( n8699 & n8701 ) | ( ~n8700 & n8701 ) ;
  assign n8703 = n8691 & n8702 ;
  assign n8704 = n8691 & ~n8703 ;
  assign n8705 = ~n8691 & n8702 ;
  assign n8706 = n8704 | n8705 ;
  assign n8707 = n8362 | n8368 ;
  assign n8708 = n8706 | n8707 ;
  assign n8709 = n8706 & n8707 ;
  assign n8710 = n8708 & ~n8709 ;
  assign n8711 = x106 & n528 ;
  assign n8712 = x105 & n523 ;
  assign n8713 = x104 & ~n522 ;
  assign n8714 = n635 & n8713 ;
  assign n8715 = n8712 | n8714 ;
  assign n8716 = n8711 | n8715 ;
  assign n8717 = n531 | n8716 ;
  assign n8718 = ( n5814 & n8716 ) | ( n5814 & n8717 ) | ( n8716 & n8717 ) ;
  assign n8719 = x11 & n8718 ;
  assign n8720 = x11 & ~n8719 ;
  assign n8721 = ( n8718 & ~n8719 ) | ( n8718 & n8720 ) | ( ~n8719 & n8720 ) ;
  assign n8722 = n8710 | n8721 ;
  assign n8723 = n8710 & n8721 ;
  assign n8724 = n8722 & ~n8723 ;
  assign n8725 = n8381 | n8387 ;
  assign n8726 = n8724 & n8725 ;
  assign n8727 = n8724 | n8725 ;
  assign n8728 = ~n8726 & n8727 ;
  assign n8729 = ( n8402 & n8478 ) | ( n8402 & ~n8728 ) | ( n8478 & ~n8728 ) ;
  assign n8730 = ( ~n8402 & n8728 ) | ( ~n8402 & n8729 ) | ( n8728 & n8729 ) ;
  assign n8731 = ( ~n8478 & n8729 ) | ( ~n8478 & n8730 ) | ( n8729 & n8730 ) ;
  assign n8732 = n8467 | n8731 ;
  assign n8733 = n8467 & n8731 ;
  assign n8734 = n8732 & ~n8733 ;
  assign n8735 = n8419 | n8425 ;
  assign n8736 = n8734 & n8735 ;
  assign n8737 = n8734 | n8735 ;
  assign n8738 = ~n8736 & n8737 ;
  assign n8739 = x114 | x115 ;
  assign n8740 = x114 & x115 ;
  assign n8741 = n8739 & ~n8740 ;
  assign n8742 = n8428 | n8431 ;
  assign n8743 = n8741 & n8742 ;
  assign n8744 = n8428 | n8433 ;
  assign n8745 = n8741 & n8744 ;
  assign n8746 = ( n7786 & n8743 ) | ( n7786 & n8745 ) | ( n8743 & n8745 ) ;
  assign n8747 = ( n7786 & n8742 ) | ( n7786 & n8744 ) | ( n8742 & n8744 ) ;
  assign n8748 = n8741 | n8747 ;
  assign n8749 = ~n8746 & n8748 ;
  assign n8750 = x114 & n131 ;
  assign n8751 = x113 & ~n156 ;
  assign n8752 = ( n135 & n8750 ) | ( n135 & n8751 ) | ( n8750 & n8751 ) ;
  assign n8753 = x0 & x115 ;
  assign n8754 = ( ~n135 & n8750 ) | ( ~n135 & n8753 ) | ( n8750 & n8753 ) ;
  assign n8755 = n8752 | n8754 ;
  assign n8756 = n139 | n8755 ;
  assign n8757 = ( n8749 & n8755 ) | ( n8749 & n8756 ) | ( n8755 & n8756 ) ;
  assign n8758 = x2 & n8757 ;
  assign n8759 = x2 & ~n8758 ;
  assign n8760 = ( n8757 & ~n8758 ) | ( n8757 & n8759 ) | ( ~n8758 & n8759 ) ;
  assign n8761 = n8738 & n8760 ;
  assign n8762 = n8738 | n8760 ;
  assign n8763 = ~n8761 & n8762 ;
  assign n8764 = n8449 | n8454 ;
  assign n8765 = n8763 & n8764 ;
  assign n8766 = n8763 | n8764 ;
  assign n8767 = ~n8765 & n8766 ;
  assign n8768 = x115 | x116 ;
  assign n8769 = x115 & x116 ;
  assign n8770 = n8768 & ~n8769 ;
  assign n8771 = n8740 | n8743 ;
  assign n8772 = n8770 & n8771 ;
  assign n8773 = n8740 | n8745 ;
  assign n8774 = n8770 & n8773 ;
  assign n8775 = ( n7786 & n8772 ) | ( n7786 & n8774 ) | ( n8772 & n8774 ) ;
  assign n8776 = ( n7786 & n8771 ) | ( n7786 & n8773 ) | ( n8771 & n8773 ) ;
  assign n8777 = n8770 | n8776 ;
  assign n8778 = ~n8775 & n8777 ;
  assign n8779 = x115 & n131 ;
  assign n8780 = x114 & ~n156 ;
  assign n8781 = ( n135 & n8779 ) | ( n135 & n8780 ) | ( n8779 & n8780 ) ;
  assign n8782 = x0 & x116 ;
  assign n8783 = ( ~n135 & n8779 ) | ( ~n135 & n8782 ) | ( n8779 & n8782 ) ;
  assign n8784 = n8781 | n8783 ;
  assign n8785 = n139 | n8784 ;
  assign n8786 = ( n8778 & n8784 ) | ( n8778 & n8785 ) | ( n8784 & n8785 ) ;
  assign n8787 = x2 & n8786 ;
  assign n8788 = x2 & ~n8787 ;
  assign n8789 = ( n8786 & ~n8787 ) | ( n8786 & n8788 ) | ( ~n8787 & n8788 ) ;
  assign n8790 = x113 & n206 ;
  assign n8791 = x112 & n201 ;
  assign n8792 = x111 & ~n200 ;
  assign n8793 = n243 & n8792 ;
  assign n8794 = n8791 | n8793 ;
  assign n8795 = n8790 | n8794 ;
  assign n8796 = n209 | n8795 ;
  assign n8797 = ( n8113 & n8795 ) | ( n8113 & n8796 ) | ( n8795 & n8796 ) ;
  assign n8798 = x5 & n8797 ;
  assign n8799 = x5 & ~n8798 ;
  assign n8800 = ( n8797 & ~n8798 ) | ( n8797 & n8799 ) | ( ~n8798 & n8799 ) ;
  assign n8801 = x92 & n2280 ;
  assign n8802 = x91 & n2275 ;
  assign n8803 = x90 & ~n2274 ;
  assign n8804 = n2481 & n8803 ;
  assign n8805 = n8802 | n8804 ;
  assign n8806 = n8801 | n8805 ;
  assign n8807 = n2283 | n8806 ;
  assign n8808 = ( n2904 & n8806 ) | ( n2904 & n8807 ) | ( n8806 & n8807 ) ;
  assign n8809 = x26 & n8808 ;
  assign n8810 = x26 & ~n8809 ;
  assign n8811 = ( n8808 & ~n8809 ) | ( n8808 & n8810 ) | ( ~n8809 & n8810 ) ;
  assign n8812 = x89 & n2775 ;
  assign n8813 = x88 & n2770 ;
  assign n8814 = x87 & ~n2769 ;
  assign n8815 = n2978 & n8814 ;
  assign n8816 = n8813 | n8815 ;
  assign n8817 = n8812 | n8816 ;
  assign n8818 = n2778 | n8817 ;
  assign n8819 = ( n2244 & n8817 ) | ( n2244 & n8818 ) | ( n8817 & n8818 ) ;
  assign n8820 = x29 & n8819 ;
  assign n8821 = x29 & ~n8820 ;
  assign n8822 = ( n8819 & ~n8820 ) | ( n8819 & n8821 ) | ( ~n8820 & n8821 ) ;
  assign n8823 = n8668 | n8671 ;
  assign n8824 = n8596 | n8600 ;
  assign n8825 = n8579 | n8582 ;
  assign n8826 = ~x51 & x52 ;
  assign n8827 = x51 & ~x52 ;
  assign n8828 = n8826 | n8827 ;
  assign n8829 = ~n8532 & n8828 ;
  assign n8830 = x64 & n8829 ;
  assign n8831 = ~x52 & x53 ;
  assign n8832 = x52 & ~x53 ;
  assign n8833 = n8831 | n8832 ;
  assign n8834 = n8532 & ~n8833 ;
  assign n8835 = x65 & n8834 ;
  assign n8836 = n8830 | n8835 ;
  assign n8837 = n8532 & n8833 ;
  assign n8838 = n142 & n8837 ;
  assign n8839 = n8836 | n8838 ;
  assign n8840 = x53 | n8839 ;
  assign n8841 = ~x53 & n8840 ;
  assign n8842 = ( ~n8839 & n8840 ) | ( ~n8839 & n8841 ) | ( n8840 & n8841 ) ;
  assign n8843 = x53 & ~n8533 ;
  assign n8844 = n8842 & n8843 ;
  assign n8845 = n8842 | n8843 ;
  assign n8846 = ~n8844 & n8845 ;
  assign n8847 = n229 & n7815 ;
  assign n8848 = x68 & n7812 ;
  assign n8849 = x67 & n7807 ;
  assign n8850 = x66 & ~n7806 ;
  assign n8851 = n8136 & n8850 ;
  assign n8852 = n8849 | n8851 ;
  assign n8853 = n8848 | n8852 ;
  assign n8854 = n8847 | n8853 ;
  assign n8855 = x50 | n8854 ;
  assign n8856 = ~x50 & n8855 ;
  assign n8857 = ( ~n8854 & n8855 ) | ( ~n8854 & n8856 ) | ( n8855 & n8856 ) ;
  assign n8858 = n8846 | n8857 ;
  assign n8859 = n8846 & n8857 ;
  assign n8860 = n8858 & ~n8859 ;
  assign n8861 = n8545 | n8860 ;
  assign n8862 = n8545 & n8860 ;
  assign n8863 = n8861 & ~n8862 ;
  assign n8864 = x71 & n6937 ;
  assign n8865 = x70 & n6932 ;
  assign n8866 = x69 & ~n6931 ;
  assign n8867 = n7216 & n8866 ;
  assign n8868 = n8865 | n8867 ;
  assign n8869 = n8864 | n8868 ;
  assign n8870 = n6940 | n8869 ;
  assign n8871 = ( n376 & n8869 ) | ( n376 & n8870 ) | ( n8869 & n8870 ) ;
  assign n8872 = x47 & ~n8871 ;
  assign n8873 = ~x47 & n8871 ;
  assign n8874 = n8872 | n8873 ;
  assign n8875 = n8863 & n8874 ;
  assign n8876 = n8863 & ~n8875 ;
  assign n8877 = ~n8863 & n8874 ;
  assign n8878 = n8876 | n8877 ;
  assign n8879 = n8559 | n8565 ;
  assign n8880 = n8878 | n8879 ;
  assign n8881 = n8878 & n8879 ;
  assign n8882 = n8880 & ~n8881 ;
  assign n8883 = x74 & n6068 ;
  assign n8884 = x73 & n6063 ;
  assign n8885 = x72 & ~n6062 ;
  assign n8886 = n6398 & n8885 ;
  assign n8887 = n8884 | n8886 ;
  assign n8888 = n8883 | n8887 ;
  assign n8889 = n6071 | n8888 ;
  assign n8890 = ( n587 & n8888 ) | ( n587 & n8889 ) | ( n8888 & n8889 ) ;
  assign n8891 = x44 & n8890 ;
  assign n8892 = x44 & ~n8891 ;
  assign n8893 = ( n8890 & ~n8891 ) | ( n8890 & n8892 ) | ( ~n8891 & n8892 ) ;
  assign n8894 = n8882 | n8893 ;
  assign n8895 = n8825 & n8894 ;
  assign n8896 = n8882 & n8893 ;
  assign n8897 = n8894 & ~n8896 ;
  assign n8898 = ~n8895 & n8897 ;
  assign n8899 = x77 & n5340 ;
  assign n8900 = x76 & n5335 ;
  assign n8901 = x75 & ~n5334 ;
  assign n8902 = n5580 & n8901 ;
  assign n8903 = n8900 | n8902 ;
  assign n8904 = n8899 | n8903 ;
  assign n8905 = n5343 | n8904 ;
  assign n8906 = ( n846 & n8904 ) | ( n846 & n8905 ) | ( n8904 & n8905 ) ;
  assign n8907 = x41 & n8906 ;
  assign n8908 = x41 & ~n8907 ;
  assign n8909 = ( n8906 & ~n8907 ) | ( n8906 & n8908 ) | ( ~n8907 & n8908 ) ;
  assign n8910 = n8898 | n8909 ;
  assign n8911 = n8825 & ~n8897 ;
  assign n8912 = n8910 | n8911 ;
  assign n8913 = ( n8898 & n8909 ) | ( n8898 & n8911 ) | ( n8909 & n8911 ) ;
  assign n8914 = n8912 & ~n8913 ;
  assign n8915 = n8824 & n8914 ;
  assign n8916 = n8824 | n8914 ;
  assign n8917 = ~n8915 & n8916 ;
  assign n8918 = x80 & n4572 ;
  assign n8919 = x79 & n4567 ;
  assign n8920 = x78 & ~n4566 ;
  assign n8921 = n4828 & n8920 ;
  assign n8922 = n8919 | n8921 ;
  assign n8923 = n8918 | n8922 ;
  assign n8924 = n4575 | n8923 ;
  assign n8925 = ( n1147 & n8923 ) | ( n1147 & n8924 ) | ( n8923 & n8924 ) ;
  assign n8926 = x38 & n8925 ;
  assign n8927 = x38 & ~n8926 ;
  assign n8928 = ( n8925 & ~n8926 ) | ( n8925 & n8927 ) | ( ~n8926 & n8927 ) ;
  assign n8929 = n8917 & n8928 ;
  assign n8930 = n8917 & ~n8929 ;
  assign n8931 = ~n8917 & n8928 ;
  assign n8932 = n8930 | n8931 ;
  assign n8933 = n8614 | n8617 ;
  assign n8934 = n8932 | n8933 ;
  assign n8935 = n8932 & n8933 ;
  assign n8936 = n8934 & ~n8935 ;
  assign n8937 = x83 & n3913 ;
  assign n8938 = x82 & n3908 ;
  assign n8939 = x81 & ~n3907 ;
  assign n8940 = n4152 & n8939 ;
  assign n8941 = n8938 | n8940 ;
  assign n8942 = n8937 | n8941 ;
  assign n8943 = n3916 | n8942 ;
  assign n8944 = ( n1510 & n8942 ) | ( n1510 & n8943 ) | ( n8942 & n8943 ) ;
  assign n8945 = x35 & n8944 ;
  assign n8946 = x35 & ~n8945 ;
  assign n8947 = ( n8944 & ~n8945 ) | ( n8944 & n8946 ) | ( ~n8945 & n8946 ) ;
  assign n8948 = n8936 & n8947 ;
  assign n8949 = n8936 | n8947 ;
  assign n8950 = ~n8948 & n8949 ;
  assign n8951 = n8631 | n8634 ;
  assign n8952 = n8950 & n8951 ;
  assign n8953 = n8951 & ~n8952 ;
  assign n8954 = ( n8950 & ~n8952 ) | ( n8950 & n8953 ) | ( ~n8952 & n8953 ) ;
  assign n8955 = x86 & n3314 ;
  assign n8956 = x85 & n3309 ;
  assign n8957 = x84 & ~n3308 ;
  assign n8958 = n3570 & n8957 ;
  assign n8959 = n8956 | n8958 ;
  assign n8960 = n8955 | n8959 ;
  assign n8961 = n3317 | n8960 ;
  assign n8962 = ( n1921 & n8960 ) | ( n1921 & n8961 ) | ( n8960 & n8961 ) ;
  assign n8963 = x32 & n8962 ;
  assign n8964 = x32 & ~n8963 ;
  assign n8965 = ( n8962 & ~n8963 ) | ( n8962 & n8964 ) | ( ~n8963 & n8964 ) ;
  assign n8966 = n8954 & n8965 ;
  assign n8967 = n8954 & ~n8966 ;
  assign n8968 = ~n8954 & n8965 ;
  assign n8969 = n8967 | n8968 ;
  assign n8970 = n8648 | n8654 ;
  assign n8971 = n8969 | n8970 ;
  assign n8972 = n8969 & n8970 ;
  assign n8973 = n8971 & ~n8972 ;
  assign n8974 = ( n8822 & n8823 ) | ( n8822 & ~n8973 ) | ( n8823 & ~n8973 ) ;
  assign n8975 = ( ~n8823 & n8973 ) | ( ~n8823 & n8974 ) | ( n8973 & n8974 ) ;
  assign n8976 = ( ~n8822 & n8974 ) | ( ~n8822 & n8975 ) | ( n8974 & n8975 ) ;
  assign n8977 = n8811 & n8976 ;
  assign n8978 = n8811 | n8976 ;
  assign n8979 = ~n8977 & n8978 ;
  assign n8980 = ( n8525 & n8526 ) | ( n8525 & n8673 ) | ( n8526 & n8673 ) ;
  assign n8981 = n8979 | n8980 ;
  assign n8982 = n8979 & n8980 ;
  assign n8983 = n8981 & ~n8982 ;
  assign n8984 = x95 & n1817 ;
  assign n8985 = x94 & n1812 ;
  assign n8986 = x93 & ~n1811 ;
  assign n8987 = n1977 & n8986 ;
  assign n8988 = n8985 | n8987 ;
  assign n8989 = n8984 | n8988 ;
  assign n8990 = n1820 | n8989 ;
  assign n8991 = ( n3479 & n8989 ) | ( n3479 & n8990 ) | ( n8989 & n8990 ) ;
  assign n8992 = x23 & n8991 ;
  assign n8993 = x23 & ~n8992 ;
  assign n8994 = ( n8991 & ~n8992 ) | ( n8991 & n8993 ) | ( ~n8992 & n8993 ) ;
  assign n8995 = n8983 & n8994 ;
  assign n8996 = n8983 & ~n8995 ;
  assign n8997 = ~n8983 & n8994 ;
  assign n8998 = n8996 | n8997 ;
  assign n8999 = n8677 | n8680 ;
  assign n9000 = n8998 | n8999 ;
  assign n9001 = n8998 & n8999 ;
  assign n9002 = n9000 & ~n9001 ;
  assign n9003 = x98 & n1421 ;
  assign n9004 = x97 & n1416 ;
  assign n9005 = x96 & ~n1415 ;
  assign n9006 = n1584 & n9005 ;
  assign n9007 = n9004 | n9006 ;
  assign n9008 = n9003 | n9007 ;
  assign n9009 = n1424 | n9008 ;
  assign n9010 = ( n4105 & n9008 ) | ( n4105 & n9009 ) | ( n9008 & n9009 ) ;
  assign n9011 = x20 & n9010 ;
  assign n9012 = x20 & ~n9011 ;
  assign n9013 = ( n9010 & ~n9011 ) | ( n9010 & n9012 ) | ( ~n9011 & n9012 ) ;
  assign n9014 = n9002 & n9013 ;
  assign n9015 = n9002 & ~n9014 ;
  assign n9016 = ~n9002 & n9013 ;
  assign n9017 = n9015 | n9016 ;
  assign n9018 = ( n8501 & n8502 ) | ( n8501 & n8682 ) | ( n8502 & n8682 ) ;
  assign n9019 = n9017 | n9018 ;
  assign n9020 = n9017 & n9018 ;
  assign n9021 = n9019 & ~n9020 ;
  assign n9022 = x101 & n1071 ;
  assign n9023 = x100 & n1066 ;
  assign n9024 = x99 & ~n1065 ;
  assign n9025 = n1189 & n9024 ;
  assign n9026 = n9023 | n9025 ;
  assign n9027 = n9022 | n9026 ;
  assign n9028 = n1074 | n9027 ;
  assign n9029 = ( n4783 & n9027 ) | ( n4783 & n9028 ) | ( n9027 & n9028 ) ;
  assign n9030 = x17 & n9029 ;
  assign n9031 = x17 & ~n9030 ;
  assign n9032 = ( n9029 & ~n9030 ) | ( n9029 & n9031 ) | ( ~n9030 & n9031 ) ;
  assign n9033 = n9021 & n9032 ;
  assign n9034 = n9021 & ~n9033 ;
  assign n9035 = ~n9021 & n9032 ;
  assign n9036 = n9034 | n9035 ;
  assign n9037 = n8686 | n8690 ;
  assign n9038 = n9036 | n9037 ;
  assign n9039 = n9036 & n9037 ;
  assign n9040 = n9038 & ~n9039 ;
  assign n9041 = x104 & n771 ;
  assign n9042 = x103 & n766 ;
  assign n9043 = x102 & ~n765 ;
  assign n9044 = n905 & n9043 ;
  assign n9045 = n9042 | n9044 ;
  assign n9046 = n9041 | n9045 ;
  assign n9047 = n774 | n9046 ;
  assign n9048 = ( n5295 & n9046 ) | ( n5295 & n9047 ) | ( n9046 & n9047 ) ;
  assign n9049 = x14 & n9048 ;
  assign n9050 = x14 & ~n9049 ;
  assign n9051 = ( n9048 & ~n9049 ) | ( n9048 & n9050 ) | ( ~n9049 & n9050 ) ;
  assign n9052 = n9040 & n9051 ;
  assign n9053 = n9040 & ~n9052 ;
  assign n9054 = ~n9040 & n9051 ;
  assign n9055 = n9053 | n9054 ;
  assign n9056 = n8703 | n8709 ;
  assign n9057 = n9055 | n9056 ;
  assign n9058 = n9055 & n9056 ;
  assign n9059 = n9057 & ~n9058 ;
  assign n9060 = x107 & n528 ;
  assign n9061 = x106 & n523 ;
  assign n9062 = x105 & ~n522 ;
  assign n9063 = n635 & n9062 ;
  assign n9064 = n9061 | n9063 ;
  assign n9065 = n9060 | n9064 ;
  assign n9066 = n531 | n9065 ;
  assign n9067 = ( n6328 & n9065 ) | ( n6328 & n9066 ) | ( n9065 & n9066 ) ;
  assign n9068 = x11 & n9067 ;
  assign n9069 = x11 & ~n9068 ;
  assign n9070 = ( n9067 & ~n9068 ) | ( n9067 & n9069 ) | ( ~n9068 & n9069 ) ;
  assign n9071 = n9059 & n9070 ;
  assign n9072 = n9059 | n9070 ;
  assign n9073 = ~n9071 & n9072 ;
  assign n9074 = n8723 | n8726 ;
  assign n9075 = n9073 & n9074 ;
  assign n9076 = n9074 & ~n9075 ;
  assign n9077 = ( n9073 & ~n9075 ) | ( n9073 & n9076 ) | ( ~n9075 & n9076 ) ;
  assign n9078 = x110 & n337 ;
  assign n9079 = x109 & n332 ;
  assign n9080 = x108 & ~n331 ;
  assign n9081 = n396 & n9080 ;
  assign n9082 = n9079 | n9081 ;
  assign n9083 = n9078 | n9082 ;
  assign n9084 = n340 | n9083 ;
  assign n9085 = ( n7189 & n9083 ) | ( n7189 & n9084 ) | ( n9083 & n9084 ) ;
  assign n9086 = x8 & n9085 ;
  assign n9087 = x8 & ~n9086 ;
  assign n9088 = ( n9085 & ~n9086 ) | ( n9085 & n9087 ) | ( ~n9086 & n9087 ) ;
  assign n9089 = n9077 & n9088 ;
  assign n9090 = n9077 & ~n9089 ;
  assign n9091 = ~n9077 & n9088 ;
  assign n9092 = n9090 | n9091 ;
  assign n9093 = ( n8402 & n8478 ) | ( n8402 & n8728 ) | ( n8478 & n8728 ) ;
  assign n9094 = n9092 | n9093 ;
  assign n9095 = n9092 & n9093 ;
  assign n9096 = n9094 & ~n9095 ;
  assign n9097 = n8733 | n8736 ;
  assign n9098 = ( n8800 & n9096 ) | ( n8800 & n9097 ) | ( n9096 & n9097 ) ;
  assign n9099 = ( n9096 & n9097 ) | ( n9096 & ~n9098 ) | ( n9097 & ~n9098 ) ;
  assign n9100 = ( n8800 & ~n9098 ) | ( n8800 & n9099 ) | ( ~n9098 & n9099 ) ;
  assign n9101 = n8789 & n9100 ;
  assign n9102 = n8789 | n9100 ;
  assign n9103 = ~n9101 & n9102 ;
  assign n9104 = n8761 | n8765 ;
  assign n9105 = n9103 & n9104 ;
  assign n9106 = n9103 | n9104 ;
  assign n9107 = ~n9105 & n9106 ;
  assign n9108 = x116 | x117 ;
  assign n9109 = x116 & x117 ;
  assign n9110 = n9108 & ~n9109 ;
  assign n9111 = n8769 | n8772 ;
  assign n9112 = n9110 & n9111 ;
  assign n9113 = n8769 | n8774 ;
  assign n9114 = n9110 & n9113 ;
  assign n9115 = ( n7786 & n9112 ) | ( n7786 & n9114 ) | ( n9112 & n9114 ) ;
  assign n9116 = ( n7786 & n9111 ) | ( n7786 & n9113 ) | ( n9111 & n9113 ) ;
  assign n9117 = n9110 | n9116 ;
  assign n9118 = ~n9115 & n9117 ;
  assign n9119 = x116 & n131 ;
  assign n9120 = x115 & ~n156 ;
  assign n9121 = ( n135 & n9119 ) | ( n135 & n9120 ) | ( n9119 & n9120 ) ;
  assign n9122 = x0 & x117 ;
  assign n9123 = ( ~n135 & n9119 ) | ( ~n135 & n9122 ) | ( n9119 & n9122 ) ;
  assign n9124 = n9121 | n9123 ;
  assign n9125 = n139 | n9124 ;
  assign n9126 = ( n9118 & n9124 ) | ( n9118 & n9125 ) | ( n9124 & n9125 ) ;
  assign n9127 = x2 & n9126 ;
  assign n9128 = x2 & ~n9127 ;
  assign n9129 = ( n9126 & ~n9127 ) | ( n9126 & n9128 ) | ( ~n9127 & n9128 ) ;
  assign n9130 = n9101 | n9105 ;
  assign n9131 = n8966 | n8972 ;
  assign n9132 = n8948 | n8952 ;
  assign n9133 = n8929 | n8935 ;
  assign n9134 = n8875 | n8881 ;
  assign n9135 = x72 & n6937 ;
  assign n9136 = x71 & n6932 ;
  assign n9137 = x70 & ~n6931 ;
  assign n9138 = n7216 & n9137 ;
  assign n9139 = n9136 | n9138 ;
  assign n9140 = n9135 | n9139 ;
  assign n9141 = ( n435 & n6940 ) | ( n435 & n9140 ) | ( n6940 & n9140 ) ;
  assign n9142 = ( x47 & ~n9140 ) | ( x47 & n9141 ) | ( ~n9140 & n9141 ) ;
  assign n9143 = ~n9141 & n9142 ;
  assign n9144 = n9140 | n9142 ;
  assign n9145 = ( ~x47 & n9143 ) | ( ~x47 & n9144 ) | ( n9143 & n9144 ) ;
  assign n9146 = n264 & n7815 ;
  assign n9147 = x69 & n7812 ;
  assign n9148 = x68 & n7807 ;
  assign n9149 = x67 & ~n7806 ;
  assign n9150 = n8136 & n9149 ;
  assign n9151 = n9148 | n9150 ;
  assign n9152 = n9147 | n9151 ;
  assign n9153 = n9146 | n9152 ;
  assign n9154 = x50 | n9153 ;
  assign n9155 = ~x50 & n9154 ;
  assign n9156 = ( ~n9153 & n9154 ) | ( ~n9153 & n9155 ) | ( n9154 & n9155 ) ;
  assign n9157 = x66 & n8834 ;
  assign n9158 = x65 & n8829 ;
  assign n9159 = ~n8532 & n8833 ;
  assign n9160 = x64 & ~n8828 ;
  assign n9161 = n9159 & n9160 ;
  assign n9162 = n9158 | n9161 ;
  assign n9163 = n9157 | n9162 ;
  assign n9164 = n153 & n8837 ;
  assign n9165 = n9163 | n9164 ;
  assign n9166 = x53 | n9165 ;
  assign n9167 = ~x53 & n9166 ;
  assign n9168 = ( ~n9165 & n9166 ) | ( ~n9165 & n9167 ) | ( n9166 & n9167 ) ;
  assign n9169 = n8844 | n9168 ;
  assign n9170 = n8844 & n9168 ;
  assign n9171 = n9169 & ~n9170 ;
  assign n9172 = n8859 | n8862 ;
  assign n9173 = ( n9156 & n9171 ) | ( n9156 & n9172 ) | ( n9171 & n9172 ) ;
  assign n9174 = ( n9171 & n9172 ) | ( n9171 & ~n9173 ) | ( n9172 & ~n9173 ) ;
  assign n9175 = ( n9156 & ~n9173 ) | ( n9156 & n9174 ) | ( ~n9173 & n9174 ) ;
  assign n9176 = n9145 | n9175 ;
  assign n9177 = n9145 & n9175 ;
  assign n9178 = n9176 & ~n9177 ;
  assign n9179 = n9134 & n9178 ;
  assign n9180 = n9134 | n9178 ;
  assign n9181 = ~n9179 & n9180 ;
  assign n9182 = x75 & n6068 ;
  assign n9183 = x74 & n6063 ;
  assign n9184 = x73 & ~n6062 ;
  assign n9185 = n6398 & n9184 ;
  assign n9186 = n9183 | n9185 ;
  assign n9187 = n9182 | n9186 ;
  assign n9188 = n6071 | n9187 ;
  assign n9189 = ( n609 & n9187 ) | ( n609 & n9188 ) | ( n9187 & n9188 ) ;
  assign n9190 = x44 & n9189 ;
  assign n9191 = x44 & ~n9190 ;
  assign n9192 = ( n9189 & ~n9190 ) | ( n9189 & n9191 ) | ( ~n9190 & n9191 ) ;
  assign n9193 = n9181 | n9192 ;
  assign n9194 = n9181 & n9192 ;
  assign n9195 = n9193 & ~n9194 ;
  assign n9196 = n8895 | n8896 ;
  assign n9197 = n9195 & n9196 ;
  assign n9198 = n9195 | n9196 ;
  assign n9199 = ~n9197 & n9198 ;
  assign n9200 = x78 & n5340 ;
  assign n9201 = x77 & n5335 ;
  assign n9202 = x76 & ~n5334 ;
  assign n9203 = n5580 & n9202 ;
  assign n9204 = n9201 | n9203 ;
  assign n9205 = n9200 | n9204 ;
  assign n9206 = n5343 | n9205 ;
  assign n9207 = ( n868 & n9205 ) | ( n868 & n9206 ) | ( n9205 & n9206 ) ;
  assign n9208 = x41 & n9207 ;
  assign n9209 = x41 & ~n9208 ;
  assign n9210 = ( n9207 & ~n9208 ) | ( n9207 & n9209 ) | ( ~n9208 & n9209 ) ;
  assign n9211 = n9199 & n9210 ;
  assign n9212 = n9199 & ~n9211 ;
  assign n9213 = ~n9199 & n9210 ;
  assign n9214 = n9212 | n9213 ;
  assign n9215 = n8913 | n8915 ;
  assign n9216 = n9214 & n9215 ;
  assign n9217 = n9214 | n9215 ;
  assign n9218 = ~n9216 & n9217 ;
  assign n9219 = x81 & n4572 ;
  assign n9220 = x80 & n4567 ;
  assign n9221 = x79 & ~n4566 ;
  assign n9222 = n4828 & n9221 ;
  assign n9223 = n9220 | n9222 ;
  assign n9224 = n9219 | n9223 ;
  assign n9225 = n4575 | n9224 ;
  assign n9226 = ( n1256 & n9224 ) | ( n1256 & n9225 ) | ( n9224 & n9225 ) ;
  assign n9227 = x38 & n9226 ;
  assign n9228 = x38 & ~n9227 ;
  assign n9229 = ( n9226 & ~n9227 ) | ( n9226 & n9228 ) | ( ~n9227 & n9228 ) ;
  assign n9230 = n9218 & n9229 ;
  assign n9231 = n9218 & ~n9230 ;
  assign n9232 = ~n9218 & n9229 ;
  assign n9233 = n9231 | n9232 ;
  assign n9234 = n9133 & n9233 ;
  assign n9235 = n9133 & ~n9234 ;
  assign n9236 = n9233 & ~n9234 ;
  assign n9237 = n9235 | n9236 ;
  assign n9238 = x84 & n3913 ;
  assign n9239 = x83 & n3908 ;
  assign n9240 = x82 & ~n3907 ;
  assign n9241 = n4152 & n9240 ;
  assign n9242 = n9239 | n9241 ;
  assign n9243 = n9238 | n9242 ;
  assign n9244 = n3916 | n9243 ;
  assign n9245 = ( n1537 & n9243 ) | ( n1537 & n9244 ) | ( n9243 & n9244 ) ;
  assign n9246 = x35 & n9245 ;
  assign n9247 = x35 & ~n9246 ;
  assign n9248 = ( n9245 & ~n9246 ) | ( n9245 & n9247 ) | ( ~n9246 & n9247 ) ;
  assign n9249 = n9237 & n9248 ;
  assign n9250 = n9237 & ~n9249 ;
  assign n9251 = ~n9237 & n9248 ;
  assign n9252 = n9250 | n9251 ;
  assign n9253 = n9132 & n9252 ;
  assign n9254 = n9132 | n9252 ;
  assign n9255 = ~n9253 & n9254 ;
  assign n9256 = x87 & n3314 ;
  assign n9257 = x86 & n3309 ;
  assign n9258 = x85 & ~n3308 ;
  assign n9259 = n3570 & n9258 ;
  assign n9260 = n9257 | n9259 ;
  assign n9261 = n9256 | n9260 ;
  assign n9262 = n3317 | n9261 ;
  assign n9263 = ( n2067 & n9261 ) | ( n2067 & n9262 ) | ( n9261 & n9262 ) ;
  assign n9264 = x32 & n9263 ;
  assign n9265 = x32 & ~n9264 ;
  assign n9266 = ( n9263 & ~n9264 ) | ( n9263 & n9265 ) | ( ~n9264 & n9265 ) ;
  assign n9267 = n9255 & n9266 ;
  assign n9268 = n9255 & ~n9267 ;
  assign n9269 = ~n9255 & n9266 ;
  assign n9270 = n9268 | n9269 ;
  assign n9271 = n9131 & n9270 ;
  assign n9272 = n9131 & ~n9271 ;
  assign n9273 = n9270 & ~n9271 ;
  assign n9274 = n9272 | n9273 ;
  assign n9275 = x90 & n2775 ;
  assign n9276 = x89 & n2770 ;
  assign n9277 = x88 & ~n2769 ;
  assign n9278 = n2978 & n9277 ;
  assign n9279 = n9276 | n9278 ;
  assign n9280 = n9275 | n9279 ;
  assign n9281 = n2778 | n9280 ;
  assign n9282 = ( n2410 & n9280 ) | ( n2410 & n9281 ) | ( n9280 & n9281 ) ;
  assign n9283 = x29 & n9282 ;
  assign n9284 = x29 & ~n9283 ;
  assign n9285 = ( n9282 & ~n9283 ) | ( n9282 & n9284 ) | ( ~n9283 & n9284 ) ;
  assign n9286 = n9274 | n9285 ;
  assign n9287 = n9274 & n9285 ;
  assign n9288 = n9286 & ~n9287 ;
  assign n9289 = ( n8822 & n8823 ) | ( n8822 & n8973 ) | ( n8823 & n8973 ) ;
  assign n9290 = n9288 | n9289 ;
  assign n9291 = n9288 & n9289 ;
  assign n9292 = n9290 & ~n9291 ;
  assign n9293 = x93 & n2280 ;
  assign n9294 = x92 & n2275 ;
  assign n9295 = x91 & ~n2274 ;
  assign n9296 = n2481 & n9295 ;
  assign n9297 = n9294 | n9296 ;
  assign n9298 = n9293 | n9297 ;
  assign n9299 = n2283 | n9298 ;
  assign n9300 = ( n2931 & n9298 ) | ( n2931 & n9299 ) | ( n9298 & n9299 ) ;
  assign n9301 = x26 & n9300 ;
  assign n9302 = x26 & ~n9301 ;
  assign n9303 = ( n9300 & ~n9301 ) | ( n9300 & n9302 ) | ( ~n9301 & n9302 ) ;
  assign n9304 = n9292 | n9303 ;
  assign n9305 = n9292 & n9303 ;
  assign n9306 = n9304 & ~n9305 ;
  assign n9307 = n8977 | n8982 ;
  assign n9308 = n9306 & n9307 ;
  assign n9309 = n9306 | n9307 ;
  assign n9310 = ~n9308 & n9309 ;
  assign n9311 = x96 & n1817 ;
  assign n9312 = x95 & n1812 ;
  assign n9313 = x94 & ~n1811 ;
  assign n9314 = n1977 & n9313 ;
  assign n9315 = n9312 | n9314 ;
  assign n9316 = n9311 | n9315 ;
  assign n9317 = n1820 | n9316 ;
  assign n9318 = ( n3509 & n9316 ) | ( n3509 & n9317 ) | ( n9316 & n9317 ) ;
  assign n9319 = x23 & n9318 ;
  assign n9320 = x23 & ~n9319 ;
  assign n9321 = ( n9318 & ~n9319 ) | ( n9318 & n9320 ) | ( ~n9319 & n9320 ) ;
  assign n9322 = n9310 | n9321 ;
  assign n9323 = n9310 & n9321 ;
  assign n9324 = n9322 & ~n9323 ;
  assign n9325 = n8995 | n9001 ;
  assign n9326 = n9324 & n9325 ;
  assign n9327 = n9324 | n9325 ;
  assign n9328 = ~n9326 & n9327 ;
  assign n9329 = x99 & n1421 ;
  assign n9330 = x98 & n1416 ;
  assign n9331 = x97 & ~n1415 ;
  assign n9332 = n1584 & n9331 ;
  assign n9333 = n9330 | n9332 ;
  assign n9334 = n9329 | n9333 ;
  assign n9335 = n1424 | n9334 ;
  assign n9336 = ( n4325 & n9334 ) | ( n4325 & n9335 ) | ( n9334 & n9335 ) ;
  assign n9337 = x20 & n9336 ;
  assign n9338 = x20 & ~n9337 ;
  assign n9339 = ( n9336 & ~n9337 ) | ( n9336 & n9338 ) | ( ~n9337 & n9338 ) ;
  assign n9340 = n9328 & n9339 ;
  assign n9341 = n9328 & ~n9340 ;
  assign n9342 = ~n9328 & n9339 ;
  assign n9343 = n9341 | n9342 ;
  assign n9344 = n9014 | n9020 ;
  assign n9345 = n9343 | n9344 ;
  assign n9346 = n9343 & n9344 ;
  assign n9347 = n9345 & ~n9346 ;
  assign n9348 = x102 & n1071 ;
  assign n9349 = x101 & n1066 ;
  assign n9350 = x100 & ~n1065 ;
  assign n9351 = n1189 & n9350 ;
  assign n9352 = n9349 | n9351 ;
  assign n9353 = n9348 | n9352 ;
  assign n9354 = n1074 | n9353 ;
  assign n9355 = ( n5025 & n9353 ) | ( n5025 & n9354 ) | ( n9353 & n9354 ) ;
  assign n9356 = x17 & n9355 ;
  assign n9357 = x17 & ~n9356 ;
  assign n9358 = ( n9355 & ~n9356 ) | ( n9355 & n9357 ) | ( ~n9356 & n9357 ) ;
  assign n9359 = n9347 & n9358 ;
  assign n9360 = n9347 & ~n9359 ;
  assign n9361 = ~n9347 & n9358 ;
  assign n9362 = n9360 | n9361 ;
  assign n9363 = n9033 | n9039 ;
  assign n9364 = n9362 | n9363 ;
  assign n9365 = n9362 & n9363 ;
  assign n9366 = n9364 & ~n9365 ;
  assign n9367 = x105 & n771 ;
  assign n9368 = x104 & n766 ;
  assign n9369 = x103 & ~n765 ;
  assign n9370 = n905 & n9369 ;
  assign n9371 = n9368 | n9370 ;
  assign n9372 = n9367 | n9371 ;
  assign n9373 = n774 | n9372 ;
  assign n9374 = ( n5788 & n9372 ) | ( n5788 & n9373 ) | ( n9372 & n9373 ) ;
  assign n9375 = x14 & n9374 ;
  assign n9376 = x14 & ~n9375 ;
  assign n9377 = ( n9374 & ~n9375 ) | ( n9374 & n9376 ) | ( ~n9375 & n9376 ) ;
  assign n9378 = n9366 & n9377 ;
  assign n9379 = n9366 & ~n9378 ;
  assign n9380 = ~n9366 & n9377 ;
  assign n9381 = n9379 | n9380 ;
  assign n9382 = n9052 | n9058 ;
  assign n9383 = n9381 | n9382 ;
  assign n9384 = n9381 & n9382 ;
  assign n9385 = n9383 & ~n9384 ;
  assign n9386 = x108 & n528 ;
  assign n9387 = x107 & n523 ;
  assign n9388 = x106 & ~n522 ;
  assign n9389 = n635 & n9388 ;
  assign n9390 = n9387 | n9389 ;
  assign n9391 = n9386 | n9390 ;
  assign n9392 = n531 | n9391 ;
  assign n9393 = ( n6358 & n9391 ) | ( n6358 & n9392 ) | ( n9391 & n9392 ) ;
  assign n9394 = x11 & n9393 ;
  assign n9395 = x11 & ~n9394 ;
  assign n9396 = ( n9393 & ~n9394 ) | ( n9393 & n9395 ) | ( ~n9394 & n9395 ) ;
  assign n9397 = n9385 & n9396 ;
  assign n9398 = n9385 | n9396 ;
  assign n9399 = ~n9397 & n9398 ;
  assign n9400 = n9071 | n9075 ;
  assign n9401 = n9399 & n9400 ;
  assign n9402 = n9400 & ~n9401 ;
  assign n9403 = ( n9399 & ~n9401 ) | ( n9399 & n9402 ) | ( ~n9401 & n9402 ) ;
  assign n9404 = x111 & n337 ;
  assign n9405 = x110 & n332 ;
  assign n9406 = x109 & ~n331 ;
  assign n9407 = n396 & n9406 ;
  assign n9408 = n9405 | n9407 ;
  assign n9409 = n9404 | n9408 ;
  assign n9410 = n340 | n9409 ;
  assign n9411 = ( n7492 & n9409 ) | ( n7492 & n9410 ) | ( n9409 & n9410 ) ;
  assign n9412 = x8 & n9411 ;
  assign n9413 = x8 & ~n9412 ;
  assign n9414 = ( n9411 & ~n9412 ) | ( n9411 & n9413 ) | ( ~n9412 & n9413 ) ;
  assign n9415 = n9403 & n9414 ;
  assign n9416 = n9403 & ~n9415 ;
  assign n9417 = ~n9403 & n9414 ;
  assign n9418 = n9416 | n9417 ;
  assign n9419 = n9089 | n9095 ;
  assign n9420 = n9418 | n9419 ;
  assign n9421 = n9418 & n9419 ;
  assign n9422 = n9420 & ~n9421 ;
  assign n9423 = x114 & n206 ;
  assign n9424 = x113 & n201 ;
  assign n9425 = x112 & ~n200 ;
  assign n9426 = n243 & n9425 ;
  assign n9427 = n9424 | n9426 ;
  assign n9428 = n9423 | n9427 ;
  assign n9429 = n209 | n9428 ;
  assign n9430 = ( n8437 & n9428 ) | ( n8437 & n9429 ) | ( n9428 & n9429 ) ;
  assign n9431 = x5 & n9430 ;
  assign n9432 = x5 & ~n9431 ;
  assign n9433 = ( n9430 & ~n9431 ) | ( n9430 & n9432 ) | ( ~n9431 & n9432 ) ;
  assign n9434 = n9422 & n9433 ;
  assign n9435 = n9422 | n9433 ;
  assign n9436 = ~n9434 & n9435 ;
  assign n9437 = n9098 & n9436 ;
  assign n9438 = n9098 & ~n9437 ;
  assign n9439 = ( n9436 & ~n9437 ) | ( n9436 & n9438 ) | ( ~n9437 & n9438 ) ;
  assign n9440 = ( n9129 & n9130 ) | ( n9129 & ~n9439 ) | ( n9130 & ~n9439 ) ;
  assign n9441 = ( ~n9130 & n9439 ) | ( ~n9130 & n9440 ) | ( n9439 & n9440 ) ;
  assign n9442 = ( ~n9129 & n9440 ) | ( ~n9129 & n9441 ) | ( n9440 & n9441 ) ;
  assign n9443 = n9434 | n9437 ;
  assign n9444 = n9397 | n9401 ;
  assign n9445 = x100 & n1421 ;
  assign n9446 = x99 & n1416 ;
  assign n9447 = x98 & ~n1415 ;
  assign n9448 = n1584 & n9447 ;
  assign n9449 = n9446 | n9448 ;
  assign n9450 = n9445 | n9449 ;
  assign n9451 = n1424 | n9450 ;
  assign n9452 = ( n4532 & n9450 ) | ( n4532 & n9451 ) | ( n9450 & n9451 ) ;
  assign n9453 = x20 & n9452 ;
  assign n9454 = x20 & ~n9453 ;
  assign n9455 = ( n9452 & ~n9453 ) | ( n9452 & n9454 ) | ( ~n9453 & n9454 ) ;
  assign n9456 = x97 & n1817 ;
  assign n9457 = x96 & n1812 ;
  assign n9458 = x95 & ~n1811 ;
  assign n9459 = n1977 & n9458 ;
  assign n9460 = n9457 | n9459 ;
  assign n9461 = n9456 | n9460 ;
  assign n9462 = n1820 | n9461 ;
  assign n9463 = ( n3707 & n9461 ) | ( n3707 & n9462 ) | ( n9461 & n9462 ) ;
  assign n9464 = x23 & n9463 ;
  assign n9465 = x23 & ~n9464 ;
  assign n9466 = ( n9463 & ~n9464 ) | ( n9463 & n9465 ) | ( ~n9464 & n9465 ) ;
  assign n9467 = n9305 | n9308 ;
  assign n9468 = n9230 | n9234 ;
  assign n9469 = n9211 | n9216 ;
  assign n9470 = n9194 | n9197 ;
  assign n9471 = n9177 | n9179 ;
  assign n9472 = x73 & n6937 ;
  assign n9473 = x72 & n6932 ;
  assign n9474 = x71 & ~n6931 ;
  assign n9475 = n7216 & n9474 ;
  assign n9476 = n9473 | n9475 ;
  assign n9477 = n9472 | n9476 ;
  assign n9478 = ( n499 & n6940 ) | ( n499 & n9477 ) | ( n6940 & n9477 ) ;
  assign n9479 = ( x47 & ~n9477 ) | ( x47 & n9478 ) | ( ~n9477 & n9478 ) ;
  assign n9480 = ~n9478 & n9479 ;
  assign n9481 = n9477 | n9479 ;
  assign n9482 = ( ~x47 & n9480 ) | ( ~x47 & n9481 ) | ( n9480 & n9481 ) ;
  assign n9483 = x53 & ~x54 ;
  assign n9484 = ~x53 & x54 ;
  assign n9485 = n9483 | n9484 ;
  assign n9486 = x64 & n9485 ;
  assign n9487 = x67 & n8834 ;
  assign n9488 = x66 & n8829 ;
  assign n9489 = x65 & ~n8828 ;
  assign n9490 = n9159 & n9489 ;
  assign n9491 = n9488 | n9490 ;
  assign n9492 = n9487 | n9491 ;
  assign n9493 = n180 & n8837 ;
  assign n9494 = n9492 | n9493 ;
  assign n9495 = x53 & ~n9494 ;
  assign n9496 = ~x53 & n9494 ;
  assign n9497 = n9495 | n9496 ;
  assign n9498 = ( n9170 & n9486 ) | ( n9170 & n9497 ) | ( n9486 & n9497 ) ;
  assign n9499 = ( n9170 & n9497 ) | ( n9170 & ~n9498 ) | ( n9497 & ~n9498 ) ;
  assign n9500 = ( n9486 & ~n9498 ) | ( n9486 & n9499 ) | ( ~n9498 & n9499 ) ;
  assign n9501 = x70 & n7812 ;
  assign n9502 = x69 & n7807 ;
  assign n9503 = x68 & ~n7806 ;
  assign n9504 = n8136 & n9503 ;
  assign n9505 = n9502 | n9504 ;
  assign n9506 = n9501 | n9505 ;
  assign n9507 = n7815 | n9506 ;
  assign n9508 = ( n310 & n9506 ) | ( n310 & n9507 ) | ( n9506 & n9507 ) ;
  assign n9509 = x50 & ~n9508 ;
  assign n9510 = ~x50 & n9508 ;
  assign n9511 = n9509 | n9510 ;
  assign n9512 = n9500 & n9511 ;
  assign n9513 = n9500 & ~n9512 ;
  assign n9514 = ~n9500 & n9511 ;
  assign n9515 = n9173 | n9514 ;
  assign n9516 = n9513 | n9515 ;
  assign n9517 = ( n9173 & n9513 ) | ( n9173 & n9514 ) | ( n9513 & n9514 ) ;
  assign n9518 = n9516 & ~n9517 ;
  assign n9519 = n9482 & n9518 ;
  assign n9520 = n9518 & ~n9519 ;
  assign n9521 = ( n9482 & ~n9519 ) | ( n9482 & n9520 ) | ( ~n9519 & n9520 ) ;
  assign n9522 = n9471 & n9521 ;
  assign n9523 = n9471 | n9521 ;
  assign n9524 = ~n9522 & n9523 ;
  assign n9525 = x76 & n6068 ;
  assign n9526 = x75 & n6063 ;
  assign n9527 = x74 & ~n6062 ;
  assign n9528 = n6398 & n9527 ;
  assign n9529 = n9526 | n9528 ;
  assign n9530 = n9525 | n9529 ;
  assign n9531 = n6071 | n9530 ;
  assign n9532 = ( n740 & n9530 ) | ( n740 & n9531 ) | ( n9530 & n9531 ) ;
  assign n9533 = x44 & n9532 ;
  assign n9534 = x44 & ~n9533 ;
  assign n9535 = ( n9532 & ~n9533 ) | ( n9532 & n9534 ) | ( ~n9533 & n9534 ) ;
  assign n9536 = n9524 & n9535 ;
  assign n9537 = n9524 & ~n9536 ;
  assign n9538 = ~n9524 & n9535 ;
  assign n9539 = n9537 | n9538 ;
  assign n9540 = n9470 & n9539 ;
  assign n9541 = n9470 | n9539 ;
  assign n9542 = ~n9540 & n9541 ;
  assign n9543 = x79 & n5340 ;
  assign n9544 = x78 & n5335 ;
  assign n9545 = x77 & ~n5334 ;
  assign n9546 = n5580 & n9545 ;
  assign n9547 = n9544 | n9546 ;
  assign n9548 = n9543 | n9547 ;
  assign n9549 = n5343 | n9548 ;
  assign n9550 = ( n961 & n9548 ) | ( n961 & n9549 ) | ( n9548 & n9549 ) ;
  assign n9551 = x41 & n9550 ;
  assign n9552 = x41 & ~n9551 ;
  assign n9553 = ( n9550 & ~n9551 ) | ( n9550 & n9552 ) | ( ~n9551 & n9552 ) ;
  assign n9554 = n9542 & n9553 ;
  assign n9555 = n9542 | n9553 ;
  assign n9556 = ~n9554 & n9555 ;
  assign n9557 = n9469 & n9556 ;
  assign n9558 = n9469 | n9556 ;
  assign n9559 = ~n9557 & n9558 ;
  assign n9560 = x82 & n4572 ;
  assign n9561 = x81 & n4567 ;
  assign n9562 = x80 & ~n4566 ;
  assign n9563 = n4828 & n9562 ;
  assign n9564 = n9561 | n9563 ;
  assign n9565 = n9560 | n9564 ;
  assign n9566 = n4575 | n9565 ;
  assign n9567 = ( n1371 & n9565 ) | ( n1371 & n9566 ) | ( n9565 & n9566 ) ;
  assign n9568 = x38 & n9567 ;
  assign n9569 = x38 & ~n9568 ;
  assign n9570 = ( n9567 & ~n9568 ) | ( n9567 & n9569 ) | ( ~n9568 & n9569 ) ;
  assign n9571 = n9559 & n9570 ;
  assign n9572 = n9559 & ~n9571 ;
  assign n9573 = ~n9559 & n9570 ;
  assign n9574 = n9572 | n9573 ;
  assign n9575 = n9468 & n9574 ;
  assign n9576 = n9468 | n9574 ;
  assign n9577 = ~n9575 & n9576 ;
  assign n9578 = x85 & n3913 ;
  assign n9579 = x84 & n3908 ;
  assign n9580 = x83 & ~n3907 ;
  assign n9581 = n4152 & n9580 ;
  assign n9582 = n9579 | n9581 ;
  assign n9583 = n9578 | n9582 ;
  assign n9584 = n3916 | n9583 ;
  assign n9585 = ( n1765 & n9583 ) | ( n1765 & n9584 ) | ( n9583 & n9584 ) ;
  assign n9586 = x35 & n9585 ;
  assign n9587 = x35 & ~n9586 ;
  assign n9588 = ( n9585 & ~n9586 ) | ( n9585 & n9587 ) | ( ~n9586 & n9587 ) ;
  assign n9589 = n9577 & n9588 ;
  assign n9590 = n9577 | n9588 ;
  assign n9591 = ~n9589 & n9590 ;
  assign n9592 = n9249 | n9253 ;
  assign n9593 = n9591 & n9592 ;
  assign n9594 = n9591 | n9592 ;
  assign n9595 = ~n9593 & n9594 ;
  assign n9596 = x88 & n3314 ;
  assign n9597 = x87 & n3309 ;
  assign n9598 = x86 & ~n3308 ;
  assign n9599 = n3570 & n9598 ;
  assign n9600 = n9597 | n9599 ;
  assign n9601 = n9596 | n9600 ;
  assign n9602 = n3317 | n9601 ;
  assign n9603 = ( n2095 & n9601 ) | ( n2095 & n9602 ) | ( n9601 & n9602 ) ;
  assign n9604 = x32 & n9603 ;
  assign n9605 = x32 & ~n9604 ;
  assign n9606 = ( n9603 & ~n9604 ) | ( n9603 & n9605 ) | ( ~n9604 & n9605 ) ;
  assign n9607 = n9595 & n9606 ;
  assign n9608 = n9595 | n9606 ;
  assign n9609 = ~n9607 & n9608 ;
  assign n9610 = n9267 | n9609 ;
  assign n9611 = n9271 | n9610 ;
  assign n9612 = ( n9267 & n9271 ) | ( n9267 & n9609 ) | ( n9271 & n9609 ) ;
  assign n9613 = n9611 & ~n9612 ;
  assign n9614 = x91 & n2775 ;
  assign n9615 = x90 & n2770 ;
  assign n9616 = x89 & ~n2769 ;
  assign n9617 = n2978 & n9616 ;
  assign n9618 = n9615 | n9617 ;
  assign n9619 = n9614 | n9618 ;
  assign n9620 = n2778 | n9619 ;
  assign n9621 = ( n2714 & n9619 ) | ( n2714 & n9620 ) | ( n9619 & n9620 ) ;
  assign n9622 = x29 & n9621 ;
  assign n9623 = x29 & ~n9622 ;
  assign n9624 = ( n9621 & ~n9622 ) | ( n9621 & n9623 ) | ( ~n9622 & n9623 ) ;
  assign n9625 = n9613 & n9624 ;
  assign n9626 = n9613 | n9624 ;
  assign n9627 = ~n9625 & n9626 ;
  assign n9628 = n9287 | n9627 ;
  assign n9629 = n9291 | n9628 ;
  assign n9630 = ( n9287 & n9291 ) | ( n9287 & n9627 ) | ( n9291 & n9627 ) ;
  assign n9631 = n9629 & ~n9630 ;
  assign n9632 = x94 & n2280 ;
  assign n9633 = x93 & n2275 ;
  assign n9634 = x92 & ~n2274 ;
  assign n9635 = n2481 & n9634 ;
  assign n9636 = n9633 | n9635 ;
  assign n9637 = n9632 | n9636 ;
  assign n9638 = n2283 | n9637 ;
  assign n9639 = ( n3271 & n9637 ) | ( n3271 & n9638 ) | ( n9637 & n9638 ) ;
  assign n9640 = x26 & n9639 ;
  assign n9641 = x26 & ~n9640 ;
  assign n9642 = ( n9639 & ~n9640 ) | ( n9639 & n9641 ) | ( ~n9640 & n9641 ) ;
  assign n9643 = n9631 & n9642 ;
  assign n9644 = n9631 | n9642 ;
  assign n9645 = ~n9643 & n9644 ;
  assign n9646 = n9467 & n9645 ;
  assign n9647 = n9467 | n9645 ;
  assign n9648 = ~n9646 & n9647 ;
  assign n9649 = n9323 | n9326 ;
  assign n9650 = ( n9466 & n9648 ) | ( n9466 & n9649 ) | ( n9648 & n9649 ) ;
  assign n9651 = ( n9648 & n9649 ) | ( n9648 & ~n9650 ) | ( n9649 & ~n9650 ) ;
  assign n9652 = ( n9466 & ~n9650 ) | ( n9466 & n9651 ) | ( ~n9650 & n9651 ) ;
  assign n9653 = n9455 & n9652 ;
  assign n9654 = n9455 | n9652 ;
  assign n9655 = ~n9653 & n9654 ;
  assign n9656 = n9340 | n9346 ;
  assign n9657 = n9655 | n9656 ;
  assign n9658 = n9655 & n9656 ;
  assign n9659 = n9657 & ~n9658 ;
  assign n9660 = x103 & n1071 ;
  assign n9661 = x102 & n1066 ;
  assign n9662 = x101 & ~n1065 ;
  assign n9663 = n1189 & n9662 ;
  assign n9664 = n9661 | n9663 ;
  assign n9665 = n9660 | n9664 ;
  assign n9666 = n1074 | n9665 ;
  assign n9667 = ( n5264 & n9665 ) | ( n5264 & n9666 ) | ( n9665 & n9666 ) ;
  assign n9668 = x17 & n9667 ;
  assign n9669 = x17 & ~n9668 ;
  assign n9670 = ( n9667 & ~n9668 ) | ( n9667 & n9669 ) | ( ~n9668 & n9669 ) ;
  assign n9671 = n9659 & n9670 ;
  assign n9672 = n9659 & ~n9671 ;
  assign n9673 = ~n9659 & n9670 ;
  assign n9674 = n9672 | n9673 ;
  assign n9675 = n9359 | n9365 ;
  assign n9676 = n9674 | n9675 ;
  assign n9677 = n9674 & n9675 ;
  assign n9678 = n9676 & ~n9677 ;
  assign n9679 = x106 & n771 ;
  assign n9680 = x105 & n766 ;
  assign n9681 = x104 & ~n765 ;
  assign n9682 = n905 & n9681 ;
  assign n9683 = n9680 | n9682 ;
  assign n9684 = n9679 | n9683 ;
  assign n9685 = n774 | n9684 ;
  assign n9686 = ( n5814 & n9684 ) | ( n5814 & n9685 ) | ( n9684 & n9685 ) ;
  assign n9687 = x14 & n9686 ;
  assign n9688 = x14 & ~n9687 ;
  assign n9689 = ( n9686 & ~n9687 ) | ( n9686 & n9688 ) | ( ~n9687 & n9688 ) ;
  assign n9690 = n9678 | n9689 ;
  assign n9691 = n9678 & n9689 ;
  assign n9692 = n9690 & ~n9691 ;
  assign n9693 = n9378 | n9692 ;
  assign n9694 = n9384 | n9693 ;
  assign n9695 = ( n9378 & n9384 ) | ( n9378 & n9692 ) | ( n9384 & n9692 ) ;
  assign n9696 = n9694 & ~n9695 ;
  assign n9697 = x109 & n528 ;
  assign n9698 = x108 & n523 ;
  assign n9699 = x107 & ~n522 ;
  assign n9700 = n635 & n9699 ;
  assign n9701 = n9698 | n9700 ;
  assign n9702 = n9697 | n9701 ;
  assign n9703 = n531 | n9702 ;
  assign n9704 = ( n6884 & n9702 ) | ( n6884 & n9703 ) | ( n9702 & n9703 ) ;
  assign n9705 = x11 & n9704 ;
  assign n9706 = x11 & ~n9705 ;
  assign n9707 = ( n9704 & ~n9705 ) | ( n9704 & n9706 ) | ( ~n9705 & n9706 ) ;
  assign n9708 = n9696 & n9707 ;
  assign n9709 = n9696 & ~n9708 ;
  assign n9710 = ~n9696 & n9707 ;
  assign n9711 = n9709 | n9710 ;
  assign n9712 = n9444 & n9711 ;
  assign n9713 = n9444 & ~n9712 ;
  assign n9714 = n9711 & ~n9712 ;
  assign n9715 = n9713 | n9714 ;
  assign n9716 = x112 & n337 ;
  assign n9717 = x111 & n332 ;
  assign n9718 = x110 & ~n331 ;
  assign n9719 = n396 & n9718 ;
  assign n9720 = n9717 | n9719 ;
  assign n9721 = n9716 | n9720 ;
  assign n9722 = n340 | n9721 ;
  assign n9723 = ( n7789 & n9721 ) | ( n7789 & n9722 ) | ( n9721 & n9722 ) ;
  assign n9724 = x8 & n9723 ;
  assign n9725 = x8 & ~n9724 ;
  assign n9726 = ( n9723 & ~n9724 ) | ( n9723 & n9725 ) | ( ~n9724 & n9725 ) ;
  assign n9727 = n9715 & n9726 ;
  assign n9728 = n9715 & ~n9727 ;
  assign n9729 = ~n9715 & n9726 ;
  assign n9730 = n9728 | n9729 ;
  assign n9731 = n9415 | n9421 ;
  assign n9732 = n9730 | n9731 ;
  assign n9733 = n9730 & n9731 ;
  assign n9734 = n9732 & ~n9733 ;
  assign n9735 = x115 & n206 ;
  assign n9736 = x114 & n201 ;
  assign n9737 = x113 & ~n200 ;
  assign n9738 = n243 & n9737 ;
  assign n9739 = n9736 | n9738 ;
  assign n9740 = n9735 | n9739 ;
  assign n9741 = n209 | n9740 ;
  assign n9742 = ( n8749 & n9740 ) | ( n8749 & n9741 ) | ( n9740 & n9741 ) ;
  assign n9743 = x5 & n9742 ;
  assign n9744 = x5 & ~n9743 ;
  assign n9745 = ( n9742 & ~n9743 ) | ( n9742 & n9744 ) | ( ~n9743 & n9744 ) ;
  assign n9746 = n9734 | n9745 ;
  assign n9747 = n9734 & n9745 ;
  assign n9748 = n9746 & ~n9747 ;
  assign n9749 = n9443 & n9748 ;
  assign n9750 = n9443 | n9748 ;
  assign n9751 = ~n9749 & n9750 ;
  assign n9752 = x117 | x118 ;
  assign n9753 = x117 & x118 ;
  assign n9754 = n9752 & ~n9753 ;
  assign n9755 = n9109 | n9112 ;
  assign n9756 = n9109 | n9114 ;
  assign n9757 = ( n7786 & n9755 ) | ( n7786 & n9756 ) | ( n9755 & n9756 ) ;
  assign n9758 = n9754 | n9757 ;
  assign n9759 = n9754 & n9757 ;
  assign n9760 = n9758 & ~n9759 ;
  assign n9761 = x117 & n131 ;
  assign n9762 = x116 & ~n156 ;
  assign n9763 = ( n135 & n9761 ) | ( n135 & n9762 ) | ( n9761 & n9762 ) ;
  assign n9764 = x0 & x118 ;
  assign n9765 = ( ~n135 & n9761 ) | ( ~n135 & n9764 ) | ( n9761 & n9764 ) ;
  assign n9766 = n9763 | n9765 ;
  assign n9767 = n139 | n9766 ;
  assign n9768 = ( n9760 & n9766 ) | ( n9760 & n9767 ) | ( n9766 & n9767 ) ;
  assign n9769 = x2 & n9768 ;
  assign n9770 = x2 & ~n9769 ;
  assign n9771 = ( n9768 & ~n9769 ) | ( n9768 & n9770 ) | ( ~n9769 & n9770 ) ;
  assign n9772 = n9751 & n9771 ;
  assign n9773 = n9751 | n9771 ;
  assign n9774 = ~n9772 & n9773 ;
  assign n9775 = ( n9129 & n9130 ) | ( n9129 & n9439 ) | ( n9130 & n9439 ) ;
  assign n9776 = n9774 | n9775 ;
  assign n9777 = n9774 & n9775 ;
  assign n9778 = n9776 & ~n9777 ;
  assign n9779 = x118 & n131 ;
  assign n9780 = x117 & ~n156 ;
  assign n9781 = ( n135 & n9779 ) | ( n135 & n9780 ) | ( n9779 & n9780 ) ;
  assign n9782 = x0 & x119 ;
  assign n9783 = ( ~n135 & n9779 ) | ( ~n135 & n9782 ) | ( n9779 & n9782 ) ;
  assign n9784 = n9781 | n9783 ;
  assign n9785 = n139 | n9784 ;
  assign n9786 = n9753 | n9759 ;
  assign n9787 = ( x118 & ~x119 ) | ( x118 & n9786 ) | ( ~x119 & n9786 ) ;
  assign n9788 = ( ~x118 & x119 ) | ( ~x118 & n9787 ) | ( x119 & n9787 ) ;
  assign n9789 = ( ~n9786 & n9787 ) | ( ~n9786 & n9788 ) | ( n9787 & n9788 ) ;
  assign n9790 = ( n9784 & n9785 ) | ( n9784 & n9789 ) | ( n9785 & n9789 ) ;
  assign n9791 = x2 & n9790 ;
  assign n9792 = x2 & ~n9791 ;
  assign n9793 = ( n9790 & ~n9791 ) | ( n9790 & n9792 ) | ( ~n9791 & n9792 ) ;
  assign n9794 = x116 & n206 ;
  assign n9795 = x115 & n201 ;
  assign n9796 = x114 & ~n200 ;
  assign n9797 = n243 & n9796 ;
  assign n9798 = n9795 | n9797 ;
  assign n9799 = n9794 | n9798 ;
  assign n9800 = n209 | n9799 ;
  assign n9801 = ( n8778 & n9799 ) | ( n8778 & n9800 ) | ( n9799 & n9800 ) ;
  assign n9802 = x5 & n9801 ;
  assign n9803 = x5 & ~n9802 ;
  assign n9804 = ( n9801 & ~n9802 ) | ( n9801 & n9803 ) | ( ~n9802 & n9803 ) ;
  assign n9805 = n9747 | n9749 ;
  assign n9806 = n9708 | n9712 ;
  assign n9807 = n9691 | n9695 ;
  assign n9808 = x86 & n3913 ;
  assign n9809 = x85 & n3908 ;
  assign n9810 = x84 & ~n3907 ;
  assign n9811 = n4152 & n9810 ;
  assign n9812 = n9809 | n9811 ;
  assign n9813 = n9808 | n9812 ;
  assign n9814 = n3916 | n9813 ;
  assign n9815 = ( n1921 & n9813 ) | ( n1921 & n9814 ) | ( n9813 & n9814 ) ;
  assign n9816 = x35 & n9815 ;
  assign n9817 = x35 & ~n9816 ;
  assign n9818 = ( n9815 & ~n9816 ) | ( n9815 & n9817 ) | ( ~n9816 & n9817 ) ;
  assign n9819 = x83 & n4572 ;
  assign n9820 = x82 & n4567 ;
  assign n9821 = x81 & ~n4566 ;
  assign n9822 = n4828 & n9821 ;
  assign n9823 = n9820 | n9822 ;
  assign n9824 = n9819 | n9823 ;
  assign n9825 = n4575 | n9824 ;
  assign n9826 = ( n1510 & n9824 ) | ( n1510 & n9825 ) | ( n9824 & n9825 ) ;
  assign n9827 = x38 & n9826 ;
  assign n9828 = x38 & ~n9827 ;
  assign n9829 = ( n9826 & ~n9827 ) | ( n9826 & n9828 ) | ( ~n9827 & n9828 ) ;
  assign n9830 = n9571 | n9575 ;
  assign n9831 = n9536 | n9540 ;
  assign n9832 = n9519 | n9522 ;
  assign n9833 = n9512 | n9517 ;
  assign n9834 = x71 & n7812 ;
  assign n9835 = x70 & n7807 ;
  assign n9836 = x69 & ~n7806 ;
  assign n9837 = n8136 & n9836 ;
  assign n9838 = n9835 | n9837 ;
  assign n9839 = n9834 | n9838 ;
  assign n9840 = n7815 | n9839 ;
  assign n9841 = ( n376 & n9839 ) | ( n376 & n9840 ) | ( n9839 & n9840 ) ;
  assign n9842 = x50 & ~n9841 ;
  assign n9843 = ~x50 & n9841 ;
  assign n9844 = n9842 | n9843 ;
  assign n9845 = ~x54 & x55 ;
  assign n9846 = x54 & ~x55 ;
  assign n9847 = n9845 | n9846 ;
  assign n9848 = ~n9485 & n9847 ;
  assign n9849 = x64 & n9848 ;
  assign n9850 = ~x55 & x56 ;
  assign n9851 = x55 & ~x56 ;
  assign n9852 = n9850 | n9851 ;
  assign n9853 = n9485 & ~n9852 ;
  assign n9854 = x65 & n9853 ;
  assign n9855 = n9849 | n9854 ;
  assign n9856 = n9485 & n9852 ;
  assign n9857 = n142 & n9856 ;
  assign n9858 = n9855 | n9857 ;
  assign n9859 = x56 | n9858 ;
  assign n9860 = ~x56 & n9859 ;
  assign n9861 = ( ~n9858 & n9859 ) | ( ~n9858 & n9860 ) | ( n9859 & n9860 ) ;
  assign n9862 = x56 & ~n9486 ;
  assign n9863 = n9861 & n9862 ;
  assign n9864 = n9861 | n9862 ;
  assign n9865 = ~n9863 & n9864 ;
  assign n9866 = n229 & n8837 ;
  assign n9867 = x68 & n8834 ;
  assign n9868 = x67 & n8829 ;
  assign n9869 = x66 & ~n8828 ;
  assign n9870 = n9159 & n9869 ;
  assign n9871 = n9868 | n9870 ;
  assign n9872 = n9867 | n9871 ;
  assign n9873 = n9866 | n9872 ;
  assign n9874 = x53 | n9873 ;
  assign n9875 = ~x53 & n9874 ;
  assign n9876 = ( ~n9873 & n9874 ) | ( ~n9873 & n9875 ) | ( n9874 & n9875 ) ;
  assign n9877 = n9865 | n9876 ;
  assign n9878 = n9865 & n9876 ;
  assign n9879 = n9877 & ~n9878 ;
  assign n9880 = n9498 | n9879 ;
  assign n9881 = n9498 & n9879 ;
  assign n9882 = n9880 & ~n9881 ;
  assign n9883 = n9844 | n9882 ;
  assign n9884 = n9844 & n9882 ;
  assign n9885 = n9883 & ~n9884 ;
  assign n9886 = n9833 & n9885 ;
  assign n9887 = n9833 | n9885 ;
  assign n9888 = ~n9886 & n9887 ;
  assign n9889 = x74 & n6937 ;
  assign n9890 = x73 & n6932 ;
  assign n9891 = x72 & ~n6931 ;
  assign n9892 = n7216 & n9891 ;
  assign n9893 = n9890 | n9892 ;
  assign n9894 = n9889 | n9893 ;
  assign n9895 = n6940 | n9894 ;
  assign n9896 = ( n587 & n9894 ) | ( n587 & n9895 ) | ( n9894 & n9895 ) ;
  assign n9897 = x47 & n9896 ;
  assign n9898 = x47 & ~n9897 ;
  assign n9899 = ( n9896 & ~n9897 ) | ( n9896 & n9898 ) | ( ~n9897 & n9898 ) ;
  assign n9900 = n9888 | n9899 ;
  assign n9901 = n9888 & n9899 ;
  assign n9902 = n9900 & ~n9901 ;
  assign n9903 = n9832 & n9902 ;
  assign n9904 = n9832 | n9902 ;
  assign n9905 = ~n9903 & n9904 ;
  assign n9906 = x77 & n6068 ;
  assign n9907 = x76 & n6063 ;
  assign n9908 = x75 & ~n6062 ;
  assign n9909 = n6398 & n9908 ;
  assign n9910 = n9907 | n9909 ;
  assign n9911 = n9906 | n9910 ;
  assign n9912 = n6071 | n9911 ;
  assign n9913 = ( n846 & n9911 ) | ( n846 & n9912 ) | ( n9911 & n9912 ) ;
  assign n9914 = x44 & n9913 ;
  assign n9915 = x44 & ~n9914 ;
  assign n9916 = ( n9913 & ~n9914 ) | ( n9913 & n9915 ) | ( ~n9914 & n9915 ) ;
  assign n9917 = n9905 | n9916 ;
  assign n9918 = n9905 & n9916 ;
  assign n9919 = n9917 & ~n9918 ;
  assign n9920 = n9831 & n9919 ;
  assign n9921 = n9831 | n9919 ;
  assign n9922 = ~n9920 & n9921 ;
  assign n9923 = x80 & n5340 ;
  assign n9924 = x79 & n5335 ;
  assign n9925 = x78 & ~n5334 ;
  assign n9926 = n5580 & n9925 ;
  assign n9927 = n9924 | n9926 ;
  assign n9928 = n9923 | n9927 ;
  assign n9929 = n5343 | n9928 ;
  assign n9930 = ( n1147 & n9928 ) | ( n1147 & n9929 ) | ( n9928 & n9929 ) ;
  assign n9931 = x41 & n9930 ;
  assign n9932 = x41 & ~n9931 ;
  assign n9933 = ( n9930 & ~n9931 ) | ( n9930 & n9932 ) | ( ~n9931 & n9932 ) ;
  assign n9934 = n9922 & n9933 ;
  assign n9935 = n9922 & ~n9934 ;
  assign n9936 = ~n9922 & n9933 ;
  assign n9937 = n9935 | n9936 ;
  assign n9938 = n9554 | n9557 ;
  assign n9939 = n9937 | n9938 ;
  assign n9940 = n9937 & n9938 ;
  assign n9941 = n9939 & ~n9940 ;
  assign n9942 = ( n9829 & n9830 ) | ( n9829 & ~n9941 ) | ( n9830 & ~n9941 ) ;
  assign n9943 = ( ~n9830 & n9941 ) | ( ~n9830 & n9942 ) | ( n9941 & n9942 ) ;
  assign n9944 = ( ~n9829 & n9942 ) | ( ~n9829 & n9943 ) | ( n9942 & n9943 ) ;
  assign n9945 = n9818 & n9944 ;
  assign n9946 = n9818 | n9944 ;
  assign n9947 = ~n9945 & n9946 ;
  assign n9948 = n9589 | n9593 ;
  assign n9949 = n9947 | n9948 ;
  assign n9950 = n9947 & n9948 ;
  assign n9951 = n9949 & ~n9950 ;
  assign n9952 = x89 & n3314 ;
  assign n9953 = x88 & n3309 ;
  assign n9954 = x87 & ~n3308 ;
  assign n9955 = n3570 & n9954 ;
  assign n9956 = n9953 | n9955 ;
  assign n9957 = n9952 | n9956 ;
  assign n9958 = n3317 | n9957 ;
  assign n9959 = ( n2244 & n9957 ) | ( n2244 & n9958 ) | ( n9957 & n9958 ) ;
  assign n9960 = x32 & n9959 ;
  assign n9961 = x32 & ~n9960 ;
  assign n9962 = ( n9959 & ~n9960 ) | ( n9959 & n9961 ) | ( ~n9960 & n9961 ) ;
  assign n9963 = n9951 & n9962 ;
  assign n9964 = n9951 & ~n9963 ;
  assign n9965 = ~n9951 & n9962 ;
  assign n9966 = n9964 | n9965 ;
  assign n9967 = n9607 | n9612 ;
  assign n9968 = n9966 | n9967 ;
  assign n9969 = n9966 & n9967 ;
  assign n9970 = n9968 & ~n9969 ;
  assign n9971 = x92 & n2775 ;
  assign n9972 = x91 & n2770 ;
  assign n9973 = x90 & ~n2769 ;
  assign n9974 = n2978 & n9973 ;
  assign n9975 = n9972 | n9974 ;
  assign n9976 = n9971 | n9975 ;
  assign n9977 = n2778 | n9976 ;
  assign n9978 = ( n2904 & n9976 ) | ( n2904 & n9977 ) | ( n9976 & n9977 ) ;
  assign n9979 = x29 & n9978 ;
  assign n9980 = x29 & ~n9979 ;
  assign n9981 = ( n9978 & ~n9979 ) | ( n9978 & n9980 ) | ( ~n9979 & n9980 ) ;
  assign n9982 = n9970 & n9981 ;
  assign n9983 = n9970 & ~n9982 ;
  assign n9984 = ~n9970 & n9981 ;
  assign n9985 = n9983 | n9984 ;
  assign n9986 = n9625 | n9630 ;
  assign n9987 = n9985 | n9986 ;
  assign n9988 = n9985 & n9986 ;
  assign n9989 = n9987 & ~n9988 ;
  assign n9990 = x95 & n2280 ;
  assign n9991 = x94 & n2275 ;
  assign n9992 = x93 & ~n2274 ;
  assign n9993 = n2481 & n9992 ;
  assign n9994 = n9991 | n9993 ;
  assign n9995 = n9990 | n9994 ;
  assign n9996 = n2283 | n9995 ;
  assign n9997 = ( n3479 & n9995 ) | ( n3479 & n9996 ) | ( n9995 & n9996 ) ;
  assign n9998 = x26 & n9997 ;
  assign n9999 = x26 & ~n9998 ;
  assign n10000 = ( n9997 & ~n9998 ) | ( n9997 & n9999 ) | ( ~n9998 & n9999 ) ;
  assign n10001 = n9989 & n10000 ;
  assign n10002 = n9989 & ~n10001 ;
  assign n10003 = ~n9989 & n10000 ;
  assign n10004 = n10002 | n10003 ;
  assign n10005 = n9643 | n9646 ;
  assign n10006 = n10004 | n10005 ;
  assign n10007 = n10004 & n10005 ;
  assign n10008 = n10006 & ~n10007 ;
  assign n10009 = x98 & n1817 ;
  assign n10010 = x97 & n1812 ;
  assign n10011 = x96 & ~n1811 ;
  assign n10012 = n1977 & n10011 ;
  assign n10013 = n10010 | n10012 ;
  assign n10014 = n10009 | n10013 ;
  assign n10015 = n1820 | n10014 ;
  assign n10016 = ( n4105 & n10014 ) | ( n4105 & n10015 ) | ( n10014 & n10015 ) ;
  assign n10017 = x23 & n10016 ;
  assign n10018 = x23 & ~n10017 ;
  assign n10019 = ( n10016 & ~n10017 ) | ( n10016 & n10018 ) | ( ~n10017 & n10018 ) ;
  assign n10020 = n10008 & n10019 ;
  assign n10021 = n10008 & ~n10020 ;
  assign n10022 = ~n10008 & n10019 ;
  assign n10023 = n10021 | n10022 ;
  assign n10024 = n9650 | n10023 ;
  assign n10025 = n9650 & n10023 ;
  assign n10026 = n10024 & ~n10025 ;
  assign n10027 = x101 & n1421 ;
  assign n10028 = x100 & n1416 ;
  assign n10029 = x99 & ~n1415 ;
  assign n10030 = n1584 & n10029 ;
  assign n10031 = n10028 | n10030 ;
  assign n10032 = n10027 | n10031 ;
  assign n10033 = n1424 | n10032 ;
  assign n10034 = ( n4783 & n10032 ) | ( n4783 & n10033 ) | ( n10032 & n10033 ) ;
  assign n10035 = x20 & n10034 ;
  assign n10036 = x20 & ~n10035 ;
  assign n10037 = ( n10034 & ~n10035 ) | ( n10034 & n10036 ) | ( ~n10035 & n10036 ) ;
  assign n10038 = n10026 & n10037 ;
  assign n10039 = n10026 & ~n10038 ;
  assign n10040 = ~n10026 & n10037 ;
  assign n10041 = n10039 | n10040 ;
  assign n10042 = n9653 | n9658 ;
  assign n10043 = n10041 | n10042 ;
  assign n10044 = n10041 & n10042 ;
  assign n10045 = n10043 & ~n10044 ;
  assign n10046 = x104 & n1071 ;
  assign n10047 = x103 & n1066 ;
  assign n10048 = x102 & ~n1065 ;
  assign n10049 = n1189 & n10048 ;
  assign n10050 = n10047 | n10049 ;
  assign n10051 = n10046 | n10050 ;
  assign n10052 = n1074 | n10051 ;
  assign n10053 = ( n5295 & n10051 ) | ( n5295 & n10052 ) | ( n10051 & n10052 ) ;
  assign n10054 = x17 & n10053 ;
  assign n10055 = x17 & ~n10054 ;
  assign n10056 = ( n10053 & ~n10054 ) | ( n10053 & n10055 ) | ( ~n10054 & n10055 ) ;
  assign n10057 = n10045 & n10056 ;
  assign n10058 = n10045 & ~n10057 ;
  assign n10059 = ~n10045 & n10056 ;
  assign n10060 = n10058 | n10059 ;
  assign n10061 = n9671 | n9677 ;
  assign n10062 = n10060 | n10061 ;
  assign n10063 = n10060 & n10061 ;
  assign n10064 = n10062 & ~n10063 ;
  assign n10065 = x107 & n771 ;
  assign n10066 = x106 & n766 ;
  assign n10067 = x105 & ~n765 ;
  assign n10068 = n905 & n10067 ;
  assign n10069 = n10066 | n10068 ;
  assign n10070 = n10065 | n10069 ;
  assign n10071 = n774 | n10070 ;
  assign n10072 = ( n6328 & n10070 ) | ( n6328 & n10071 ) | ( n10070 & n10071 ) ;
  assign n10073 = x14 & n10072 ;
  assign n10074 = x14 & ~n10073 ;
  assign n10075 = ( n10072 & ~n10073 ) | ( n10072 & n10074 ) | ( ~n10073 & n10074 ) ;
  assign n10076 = n10064 | n10075 ;
  assign n10077 = n9807 & n10076 ;
  assign n10078 = n10064 & n10075 ;
  assign n10079 = n10076 & ~n10078 ;
  assign n10080 = ~n10077 & n10079 ;
  assign n10081 = x110 & n528 ;
  assign n10082 = x109 & n523 ;
  assign n10083 = x108 & ~n522 ;
  assign n10084 = n635 & n10083 ;
  assign n10085 = n10082 | n10084 ;
  assign n10086 = n10081 | n10085 ;
  assign n10087 = n531 | n10086 ;
  assign n10088 = ( n7189 & n10086 ) | ( n7189 & n10087 ) | ( n10086 & n10087 ) ;
  assign n10089 = x11 & n10088 ;
  assign n10090 = x11 & ~n10089 ;
  assign n10091 = ( n10088 & ~n10089 ) | ( n10088 & n10090 ) | ( ~n10089 & n10090 ) ;
  assign n10092 = n10080 | n10091 ;
  assign n10093 = n9807 & ~n10079 ;
  assign n10094 = n10092 | n10093 ;
  assign n10095 = ( n10080 & n10091 ) | ( n10080 & n10093 ) | ( n10091 & n10093 ) ;
  assign n10096 = n10094 & ~n10095 ;
  assign n10097 = n9806 & n10096 ;
  assign n10098 = n9806 | n10096 ;
  assign n10099 = ~n10097 & n10098 ;
  assign n10100 = x113 & n337 ;
  assign n10101 = x112 & n332 ;
  assign n10102 = x111 & ~n331 ;
  assign n10103 = n396 & n10102 ;
  assign n10104 = n10101 | n10103 ;
  assign n10105 = n10100 | n10104 ;
  assign n10106 = n340 | n10105 ;
  assign n10107 = ( n8113 & n10105 ) | ( n8113 & n10106 ) | ( n10105 & n10106 ) ;
  assign n10108 = x8 & n10107 ;
  assign n10109 = x8 & ~n10108 ;
  assign n10110 = ( n10107 & ~n10108 ) | ( n10107 & n10109 ) | ( ~n10108 & n10109 ) ;
  assign n10111 = n10099 | n10110 ;
  assign n10112 = n10099 & n10110 ;
  assign n10113 = n10111 & ~n10112 ;
  assign n10114 = n9727 | n9733 ;
  assign n10115 = n10113 & n10114 ;
  assign n10116 = n10113 | n10114 ;
  assign n10117 = ~n10115 & n10116 ;
  assign n10118 = ( n9804 & n9805 ) | ( n9804 & ~n10117 ) | ( n9805 & ~n10117 ) ;
  assign n10119 = ( ~n9805 & n10117 ) | ( ~n9805 & n10118 ) | ( n10117 & n10118 ) ;
  assign n10120 = ( ~n9804 & n10118 ) | ( ~n9804 & n10119 ) | ( n10118 & n10119 ) ;
  assign n10121 = n9793 & n10120 ;
  assign n10122 = n9793 | n10120 ;
  assign n10123 = ~n10121 & n10122 ;
  assign n10124 = n9772 | n9777 ;
  assign n10125 = n10123 & n10124 ;
  assign n10126 = n10123 | n10124 ;
  assign n10127 = ~n10125 & n10126 ;
  assign n10128 = n9982 | n9988 ;
  assign n10129 = x87 & n3913 ;
  assign n10130 = x86 & n3908 ;
  assign n10131 = x85 & ~n3907 ;
  assign n10132 = n4152 & n10131 ;
  assign n10133 = n10130 | n10132 ;
  assign n10134 = n10129 | n10133 ;
  assign n10135 = n3916 | n10134 ;
  assign n10136 = ( n2067 & n10134 ) | ( n2067 & n10135 ) | ( n10134 & n10135 ) ;
  assign n10137 = x35 & n10136 ;
  assign n10138 = x35 & ~n10137 ;
  assign n10139 = ( n10136 & ~n10137 ) | ( n10136 & n10138 ) | ( ~n10137 & n10138 ) ;
  assign n10256 = ( n9829 & n9830 ) | ( n9829 & n9941 ) | ( n9830 & n9941 ) ;
  assign n10140 = n9934 | n9940 ;
  assign n10141 = x72 & n7812 ;
  assign n10142 = x71 & n7807 ;
  assign n10143 = x70 & ~n7806 ;
  assign n10144 = n8136 & n10143 ;
  assign n10145 = n10142 | n10144 ;
  assign n10146 = n10141 | n10145 ;
  assign n10147 = ( n435 & n7815 ) | ( n435 & n10146 ) | ( n7815 & n10146 ) ;
  assign n10148 = ( x50 & ~n10146 ) | ( x50 & n10147 ) | ( ~n10146 & n10147 ) ;
  assign n10149 = ~n10147 & n10148 ;
  assign n10150 = n10146 | n10148 ;
  assign n10151 = ( ~x50 & n10149 ) | ( ~x50 & n10150 ) | ( n10149 & n10150 ) ;
  assign n10152 = n264 & n8837 ;
  assign n10153 = x69 & n8834 ;
  assign n10154 = x68 & n8829 ;
  assign n10155 = x67 & ~n8828 ;
  assign n10156 = n9159 & n10155 ;
  assign n10157 = n10154 | n10156 ;
  assign n10158 = n10153 | n10157 ;
  assign n10159 = n10152 | n10158 ;
  assign n10160 = x53 | n10159 ;
  assign n10161 = ~x53 & n10160 ;
  assign n10162 = ( ~n10159 & n10160 ) | ( ~n10159 & n10161 ) | ( n10160 & n10161 ) ;
  assign n10163 = x66 & n9853 ;
  assign n10164 = x65 & n9848 ;
  assign n10165 = ~n9485 & n9852 ;
  assign n10166 = x64 & ~n9847 ;
  assign n10167 = n10165 & n10166 ;
  assign n10168 = n10164 | n10167 ;
  assign n10169 = n10163 | n10168 ;
  assign n10170 = n153 & n9856 ;
  assign n10171 = n10169 | n10170 ;
  assign n10172 = x56 | n10171 ;
  assign n10173 = ~x56 & n10172 ;
  assign n10174 = ( ~n10171 & n10172 ) | ( ~n10171 & n10173 ) | ( n10172 & n10173 ) ;
  assign n10175 = n9863 | n10174 ;
  assign n10176 = n9863 & n10174 ;
  assign n10177 = n10175 & ~n10176 ;
  assign n10178 = n9878 | n9881 ;
  assign n10179 = ( n10162 & n10177 ) | ( n10162 & n10178 ) | ( n10177 & n10178 ) ;
  assign n10180 = ( n10177 & n10178 ) | ( n10177 & ~n10179 ) | ( n10178 & ~n10179 ) ;
  assign n10181 = ( n10162 & ~n10179 ) | ( n10162 & n10180 ) | ( ~n10179 & n10180 ) ;
  assign n10182 = n10151 | n10181 ;
  assign n10183 = n10151 & n10181 ;
  assign n10184 = n10182 & ~n10183 ;
  assign n10185 = n9884 | n9886 ;
  assign n10186 = n10184 & n10185 ;
  assign n10187 = n10184 | n10185 ;
  assign n10188 = ~n10186 & n10187 ;
  assign n10189 = x75 & n6937 ;
  assign n10190 = x74 & n6932 ;
  assign n10191 = x73 & ~n6931 ;
  assign n10192 = n7216 & n10191 ;
  assign n10193 = n10190 | n10192 ;
  assign n10194 = n10189 | n10193 ;
  assign n10195 = n6940 | n10194 ;
  assign n10196 = ( n609 & n10194 ) | ( n609 & n10195 ) | ( n10194 & n10195 ) ;
  assign n10197 = x47 & n10196 ;
  assign n10198 = x47 & ~n10197 ;
  assign n10199 = ( n10196 & ~n10197 ) | ( n10196 & n10198 ) | ( ~n10197 & n10198 ) ;
  assign n10200 = n10188 | n10199 ;
  assign n10201 = n10188 & n10199 ;
  assign n10202 = n10200 & ~n10201 ;
  assign n10203 = n9901 | n9903 ;
  assign n10204 = n10202 & n10203 ;
  assign n10205 = n10202 | n10203 ;
  assign n10206 = ~n10204 & n10205 ;
  assign n10207 = x78 & n6068 ;
  assign n10208 = x77 & n6063 ;
  assign n10209 = x76 & ~n6062 ;
  assign n10210 = n6398 & n10209 ;
  assign n10211 = n10208 | n10210 ;
  assign n10212 = n10207 | n10211 ;
  assign n10213 = n6071 | n10212 ;
  assign n10214 = ( n868 & n10212 ) | ( n868 & n10213 ) | ( n10212 & n10213 ) ;
  assign n10215 = x44 & n10214 ;
  assign n10216 = x44 & ~n10215 ;
  assign n10217 = ( n10214 & ~n10215 ) | ( n10214 & n10216 ) | ( ~n10215 & n10216 ) ;
  assign n10218 = n10206 & n10217 ;
  assign n10219 = n10206 & ~n10218 ;
  assign n10220 = ~n10206 & n10217 ;
  assign n10221 = n10219 | n10220 ;
  assign n10222 = n9918 | n9920 ;
  assign n10223 = n10221 & n10222 ;
  assign n10224 = n10221 | n10222 ;
  assign n10225 = ~n10223 & n10224 ;
  assign n10226 = x81 & n5340 ;
  assign n10227 = x80 & n5335 ;
  assign n10228 = x79 & ~n5334 ;
  assign n10229 = n5580 & n10228 ;
  assign n10230 = n10227 | n10229 ;
  assign n10231 = n10226 | n10230 ;
  assign n10232 = n5343 | n10231 ;
  assign n10233 = ( n1256 & n10231 ) | ( n1256 & n10232 ) | ( n10231 & n10232 ) ;
  assign n10234 = x41 & n10233 ;
  assign n10235 = x41 & ~n10234 ;
  assign n10236 = ( n10233 & ~n10234 ) | ( n10233 & n10235 ) | ( ~n10234 & n10235 ) ;
  assign n10237 = n10225 & n10236 ;
  assign n10238 = n10225 & ~n10237 ;
  assign n10239 = ~n10225 & n10236 ;
  assign n10240 = n10238 | n10239 ;
  assign n10241 = n10140 & n10240 ;
  assign n10242 = n10140 & ~n10241 ;
  assign n10243 = n10240 & ~n10241 ;
  assign n10244 = n10242 | n10243 ;
  assign n10245 = x84 & n4572 ;
  assign n10246 = x83 & n4567 ;
  assign n10247 = x82 & ~n4566 ;
  assign n10248 = n4828 & n10247 ;
  assign n10249 = n10246 | n10248 ;
  assign n10250 = n10245 | n10249 ;
  assign n10251 = n4575 | n10250 ;
  assign n10252 = ( n1537 & n10250 ) | ( n1537 & n10251 ) | ( n10250 & n10251 ) ;
  assign n10253 = x38 & n10252 ;
  assign n10254 = x38 & ~n10253 ;
  assign n10255 = ( n10252 & ~n10253 ) | ( n10252 & n10254 ) | ( ~n10253 & n10254 ) ;
  assign n10257 = ( n10244 & ~n10255 ) | ( n10244 & n10256 ) | ( ~n10255 & n10256 ) ;
  assign n10258 = ( ~n10244 & n10255 ) | ( ~n10244 & n10257 ) | ( n10255 & n10257 ) ;
  assign n10259 = ( ~n10256 & n10257 ) | ( ~n10256 & n10258 ) | ( n10257 & n10258 ) ;
  assign n10260 = n10139 & n10259 ;
  assign n10261 = n10139 | n10259 ;
  assign n10262 = ~n10260 & n10261 ;
  assign n10263 = n9945 | n9950 ;
  assign n10264 = n10262 | n10263 ;
  assign n10265 = n10262 & n10263 ;
  assign n10266 = n10264 & ~n10265 ;
  assign n10267 = x90 & n3314 ;
  assign n10268 = x89 & n3309 ;
  assign n10269 = x88 & ~n3308 ;
  assign n10270 = n3570 & n10269 ;
  assign n10271 = n10268 | n10270 ;
  assign n10272 = n10267 | n10271 ;
  assign n10273 = n3317 | n10272 ;
  assign n10274 = ( n2410 & n10272 ) | ( n2410 & n10273 ) | ( n10272 & n10273 ) ;
  assign n10275 = x32 & n10274 ;
  assign n10276 = x32 & ~n10275 ;
  assign n10277 = ( n10274 & ~n10275 ) | ( n10274 & n10276 ) | ( ~n10275 & n10276 ) ;
  assign n10278 = n10266 & n10277 ;
  assign n10279 = n10266 | n10277 ;
  assign n10280 = ~n10278 & n10279 ;
  assign n10281 = n9963 | n9969 ;
  assign n10282 = n10280 | n10281 ;
  assign n10283 = n10280 & n10281 ;
  assign n10284 = n10282 & ~n10283 ;
  assign n10285 = x93 & n2775 ;
  assign n10286 = x92 & n2770 ;
  assign n10287 = x91 & ~n2769 ;
  assign n10288 = n2978 & n10287 ;
  assign n10289 = n10286 | n10288 ;
  assign n10290 = n10285 | n10289 ;
  assign n10291 = n2778 | n10290 ;
  assign n10292 = ( n2931 & n10290 ) | ( n2931 & n10291 ) | ( n10290 & n10291 ) ;
  assign n10293 = x29 & n10292 ;
  assign n10294 = x29 & ~n10293 ;
  assign n10295 = ( n10292 & ~n10293 ) | ( n10292 & n10294 ) | ( ~n10293 & n10294 ) ;
  assign n10296 = n10284 | n10295 ;
  assign n10297 = n10284 & n10295 ;
  assign n10298 = n10296 & ~n10297 ;
  assign n10299 = n10128 & n10298 ;
  assign n10300 = n10128 | n10298 ;
  assign n10301 = ~n10299 & n10300 ;
  assign n10302 = x96 & n2280 ;
  assign n10303 = x95 & n2275 ;
  assign n10304 = x94 & ~n2274 ;
  assign n10305 = n2481 & n10304 ;
  assign n10306 = n10303 | n10305 ;
  assign n10307 = n10302 | n10306 ;
  assign n10308 = n2283 | n10307 ;
  assign n10309 = ( n3509 & n10307 ) | ( n3509 & n10308 ) | ( n10307 & n10308 ) ;
  assign n10310 = x26 & n10309 ;
  assign n10311 = x26 & ~n10310 ;
  assign n10312 = ( n10309 & ~n10310 ) | ( n10309 & n10311 ) | ( ~n10310 & n10311 ) ;
  assign n10313 = n10301 | n10312 ;
  assign n10314 = n10301 & n10312 ;
  assign n10315 = n10313 & ~n10314 ;
  assign n10316 = n10001 | n10007 ;
  assign n10317 = n10315 & n10316 ;
  assign n10318 = n10315 | n10316 ;
  assign n10319 = ~n10317 & n10318 ;
  assign n10320 = x99 & n1817 ;
  assign n10321 = x98 & n1812 ;
  assign n10322 = x97 & ~n1811 ;
  assign n10323 = n1977 & n10322 ;
  assign n10324 = n10321 | n10323 ;
  assign n10325 = n10320 | n10324 ;
  assign n10326 = n1820 | n10325 ;
  assign n10327 = ( n4325 & n10325 ) | ( n4325 & n10326 ) | ( n10325 & n10326 ) ;
  assign n10328 = x23 & n10327 ;
  assign n10329 = x23 & ~n10328 ;
  assign n10330 = ( n10327 & ~n10328 ) | ( n10327 & n10329 ) | ( ~n10328 & n10329 ) ;
  assign n10331 = n10319 & n10330 ;
  assign n10332 = n10319 & ~n10331 ;
  assign n10333 = ~n10319 & n10330 ;
  assign n10334 = n10332 | n10333 ;
  assign n10335 = n10020 | n10025 ;
  assign n10336 = n10334 | n10335 ;
  assign n10337 = n10334 & n10335 ;
  assign n10338 = n10336 & ~n10337 ;
  assign n10339 = x102 & n1421 ;
  assign n10340 = x101 & n1416 ;
  assign n10341 = x100 & ~n1415 ;
  assign n10342 = n1584 & n10341 ;
  assign n10343 = n10340 | n10342 ;
  assign n10344 = n10339 | n10343 ;
  assign n10345 = n1424 | n10344 ;
  assign n10346 = ( n5025 & n10344 ) | ( n5025 & n10345 ) | ( n10344 & n10345 ) ;
  assign n10347 = x20 & n10346 ;
  assign n10348 = x20 & ~n10347 ;
  assign n10349 = ( n10346 & ~n10347 ) | ( n10346 & n10348 ) | ( ~n10347 & n10348 ) ;
  assign n10350 = n10338 & n10349 ;
  assign n10351 = n10338 & ~n10350 ;
  assign n10352 = ~n10338 & n10349 ;
  assign n10353 = n10351 | n10352 ;
  assign n10354 = n10038 | n10044 ;
  assign n10355 = n10353 | n10354 ;
  assign n10356 = n10353 & n10354 ;
  assign n10357 = n10355 & ~n10356 ;
  assign n10358 = x105 & n1071 ;
  assign n10359 = x104 & n1066 ;
  assign n10360 = x103 & ~n1065 ;
  assign n10361 = n1189 & n10360 ;
  assign n10362 = n10359 | n10361 ;
  assign n10363 = n10358 | n10362 ;
  assign n10364 = n1074 | n10363 ;
  assign n10365 = ( n5788 & n10363 ) | ( n5788 & n10364 ) | ( n10363 & n10364 ) ;
  assign n10366 = x17 & n10365 ;
  assign n10367 = x17 & ~n10366 ;
  assign n10368 = ( n10365 & ~n10366 ) | ( n10365 & n10367 ) | ( ~n10366 & n10367 ) ;
  assign n10369 = n10357 & n10368 ;
  assign n10370 = n10357 & ~n10369 ;
  assign n10371 = ~n10357 & n10368 ;
  assign n10372 = n10370 | n10371 ;
  assign n10373 = n10057 | n10063 ;
  assign n10374 = n10372 | n10373 ;
  assign n10375 = n10372 & n10373 ;
  assign n10376 = n10374 & ~n10375 ;
  assign n10377 = x108 & n771 ;
  assign n10378 = x107 & n766 ;
  assign n10379 = x106 & ~n765 ;
  assign n10380 = n905 & n10379 ;
  assign n10381 = n10378 | n10380 ;
  assign n10382 = n10377 | n10381 ;
  assign n10383 = n774 | n10382 ;
  assign n10384 = ( n6358 & n10382 ) | ( n6358 & n10383 ) | ( n10382 & n10383 ) ;
  assign n10385 = x14 & n10384 ;
  assign n10386 = x14 & ~n10385 ;
  assign n10387 = ( n10384 & ~n10385 ) | ( n10384 & n10386 ) | ( ~n10385 & n10386 ) ;
  assign n10388 = n10376 & n10387 ;
  assign n10389 = n10376 | n10387 ;
  assign n10390 = ~n10388 & n10389 ;
  assign n10391 = n10077 | n10078 ;
  assign n10392 = n10390 & n10391 ;
  assign n10393 = n10391 & ~n10392 ;
  assign n10394 = ( n10390 & ~n10392 ) | ( n10390 & n10393 ) | ( ~n10392 & n10393 ) ;
  assign n10395 = x111 & n528 ;
  assign n10396 = x110 & n523 ;
  assign n10397 = x109 & ~n522 ;
  assign n10398 = n635 & n10397 ;
  assign n10399 = n10396 | n10398 ;
  assign n10400 = n10395 | n10399 ;
  assign n10401 = n531 | n10400 ;
  assign n10402 = ( n7492 & n10400 ) | ( n7492 & n10401 ) | ( n10400 & n10401 ) ;
  assign n10403 = x11 & n10402 ;
  assign n10404 = x11 & ~n10403 ;
  assign n10405 = ( n10402 & ~n10403 ) | ( n10402 & n10404 ) | ( ~n10403 & n10404 ) ;
  assign n10406 = n10394 & n10405 ;
  assign n10407 = n10394 & ~n10406 ;
  assign n10408 = ~n10394 & n10405 ;
  assign n10409 = n10407 | n10408 ;
  assign n10410 = n10095 | n10097 ;
  assign n10411 = n10409 & n10410 ;
  assign n10412 = n10409 | n10410 ;
  assign n10413 = ~n10411 & n10412 ;
  assign n10414 = x114 & n337 ;
  assign n10415 = x113 & n332 ;
  assign n10416 = x112 & ~n331 ;
  assign n10417 = n396 & n10416 ;
  assign n10418 = n10415 | n10417 ;
  assign n10419 = n10414 | n10418 ;
  assign n10420 = n340 | n10419 ;
  assign n10421 = ( n8437 & n10419 ) | ( n8437 & n10420 ) | ( n10419 & n10420 ) ;
  assign n10422 = x8 & n10421 ;
  assign n10423 = x8 & ~n10422 ;
  assign n10424 = ( n10421 & ~n10422 ) | ( n10421 & n10423 ) | ( ~n10422 & n10423 ) ;
  assign n10425 = ~n10413 & n10424 ;
  assign n10426 = n10413 & ~n10424 ;
  assign n10427 = n10425 | n10426 ;
  assign n10428 = n10112 | n10115 ;
  assign n10429 = n10427 & ~n10428 ;
  assign n10430 = ~n10427 & n10428 ;
  assign n10431 = x117 & n206 ;
  assign n10432 = x116 & n201 ;
  assign n10433 = x115 & ~n200 ;
  assign n10434 = n243 & n10433 ;
  assign n10435 = n10432 | n10434 ;
  assign n10436 = n10431 | n10435 ;
  assign n10437 = n209 | n10436 ;
  assign n10438 = ( n9118 & n10436 ) | ( n9118 & n10437 ) | ( n10436 & n10437 ) ;
  assign n10439 = x5 & n10438 ;
  assign n10440 = x5 & ~n10439 ;
  assign n10441 = ( n10438 & ~n10439 ) | ( n10438 & n10440 ) | ( ~n10439 & n10440 ) ;
  assign n10442 = n10430 | n10441 ;
  assign n10443 = n10429 | n10442 ;
  assign n10444 = ( n10429 & n10430 ) | ( n10429 & n10441 ) | ( n10430 & n10441 ) ;
  assign n10445 = n10443 & ~n10444 ;
  assign n10446 = ( n9804 & n9805 ) | ( n9804 & n10117 ) | ( n9805 & n10117 ) ;
  assign n10447 = n10445 | n10446 ;
  assign n10448 = n10445 & n10446 ;
  assign n10449 = n10447 & ~n10448 ;
  assign n10450 = x118 | x119 ;
  assign n10451 = x119 | x120 ;
  assign n10452 = x119 & x120 ;
  assign n10453 = n10451 & ~n10452 ;
  assign n10454 = n10450 & n10453 ;
  assign n10455 = x118 & x119 ;
  assign n10456 = n10453 & n10455 ;
  assign n10457 = ( n9786 & n10454 ) | ( n9786 & n10456 ) | ( n10454 & n10456 ) ;
  assign n10458 = ( n9786 & n10450 ) | ( n9786 & n10455 ) | ( n10450 & n10455 ) ;
  assign n10459 = n10453 | n10458 ;
  assign n10460 = ~n10457 & n10459 ;
  assign n10461 = x119 & n131 ;
  assign n10462 = x118 & ~n156 ;
  assign n10463 = ( n135 & n10461 ) | ( n135 & n10462 ) | ( n10461 & n10462 ) ;
  assign n10464 = x0 & x120 ;
  assign n10465 = ( ~n135 & n10461 ) | ( ~n135 & n10464 ) | ( n10461 & n10464 ) ;
  assign n10466 = n10463 | n10465 ;
  assign n10467 = n139 | n10466 ;
  assign n10468 = ( n10460 & n10466 ) | ( n10460 & n10467 ) | ( n10466 & n10467 ) ;
  assign n10469 = x2 & n10468 ;
  assign n10470 = x2 & ~n10469 ;
  assign n10471 = ( n10468 & ~n10469 ) | ( n10468 & n10470 ) | ( ~n10469 & n10470 ) ;
  assign n10472 = n10449 & n10471 ;
  assign n10473 = n10449 & ~n10472 ;
  assign n10474 = ~n10449 & n10471 ;
  assign n10475 = n10473 | n10474 ;
  assign n10476 = n10121 | n10125 ;
  assign n10477 = n10475 & n10476 ;
  assign n10478 = n10475 | n10476 ;
  assign n10479 = ~n10477 & n10478 ;
  assign n10480 = n10444 | n10448 ;
  assign n10481 = n10388 | n10392 ;
  assign n10482 = n10331 | n10337 ;
  assign n10483 = x100 & n1817 ;
  assign n10484 = x99 & n1812 ;
  assign n10485 = x98 & ~n1811 ;
  assign n10486 = n1977 & n10485 ;
  assign n10487 = n10484 | n10486 ;
  assign n10488 = n10483 | n10487 ;
  assign n10489 = n1820 | n10488 ;
  assign n10490 = ( n4532 & n10488 ) | ( n4532 & n10489 ) | ( n10488 & n10489 ) ;
  assign n10491 = x23 & n10490 ;
  assign n10492 = x23 & ~n10491 ;
  assign n10493 = ( n10490 & ~n10491 ) | ( n10490 & n10492 ) | ( ~n10491 & n10492 ) ;
  assign n10494 = x97 & n2280 ;
  assign n10495 = x96 & n2275 ;
  assign n10496 = x95 & ~n2274 ;
  assign n10497 = n2481 & n10496 ;
  assign n10498 = n10495 | n10497 ;
  assign n10499 = n10494 | n10498 ;
  assign n10500 = n2283 | n10499 ;
  assign n10501 = ( n3707 & n10499 ) | ( n3707 & n10500 ) | ( n10499 & n10500 ) ;
  assign n10502 = x26 & n10501 ;
  assign n10503 = x26 & ~n10502 ;
  assign n10504 = ( n10501 & ~n10502 ) | ( n10501 & n10503 ) | ( ~n10502 & n10503 ) ;
  assign n10505 = n10314 | n10317 ;
  assign n10506 = n10278 | n10283 ;
  assign n10507 = x85 & n4572 ;
  assign n10508 = x84 & n4567 ;
  assign n10509 = x83 & ~n4566 ;
  assign n10510 = n4828 & n10509 ;
  assign n10511 = n10508 | n10510 ;
  assign n10512 = n10507 | n10511 ;
  assign n10513 = n4575 | n10512 ;
  assign n10514 = ( n1765 & n10512 ) | ( n1765 & n10513 ) | ( n10512 & n10513 ) ;
  assign n10515 = x38 & n10514 ;
  assign n10516 = x38 & ~n10515 ;
  assign n10517 = ( n10514 & ~n10515 ) | ( n10514 & n10516 ) | ( ~n10515 & n10516 ) ;
  assign n10518 = n10237 | n10241 ;
  assign n10519 = n10183 | n10186 ;
  assign n10520 = x70 & n8834 ;
  assign n10521 = x69 & n8829 ;
  assign n10522 = x68 & ~n8828 ;
  assign n10523 = n9159 & n10522 ;
  assign n10524 = n10521 | n10523 ;
  assign n10525 = n10520 | n10524 ;
  assign n10526 = n8837 | n10525 ;
  assign n10527 = ( n310 & n10525 ) | ( n310 & n10526 ) | ( n10525 & n10526 ) ;
  assign n10528 = x53 & ~n10527 ;
  assign n10529 = ~x53 & n10527 ;
  assign n10530 = n10528 | n10529 ;
  assign n10531 = x56 & ~x57 ;
  assign n10532 = ~x56 & x57 ;
  assign n10533 = n10531 | n10532 ;
  assign n10534 = x64 & n10533 ;
  assign n10535 = x67 & n9853 ;
  assign n10536 = x66 & n9848 ;
  assign n10537 = x65 & ~n9847 ;
  assign n10538 = n10165 & n10537 ;
  assign n10539 = n10536 | n10538 ;
  assign n10540 = n10535 | n10539 ;
  assign n10541 = n180 & n9856 ;
  assign n10542 = n10540 | n10541 ;
  assign n10543 = x56 & ~n10542 ;
  assign n10544 = ~x56 & n10542 ;
  assign n10545 = n10543 | n10544 ;
  assign n10546 = ( n10176 & n10534 ) | ( n10176 & n10545 ) | ( n10534 & n10545 ) ;
  assign n10547 = ( n10176 & n10545 ) | ( n10176 & ~n10546 ) | ( n10545 & ~n10546 ) ;
  assign n10548 = ( n10534 & ~n10546 ) | ( n10534 & n10547 ) | ( ~n10546 & n10547 ) ;
  assign n10549 = ( n10179 & n10530 ) | ( n10179 & ~n10548 ) | ( n10530 & ~n10548 ) ;
  assign n10550 = ( ~n10179 & n10548 ) | ( ~n10179 & n10549 ) | ( n10548 & n10549 ) ;
  assign n10551 = ( ~n10530 & n10549 ) | ( ~n10530 & n10550 ) | ( n10549 & n10550 ) ;
  assign n10552 = x73 & n7812 ;
  assign n10553 = x72 & n7807 ;
  assign n10554 = x71 & ~n7806 ;
  assign n10555 = n8136 & n10554 ;
  assign n10556 = n10553 | n10555 ;
  assign n10557 = n10552 | n10556 ;
  assign n10558 = ( n499 & n7815 ) | ( n499 & n10557 ) | ( n7815 & n10557 ) ;
  assign n10559 = ( x50 & ~n10557 ) | ( x50 & n10558 ) | ( ~n10557 & n10558 ) ;
  assign n10560 = ~n10558 & n10559 ;
  assign n10561 = n10557 | n10559 ;
  assign n10562 = ( ~x50 & n10560 ) | ( ~x50 & n10561 ) | ( n10560 & n10561 ) ;
  assign n10563 = n10551 & n10562 ;
  assign n10564 = n10551 | n10562 ;
  assign n10565 = ~n10563 & n10564 ;
  assign n10566 = n10519 & n10565 ;
  assign n10567 = n10519 | n10565 ;
  assign n10568 = ~n10566 & n10567 ;
  assign n10569 = x76 & n6937 ;
  assign n10570 = x75 & n6932 ;
  assign n10571 = x74 & ~n6931 ;
  assign n10572 = n7216 & n10571 ;
  assign n10573 = n10570 | n10572 ;
  assign n10574 = n10569 | n10573 ;
  assign n10575 = n6940 | n10574 ;
  assign n10576 = ( n740 & n10574 ) | ( n740 & n10575 ) | ( n10574 & n10575 ) ;
  assign n10577 = x47 & n10576 ;
  assign n10578 = x47 & ~n10577 ;
  assign n10579 = ( n10576 & ~n10577 ) | ( n10576 & n10578 ) | ( ~n10577 & n10578 ) ;
  assign n10580 = n10568 | n10579 ;
  assign n10581 = n10568 & n10579 ;
  assign n10582 = n10580 & ~n10581 ;
  assign n10583 = n10201 | n10204 ;
  assign n10584 = n10582 & n10583 ;
  assign n10585 = n10582 | n10583 ;
  assign n10586 = ~n10584 & n10585 ;
  assign n10587 = x79 & n6068 ;
  assign n10588 = x78 & n6063 ;
  assign n10589 = x77 & ~n6062 ;
  assign n10590 = n6398 & n10589 ;
  assign n10591 = n10588 | n10590 ;
  assign n10592 = n10587 | n10591 ;
  assign n10593 = n6071 | n10592 ;
  assign n10594 = ( n961 & n10592 ) | ( n961 & n10593 ) | ( n10592 & n10593 ) ;
  assign n10595 = x44 & n10594 ;
  assign n10596 = x44 & ~n10595 ;
  assign n10597 = ( n10594 & ~n10595 ) | ( n10594 & n10596 ) | ( ~n10595 & n10596 ) ;
  assign n10598 = n10586 & n10597 ;
  assign n10599 = n10586 | n10597 ;
  assign n10600 = ~n10598 & n10599 ;
  assign n10601 = n10218 | n10600 ;
  assign n10602 = n10223 | n10601 ;
  assign n10603 = ( n10218 & n10223 ) | ( n10218 & n10600 ) | ( n10223 & n10600 ) ;
  assign n10604 = n10602 & ~n10603 ;
  assign n10605 = x82 & n5340 ;
  assign n10606 = x81 & n5335 ;
  assign n10607 = x80 & ~n5334 ;
  assign n10608 = n5580 & n10607 ;
  assign n10609 = n10606 | n10608 ;
  assign n10610 = n10605 | n10609 ;
  assign n10611 = n5343 | n10610 ;
  assign n10612 = ( n1371 & n10610 ) | ( n1371 & n10611 ) | ( n10610 & n10611 ) ;
  assign n10613 = x41 & n10612 ;
  assign n10614 = x41 & ~n10613 ;
  assign n10615 = ( n10612 & ~n10613 ) | ( n10612 & n10614 ) | ( ~n10613 & n10614 ) ;
  assign n10616 = ( n10518 & n10604 ) | ( n10518 & n10615 ) | ( n10604 & n10615 ) ;
  assign n10617 = ( n10604 & n10615 ) | ( n10604 & ~n10616 ) | ( n10615 & ~n10616 ) ;
  assign n10618 = ( n10518 & ~n10616 ) | ( n10518 & n10617 ) | ( ~n10616 & n10617 ) ;
  assign n10619 = n10517 & n10618 ;
  assign n10620 = n10517 | n10618 ;
  assign n10621 = ~n10619 & n10620 ;
  assign n10622 = ( n10244 & n10255 ) | ( n10244 & n10256 ) | ( n10255 & n10256 ) ;
  assign n10623 = n10621 | n10622 ;
  assign n10624 = n10621 & n10622 ;
  assign n10625 = n10623 & ~n10624 ;
  assign n10626 = x88 & n3913 ;
  assign n10627 = x87 & n3908 ;
  assign n10628 = x86 & ~n3907 ;
  assign n10629 = n4152 & n10628 ;
  assign n10630 = n10627 | n10629 ;
  assign n10631 = n10626 | n10630 ;
  assign n10632 = n3916 | n10631 ;
  assign n10633 = ( n2095 & n10631 ) | ( n2095 & n10632 ) | ( n10631 & n10632 ) ;
  assign n10634 = x35 & n10633 ;
  assign n10635 = x35 & ~n10634 ;
  assign n10636 = ( n10633 & ~n10634 ) | ( n10633 & n10635 ) | ( ~n10634 & n10635 ) ;
  assign n10637 = n10625 & n10636 ;
  assign n10638 = n10625 & ~n10637 ;
  assign n10639 = ~n10625 & n10636 ;
  assign n10640 = n10638 | n10639 ;
  assign n10641 = n10260 | n10265 ;
  assign n10642 = n10640 | n10641 ;
  assign n10643 = n10640 & n10641 ;
  assign n10644 = n10642 & ~n10643 ;
  assign n10645 = x91 & n3314 ;
  assign n10646 = x90 & n3309 ;
  assign n10647 = x89 & ~n3308 ;
  assign n10648 = n3570 & n10647 ;
  assign n10649 = n10646 | n10648 ;
  assign n10650 = n10645 | n10649 ;
  assign n10651 = n3317 | n10650 ;
  assign n10652 = ( n2714 & n10650 ) | ( n2714 & n10651 ) | ( n10650 & n10651 ) ;
  assign n10653 = x32 & n10652 ;
  assign n10654 = x32 & ~n10653 ;
  assign n10655 = ( n10652 & ~n10653 ) | ( n10652 & n10654 ) | ( ~n10653 & n10654 ) ;
  assign n10656 = n10644 | n10655 ;
  assign n10657 = n10644 & n10655 ;
  assign n10658 = n10656 & ~n10657 ;
  assign n10659 = n10506 & n10658 ;
  assign n10660 = n10506 | n10658 ;
  assign n10661 = ~n10659 & n10660 ;
  assign n10662 = x94 & n2775 ;
  assign n10663 = x93 & n2770 ;
  assign n10664 = x92 & ~n2769 ;
  assign n10665 = n2978 & n10664 ;
  assign n10666 = n10663 | n10665 ;
  assign n10667 = n10662 | n10666 ;
  assign n10668 = n2778 | n10667 ;
  assign n10669 = ( n3271 & n10667 ) | ( n3271 & n10668 ) | ( n10667 & n10668 ) ;
  assign n10670 = x29 & n10669 ;
  assign n10671 = x29 & ~n10670 ;
  assign n10672 = ( n10669 & ~n10670 ) | ( n10669 & n10671 ) | ( ~n10670 & n10671 ) ;
  assign n10673 = n10661 & n10672 ;
  assign n10674 = n10661 | n10672 ;
  assign n10675 = ~n10673 & n10674 ;
  assign n10676 = n10297 | n10299 ;
  assign n10677 = n10675 & n10676 ;
  assign n10678 = n10675 | n10676 ;
  assign n10679 = ~n10677 & n10678 ;
  assign n10680 = ( n10504 & n10505 ) | ( n10504 & ~n10679 ) | ( n10505 & ~n10679 ) ;
  assign n10681 = ( ~n10505 & n10679 ) | ( ~n10505 & n10680 ) | ( n10679 & n10680 ) ;
  assign n10682 = ( ~n10504 & n10680 ) | ( ~n10504 & n10681 ) | ( n10680 & n10681 ) ;
  assign n10683 = n10493 & n10682 ;
  assign n10684 = n10493 | n10682 ;
  assign n10685 = ~n10683 & n10684 ;
  assign n10686 = n10482 | n10685 ;
  assign n10687 = n10482 & n10685 ;
  assign n10688 = n10686 & ~n10687 ;
  assign n10689 = x103 & n1421 ;
  assign n10690 = x102 & n1416 ;
  assign n10691 = x101 & ~n1415 ;
  assign n10692 = n1584 & n10691 ;
  assign n10693 = n10690 | n10692 ;
  assign n10694 = n10689 | n10693 ;
  assign n10695 = n1424 | n10694 ;
  assign n10696 = ( n5264 & n10694 ) | ( n5264 & n10695 ) | ( n10694 & n10695 ) ;
  assign n10697 = x20 & n10696 ;
  assign n10698 = x20 & ~n10697 ;
  assign n10699 = ( n10696 & ~n10697 ) | ( n10696 & n10698 ) | ( ~n10697 & n10698 ) ;
  assign n10700 = n10688 & n10699 ;
  assign n10701 = n10688 & ~n10700 ;
  assign n10702 = ~n10688 & n10699 ;
  assign n10703 = n10701 | n10702 ;
  assign n10704 = n10350 | n10356 ;
  assign n10705 = n10703 | n10704 ;
  assign n10706 = n10703 & n10704 ;
  assign n10707 = n10705 & ~n10706 ;
  assign n10708 = x106 & n1071 ;
  assign n10709 = x105 & n1066 ;
  assign n10710 = x104 & ~n1065 ;
  assign n10711 = n1189 & n10710 ;
  assign n10712 = n10709 | n10711 ;
  assign n10713 = n10708 | n10712 ;
  assign n10714 = n1074 | n10713 ;
  assign n10715 = ( n5814 & n10713 ) | ( n5814 & n10714 ) | ( n10713 & n10714 ) ;
  assign n10716 = x17 & n10715 ;
  assign n10717 = x17 & ~n10716 ;
  assign n10718 = ( n10715 & ~n10716 ) | ( n10715 & n10717 ) | ( ~n10716 & n10717 ) ;
  assign n10719 = n10707 | n10718 ;
  assign n10720 = n10707 & n10718 ;
  assign n10721 = n10719 & ~n10720 ;
  assign n10722 = n10369 | n10375 ;
  assign n10723 = n10721 & n10722 ;
  assign n10724 = n10721 | n10722 ;
  assign n10725 = ~n10723 & n10724 ;
  assign n10726 = x109 & n771 ;
  assign n10727 = x108 & n766 ;
  assign n10728 = x107 & ~n765 ;
  assign n10729 = n905 & n10728 ;
  assign n10730 = n10727 | n10729 ;
  assign n10731 = n10726 | n10730 ;
  assign n10732 = n774 | n10731 ;
  assign n10733 = ( n6884 & n10731 ) | ( n6884 & n10732 ) | ( n10731 & n10732 ) ;
  assign n10734 = x14 & n10733 ;
  assign n10735 = x14 & ~n10734 ;
  assign n10736 = ( n10733 & ~n10734 ) | ( n10733 & n10735 ) | ( ~n10734 & n10735 ) ;
  assign n10737 = n10725 & n10736 ;
  assign n10738 = n10725 & ~n10737 ;
  assign n10739 = ~n10725 & n10736 ;
  assign n10740 = n10738 | n10739 ;
  assign n10741 = n10481 & n10740 ;
  assign n10742 = n10481 | n10740 ;
  assign n10743 = ~n10741 & n10742 ;
  assign n10744 = x112 & n528 ;
  assign n10745 = x111 & n523 ;
  assign n10746 = x110 & ~n522 ;
  assign n10747 = n635 & n10746 ;
  assign n10748 = n10745 | n10747 ;
  assign n10749 = n10744 | n10748 ;
  assign n10750 = n531 | n10749 ;
  assign n10751 = ( n7789 & n10749 ) | ( n7789 & n10750 ) | ( n10749 & n10750 ) ;
  assign n10752 = x11 & n10751 ;
  assign n10753 = x11 & ~n10752 ;
  assign n10754 = ( n10751 & ~n10752 ) | ( n10751 & n10753 ) | ( ~n10752 & n10753 ) ;
  assign n10755 = n10743 & n10754 ;
  assign n10756 = n10743 & ~n10755 ;
  assign n10757 = ~n10743 & n10754 ;
  assign n10758 = n10756 | n10757 ;
  assign n10759 = n10406 | n10411 ;
  assign n10760 = n10758 & n10759 ;
  assign n10761 = n10758 | n10759 ;
  assign n10762 = ~n10760 & n10761 ;
  assign n10763 = x115 & n337 ;
  assign n10764 = x114 & n332 ;
  assign n10765 = x113 & ~n331 ;
  assign n10766 = n396 & n10765 ;
  assign n10767 = n10764 | n10766 ;
  assign n10768 = n10763 | n10767 ;
  assign n10769 = n340 | n10768 ;
  assign n10770 = ( n8749 & n10768 ) | ( n8749 & n10769 ) | ( n10768 & n10769 ) ;
  assign n10771 = x8 & n10770 ;
  assign n10772 = x8 & ~n10771 ;
  assign n10773 = ( n10770 & ~n10771 ) | ( n10770 & n10772 ) | ( ~n10771 & n10772 ) ;
  assign n10774 = n10762 & n10773 ;
  assign n10775 = n10762 & ~n10774 ;
  assign n10776 = ~n10762 & n10773 ;
  assign n10777 = n10775 | n10776 ;
  assign n10778 = ( n10413 & n10424 ) | ( n10413 & n10428 ) | ( n10424 & n10428 ) ;
  assign n10779 = n10777 & n10778 ;
  assign n10780 = n10777 | n10778 ;
  assign n10781 = ~n10779 & n10780 ;
  assign n10782 = x118 & n206 ;
  assign n10783 = x117 & n201 ;
  assign n10784 = x116 & ~n200 ;
  assign n10785 = n243 & n10784 ;
  assign n10786 = n10783 | n10785 ;
  assign n10787 = n10782 | n10786 ;
  assign n10788 = n209 | n10787 ;
  assign n10789 = ( n9760 & n10787 ) | ( n9760 & n10788 ) | ( n10787 & n10788 ) ;
  assign n10790 = x5 & n10789 ;
  assign n10791 = x5 & ~n10790 ;
  assign n10792 = ( n10789 & ~n10790 ) | ( n10789 & n10791 ) | ( ~n10790 & n10791 ) ;
  assign n10793 = n10781 & n10792 ;
  assign n10794 = n10781 & ~n10793 ;
  assign n10795 = ~n10781 & n10792 ;
  assign n10796 = n10794 | n10795 ;
  assign n10797 = n10480 & n10796 ;
  assign n10798 = n10480 & ~n10797 ;
  assign n10799 = n10796 & ~n10797 ;
  assign n10800 = n10798 | n10799 ;
  assign n10801 = x120 | x121 ;
  assign n10802 = x120 & x121 ;
  assign n10803 = n10801 & ~n10802 ;
  assign n10804 = n10452 | n10454 ;
  assign n10805 = n10803 & n10804 ;
  assign n10806 = n10452 | n10456 ;
  assign n10807 = n10803 & n10806 ;
  assign n10808 = ( n9786 & n10805 ) | ( n9786 & n10807 ) | ( n10805 & n10807 ) ;
  assign n10809 = ( n9786 & n10804 ) | ( n9786 & n10806 ) | ( n10804 & n10806 ) ;
  assign n10810 = n10803 | n10809 ;
  assign n10811 = ~n10808 & n10810 ;
  assign n10812 = x120 & n131 ;
  assign n10813 = x119 & ~n156 ;
  assign n10814 = ( n135 & n10812 ) | ( n135 & n10813 ) | ( n10812 & n10813 ) ;
  assign n10815 = x0 & x121 ;
  assign n10816 = ( ~n135 & n10812 ) | ( ~n135 & n10815 ) | ( n10812 & n10815 ) ;
  assign n10817 = n10814 | n10816 ;
  assign n10818 = n139 | n10817 ;
  assign n10819 = ( n10811 & n10817 ) | ( n10811 & n10818 ) | ( n10817 & n10818 ) ;
  assign n10820 = x2 & n10819 ;
  assign n10821 = x2 & ~n10820 ;
  assign n10822 = ( n10819 & ~n10820 ) | ( n10819 & n10821 ) | ( ~n10820 & n10821 ) ;
  assign n10823 = n10800 & n10822 ;
  assign n10824 = n10800 & ~n10823 ;
  assign n10825 = ~n10800 & n10822 ;
  assign n10826 = n10824 | n10825 ;
  assign n10827 = n10472 | n10477 ;
  assign n10828 = n10826 & n10827 ;
  assign n10829 = n10826 | n10827 ;
  assign n10830 = ~n10828 & n10829 ;
  assign n10831 = n10793 | n10797 ;
  assign n10832 = n10774 | n10779 ;
  assign n10833 = n10755 | n10760 ;
  assign n10834 = n10737 | n10741 ;
  assign n10835 = x95 & n2775 ;
  assign n10836 = x94 & n2770 ;
  assign n10837 = x93 & ~n2769 ;
  assign n10838 = n2978 & n10837 ;
  assign n10839 = n10836 | n10838 ;
  assign n10840 = n10835 | n10839 ;
  assign n10841 = n2778 | n10840 ;
  assign n10842 = ( n3479 & n10840 ) | ( n3479 & n10841 ) | ( n10840 & n10841 ) ;
  assign n10843 = x29 & n10842 ;
  assign n10844 = x29 & ~n10843 ;
  assign n10845 = ( n10842 & ~n10843 ) | ( n10842 & n10844 ) | ( ~n10843 & n10844 ) ;
  assign n10846 = x92 & n3314 ;
  assign n10847 = x91 & n3309 ;
  assign n10848 = x90 & ~n3308 ;
  assign n10849 = n3570 & n10848 ;
  assign n10850 = n10847 | n10849 ;
  assign n10851 = n10846 | n10850 ;
  assign n10852 = n3317 | n10851 ;
  assign n10853 = ( n2904 & n10851 ) | ( n2904 & n10852 ) | ( n10851 & n10852 ) ;
  assign n10854 = x32 & n10853 ;
  assign n10855 = x32 & ~n10854 ;
  assign n10856 = ( n10853 & ~n10854 ) | ( n10853 & n10855 ) | ( ~n10854 & n10855 ) ;
  assign n10857 = x71 & n8834 ;
  assign n10858 = x70 & n8829 ;
  assign n10859 = x69 & ~n8828 ;
  assign n10860 = n9159 & n10859 ;
  assign n10861 = n10858 | n10860 ;
  assign n10862 = n10857 | n10861 ;
  assign n10863 = n8837 | n10862 ;
  assign n10864 = ( n376 & n10862 ) | ( n376 & n10863 ) | ( n10862 & n10863 ) ;
  assign n10865 = x53 & ~n10864 ;
  assign n10866 = ~x53 & n10864 ;
  assign n10867 = n10865 | n10866 ;
  assign n10868 = ~x57 & x58 ;
  assign n10869 = x57 & ~x58 ;
  assign n10870 = n10868 | n10869 ;
  assign n10871 = ~n10533 & n10870 ;
  assign n10872 = x64 & n10871 ;
  assign n10873 = ~x58 & x59 ;
  assign n10874 = x58 & ~x59 ;
  assign n10875 = n10873 | n10874 ;
  assign n10876 = n10533 & ~n10875 ;
  assign n10877 = x65 & n10876 ;
  assign n10878 = n10872 | n10877 ;
  assign n10879 = n10533 & n10875 ;
  assign n10880 = n142 & n10879 ;
  assign n10881 = n10878 | n10880 ;
  assign n10882 = x59 | n10881 ;
  assign n10883 = ~x59 & n10882 ;
  assign n10884 = ( ~n10881 & n10882 ) | ( ~n10881 & n10883 ) | ( n10882 & n10883 ) ;
  assign n10885 = x59 & ~n10534 ;
  assign n10886 = n10884 & n10885 ;
  assign n10887 = n10884 | n10885 ;
  assign n10888 = ~n10886 & n10887 ;
  assign n10889 = n229 & n9856 ;
  assign n10890 = x68 & n9853 ;
  assign n10891 = x67 & n9848 ;
  assign n10892 = x66 & ~n9847 ;
  assign n10893 = n10165 & n10892 ;
  assign n10894 = n10891 | n10893 ;
  assign n10895 = n10890 | n10894 ;
  assign n10896 = n10889 | n10895 ;
  assign n10897 = x56 | n10896 ;
  assign n10898 = ~x56 & n10897 ;
  assign n10899 = ( ~n10896 & n10897 ) | ( ~n10896 & n10898 ) | ( n10897 & n10898 ) ;
  assign n10900 = n10888 | n10899 ;
  assign n10901 = n10888 & n10899 ;
  assign n10902 = n10900 & ~n10901 ;
  assign n10903 = n10546 | n10902 ;
  assign n10904 = n10546 & n10902 ;
  assign n10905 = n10903 & ~n10904 ;
  assign n10906 = n10867 | n10905 ;
  assign n10907 = n10867 & n10905 ;
  assign n10908 = n10906 & ~n10907 ;
  assign n10909 = ( n10179 & n10530 ) | ( n10179 & n10548 ) | ( n10530 & n10548 ) ;
  assign n10910 = n10908 | n10909 ;
  assign n10911 = n10908 & n10909 ;
  assign n10912 = n10910 & ~n10911 ;
  assign n10913 = x74 & n7812 ;
  assign n10914 = x73 & n7807 ;
  assign n10915 = x72 & ~n7806 ;
  assign n10916 = n8136 & n10915 ;
  assign n10917 = n10914 | n10916 ;
  assign n10918 = n10913 | n10917 ;
  assign n10919 = n7815 | n10918 ;
  assign n10920 = ( n587 & n10918 ) | ( n587 & n10919 ) | ( n10918 & n10919 ) ;
  assign n10921 = x50 & n10920 ;
  assign n10922 = x50 & ~n10921 ;
  assign n10923 = ( n10920 & ~n10921 ) | ( n10920 & n10922 ) | ( ~n10921 & n10922 ) ;
  assign n10924 = n10912 & n10923 ;
  assign n10925 = n10912 & ~n10924 ;
  assign n10926 = ~n10912 & n10923 ;
  assign n10927 = n10925 | n10926 ;
  assign n10928 = n10563 | n10566 ;
  assign n10929 = n10927 | n10928 ;
  assign n10930 = n10927 & n10928 ;
  assign n10931 = n10929 & ~n10930 ;
  assign n10932 = x77 & n6937 ;
  assign n10933 = x76 & n6932 ;
  assign n10934 = x75 & ~n6931 ;
  assign n10935 = n7216 & n10934 ;
  assign n10936 = n10933 | n10935 ;
  assign n10937 = n10932 | n10936 ;
  assign n10938 = n6940 | n10937 ;
  assign n10939 = ( n846 & n10937 ) | ( n846 & n10938 ) | ( n10937 & n10938 ) ;
  assign n10940 = x47 & n10939 ;
  assign n10941 = x47 & ~n10940 ;
  assign n10942 = ( n10939 & ~n10940 ) | ( n10939 & n10941 ) | ( ~n10940 & n10941 ) ;
  assign n10943 = n10931 & n10942 ;
  assign n10944 = n10931 | n10942 ;
  assign n10945 = ~n10943 & n10944 ;
  assign n10946 = n10581 | n10584 ;
  assign n10947 = n10945 & n10946 ;
  assign n10948 = n10946 & ~n10947 ;
  assign n10949 = ( n10945 & ~n10947 ) | ( n10945 & n10948 ) | ( ~n10947 & n10948 ) ;
  assign n10950 = x80 & n6068 ;
  assign n10951 = x79 & n6063 ;
  assign n10952 = x78 & ~n6062 ;
  assign n10953 = n6398 & n10952 ;
  assign n10954 = n10951 | n10953 ;
  assign n10955 = n10950 | n10954 ;
  assign n10956 = n6071 | n10955 ;
  assign n10957 = ( n1147 & n10955 ) | ( n1147 & n10956 ) | ( n10955 & n10956 ) ;
  assign n10958 = x44 & n10957 ;
  assign n10959 = x44 & ~n10958 ;
  assign n10960 = ( n10957 & ~n10958 ) | ( n10957 & n10959 ) | ( ~n10958 & n10959 ) ;
  assign n10961 = n10949 & n10960 ;
  assign n10962 = n10949 & ~n10961 ;
  assign n10963 = ~n10949 & n10960 ;
  assign n10964 = n10962 | n10963 ;
  assign n10965 = n10598 | n10603 ;
  assign n10966 = n10964 | n10965 ;
  assign n10967 = n10964 & n10965 ;
  assign n10968 = n10966 & ~n10967 ;
  assign n10969 = x83 & n5340 ;
  assign n10970 = x82 & n5335 ;
  assign n10971 = x81 & ~n5334 ;
  assign n10972 = n5580 & n10971 ;
  assign n10973 = n10970 | n10972 ;
  assign n10974 = n10969 | n10973 ;
  assign n10975 = n5343 | n10974 ;
  assign n10976 = ( n1510 & n10974 ) | ( n1510 & n10975 ) | ( n10974 & n10975 ) ;
  assign n10977 = x41 & n10976 ;
  assign n10978 = x41 & ~n10977 ;
  assign n10979 = ( n10976 & ~n10977 ) | ( n10976 & n10978 ) | ( ~n10977 & n10978 ) ;
  assign n10980 = n10968 & n10979 ;
  assign n10981 = n10968 | n10979 ;
  assign n10982 = ~n10980 & n10981 ;
  assign n10983 = n10616 & n10982 ;
  assign n10984 = n10616 & ~n10983 ;
  assign n10985 = ( n10982 & ~n10983 ) | ( n10982 & n10984 ) | ( ~n10983 & n10984 ) ;
  assign n10986 = x86 & n4572 ;
  assign n10987 = x85 & n4567 ;
  assign n10988 = x84 & ~n4566 ;
  assign n10989 = n4828 & n10988 ;
  assign n10990 = n10987 | n10989 ;
  assign n10991 = n10986 | n10990 ;
  assign n10992 = n4575 | n10991 ;
  assign n10993 = ( n1921 & n10991 ) | ( n1921 & n10992 ) | ( n10991 & n10992 ) ;
  assign n10994 = x38 & n10993 ;
  assign n10995 = x38 & ~n10994 ;
  assign n10996 = ( n10993 & ~n10994 ) | ( n10993 & n10995 ) | ( ~n10994 & n10995 ) ;
  assign n10997 = n10985 & n10996 ;
  assign n10998 = n10985 & ~n10997 ;
  assign n10999 = ~n10985 & n10996 ;
  assign n11000 = n10998 | n10999 ;
  assign n11001 = n10619 | n10624 ;
  assign n11002 = n11000 | n11001 ;
  assign n11003 = n11000 & n11001 ;
  assign n11004 = n11002 & ~n11003 ;
  assign n11005 = x89 & n3913 ;
  assign n11006 = x88 & n3908 ;
  assign n11007 = x87 & ~n3907 ;
  assign n11008 = n4152 & n11007 ;
  assign n11009 = n11006 | n11008 ;
  assign n11010 = n11005 | n11009 ;
  assign n11011 = n3916 | n11010 ;
  assign n11012 = ( n2244 & n11010 ) | ( n2244 & n11011 ) | ( n11010 & n11011 ) ;
  assign n11013 = x35 & n11012 ;
  assign n11014 = x35 & ~n11013 ;
  assign n11015 = ( n11012 & ~n11013 ) | ( n11012 & n11014 ) | ( ~n11013 & n11014 ) ;
  assign n11016 = n11004 & n11015 ;
  assign n11017 = n11004 & ~n11016 ;
  assign n11018 = ~n11004 & n11015 ;
  assign n11019 = n11017 | n11018 ;
  assign n11020 = n10637 | n10643 ;
  assign n11021 = n11019 | n11020 ;
  assign n11022 = n11019 & n11020 ;
  assign n11023 = n11021 & ~n11022 ;
  assign n11024 = n10657 | n10659 ;
  assign n11025 = ( n10856 & n11023 ) | ( n10856 & n11024 ) | ( n11023 & n11024 ) ;
  assign n11026 = ( n11023 & n11024 ) | ( n11023 & ~n11025 ) | ( n11024 & ~n11025 ) ;
  assign n11027 = ( n10856 & ~n11025 ) | ( n10856 & n11026 ) | ( ~n11025 & n11026 ) ;
  assign n11028 = n10845 & n11027 ;
  assign n11029 = n10845 | n11027 ;
  assign n11030 = ~n11028 & n11029 ;
  assign n11031 = n10673 | n10677 ;
  assign n11032 = n11030 | n11031 ;
  assign n11033 = n11030 & n11031 ;
  assign n11034 = n11032 & ~n11033 ;
  assign n11035 = x98 & n2280 ;
  assign n11036 = x97 & n2275 ;
  assign n11037 = x96 & ~n2274 ;
  assign n11038 = n2481 & n11037 ;
  assign n11039 = n11036 | n11038 ;
  assign n11040 = n11035 | n11039 ;
  assign n11041 = n2283 | n11040 ;
  assign n11042 = ( n4105 & n11040 ) | ( n4105 & n11041 ) | ( n11040 & n11041 ) ;
  assign n11043 = x26 & n11042 ;
  assign n11044 = x26 & ~n11043 ;
  assign n11045 = ( n11042 & ~n11043 ) | ( n11042 & n11044 ) | ( ~n11043 & n11044 ) ;
  assign n11046 = n11034 & n11045 ;
  assign n11047 = n11034 & ~n11046 ;
  assign n11048 = ~n11034 & n11045 ;
  assign n11049 = n11047 | n11048 ;
  assign n11050 = ( n10504 & n10505 ) | ( n10504 & n10679 ) | ( n10505 & n10679 ) ;
  assign n11051 = n11049 | n11050 ;
  assign n11052 = n11049 & n11050 ;
  assign n11053 = n11051 & ~n11052 ;
  assign n11054 = x101 & n1817 ;
  assign n11055 = x100 & n1812 ;
  assign n11056 = x99 & ~n1811 ;
  assign n11057 = n1977 & n11056 ;
  assign n11058 = n11055 | n11057 ;
  assign n11059 = n11054 | n11058 ;
  assign n11060 = n1820 | n11059 ;
  assign n11061 = ( n4783 & n11059 ) | ( n4783 & n11060 ) | ( n11059 & n11060 ) ;
  assign n11062 = x23 & n11061 ;
  assign n11063 = x23 & ~n11062 ;
  assign n11064 = ( n11061 & ~n11062 ) | ( n11061 & n11063 ) | ( ~n11062 & n11063 ) ;
  assign n11065 = n11053 & n11064 ;
  assign n11066 = n11053 & ~n11065 ;
  assign n11067 = ~n11053 & n11064 ;
  assign n11068 = n11066 | n11067 ;
  assign n11069 = n10683 | n10687 ;
  assign n11070 = n11068 | n11069 ;
  assign n11071 = n11068 & n11069 ;
  assign n11072 = n11070 & ~n11071 ;
  assign n11073 = x104 & n1421 ;
  assign n11074 = x103 & n1416 ;
  assign n11075 = x102 & ~n1415 ;
  assign n11076 = n1584 & n11075 ;
  assign n11077 = n11074 | n11076 ;
  assign n11078 = n11073 | n11077 ;
  assign n11079 = n1424 | n11078 ;
  assign n11080 = ( n5295 & n11078 ) | ( n5295 & n11079 ) | ( n11078 & n11079 ) ;
  assign n11081 = x20 & n11080 ;
  assign n11082 = x20 & ~n11081 ;
  assign n11083 = ( n11080 & ~n11081 ) | ( n11080 & n11082 ) | ( ~n11081 & n11082 ) ;
  assign n11084 = n11072 & n11083 ;
  assign n11085 = n11072 & ~n11084 ;
  assign n11086 = ~n11072 & n11083 ;
  assign n11087 = n11085 | n11086 ;
  assign n11088 = n10700 | n10706 ;
  assign n11089 = n11087 | n11088 ;
  assign n11090 = n11087 & n11088 ;
  assign n11091 = n11089 & ~n11090 ;
  assign n11092 = x107 & n1071 ;
  assign n11093 = x106 & n1066 ;
  assign n11094 = x105 & ~n1065 ;
  assign n11095 = n1189 & n11094 ;
  assign n11096 = n11093 | n11095 ;
  assign n11097 = n11092 | n11096 ;
  assign n11098 = n1074 | n11097 ;
  assign n11099 = ( n6328 & n11097 ) | ( n6328 & n11098 ) | ( n11097 & n11098 ) ;
  assign n11100 = x17 & n11099 ;
  assign n11101 = x17 & ~n11100 ;
  assign n11102 = ( n11099 & ~n11100 ) | ( n11099 & n11101 ) | ( ~n11100 & n11101 ) ;
  assign n11103 = n11091 & n11102 ;
  assign n11104 = n11091 | n11102 ;
  assign n11105 = ~n11103 & n11104 ;
  assign n11106 = n10720 | n10723 ;
  assign n11107 = n11105 & n11106 ;
  assign n11108 = n11106 & ~n11107 ;
  assign n11109 = ( n11105 & ~n11107 ) | ( n11105 & n11108 ) | ( ~n11107 & n11108 ) ;
  assign n11110 = x110 & n771 ;
  assign n11111 = x109 & n766 ;
  assign n11112 = x108 & ~n765 ;
  assign n11113 = n905 & n11112 ;
  assign n11114 = n11111 | n11113 ;
  assign n11115 = n11110 | n11114 ;
  assign n11116 = n774 | n11115 ;
  assign n11117 = ( n7189 & n11115 ) | ( n7189 & n11116 ) | ( n11115 & n11116 ) ;
  assign n11118 = x14 & n11117 ;
  assign n11119 = x14 & ~n11118 ;
  assign n11120 = ( n11117 & ~n11118 ) | ( n11117 & n11119 ) | ( ~n11118 & n11119 ) ;
  assign n11121 = n11109 | n11120 ;
  assign n11122 = n11109 & n11120 ;
  assign n11123 = n11121 & ~n11122 ;
  assign n11124 = n10834 & n11123 ;
  assign n11125 = n10834 | n11123 ;
  assign n11126 = ~n11124 & n11125 ;
  assign n11127 = x113 & n528 ;
  assign n11128 = x112 & n523 ;
  assign n11129 = x111 & ~n522 ;
  assign n11130 = n635 & n11129 ;
  assign n11131 = n11128 | n11130 ;
  assign n11132 = n11127 | n11131 ;
  assign n11133 = n531 | n11132 ;
  assign n11134 = ( n8113 & n11132 ) | ( n8113 & n11133 ) | ( n11132 & n11133 ) ;
  assign n11135 = x11 & n11134 ;
  assign n11136 = x11 & ~n11135 ;
  assign n11137 = ( n11134 & ~n11135 ) | ( n11134 & n11136 ) | ( ~n11135 & n11136 ) ;
  assign n11138 = n11126 | n11137 ;
  assign n11139 = n11126 & n11137 ;
  assign n11140 = n11138 & ~n11139 ;
  assign n11141 = n10833 & n11140 ;
  assign n11142 = n10833 | n11140 ;
  assign n11143 = ~n11141 & n11142 ;
  assign n11144 = x116 & n337 ;
  assign n11145 = x115 & n332 ;
  assign n11146 = x114 & ~n331 ;
  assign n11147 = n396 & n11146 ;
  assign n11148 = n11145 | n11147 ;
  assign n11149 = n11144 | n11148 ;
  assign n11150 = n340 | n11149 ;
  assign n11151 = ( n8778 & n11149 ) | ( n8778 & n11150 ) | ( n11149 & n11150 ) ;
  assign n11152 = x8 & n11151 ;
  assign n11153 = x8 & ~n11152 ;
  assign n11154 = ( n11151 & ~n11152 ) | ( n11151 & n11153 ) | ( ~n11152 & n11153 ) ;
  assign n11155 = n11143 | n11154 ;
  assign n11156 = n11143 & n11154 ;
  assign n11157 = n11155 & ~n11156 ;
  assign n11158 = n10832 & n11157 ;
  assign n11159 = n10832 | n11157 ;
  assign n11160 = ~n11158 & n11159 ;
  assign n11161 = x119 & n206 ;
  assign n11162 = x118 & n201 ;
  assign n11163 = x117 & ~n200 ;
  assign n11164 = n243 & n11163 ;
  assign n11165 = n11162 | n11164 ;
  assign n11166 = n11161 | n11165 ;
  assign n11167 = n209 | n11166 ;
  assign n11168 = ( n9789 & n11166 ) | ( n9789 & n11167 ) | ( n11166 & n11167 ) ;
  assign n11169 = x5 & n11168 ;
  assign n11170 = x5 & ~n11169 ;
  assign n11171 = ( n11168 & ~n11169 ) | ( n11168 & n11170 ) | ( ~n11169 & n11170 ) ;
  assign n11172 = n11160 | n11171 ;
  assign n11173 = n11160 & n11171 ;
  assign n11174 = n11172 & ~n11173 ;
  assign n11175 = n10831 & n11174 ;
  assign n11176 = n10831 | n11174 ;
  assign n11177 = ~n11175 & n11176 ;
  assign n11178 = x121 | x122 ;
  assign n11179 = x121 & x122 ;
  assign n11180 = n11178 & ~n11179 ;
  assign n11181 = n10802 | n10805 ;
  assign n11182 = n11180 & n11181 ;
  assign n11183 = n10802 | n10807 ;
  assign n11184 = n11180 & n11183 ;
  assign n11185 = ( n9786 & n11182 ) | ( n9786 & n11184 ) | ( n11182 & n11184 ) ;
  assign n11186 = ( n9786 & n11181 ) | ( n9786 & n11183 ) | ( n11181 & n11183 ) ;
  assign n11187 = n11180 | n11186 ;
  assign n11188 = ~n11185 & n11187 ;
  assign n11189 = x121 & n131 ;
  assign n11190 = x120 & ~n156 ;
  assign n11191 = ( n135 & n11189 ) | ( n135 & n11190 ) | ( n11189 & n11190 ) ;
  assign n11192 = x0 & x122 ;
  assign n11193 = ( ~n135 & n11189 ) | ( ~n135 & n11192 ) | ( n11189 & n11192 ) ;
  assign n11194 = n11191 | n11193 ;
  assign n11195 = n139 | n11194 ;
  assign n11196 = ( n11188 & n11194 ) | ( n11188 & n11195 ) | ( n11194 & n11195 ) ;
  assign n11197 = x2 & n11196 ;
  assign n11198 = x2 & ~n11197 ;
  assign n11199 = ( n11196 & ~n11197 ) | ( n11196 & n11198 ) | ( ~n11197 & n11198 ) ;
  assign n11200 = n11177 & n11199 ;
  assign n11201 = n11177 & ~n11200 ;
  assign n11202 = ~n11177 & n11199 ;
  assign n11203 = n11201 | n11202 ;
  assign n11204 = n10823 | n10828 ;
  assign n11205 = n11203 & n11204 ;
  assign n11206 = n11203 | n11204 ;
  assign n11207 = ~n11205 & n11206 ;
  assign n11208 = n11200 | n11205 ;
  assign n11209 = x122 | x123 ;
  assign n11210 = x122 & x123 ;
  assign n11211 = n11209 & ~n11210 ;
  assign n11212 = n11179 | n11182 ;
  assign n11213 = n11211 & n11212 ;
  assign n11214 = n11179 | n11184 ;
  assign n11215 = n11211 & n11214 ;
  assign n11216 = ( n9786 & n11213 ) | ( n9786 & n11215 ) | ( n11213 & n11215 ) ;
  assign n11217 = ( n9786 & n11212 ) | ( n9786 & n11214 ) | ( n11212 & n11214 ) ;
  assign n11218 = n11211 | n11217 ;
  assign n11219 = ~n11216 & n11218 ;
  assign n11220 = x122 & n131 ;
  assign n11221 = x121 & ~n156 ;
  assign n11222 = ( n135 & n11220 ) | ( n135 & n11221 ) | ( n11220 & n11221 ) ;
  assign n11223 = x0 & x123 ;
  assign n11224 = ( ~n135 & n11220 ) | ( ~n135 & n11223 ) | ( n11220 & n11223 ) ;
  assign n11225 = n11222 | n11224 ;
  assign n11226 = n139 | n11225 ;
  assign n11227 = ( n11219 & n11225 ) | ( n11219 & n11226 ) | ( n11225 & n11226 ) ;
  assign n11228 = x2 & n11227 ;
  assign n11229 = x2 & ~n11228 ;
  assign n11230 = ( n11227 & ~n11228 ) | ( n11227 & n11229 ) | ( ~n11228 & n11229 ) ;
  assign n11231 = n11156 | n11158 ;
  assign n11232 = x111 & n771 ;
  assign n11233 = x110 & n766 ;
  assign n11234 = x109 & ~n765 ;
  assign n11235 = n905 & n11234 ;
  assign n11236 = n11233 | n11235 ;
  assign n11237 = n11232 | n11236 ;
  assign n11238 = n774 | n11237 ;
  assign n11239 = ( n7492 & n11237 ) | ( n7492 & n11238 ) | ( n11237 & n11238 ) ;
  assign n11240 = x14 & n11239 ;
  assign n11241 = x14 & ~n11240 ;
  assign n11242 = ( n11239 & ~n11240 ) | ( n11239 & n11241 ) | ( ~n11240 & n11241 ) ;
  assign n11243 = x108 & n1071 ;
  assign n11244 = x107 & n1066 ;
  assign n11245 = x106 & ~n1065 ;
  assign n11246 = n1189 & n11245 ;
  assign n11247 = n11244 | n11246 ;
  assign n11248 = n11243 | n11247 ;
  assign n11249 = n1074 | n11248 ;
  assign n11250 = ( n6358 & n11248 ) | ( n6358 & n11249 ) | ( n11248 & n11249 ) ;
  assign n11251 = x17 & n11250 ;
  assign n11252 = x17 & ~n11251 ;
  assign n11253 = ( n11250 & ~n11251 ) | ( n11250 & n11252 ) | ( ~n11251 & n11252 ) ;
  assign n11254 = n11103 | n11107 ;
  assign n11255 = n11028 | n11033 ;
  assign n11256 = x87 & n4572 ;
  assign n11257 = x86 & n4567 ;
  assign n11258 = x85 & ~n4566 ;
  assign n11259 = n4828 & n11258 ;
  assign n11260 = n11257 | n11259 ;
  assign n11261 = n11256 | n11260 ;
  assign n11262 = n4575 | n11261 ;
  assign n11263 = ( n2067 & n11261 ) | ( n2067 & n11262 ) | ( n11261 & n11262 ) ;
  assign n11264 = x38 & n11263 ;
  assign n11265 = x38 & ~n11264 ;
  assign n11266 = ( n11263 & ~n11264 ) | ( n11263 & n11265 ) | ( ~n11264 & n11265 ) ;
  assign n11267 = x84 & n5340 ;
  assign n11268 = x83 & n5335 ;
  assign n11269 = x82 & ~n5334 ;
  assign n11270 = n5580 & n11269 ;
  assign n11271 = n11268 | n11270 ;
  assign n11272 = n11267 | n11271 ;
  assign n11273 = n5343 | n11272 ;
  assign n11274 = ( n1537 & n11272 ) | ( n1537 & n11273 ) | ( n11272 & n11273 ) ;
  assign n11275 = x41 & n11274 ;
  assign n11276 = x41 & ~n11275 ;
  assign n11277 = ( n11274 & ~n11275 ) | ( n11274 & n11276 ) | ( ~n11275 & n11276 ) ;
  assign n11278 = n10980 | n10983 ;
  assign n11279 = n10961 | n10967 ;
  assign n11280 = n10943 | n10947 ;
  assign n11281 = x72 & n8834 ;
  assign n11282 = x71 & n8829 ;
  assign n11283 = x70 & ~n8828 ;
  assign n11284 = n9159 & n11283 ;
  assign n11285 = n11282 | n11284 ;
  assign n11286 = n11281 | n11285 ;
  assign n11287 = ( n435 & n8837 ) | ( n435 & n11286 ) | ( n8837 & n11286 ) ;
  assign n11288 = ( x53 & ~n11286 ) | ( x53 & n11287 ) | ( ~n11286 & n11287 ) ;
  assign n11289 = ~n11287 & n11288 ;
  assign n11290 = n11286 | n11288 ;
  assign n11291 = ( ~x53 & n11289 ) | ( ~x53 & n11290 ) | ( n11289 & n11290 ) ;
  assign n11292 = n264 & n9856 ;
  assign n11293 = x69 & n9853 ;
  assign n11294 = x68 & n9848 ;
  assign n11295 = x67 & ~n9847 ;
  assign n11296 = n10165 & n11295 ;
  assign n11297 = n11294 | n11296 ;
  assign n11298 = n11293 | n11297 ;
  assign n11299 = n11292 | n11298 ;
  assign n11300 = x56 | n11299 ;
  assign n11301 = ~x56 & n11300 ;
  assign n11302 = ( ~n11299 & n11300 ) | ( ~n11299 & n11301 ) | ( n11300 & n11301 ) ;
  assign n11303 = x66 & n10876 ;
  assign n11304 = x65 & n10871 ;
  assign n11305 = ~n10533 & n10875 ;
  assign n11306 = x64 & ~n10870 ;
  assign n11307 = n11305 & n11306 ;
  assign n11308 = n11304 | n11307 ;
  assign n11309 = n11303 | n11308 ;
  assign n11310 = n153 & n10879 ;
  assign n11311 = n11309 | n11310 ;
  assign n11312 = x59 | n11311 ;
  assign n11313 = ~x59 & n11312 ;
  assign n11314 = ( ~n11311 & n11312 ) | ( ~n11311 & n11313 ) | ( n11312 & n11313 ) ;
  assign n11315 = n10886 | n11314 ;
  assign n11316 = n10886 & n11314 ;
  assign n11317 = n11315 & ~n11316 ;
  assign n11318 = n10901 | n10904 ;
  assign n11319 = ( n11302 & n11317 ) | ( n11302 & n11318 ) | ( n11317 & n11318 ) ;
  assign n11320 = ( n11317 & n11318 ) | ( n11317 & ~n11319 ) | ( n11318 & ~n11319 ) ;
  assign n11321 = ( n11302 & ~n11319 ) | ( n11302 & n11320 ) | ( ~n11319 & n11320 ) ;
  assign n11322 = n11291 | n11321 ;
  assign n11323 = n11291 & n11321 ;
  assign n11324 = n11322 & ~n11323 ;
  assign n11325 = n10907 | n10911 ;
  assign n11326 = n11324 & n11325 ;
  assign n11327 = n11324 | n11325 ;
  assign n11328 = ~n11326 & n11327 ;
  assign n11329 = x75 & n7812 ;
  assign n11330 = x74 & n7807 ;
  assign n11331 = x73 & ~n7806 ;
  assign n11332 = n8136 & n11331 ;
  assign n11333 = n11330 | n11332 ;
  assign n11334 = n11329 | n11333 ;
  assign n11335 = n7815 | n11334 ;
  assign n11336 = ( n609 & n11334 ) | ( n609 & n11335 ) | ( n11334 & n11335 ) ;
  assign n11337 = x50 & n11336 ;
  assign n11338 = x50 & ~n11337 ;
  assign n11339 = ( n11336 & ~n11337 ) | ( n11336 & n11338 ) | ( ~n11337 & n11338 ) ;
  assign n11340 = n11328 | n11339 ;
  assign n11341 = n11328 & n11339 ;
  assign n11342 = n11340 & ~n11341 ;
  assign n11343 = n10924 | n10930 ;
  assign n11344 = n11342 & n11343 ;
  assign n11345 = n11342 | n11343 ;
  assign n11346 = ~n11344 & n11345 ;
  assign n11347 = x78 & n6937 ;
  assign n11348 = x77 & n6932 ;
  assign n11349 = x76 & ~n6931 ;
  assign n11350 = n7216 & n11349 ;
  assign n11351 = n11348 | n11350 ;
  assign n11352 = n11347 | n11351 ;
  assign n11353 = n6940 | n11352 ;
  assign n11354 = ( n868 & n11352 ) | ( n868 & n11353 ) | ( n11352 & n11353 ) ;
  assign n11355 = x47 & n11354 ;
  assign n11356 = x47 & ~n11355 ;
  assign n11357 = ( n11354 & ~n11355 ) | ( n11354 & n11356 ) | ( ~n11355 & n11356 ) ;
  assign n11358 = n11346 & n11357 ;
  assign n11359 = n11346 & ~n11358 ;
  assign n11360 = ~n11346 & n11357 ;
  assign n11361 = n11359 | n11360 ;
  assign n11362 = n11280 & n11361 ;
  assign n11363 = n11280 | n11361 ;
  assign n11364 = ~n11362 & n11363 ;
  assign n11365 = x81 & n6068 ;
  assign n11366 = x80 & n6063 ;
  assign n11367 = x79 & ~n6062 ;
  assign n11368 = n6398 & n11367 ;
  assign n11369 = n11366 | n11368 ;
  assign n11370 = n11365 | n11369 ;
  assign n11371 = n6071 | n11370 ;
  assign n11372 = ( n1256 & n11370 ) | ( n1256 & n11371 ) | ( n11370 & n11371 ) ;
  assign n11373 = x44 & n11372 ;
  assign n11374 = x44 & ~n11373 ;
  assign n11375 = ( n11372 & ~n11373 ) | ( n11372 & n11374 ) | ( ~n11373 & n11374 ) ;
  assign n11376 = n11364 & n11375 ;
  assign n11377 = n11364 & ~n11376 ;
  assign n11378 = ~n11364 & n11375 ;
  assign n11379 = n11377 | n11378 ;
  assign n11380 = n11279 & n11379 ;
  assign n11381 = n11279 & ~n11380 ;
  assign n11382 = n11379 & ~n11380 ;
  assign n11383 = n11381 | n11382 ;
  assign n11384 = ( n11277 & n11278 ) | ( n11277 & ~n11383 ) | ( n11278 & ~n11383 ) ;
  assign n11385 = ( ~n11278 & n11383 ) | ( ~n11278 & n11384 ) | ( n11383 & n11384 ) ;
  assign n11386 = ( ~n11277 & n11384 ) | ( ~n11277 & n11385 ) | ( n11384 & n11385 ) ;
  assign n11387 = n11266 & n11386 ;
  assign n11388 = n11266 | n11386 ;
  assign n11389 = ~n11387 & n11388 ;
  assign n11390 = n10997 | n11003 ;
  assign n11391 = n11389 | n11390 ;
  assign n11392 = n11389 & n11390 ;
  assign n11393 = n11391 & ~n11392 ;
  assign n11394 = x90 & n3913 ;
  assign n11395 = x89 & n3908 ;
  assign n11396 = x88 & ~n3907 ;
  assign n11397 = n4152 & n11396 ;
  assign n11398 = n11395 | n11397 ;
  assign n11399 = n11394 | n11398 ;
  assign n11400 = n3916 | n11399 ;
  assign n11401 = ( n2410 & n11399 ) | ( n2410 & n11400 ) | ( n11399 & n11400 ) ;
  assign n11402 = x35 & n11401 ;
  assign n11403 = x35 & ~n11402 ;
  assign n11404 = ( n11401 & ~n11402 ) | ( n11401 & n11403 ) | ( ~n11402 & n11403 ) ;
  assign n11405 = n11393 & n11404 ;
  assign n11406 = n11393 & ~n11405 ;
  assign n11407 = ~n11393 & n11404 ;
  assign n11408 = n11406 | n11407 ;
  assign n11409 = n11016 | n11022 ;
  assign n11410 = n11408 | n11409 ;
  assign n11411 = n11408 & n11409 ;
  assign n11412 = n11410 & ~n11411 ;
  assign n11413 = x93 & n3314 ;
  assign n11414 = x92 & n3309 ;
  assign n11415 = x91 & ~n3308 ;
  assign n11416 = n3570 & n11415 ;
  assign n11417 = n11414 | n11416 ;
  assign n11418 = n11413 | n11417 ;
  assign n11419 = n3317 | n11418 ;
  assign n11420 = ( n2931 & n11418 ) | ( n2931 & n11419 ) | ( n11418 & n11419 ) ;
  assign n11421 = x32 & n11420 ;
  assign n11422 = x32 & ~n11421 ;
  assign n11423 = ( n11420 & ~n11421 ) | ( n11420 & n11422 ) | ( ~n11421 & n11422 ) ;
  assign n11424 = n11412 & n11423 ;
  assign n11425 = n11412 | n11423 ;
  assign n11426 = ~n11424 & n11425 ;
  assign n11427 = n11025 & n11426 ;
  assign n11428 = n11025 & ~n11427 ;
  assign n11429 = ( n11426 & ~n11427 ) | ( n11426 & n11428 ) | ( ~n11427 & n11428 ) ;
  assign n11430 = x96 & n2775 ;
  assign n11431 = x95 & n2770 ;
  assign n11432 = x94 & ~n2769 ;
  assign n11433 = n2978 & n11432 ;
  assign n11434 = n11431 | n11433 ;
  assign n11435 = n11430 | n11434 ;
  assign n11436 = n2778 | n11435 ;
  assign n11437 = ( n3509 & n11435 ) | ( n3509 & n11436 ) | ( n11435 & n11436 ) ;
  assign n11438 = x29 & n11437 ;
  assign n11439 = x29 & ~n11438 ;
  assign n11440 = ( n11437 & ~n11438 ) | ( n11437 & n11439 ) | ( ~n11438 & n11439 ) ;
  assign n11441 = n11429 | n11440 ;
  assign n11442 = n11429 & n11440 ;
  assign n11443 = n11441 & ~n11442 ;
  assign n11444 = n11255 & n11443 ;
  assign n11445 = n11255 | n11443 ;
  assign n11446 = ~n11444 & n11445 ;
  assign n11447 = x99 & n2280 ;
  assign n11448 = x98 & n2275 ;
  assign n11449 = x97 & ~n2274 ;
  assign n11450 = n2481 & n11449 ;
  assign n11451 = n11448 | n11450 ;
  assign n11452 = n11447 | n11451 ;
  assign n11453 = n2283 | n11452 ;
  assign n11454 = ( n4325 & n11452 ) | ( n4325 & n11453 ) | ( n11452 & n11453 ) ;
  assign n11455 = x26 & n11454 ;
  assign n11456 = x26 & ~n11455 ;
  assign n11457 = ( n11454 & ~n11455 ) | ( n11454 & n11456 ) | ( ~n11455 & n11456 ) ;
  assign n11458 = n11446 & n11457 ;
  assign n11459 = n11446 & ~n11458 ;
  assign n11460 = ~n11446 & n11457 ;
  assign n11461 = n11459 | n11460 ;
  assign n11462 = n11046 | n11052 ;
  assign n11463 = n11461 | n11462 ;
  assign n11464 = n11461 & n11462 ;
  assign n11465 = n11463 & ~n11464 ;
  assign n11466 = x102 & n1817 ;
  assign n11467 = x101 & n1812 ;
  assign n11468 = x100 & ~n1811 ;
  assign n11469 = n1977 & n11468 ;
  assign n11470 = n11467 | n11469 ;
  assign n11471 = n11466 | n11470 ;
  assign n11472 = n1820 | n11471 ;
  assign n11473 = ( n5025 & n11471 ) | ( n5025 & n11472 ) | ( n11471 & n11472 ) ;
  assign n11474 = x23 & n11473 ;
  assign n11475 = x23 & ~n11474 ;
  assign n11476 = ( n11473 & ~n11474 ) | ( n11473 & n11475 ) | ( ~n11474 & n11475 ) ;
  assign n11477 = n11465 & n11476 ;
  assign n11478 = n11465 & ~n11477 ;
  assign n11479 = ~n11465 & n11476 ;
  assign n11480 = n11478 | n11479 ;
  assign n11481 = n11065 | n11071 ;
  assign n11482 = n11480 | n11481 ;
  assign n11483 = n11480 & n11481 ;
  assign n11484 = n11482 & ~n11483 ;
  assign n11485 = x105 & n1421 ;
  assign n11486 = x104 & n1416 ;
  assign n11487 = x103 & ~n1415 ;
  assign n11488 = n1584 & n11487 ;
  assign n11489 = n11486 | n11488 ;
  assign n11490 = n11485 | n11489 ;
  assign n11491 = n1424 | n11490 ;
  assign n11492 = ( n5788 & n11490 ) | ( n5788 & n11491 ) | ( n11490 & n11491 ) ;
  assign n11493 = x20 & n11492 ;
  assign n11494 = x20 & ~n11493 ;
  assign n11495 = ( n11492 & ~n11493 ) | ( n11492 & n11494 ) | ( ~n11493 & n11494 ) ;
  assign n11496 = n11484 & n11495 ;
  assign n11497 = n11484 | n11495 ;
  assign n11498 = ~n11496 & n11497 ;
  assign n11499 = n11084 | n11090 ;
  assign n11500 = n11498 | n11499 ;
  assign n11501 = ( n11084 & n11090 ) | ( n11084 & n11498 ) | ( n11090 & n11498 ) ;
  assign n11502 = n11500 & ~n11501 ;
  assign n11503 = ( n11253 & n11254 ) | ( n11253 & ~n11502 ) | ( n11254 & ~n11502 ) ;
  assign n11504 = ( ~n11254 & n11502 ) | ( ~n11254 & n11503 ) | ( n11502 & n11503 ) ;
  assign n11505 = ( ~n11253 & n11503 ) | ( ~n11253 & n11504 ) | ( n11503 & n11504 ) ;
  assign n11506 = n11242 & n11505 ;
  assign n11507 = n11242 | n11505 ;
  assign n11508 = ~n11506 & n11507 ;
  assign n11509 = n11122 | n11124 ;
  assign n11510 = n11508 & n11509 ;
  assign n11511 = n11508 | n11509 ;
  assign n11512 = ~n11510 & n11511 ;
  assign n11513 = x114 & n528 ;
  assign n11514 = x113 & n523 ;
  assign n11515 = x112 & ~n522 ;
  assign n11516 = n635 & n11515 ;
  assign n11517 = n11514 | n11516 ;
  assign n11518 = n11513 | n11517 ;
  assign n11519 = n531 | n11518 ;
  assign n11520 = ( n8437 & n11518 ) | ( n8437 & n11519 ) | ( n11518 & n11519 ) ;
  assign n11521 = x11 & n11520 ;
  assign n11522 = x11 & ~n11521 ;
  assign n11523 = ( n11520 & ~n11521 ) | ( n11520 & n11522 ) | ( ~n11521 & n11522 ) ;
  assign n11524 = n11512 & n11523 ;
  assign n11525 = n11512 & ~n11524 ;
  assign n11526 = ~n11512 & n11523 ;
  assign n11527 = n11525 | n11526 ;
  assign n11528 = n11139 | n11141 ;
  assign n11529 = n11527 & n11528 ;
  assign n11530 = n11527 | n11528 ;
  assign n11531 = ~n11529 & n11530 ;
  assign n11532 = x117 & n337 ;
  assign n11533 = x116 & n332 ;
  assign n11534 = x115 & ~n331 ;
  assign n11535 = n396 & n11534 ;
  assign n11536 = n11533 | n11535 ;
  assign n11537 = n11532 | n11536 ;
  assign n11538 = n340 | n11537 ;
  assign n11539 = ( n9118 & n11537 ) | ( n9118 & n11538 ) | ( n11537 & n11538 ) ;
  assign n11540 = x8 & n11539 ;
  assign n11541 = x8 & ~n11540 ;
  assign n11542 = ( n11539 & ~n11540 ) | ( n11539 & n11541 ) | ( ~n11540 & n11541 ) ;
  assign n11543 = n11531 & n11542 ;
  assign n11544 = n11531 & ~n11543 ;
  assign n11545 = ~n11531 & n11542 ;
  assign n11546 = n11544 | n11545 ;
  assign n11547 = n11231 & n11546 ;
  assign n11548 = n11231 & ~n11547 ;
  assign n11549 = n11546 & ~n11547 ;
  assign n11550 = n11548 | n11549 ;
  assign n11551 = x120 & n206 ;
  assign n11552 = x119 & n201 ;
  assign n11553 = x118 & ~n200 ;
  assign n11554 = n243 & n11553 ;
  assign n11555 = n11552 | n11554 ;
  assign n11556 = n11551 | n11555 ;
  assign n11557 = n209 | n11556 ;
  assign n11558 = ( n10460 & n11556 ) | ( n10460 & n11557 ) | ( n11556 & n11557 ) ;
  assign n11559 = x5 & n11558 ;
  assign n11560 = x5 & ~n11559 ;
  assign n11561 = ( n11558 & ~n11559 ) | ( n11558 & n11560 ) | ( ~n11559 & n11560 ) ;
  assign n11562 = ( n11230 & n11550 ) | ( n11230 & ~n11561 ) | ( n11550 & ~n11561 ) ;
  assign n11563 = ( ~n11550 & n11561 ) | ( ~n11550 & n11562 ) | ( n11561 & n11562 ) ;
  assign n11564 = ( ~n11230 & n11562 ) | ( ~n11230 & n11563 ) | ( n11562 & n11563 ) ;
  assign n11565 = n11173 | n11175 ;
  assign n11566 = n11564 & n11565 ;
  assign n11567 = n11565 & ~n11566 ;
  assign n11568 = ( n11564 & ~n11566 ) | ( n11564 & n11567 ) | ( ~n11566 & n11567 ) ;
  assign n11569 = n11208 & n11568 ;
  assign n11570 = n11208 | n11568 ;
  assign n11571 = ~n11569 & n11570 ;
  assign n11572 = n11543 | n11547 ;
  assign n11573 = n11524 | n11529 ;
  assign n11574 = n11506 | n11510 ;
  assign n11575 = n11496 | n11501 ;
  assign n11576 = n11458 | n11464 ;
  assign n11577 = x100 & n2280 ;
  assign n11578 = x99 & n2275 ;
  assign n11579 = x98 & ~n2274 ;
  assign n11580 = n2481 & n11579 ;
  assign n11581 = n11578 | n11580 ;
  assign n11582 = n11577 | n11581 ;
  assign n11583 = n2283 | n11582 ;
  assign n11584 = ( n4532 & n11582 ) | ( n4532 & n11583 ) | ( n11582 & n11583 ) ;
  assign n11585 = x26 & n11584 ;
  assign n11586 = x26 & ~n11585 ;
  assign n11587 = ( n11584 & ~n11585 ) | ( n11584 & n11586 ) | ( ~n11585 & n11586 ) ;
  assign n11588 = x97 & n2775 ;
  assign n11589 = x96 & n2770 ;
  assign n11590 = x95 & ~n2769 ;
  assign n11591 = n2978 & n11590 ;
  assign n11592 = n11589 | n11591 ;
  assign n11593 = n11588 | n11592 ;
  assign n11594 = n2778 | n11593 ;
  assign n11595 = ( n3707 & n11593 ) | ( n3707 & n11594 ) | ( n11593 & n11594 ) ;
  assign n11596 = x29 & n11595 ;
  assign n11597 = x29 & ~n11596 ;
  assign n11598 = ( n11595 & ~n11596 ) | ( n11595 & n11597 ) | ( ~n11596 & n11597 ) ;
  assign n11599 = n11442 | n11444 ;
  assign n11600 = n11424 | n11427 ;
  assign n11601 = x85 & n5340 ;
  assign n11602 = x84 & n5335 ;
  assign n11603 = x83 & ~n5334 ;
  assign n11604 = n5580 & n11603 ;
  assign n11605 = n11602 | n11604 ;
  assign n11606 = n11601 | n11605 ;
  assign n11607 = n5343 | n11606 ;
  assign n11608 = ( n1765 & n11606 ) | ( n1765 & n11607 ) | ( n11606 & n11607 ) ;
  assign n11609 = x41 & n11608 ;
  assign n11610 = x41 & ~n11609 ;
  assign n11611 = ( n11608 & ~n11609 ) | ( n11608 & n11610 ) | ( ~n11609 & n11610 ) ;
  assign n11612 = n11376 | n11380 ;
  assign n11613 = n11323 | n11326 ;
  assign n11614 = x70 & n9853 ;
  assign n11615 = x69 & n9848 ;
  assign n11616 = x68 & ~n9847 ;
  assign n11617 = n10165 & n11616 ;
  assign n11618 = n11615 | n11617 ;
  assign n11619 = n11614 | n11618 ;
  assign n11620 = n9856 | n11619 ;
  assign n11621 = ( n310 & n11619 ) | ( n310 & n11620 ) | ( n11619 & n11620 ) ;
  assign n11622 = x56 & ~n11621 ;
  assign n11623 = ~x56 & n11621 ;
  assign n11624 = n11622 | n11623 ;
  assign n11625 = x59 & ~x60 ;
  assign n11626 = ~x59 & x60 ;
  assign n11627 = n11625 | n11626 ;
  assign n11628 = x64 & n11627 ;
  assign n11629 = x67 & n10876 ;
  assign n11630 = x66 & n10871 ;
  assign n11631 = x65 & ~n10870 ;
  assign n11632 = n11305 & n11631 ;
  assign n11633 = n11630 | n11632 ;
  assign n11634 = n11629 | n11633 ;
  assign n11635 = n180 & n10879 ;
  assign n11636 = n11634 | n11635 ;
  assign n11637 = x59 & ~n11636 ;
  assign n11638 = ~x59 & n11636 ;
  assign n11639 = n11637 | n11638 ;
  assign n11640 = ( n11316 & n11628 ) | ( n11316 & n11639 ) | ( n11628 & n11639 ) ;
  assign n11641 = ( n11316 & n11639 ) | ( n11316 & ~n11640 ) | ( n11639 & ~n11640 ) ;
  assign n11642 = ( n11628 & ~n11640 ) | ( n11628 & n11641 ) | ( ~n11640 & n11641 ) ;
  assign n11643 = ( n11319 & n11624 ) | ( n11319 & ~n11642 ) | ( n11624 & ~n11642 ) ;
  assign n11644 = ( ~n11319 & n11642 ) | ( ~n11319 & n11643 ) | ( n11642 & n11643 ) ;
  assign n11645 = ( ~n11624 & n11643 ) | ( ~n11624 & n11644 ) | ( n11643 & n11644 ) ;
  assign n11646 = x73 & n8834 ;
  assign n11647 = x72 & n8829 ;
  assign n11648 = x71 & ~n8828 ;
  assign n11649 = n9159 & n11648 ;
  assign n11650 = n11647 | n11649 ;
  assign n11651 = n11646 | n11650 ;
  assign n11652 = ( n499 & n8837 ) | ( n499 & n11651 ) | ( n8837 & n11651 ) ;
  assign n11653 = ( x53 & ~n11651 ) | ( x53 & n11652 ) | ( ~n11651 & n11652 ) ;
  assign n11654 = ~n11652 & n11653 ;
  assign n11655 = n11651 | n11653 ;
  assign n11656 = ( ~x53 & n11654 ) | ( ~x53 & n11655 ) | ( n11654 & n11655 ) ;
  assign n11657 = n11645 & n11656 ;
  assign n11658 = n11645 | n11656 ;
  assign n11659 = ~n11657 & n11658 ;
  assign n11660 = n11613 & n11659 ;
  assign n11661 = n11613 | n11659 ;
  assign n11662 = ~n11660 & n11661 ;
  assign n11663 = x76 & n7812 ;
  assign n11664 = x75 & n7807 ;
  assign n11665 = x74 & ~n7806 ;
  assign n11666 = n8136 & n11665 ;
  assign n11667 = n11664 | n11666 ;
  assign n11668 = n11663 | n11667 ;
  assign n11669 = n7815 | n11668 ;
  assign n11670 = ( n740 & n11668 ) | ( n740 & n11669 ) | ( n11668 & n11669 ) ;
  assign n11671 = x50 & n11670 ;
  assign n11672 = x50 & ~n11671 ;
  assign n11673 = ( n11670 & ~n11671 ) | ( n11670 & n11672 ) | ( ~n11671 & n11672 ) ;
  assign n11674 = n11662 | n11673 ;
  assign n11675 = n11662 & n11673 ;
  assign n11676 = n11674 & ~n11675 ;
  assign n11677 = n11341 | n11344 ;
  assign n11678 = n11676 & n11677 ;
  assign n11679 = n11676 | n11677 ;
  assign n11680 = ~n11678 & n11679 ;
  assign n11681 = x79 & n6937 ;
  assign n11682 = x78 & n6932 ;
  assign n11683 = x77 & ~n6931 ;
  assign n11684 = n7216 & n11683 ;
  assign n11685 = n11682 | n11684 ;
  assign n11686 = n11681 | n11685 ;
  assign n11687 = n6940 | n11686 ;
  assign n11688 = ( n961 & n11686 ) | ( n961 & n11687 ) | ( n11686 & n11687 ) ;
  assign n11689 = x47 & n11688 ;
  assign n11690 = x47 & ~n11689 ;
  assign n11691 = ( n11688 & ~n11689 ) | ( n11688 & n11690 ) | ( ~n11689 & n11690 ) ;
  assign n11692 = n11680 & n11691 ;
  assign n11693 = n11680 | n11691 ;
  assign n11694 = ~n11692 & n11693 ;
  assign n11695 = n11358 | n11694 ;
  assign n11696 = n11362 | n11695 ;
  assign n11697 = ( n11358 & n11362 ) | ( n11358 & n11694 ) | ( n11362 & n11694 ) ;
  assign n11698 = n11696 & ~n11697 ;
  assign n11699 = x82 & n6068 ;
  assign n11700 = x81 & n6063 ;
  assign n11701 = x80 & ~n6062 ;
  assign n11702 = n6398 & n11701 ;
  assign n11703 = n11700 | n11702 ;
  assign n11704 = n11699 | n11703 ;
  assign n11705 = n6071 | n11704 ;
  assign n11706 = ( n1371 & n11704 ) | ( n1371 & n11705 ) | ( n11704 & n11705 ) ;
  assign n11707 = x44 & n11706 ;
  assign n11708 = x44 & ~n11707 ;
  assign n11709 = ( n11706 & ~n11707 ) | ( n11706 & n11708 ) | ( ~n11707 & n11708 ) ;
  assign n11710 = ( n11612 & n11698 ) | ( n11612 & n11709 ) | ( n11698 & n11709 ) ;
  assign n11711 = ( n11698 & n11709 ) | ( n11698 & ~n11710 ) | ( n11709 & ~n11710 ) ;
  assign n11712 = ( n11612 & ~n11710 ) | ( n11612 & n11711 ) | ( ~n11710 & n11711 ) ;
  assign n11713 = n11611 & n11712 ;
  assign n11714 = n11611 | n11712 ;
  assign n11715 = ~n11713 & n11714 ;
  assign n11716 = ( n11277 & n11278 ) | ( n11277 & n11383 ) | ( n11278 & n11383 ) ;
  assign n11717 = n11715 | n11716 ;
  assign n11718 = n11715 & n11716 ;
  assign n11719 = n11717 & ~n11718 ;
  assign n11720 = x88 & n4572 ;
  assign n11721 = x87 & n4567 ;
  assign n11722 = x86 & ~n4566 ;
  assign n11723 = n4828 & n11722 ;
  assign n11724 = n11721 | n11723 ;
  assign n11725 = n11720 | n11724 ;
  assign n11726 = n4575 | n11725 ;
  assign n11727 = ( n2095 & n11725 ) | ( n2095 & n11726 ) | ( n11725 & n11726 ) ;
  assign n11728 = x38 & n11727 ;
  assign n11729 = x38 & ~n11728 ;
  assign n11730 = ( n11727 & ~n11728 ) | ( n11727 & n11729 ) | ( ~n11728 & n11729 ) ;
  assign n11731 = n11719 & n11730 ;
  assign n11732 = n11719 & ~n11731 ;
  assign n11733 = ~n11719 & n11730 ;
  assign n11734 = n11732 | n11733 ;
  assign n11735 = n11387 | n11392 ;
  assign n11736 = n11734 | n11735 ;
  assign n11737 = n11734 & n11735 ;
  assign n11738 = n11736 & ~n11737 ;
  assign n11739 = x91 & n3913 ;
  assign n11740 = x90 & n3908 ;
  assign n11741 = x89 & ~n3907 ;
  assign n11742 = n4152 & n11741 ;
  assign n11743 = n11740 | n11742 ;
  assign n11744 = n11739 | n11743 ;
  assign n11745 = n3916 | n11744 ;
  assign n11746 = ( n2714 & n11744 ) | ( n2714 & n11745 ) | ( n11744 & n11745 ) ;
  assign n11747 = x35 & n11746 ;
  assign n11748 = x35 & ~n11747 ;
  assign n11749 = ( n11746 & ~n11747 ) | ( n11746 & n11748 ) | ( ~n11747 & n11748 ) ;
  assign n11750 = n11738 & n11749 ;
  assign n11751 = n11738 & ~n11750 ;
  assign n11752 = ~n11738 & n11749 ;
  assign n11753 = n11751 | n11752 ;
  assign n11754 = n11405 | n11411 ;
  assign n11755 = n11753 | n11754 ;
  assign n11756 = n11753 & n11754 ;
  assign n11757 = n11755 & ~n11756 ;
  assign n11758 = x94 & n3314 ;
  assign n11759 = x93 & n3309 ;
  assign n11760 = x92 & ~n3308 ;
  assign n11761 = n3570 & n11760 ;
  assign n11762 = n11759 | n11761 ;
  assign n11763 = n11758 | n11762 ;
  assign n11764 = n3317 | n11763 ;
  assign n11765 = ( n3271 & n11763 ) | ( n3271 & n11764 ) | ( n11763 & n11764 ) ;
  assign n11766 = x32 & n11765 ;
  assign n11767 = x32 & ~n11766 ;
  assign n11768 = ( n11765 & ~n11766 ) | ( n11765 & n11767 ) | ( ~n11766 & n11767 ) ;
  assign n11769 = n11757 | n11768 ;
  assign n11770 = n11757 & n11768 ;
  assign n11771 = n11769 & ~n11770 ;
  assign n11772 = n11600 & n11771 ;
  assign n11773 = n11600 | n11771 ;
  assign n11774 = ~n11772 & n11773 ;
  assign n11775 = ( n11598 & n11599 ) | ( n11598 & ~n11774 ) | ( n11599 & ~n11774 ) ;
  assign n11776 = ( ~n11599 & n11774 ) | ( ~n11599 & n11775 ) | ( n11774 & n11775 ) ;
  assign n11777 = ( ~n11598 & n11775 ) | ( ~n11598 & n11776 ) | ( n11775 & n11776 ) ;
  assign n11778 = n11587 & n11777 ;
  assign n11779 = n11587 | n11777 ;
  assign n11780 = ~n11778 & n11779 ;
  assign n11781 = n11576 | n11780 ;
  assign n11782 = n11576 & n11780 ;
  assign n11783 = n11781 & ~n11782 ;
  assign n11784 = x103 & n1817 ;
  assign n11785 = x102 & n1812 ;
  assign n11786 = x101 & ~n1811 ;
  assign n11787 = n1977 & n11786 ;
  assign n11788 = n11785 | n11787 ;
  assign n11789 = n11784 | n11788 ;
  assign n11790 = n1820 | n11789 ;
  assign n11791 = ( n5264 & n11789 ) | ( n5264 & n11790 ) | ( n11789 & n11790 ) ;
  assign n11792 = x23 & n11791 ;
  assign n11793 = x23 & ~n11792 ;
  assign n11794 = ( n11791 & ~n11792 ) | ( n11791 & n11793 ) | ( ~n11792 & n11793 ) ;
  assign n11795 = n11783 & n11794 ;
  assign n11796 = n11783 & ~n11795 ;
  assign n11797 = ~n11783 & n11794 ;
  assign n11798 = n11796 | n11797 ;
  assign n11799 = n11477 | n11483 ;
  assign n11800 = n11798 | n11799 ;
  assign n11801 = n11798 & n11799 ;
  assign n11802 = n11800 & ~n11801 ;
  assign n11803 = x106 & n1421 ;
  assign n11804 = x105 & n1416 ;
  assign n11805 = x104 & ~n1415 ;
  assign n11806 = n1584 & n11805 ;
  assign n11807 = n11804 | n11806 ;
  assign n11808 = n11803 | n11807 ;
  assign n11809 = n1424 | n11808 ;
  assign n11810 = ( n5814 & n11808 ) | ( n5814 & n11809 ) | ( n11808 & n11809 ) ;
  assign n11811 = x20 & n11810 ;
  assign n11812 = x20 & ~n11811 ;
  assign n11813 = ( n11810 & ~n11811 ) | ( n11810 & n11812 ) | ( ~n11811 & n11812 ) ;
  assign n11814 = n11802 | n11813 ;
  assign n11815 = n11802 & n11813 ;
  assign n11816 = n11814 & ~n11815 ;
  assign n11817 = n11575 & n11816 ;
  assign n11818 = n11575 | n11816 ;
  assign n11819 = ~n11817 & n11818 ;
  assign n11820 = x109 & n1071 ;
  assign n11821 = x108 & n1066 ;
  assign n11822 = x107 & ~n1065 ;
  assign n11823 = n1189 & n11822 ;
  assign n11824 = n11821 | n11823 ;
  assign n11825 = n11820 | n11824 ;
  assign n11826 = n1074 | n11825 ;
  assign n11827 = ( n6884 & n11825 ) | ( n6884 & n11826 ) | ( n11825 & n11826 ) ;
  assign n11828 = x17 & n11827 ;
  assign n11829 = x17 & ~n11828 ;
  assign n11830 = ( n11827 & ~n11828 ) | ( n11827 & n11829 ) | ( ~n11828 & n11829 ) ;
  assign n11831 = n11819 & n11830 ;
  assign n11832 = n11819 & ~n11831 ;
  assign n11833 = ~n11819 & n11830 ;
  assign n11834 = n11832 | n11833 ;
  assign n11835 = ( n11253 & n11254 ) | ( n11253 & n11502 ) | ( n11254 & n11502 ) ;
  assign n11836 = n11834 & n11835 ;
  assign n11837 = n11834 | n11835 ;
  assign n11838 = ~n11836 & n11837 ;
  assign n11839 = x112 & n771 ;
  assign n11840 = x111 & n766 ;
  assign n11841 = x110 & ~n765 ;
  assign n11842 = n905 & n11841 ;
  assign n11843 = n11840 | n11842 ;
  assign n11844 = n11839 | n11843 ;
  assign n11845 = n774 | n11844 ;
  assign n11846 = ( n7789 & n11844 ) | ( n7789 & n11845 ) | ( n11844 & n11845 ) ;
  assign n11847 = x14 & n11846 ;
  assign n11848 = x14 & ~n11847 ;
  assign n11849 = ( n11846 & ~n11847 ) | ( n11846 & n11848 ) | ( ~n11847 & n11848 ) ;
  assign n11850 = n11838 & n11849 ;
  assign n11851 = n11838 & ~n11850 ;
  assign n11852 = ~n11838 & n11849 ;
  assign n11853 = n11851 | n11852 ;
  assign n11854 = n11574 & n11853 ;
  assign n11855 = n11574 | n11853 ;
  assign n11856 = ~n11854 & n11855 ;
  assign n11857 = x115 & n528 ;
  assign n11858 = x114 & n523 ;
  assign n11859 = x113 & ~n522 ;
  assign n11860 = n635 & n11859 ;
  assign n11861 = n11858 | n11860 ;
  assign n11862 = n11857 | n11861 ;
  assign n11863 = n531 | n11862 ;
  assign n11864 = ( n8749 & n11862 ) | ( n8749 & n11863 ) | ( n11862 & n11863 ) ;
  assign n11865 = x11 & n11864 ;
  assign n11866 = x11 & ~n11865 ;
  assign n11867 = ( n11864 & ~n11865 ) | ( n11864 & n11866 ) | ( ~n11865 & n11866 ) ;
  assign n11868 = n11856 & n11867 ;
  assign n11869 = n11856 & ~n11868 ;
  assign n11870 = ~n11856 & n11867 ;
  assign n11871 = n11869 | n11870 ;
  assign n11872 = n11573 & n11871 ;
  assign n11873 = n11573 | n11871 ;
  assign n11874 = ~n11872 & n11873 ;
  assign n11875 = x118 & n337 ;
  assign n11876 = x117 & n332 ;
  assign n11877 = x116 & ~n331 ;
  assign n11878 = n396 & n11877 ;
  assign n11879 = n11876 | n11878 ;
  assign n11880 = n11875 | n11879 ;
  assign n11881 = n340 | n11880 ;
  assign n11882 = ( n9760 & n11880 ) | ( n9760 & n11881 ) | ( n11880 & n11881 ) ;
  assign n11883 = x8 & n11882 ;
  assign n11884 = x8 & ~n11883 ;
  assign n11885 = ( n11882 & ~n11883 ) | ( n11882 & n11884 ) | ( ~n11883 & n11884 ) ;
  assign n11886 = n11874 & n11885 ;
  assign n11887 = n11874 | n11885 ;
  assign n11888 = ~n11886 & n11887 ;
  assign n11889 = n11572 & n11888 ;
  assign n11890 = n11572 | n11888 ;
  assign n11891 = ~n11889 & n11890 ;
  assign n11892 = x121 & n206 ;
  assign n11893 = x120 & n201 ;
  assign n11894 = x119 & ~n200 ;
  assign n11895 = n243 & n11894 ;
  assign n11896 = n11893 | n11895 ;
  assign n11897 = n11892 | n11896 ;
  assign n11898 = n209 | n11897 ;
  assign n11899 = ( n10811 & n11897 ) | ( n10811 & n11898 ) | ( n11897 & n11898 ) ;
  assign n11900 = x5 & n11899 ;
  assign n11901 = x5 & ~n11900 ;
  assign n11902 = ( n11899 & ~n11900 ) | ( n11899 & n11901 ) | ( ~n11900 & n11901 ) ;
  assign n11903 = n11891 & n11902 ;
  assign n11904 = n11891 | n11902 ;
  assign n11905 = ~n11903 & n11904 ;
  assign n11906 = x123 | x124 ;
  assign n11907 = x123 & x124 ;
  assign n11908 = n11906 & ~n11907 ;
  assign n11909 = n11210 | n11213 ;
  assign n11910 = n11908 & n11909 ;
  assign n11911 = n11210 | n11215 ;
  assign n11912 = n11908 & n11911 ;
  assign n11913 = ( n9786 & n11910 ) | ( n9786 & n11912 ) | ( n11910 & n11912 ) ;
  assign n11914 = ( n9786 & n11909 ) | ( n9786 & n11911 ) | ( n11909 & n11911 ) ;
  assign n11915 = n11908 | n11914 ;
  assign n11916 = ~n11913 & n11915 ;
  assign n11917 = x123 & n131 ;
  assign n11918 = x122 & ~n156 ;
  assign n11919 = ( n135 & n11917 ) | ( n135 & n11918 ) | ( n11917 & n11918 ) ;
  assign n11920 = x0 & x124 ;
  assign n11921 = ( ~n135 & n11917 ) | ( ~n135 & n11920 ) | ( n11917 & n11920 ) ;
  assign n11922 = n11919 | n11921 ;
  assign n11923 = n139 | n11922 ;
  assign n11924 = ( n11916 & n11922 ) | ( n11916 & n11923 ) | ( n11922 & n11923 ) ;
  assign n11925 = x2 & n11924 ;
  assign n11926 = x2 & ~n11925 ;
  assign n11927 = ( n11924 & ~n11925 ) | ( n11924 & n11926 ) | ( ~n11925 & n11926 ) ;
  assign n11928 = n11905 & n11927 ;
  assign n11929 = n11905 | n11927 ;
  assign n11930 = ~n11928 & n11929 ;
  assign n11931 = ( n11230 & n11561 ) | ( n11230 & ~n11564 ) | ( n11561 & ~n11564 ) ;
  assign n11932 = n11930 & n11931 ;
  assign n11933 = n11930 | n11931 ;
  assign n11934 = ~n11932 & n11933 ;
  assign n11935 = n11566 | n11569 ;
  assign n11936 = n11934 & n11935 ;
  assign n11937 = n11934 | n11935 ;
  assign n11938 = ~n11936 & n11937 ;
  assign n11939 = n11903 | n11928 ;
  assign n11940 = n11868 | n11872 ;
  assign n11941 = n11850 | n11854 ;
  assign n11942 = n11831 | n11836 ;
  assign n11943 = x98 & n2775 ;
  assign n11944 = x97 & n2770 ;
  assign n11945 = x96 & ~n2769 ;
  assign n11946 = n2978 & n11945 ;
  assign n11947 = n11944 | n11946 ;
  assign n11948 = n11943 | n11947 ;
  assign n11949 = n2778 | n11948 ;
  assign n11950 = ( n4105 & n11948 ) | ( n4105 & n11949 ) | ( n11948 & n11949 ) ;
  assign n11951 = x29 & n11950 ;
  assign n11952 = x29 & ~n11951 ;
  assign n11953 = ( n11950 & ~n11951 ) | ( n11950 & n11952 ) | ( ~n11951 & n11952 ) ;
  assign n11954 = x95 & n3314 ;
  assign n11955 = x94 & n3309 ;
  assign n11956 = x93 & ~n3308 ;
  assign n11957 = n3570 & n11956 ;
  assign n11958 = n11955 | n11957 ;
  assign n11959 = n11954 | n11958 ;
  assign n11960 = n3317 | n11959 ;
  assign n11961 = ( n3479 & n11959 ) | ( n3479 & n11960 ) | ( n11959 & n11960 ) ;
  assign n11962 = x32 & n11961 ;
  assign n11963 = x32 & ~n11962 ;
  assign n11964 = ( n11961 & ~n11962 ) | ( n11961 & n11963 ) | ( ~n11962 & n11963 ) ;
  assign n11965 = x71 & n9853 ;
  assign n11966 = x70 & n9848 ;
  assign n11967 = x69 & ~n9847 ;
  assign n11968 = n10165 & n11967 ;
  assign n11969 = n11966 | n11968 ;
  assign n11970 = n11965 | n11969 ;
  assign n11971 = n9856 | n11970 ;
  assign n11972 = ( n376 & n11970 ) | ( n376 & n11971 ) | ( n11970 & n11971 ) ;
  assign n11973 = x56 & ~n11972 ;
  assign n11974 = ~x56 & n11972 ;
  assign n11975 = n11973 | n11974 ;
  assign n11976 = ~x60 & x61 ;
  assign n11977 = x60 & ~x61 ;
  assign n11978 = n11976 | n11977 ;
  assign n11979 = ~n11627 & n11978 ;
  assign n11980 = x64 & n11979 ;
  assign n11981 = ~x61 & x62 ;
  assign n11982 = x61 & ~x62 ;
  assign n11983 = n11981 | n11982 ;
  assign n11984 = n11627 & ~n11983 ;
  assign n11985 = x65 & n11984 ;
  assign n11986 = n11980 | n11985 ;
  assign n11987 = n11627 & n11983 ;
  assign n11988 = n142 & n11987 ;
  assign n11989 = n11986 | n11988 ;
  assign n11990 = x62 | n11989 ;
  assign n11991 = ~x62 & n11990 ;
  assign n11992 = ( ~n11989 & n11990 ) | ( ~n11989 & n11991 ) | ( n11990 & n11991 ) ;
  assign n11993 = x62 & ~n11628 ;
  assign n11994 = n11992 & n11993 ;
  assign n11995 = n11992 | n11993 ;
  assign n11996 = ~n11994 & n11995 ;
  assign n11997 = n229 & n10879 ;
  assign n11998 = x68 & n10876 ;
  assign n11999 = x67 & n10871 ;
  assign n12000 = x66 & ~n10870 ;
  assign n12001 = n11305 & n12000 ;
  assign n12002 = n11999 | n12001 ;
  assign n12003 = n11998 | n12002 ;
  assign n12004 = n11997 | n12003 ;
  assign n12005 = x59 | n12004 ;
  assign n12006 = ~x59 & n12005 ;
  assign n12007 = ( ~n12004 & n12005 ) | ( ~n12004 & n12006 ) | ( n12005 & n12006 ) ;
  assign n12008 = n11996 | n12007 ;
  assign n12009 = n11996 & n12007 ;
  assign n12010 = n12008 & ~n12009 ;
  assign n12011 = n11640 | n12010 ;
  assign n12012 = n11640 & n12010 ;
  assign n12013 = n12011 & ~n12012 ;
  assign n12014 = n11975 | n12013 ;
  assign n12015 = n11975 & n12013 ;
  assign n12016 = n12014 & ~n12015 ;
  assign n12017 = ( n11319 & n11624 ) | ( n11319 & n11642 ) | ( n11624 & n11642 ) ;
  assign n12018 = n12016 | n12017 ;
  assign n12019 = n12016 & n12017 ;
  assign n12020 = n12018 & ~n12019 ;
  assign n12021 = x74 & n8834 ;
  assign n12022 = x73 & n8829 ;
  assign n12023 = x72 & ~n8828 ;
  assign n12024 = n9159 & n12023 ;
  assign n12025 = n12022 | n12024 ;
  assign n12026 = n12021 | n12025 ;
  assign n12027 = n8837 | n12026 ;
  assign n12028 = ( n587 & n12026 ) | ( n587 & n12027 ) | ( n12026 & n12027 ) ;
  assign n12029 = x53 & n12028 ;
  assign n12030 = x53 & ~n12029 ;
  assign n12031 = ( n12028 & ~n12029 ) | ( n12028 & n12030 ) | ( ~n12029 & n12030 ) ;
  assign n12032 = n12020 & n12031 ;
  assign n12033 = n12020 & ~n12032 ;
  assign n12034 = ~n12020 & n12031 ;
  assign n12035 = n12033 | n12034 ;
  assign n12036 = n11657 | n11660 ;
  assign n12037 = n12035 | n12036 ;
  assign n12038 = n12035 & n12036 ;
  assign n12039 = n12037 & ~n12038 ;
  assign n12040 = x77 & n7812 ;
  assign n12041 = x76 & n7807 ;
  assign n12042 = x75 & ~n7806 ;
  assign n12043 = n8136 & n12042 ;
  assign n12044 = n12041 | n12043 ;
  assign n12045 = n12040 | n12044 ;
  assign n12046 = n7815 | n12045 ;
  assign n12047 = ( n846 & n12045 ) | ( n846 & n12046 ) | ( n12045 & n12046 ) ;
  assign n12048 = x50 & n12047 ;
  assign n12049 = x50 & ~n12048 ;
  assign n12050 = ( n12047 & ~n12048 ) | ( n12047 & n12049 ) | ( ~n12048 & n12049 ) ;
  assign n12051 = n12039 & n12050 ;
  assign n12052 = n12039 | n12050 ;
  assign n12053 = ~n12051 & n12052 ;
  assign n12054 = n11675 | n11678 ;
  assign n12055 = n12053 & n12054 ;
  assign n12056 = n12054 & ~n12055 ;
  assign n12057 = ( n12053 & ~n12055 ) | ( n12053 & n12056 ) | ( ~n12055 & n12056 ) ;
  assign n12058 = x80 & n6937 ;
  assign n12059 = x79 & n6932 ;
  assign n12060 = x78 & ~n6931 ;
  assign n12061 = n7216 & n12060 ;
  assign n12062 = n12059 | n12061 ;
  assign n12063 = n12058 | n12062 ;
  assign n12064 = n6940 | n12063 ;
  assign n12065 = ( n1147 & n12063 ) | ( n1147 & n12064 ) | ( n12063 & n12064 ) ;
  assign n12066 = x47 & n12065 ;
  assign n12067 = x47 & ~n12066 ;
  assign n12068 = ( n12065 & ~n12066 ) | ( n12065 & n12067 ) | ( ~n12066 & n12067 ) ;
  assign n12069 = n12057 & n12068 ;
  assign n12070 = n12057 & ~n12069 ;
  assign n12071 = ~n12057 & n12068 ;
  assign n12072 = n12070 | n12071 ;
  assign n12073 = n11692 | n11697 ;
  assign n12074 = n12072 | n12073 ;
  assign n12075 = n12072 & n12073 ;
  assign n12076 = n12074 & ~n12075 ;
  assign n12077 = x83 & n6068 ;
  assign n12078 = x82 & n6063 ;
  assign n12079 = x81 & ~n6062 ;
  assign n12080 = n6398 & n12079 ;
  assign n12081 = n12078 | n12080 ;
  assign n12082 = n12077 | n12081 ;
  assign n12083 = n6071 | n12082 ;
  assign n12084 = ( n1510 & n12082 ) | ( n1510 & n12083 ) | ( n12082 & n12083 ) ;
  assign n12085 = x44 & n12084 ;
  assign n12086 = x44 & ~n12085 ;
  assign n12087 = ( n12084 & ~n12085 ) | ( n12084 & n12086 ) | ( ~n12085 & n12086 ) ;
  assign n12088 = n12076 & n12087 ;
  assign n12089 = n12076 | n12087 ;
  assign n12090 = ~n12088 & n12089 ;
  assign n12091 = n11710 & n12090 ;
  assign n12092 = n11710 & ~n12091 ;
  assign n12093 = ( n12090 & ~n12091 ) | ( n12090 & n12092 ) | ( ~n12091 & n12092 ) ;
  assign n12094 = x86 & n5340 ;
  assign n12095 = x85 & n5335 ;
  assign n12096 = x84 & ~n5334 ;
  assign n12097 = n5580 & n12096 ;
  assign n12098 = n12095 | n12097 ;
  assign n12099 = n12094 | n12098 ;
  assign n12100 = n5343 | n12099 ;
  assign n12101 = ( n1921 & n12099 ) | ( n1921 & n12100 ) | ( n12099 & n12100 ) ;
  assign n12102 = x41 & n12101 ;
  assign n12103 = x41 & ~n12102 ;
  assign n12104 = ( n12101 & ~n12102 ) | ( n12101 & n12103 ) | ( ~n12102 & n12103 ) ;
  assign n12105 = n12093 & n12104 ;
  assign n12106 = n12093 & ~n12105 ;
  assign n12107 = ~n12093 & n12104 ;
  assign n12108 = n12106 | n12107 ;
  assign n12109 = n11713 | n11718 ;
  assign n12110 = n12108 | n12109 ;
  assign n12111 = n12108 & n12109 ;
  assign n12112 = n12110 & ~n12111 ;
  assign n12113 = x89 & n4572 ;
  assign n12114 = x88 & n4567 ;
  assign n12115 = x87 & ~n4566 ;
  assign n12116 = n4828 & n12115 ;
  assign n12117 = n12114 | n12116 ;
  assign n12118 = n12113 | n12117 ;
  assign n12119 = n4575 | n12118 ;
  assign n12120 = ( n2244 & n12118 ) | ( n2244 & n12119 ) | ( n12118 & n12119 ) ;
  assign n12121 = x38 & n12120 ;
  assign n12122 = x38 & ~n12121 ;
  assign n12123 = ( n12120 & ~n12121 ) | ( n12120 & n12122 ) | ( ~n12121 & n12122 ) ;
  assign n12124 = n12112 & n12123 ;
  assign n12125 = n12112 & ~n12124 ;
  assign n12126 = ~n12112 & n12123 ;
  assign n12127 = n12125 | n12126 ;
  assign n12128 = n11731 | n11737 ;
  assign n12129 = n12127 | n12128 ;
  assign n12130 = n12127 & n12128 ;
  assign n12131 = n12129 & ~n12130 ;
  assign n12132 = x92 & n3913 ;
  assign n12133 = x91 & n3908 ;
  assign n12134 = x90 & ~n3907 ;
  assign n12135 = n4152 & n12134 ;
  assign n12136 = n12133 | n12135 ;
  assign n12137 = n12132 | n12136 ;
  assign n12138 = n3916 | n12137 ;
  assign n12139 = ( n2904 & n12137 ) | ( n2904 & n12138 ) | ( n12137 & n12138 ) ;
  assign n12140 = x35 & n12139 ;
  assign n12141 = x35 & ~n12140 ;
  assign n12142 = ( n12139 & ~n12140 ) | ( n12139 & n12141 ) | ( ~n12140 & n12141 ) ;
  assign n12143 = n12131 & n12142 ;
  assign n12144 = n12131 & ~n12143 ;
  assign n12145 = ~n12131 & n12142 ;
  assign n12146 = n12144 | n12145 ;
  assign n12147 = n11750 | n11756 ;
  assign n12148 = n12146 | n12147 ;
  assign n12149 = n12146 & n12147 ;
  assign n12150 = n12148 & ~n12149 ;
  assign n12151 = n11770 | n11772 ;
  assign n12152 = ( n11964 & n12150 ) | ( n11964 & n12151 ) | ( n12150 & n12151 ) ;
  assign n12153 = ( n12150 & n12151 ) | ( n12150 & ~n12152 ) | ( n12151 & ~n12152 ) ;
  assign n12154 = ( n11964 & ~n12152 ) | ( n11964 & n12153 ) | ( ~n12152 & n12153 ) ;
  assign n12155 = n11953 & n12154 ;
  assign n12156 = n11953 | n12154 ;
  assign n12157 = ~n12155 & n12156 ;
  assign n12158 = ( n11598 & n11599 ) | ( n11598 & n11774 ) | ( n11599 & n11774 ) ;
  assign n12159 = n12157 | n12158 ;
  assign n12160 = n12157 & n12158 ;
  assign n12161 = n12159 & ~n12160 ;
  assign n12162 = x101 & n2280 ;
  assign n12163 = x100 & n2275 ;
  assign n12164 = x99 & ~n2274 ;
  assign n12165 = n2481 & n12164 ;
  assign n12166 = n12163 | n12165 ;
  assign n12167 = n12162 | n12166 ;
  assign n12168 = n2283 | n12167 ;
  assign n12169 = ( n4783 & n12167 ) | ( n4783 & n12168 ) | ( n12167 & n12168 ) ;
  assign n12170 = x26 & n12169 ;
  assign n12171 = x26 & ~n12170 ;
  assign n12172 = ( n12169 & ~n12170 ) | ( n12169 & n12171 ) | ( ~n12170 & n12171 ) ;
  assign n12173 = n12161 & n12172 ;
  assign n12174 = n12161 & ~n12173 ;
  assign n12175 = ~n12161 & n12172 ;
  assign n12176 = n12174 | n12175 ;
  assign n12177 = n11778 | n11782 ;
  assign n12178 = n12176 | n12177 ;
  assign n12179 = n12176 & n12177 ;
  assign n12180 = n12178 & ~n12179 ;
  assign n12181 = x104 & n1817 ;
  assign n12182 = x103 & n1812 ;
  assign n12183 = x102 & ~n1811 ;
  assign n12184 = n1977 & n12183 ;
  assign n12185 = n12182 | n12184 ;
  assign n12186 = n12181 | n12185 ;
  assign n12187 = n1820 | n12186 ;
  assign n12188 = ( n5295 & n12186 ) | ( n5295 & n12187 ) | ( n12186 & n12187 ) ;
  assign n12189 = x23 & n12188 ;
  assign n12190 = x23 & ~n12189 ;
  assign n12191 = ( n12188 & ~n12189 ) | ( n12188 & n12190 ) | ( ~n12189 & n12190 ) ;
  assign n12192 = n12180 & n12191 ;
  assign n12193 = n12180 & ~n12192 ;
  assign n12194 = ~n12180 & n12191 ;
  assign n12195 = n12193 | n12194 ;
  assign n12196 = n11795 | n11801 ;
  assign n12197 = n12195 | n12196 ;
  assign n12198 = n12195 & n12196 ;
  assign n12199 = n12197 & ~n12198 ;
  assign n12200 = x107 & n1421 ;
  assign n12201 = x106 & n1416 ;
  assign n12202 = x105 & ~n1415 ;
  assign n12203 = n1584 & n12202 ;
  assign n12204 = n12201 | n12203 ;
  assign n12205 = n12200 | n12204 ;
  assign n12206 = n1424 | n12205 ;
  assign n12207 = ( n6328 & n12205 ) | ( n6328 & n12206 ) | ( n12205 & n12206 ) ;
  assign n12208 = x20 & n12207 ;
  assign n12209 = x20 & ~n12208 ;
  assign n12210 = ( n12207 & ~n12208 ) | ( n12207 & n12209 ) | ( ~n12208 & n12209 ) ;
  assign n12211 = n12199 & n12210 ;
  assign n12212 = n12199 | n12210 ;
  assign n12213 = ~n12211 & n12212 ;
  assign n12214 = n11815 | n11817 ;
  assign n12215 = n12213 & n12214 ;
  assign n12216 = n12214 & ~n12215 ;
  assign n12217 = ( n12213 & ~n12215 ) | ( n12213 & n12216 ) | ( ~n12215 & n12216 ) ;
  assign n12218 = x110 & n1071 ;
  assign n12219 = x109 & n1066 ;
  assign n12220 = x108 & ~n1065 ;
  assign n12221 = n1189 & n12220 ;
  assign n12222 = n12219 | n12221 ;
  assign n12223 = n12218 | n12222 ;
  assign n12224 = n1074 | n12223 ;
  assign n12225 = ( n7189 & n12223 ) | ( n7189 & n12224 ) | ( n12223 & n12224 ) ;
  assign n12226 = x17 & n12225 ;
  assign n12227 = x17 & ~n12226 ;
  assign n12228 = ( n12225 & ~n12226 ) | ( n12225 & n12227 ) | ( ~n12226 & n12227 ) ;
  assign n12229 = n12217 | n12228 ;
  assign n12230 = n12217 & n12228 ;
  assign n12231 = n12229 & ~n12230 ;
  assign n12232 = n11942 & n12231 ;
  assign n12233 = n11942 | n12231 ;
  assign n12234 = ~n12232 & n12233 ;
  assign n12235 = x113 & n771 ;
  assign n12236 = x112 & n766 ;
  assign n12237 = x111 & ~n765 ;
  assign n12238 = n905 & n12237 ;
  assign n12239 = n12236 | n12238 ;
  assign n12240 = n12235 | n12239 ;
  assign n12241 = n774 | n12240 ;
  assign n12242 = ( n8113 & n12240 ) | ( n8113 & n12241 ) | ( n12240 & n12241 ) ;
  assign n12243 = x14 & n12242 ;
  assign n12244 = x14 & ~n12243 ;
  assign n12245 = ( n12242 & ~n12243 ) | ( n12242 & n12244 ) | ( ~n12243 & n12244 ) ;
  assign n12246 = n12234 | n12245 ;
  assign n12247 = n12234 & n12245 ;
  assign n12248 = n12246 & ~n12247 ;
  assign n12249 = n11941 & n12248 ;
  assign n12250 = n11941 | n12248 ;
  assign n12251 = ~n12249 & n12250 ;
  assign n12252 = x116 & n528 ;
  assign n12253 = x115 & n523 ;
  assign n12254 = x114 & ~n522 ;
  assign n12255 = n635 & n12254 ;
  assign n12256 = n12253 | n12255 ;
  assign n12257 = n12252 | n12256 ;
  assign n12258 = n531 | n12257 ;
  assign n12259 = ( n8778 & n12257 ) | ( n8778 & n12258 ) | ( n12257 & n12258 ) ;
  assign n12260 = x11 & n12259 ;
  assign n12261 = x11 & ~n12260 ;
  assign n12262 = ( n12259 & ~n12260 ) | ( n12259 & n12261 ) | ( ~n12260 & n12261 ) ;
  assign n12263 = n12251 | n12262 ;
  assign n12264 = n12251 & n12262 ;
  assign n12265 = n12263 & ~n12264 ;
  assign n12266 = n11940 & n12265 ;
  assign n12267 = n11940 | n12265 ;
  assign n12268 = ~n12266 & n12267 ;
  assign n12269 = x119 & n337 ;
  assign n12270 = x118 & n332 ;
  assign n12271 = x117 & ~n331 ;
  assign n12272 = n396 & n12271 ;
  assign n12273 = n12270 | n12272 ;
  assign n12274 = n12269 | n12273 ;
  assign n12275 = n340 | n12274 ;
  assign n12276 = ( n9789 & n12274 ) | ( n9789 & n12275 ) | ( n12274 & n12275 ) ;
  assign n12277 = x8 & n12276 ;
  assign n12278 = x8 & ~n12277 ;
  assign n12279 = ( n12276 & ~n12277 ) | ( n12276 & n12278 ) | ( ~n12277 & n12278 ) ;
  assign n12280 = n12268 & n12279 ;
  assign n12281 = n12268 & ~n12280 ;
  assign n12282 = ~n12268 & n12279 ;
  assign n12283 = n12281 | n12282 ;
  assign n12284 = n11886 | n11889 ;
  assign n12285 = n12283 | n12284 ;
  assign n12286 = n12283 & n12284 ;
  assign n12287 = n12285 & ~n12286 ;
  assign n12288 = x122 & n206 ;
  assign n12289 = x121 & n201 ;
  assign n12290 = x120 & ~n200 ;
  assign n12291 = n243 & n12290 ;
  assign n12292 = n12289 | n12291 ;
  assign n12293 = n12288 | n12292 ;
  assign n12294 = n209 | n12293 ;
  assign n12295 = ( n11188 & n12293 ) | ( n11188 & n12294 ) | ( n12293 & n12294 ) ;
  assign n12296 = x5 & n12295 ;
  assign n12297 = x5 & ~n12296 ;
  assign n12298 = ( n12295 & ~n12296 ) | ( n12295 & n12297 ) | ( ~n12296 & n12297 ) ;
  assign n12299 = n12287 | n12298 ;
  assign n12300 = x124 | x125 ;
  assign n12301 = x124 & x125 ;
  assign n12302 = n12300 & ~n12301 ;
  assign n12303 = n11907 | n11910 ;
  assign n12304 = n12302 & n12303 ;
  assign n12305 = n11907 | n11912 ;
  assign n12306 = n12302 & n12305 ;
  assign n12307 = ( n9786 & n12304 ) | ( n9786 & n12306 ) | ( n12304 & n12306 ) ;
  assign n12308 = ( n9786 & n12303 ) | ( n9786 & n12305 ) | ( n12303 & n12305 ) ;
  assign n12309 = n12302 | n12308 ;
  assign n12310 = ~n12307 & n12309 ;
  assign n12311 = x124 & n131 ;
  assign n12312 = x123 & ~n156 ;
  assign n12313 = ( n135 & n12311 ) | ( n135 & n12312 ) | ( n12311 & n12312 ) ;
  assign n12314 = x0 & x125 ;
  assign n12315 = ( ~n135 & n12311 ) | ( ~n135 & n12314 ) | ( n12311 & n12314 ) ;
  assign n12316 = n12313 | n12315 ;
  assign n12317 = n139 | n12316 ;
  assign n12318 = ( n12310 & n12316 ) | ( n12310 & n12317 ) | ( n12316 & n12317 ) ;
  assign n12319 = x2 & n12318 ;
  assign n12320 = x2 & ~n12319 ;
  assign n12321 = ( n12318 & ~n12319 ) | ( n12318 & n12320 ) | ( ~n12319 & n12320 ) ;
  assign n12322 = ( n12298 & ~n12299 ) | ( n12298 & n12321 ) | ( ~n12299 & n12321 ) ;
  assign n12323 = ( n12287 & ~n12299 ) | ( n12287 & n12322 ) | ( ~n12299 & n12322 ) ;
  assign n12324 = n11939 | n12323 ;
  assign n12325 = ( n12287 & n12298 ) | ( n12287 & n12321 ) | ( n12298 & n12321 ) ;
  assign n12326 = n12299 & ~n12325 ;
  assign n12327 = n12324 | n12326 ;
  assign n12328 = ( n11939 & n12323 ) | ( n11939 & n12326 ) | ( n12323 & n12326 ) ;
  assign n12329 = n12327 & ~n12328 ;
  assign n12330 = n11932 | n11936 ;
  assign n12331 = n12329 & n12330 ;
  assign n12332 = n12329 | n12330 ;
  assign n12333 = ~n12331 & n12332 ;
  assign n12334 = n12280 | n12286 ;
  assign n12335 = x117 & n528 ;
  assign n12336 = x116 & n523 ;
  assign n12337 = x115 & ~n522 ;
  assign n12338 = n635 & n12337 ;
  assign n12339 = n12336 | n12338 ;
  assign n12340 = n12335 | n12339 ;
  assign n12341 = n531 | n12340 ;
  assign n12342 = ( n9118 & n12340 ) | ( n9118 & n12341 ) | ( n12340 & n12341 ) ;
  assign n12343 = x11 & n12342 ;
  assign n12344 = x11 & ~n12343 ;
  assign n12345 = ( n12342 & ~n12343 ) | ( n12342 & n12344 ) | ( ~n12343 & n12344 ) ;
  assign n12346 = x114 & n771 ;
  assign n12347 = x113 & n766 ;
  assign n12348 = x112 & ~n765 ;
  assign n12349 = n905 & n12348 ;
  assign n12350 = n12347 | n12349 ;
  assign n12351 = n12346 | n12350 ;
  assign n12352 = n774 | n12351 ;
  assign n12353 = ( n8437 & n12351 ) | ( n8437 & n12352 ) | ( n12351 & n12352 ) ;
  assign n12354 = x14 & n12353 ;
  assign n12355 = x14 & ~n12354 ;
  assign n12356 = ( n12353 & ~n12354 ) | ( n12353 & n12355 ) | ( ~n12354 & n12355 ) ;
  assign n12357 = n12211 | n12215 ;
  assign n12358 = x108 & n1421 ;
  assign n12359 = x107 & n1416 ;
  assign n12360 = x106 & ~n1415 ;
  assign n12361 = n1584 & n12360 ;
  assign n12362 = n12359 | n12361 ;
  assign n12363 = n12358 | n12362 ;
  assign n12364 = n1424 | n12363 ;
  assign n12365 = ( n6358 & n12363 ) | ( n6358 & n12364 ) | ( n12363 & n12364 ) ;
  assign n12366 = x20 & n12365 ;
  assign n12367 = x20 & ~n12366 ;
  assign n12368 = ( n12365 & ~n12366 ) | ( n12365 & n12367 ) | ( ~n12366 & n12367 ) ;
  assign n12369 = x105 & n1817 ;
  assign n12370 = x104 & n1812 ;
  assign n12371 = x103 & ~n1811 ;
  assign n12372 = n1977 & n12371 ;
  assign n12373 = n12370 | n12372 ;
  assign n12374 = n12369 | n12373 ;
  assign n12375 = n1820 | n12374 ;
  assign n12376 = ( n5788 & n12374 ) | ( n5788 & n12375 ) | ( n12374 & n12375 ) ;
  assign n12377 = x23 & n12376 ;
  assign n12378 = x23 & ~n12377 ;
  assign n12379 = ( n12376 & ~n12377 ) | ( n12376 & n12378 ) | ( ~n12377 & n12378 ) ;
  assign n12380 = n12192 | n12198 ;
  assign n12381 = x87 & n5340 ;
  assign n12382 = x86 & n5335 ;
  assign n12383 = x85 & ~n5334 ;
  assign n12384 = n5580 & n12383 ;
  assign n12385 = n12382 | n12384 ;
  assign n12386 = n12381 | n12385 ;
  assign n12387 = n5343 | n12386 ;
  assign n12388 = ( n2067 & n12386 ) | ( n2067 & n12387 ) | ( n12386 & n12387 ) ;
  assign n12389 = x41 & n12388 ;
  assign n12390 = x41 & ~n12389 ;
  assign n12391 = ( n12388 & ~n12389 ) | ( n12388 & n12390 ) | ( ~n12389 & n12390 ) ;
  assign n12392 = x84 & n6068 ;
  assign n12393 = x83 & n6063 ;
  assign n12394 = x82 & ~n6062 ;
  assign n12395 = n6398 & n12394 ;
  assign n12396 = n12393 | n12395 ;
  assign n12397 = n12392 | n12396 ;
  assign n12398 = n6071 | n12397 ;
  assign n12399 = ( n1537 & n12397 ) | ( n1537 & n12398 ) | ( n12397 & n12398 ) ;
  assign n12400 = x44 & n12399 ;
  assign n12401 = x44 & ~n12400 ;
  assign n12402 = ( n12399 & ~n12400 ) | ( n12399 & n12401 ) | ( ~n12400 & n12401 ) ;
  assign n12403 = n12088 | n12091 ;
  assign n12404 = n12069 | n12075 ;
  assign n12405 = n12051 | n12055 ;
  assign n12406 = x72 & n9853 ;
  assign n12407 = x71 & n9848 ;
  assign n12408 = x70 & ~n9847 ;
  assign n12409 = n10165 & n12408 ;
  assign n12410 = n12407 | n12409 ;
  assign n12411 = n12406 | n12410 ;
  assign n12412 = ( n435 & n9856 ) | ( n435 & n12411 ) | ( n9856 & n12411 ) ;
  assign n12413 = ( x56 & ~n12411 ) | ( x56 & n12412 ) | ( ~n12411 & n12412 ) ;
  assign n12414 = ~n12412 & n12413 ;
  assign n12415 = n12411 | n12413 ;
  assign n12416 = ( ~x56 & n12414 ) | ( ~x56 & n12415 ) | ( n12414 & n12415 ) ;
  assign n12417 = n264 & n10879 ;
  assign n12418 = x69 & n10876 ;
  assign n12419 = x68 & n10871 ;
  assign n12420 = x67 & ~n10870 ;
  assign n12421 = n11305 & n12420 ;
  assign n12422 = n12419 | n12421 ;
  assign n12423 = n12418 | n12422 ;
  assign n12424 = n12417 | n12423 ;
  assign n12425 = x59 | n12424 ;
  assign n12426 = ~x59 & n12425 ;
  assign n12427 = ( ~n12424 & n12425 ) | ( ~n12424 & n12426 ) | ( n12425 & n12426 ) ;
  assign n12428 = x66 & n11984 ;
  assign n12429 = x65 & n11979 ;
  assign n12430 = ~n11627 & n11983 ;
  assign n12431 = x64 & ~n11978 ;
  assign n12432 = n12430 & n12431 ;
  assign n12433 = n12429 | n12432 ;
  assign n12434 = n12428 | n12433 ;
  assign n12435 = n153 & n11987 ;
  assign n12436 = n12434 | n12435 ;
  assign n12437 = x62 | n12436 ;
  assign n12438 = ~x62 & n12437 ;
  assign n12439 = ( ~n12436 & n12437 ) | ( ~n12436 & n12438 ) | ( n12437 & n12438 ) ;
  assign n12440 = n11994 | n12439 ;
  assign n12441 = n11994 & n12439 ;
  assign n12442 = n12440 & ~n12441 ;
  assign n12443 = n12009 | n12012 ;
  assign n12444 = ( n12427 & n12442 ) | ( n12427 & n12443 ) | ( n12442 & n12443 ) ;
  assign n12445 = ( n12442 & n12443 ) | ( n12442 & ~n12444 ) | ( n12443 & ~n12444 ) ;
  assign n12446 = ( n12427 & ~n12444 ) | ( n12427 & n12445 ) | ( ~n12444 & n12445 ) ;
  assign n12447 = n12416 | n12446 ;
  assign n12448 = n12416 & n12446 ;
  assign n12449 = n12447 & ~n12448 ;
  assign n12450 = n12015 | n12019 ;
  assign n12451 = n12449 & n12450 ;
  assign n12452 = n12449 | n12450 ;
  assign n12453 = ~n12451 & n12452 ;
  assign n12454 = x75 & n8834 ;
  assign n12455 = x74 & n8829 ;
  assign n12456 = x73 & ~n8828 ;
  assign n12457 = n9159 & n12456 ;
  assign n12458 = n12455 | n12457 ;
  assign n12459 = n12454 | n12458 ;
  assign n12460 = n8837 | n12459 ;
  assign n12461 = ( n609 & n12459 ) | ( n609 & n12460 ) | ( n12459 & n12460 ) ;
  assign n12462 = x53 & n12461 ;
  assign n12463 = x53 & ~n12462 ;
  assign n12464 = ( n12461 & ~n12462 ) | ( n12461 & n12463 ) | ( ~n12462 & n12463 ) ;
  assign n12465 = n12453 | n12464 ;
  assign n12466 = n12453 & n12464 ;
  assign n12467 = n12465 & ~n12466 ;
  assign n12468 = n12032 | n12038 ;
  assign n12469 = n12467 & n12468 ;
  assign n12470 = n12467 | n12468 ;
  assign n12471 = ~n12469 & n12470 ;
  assign n12472 = x78 & n7812 ;
  assign n12473 = x77 & n7807 ;
  assign n12474 = x76 & ~n7806 ;
  assign n12475 = n8136 & n12474 ;
  assign n12476 = n12473 | n12475 ;
  assign n12477 = n12472 | n12476 ;
  assign n12478 = n7815 | n12477 ;
  assign n12479 = ( n868 & n12477 ) | ( n868 & n12478 ) | ( n12477 & n12478 ) ;
  assign n12480 = x50 & n12479 ;
  assign n12481 = x50 & ~n12480 ;
  assign n12482 = ( n12479 & ~n12480 ) | ( n12479 & n12481 ) | ( ~n12480 & n12481 ) ;
  assign n12483 = n12471 & n12482 ;
  assign n12484 = n12471 & ~n12483 ;
  assign n12485 = ~n12471 & n12482 ;
  assign n12486 = n12484 | n12485 ;
  assign n12487 = n12405 & n12486 ;
  assign n12488 = n12405 | n12486 ;
  assign n12489 = ~n12487 & n12488 ;
  assign n12490 = x81 & n6937 ;
  assign n12491 = x80 & n6932 ;
  assign n12492 = x79 & ~n6931 ;
  assign n12493 = n7216 & n12492 ;
  assign n12494 = n12491 | n12493 ;
  assign n12495 = n12490 | n12494 ;
  assign n12496 = n6940 | n12495 ;
  assign n12497 = ( n1256 & n12495 ) | ( n1256 & n12496 ) | ( n12495 & n12496 ) ;
  assign n12498 = x47 & n12497 ;
  assign n12499 = x47 & ~n12498 ;
  assign n12500 = ( n12497 & ~n12498 ) | ( n12497 & n12499 ) | ( ~n12498 & n12499 ) ;
  assign n12501 = n12489 & n12500 ;
  assign n12502 = n12489 & ~n12501 ;
  assign n12503 = ~n12489 & n12500 ;
  assign n12504 = n12502 | n12503 ;
  assign n12505 = n12404 & n12504 ;
  assign n12506 = n12404 & ~n12505 ;
  assign n12507 = n12504 & ~n12505 ;
  assign n12508 = n12506 | n12507 ;
  assign n12509 = ( n12402 & n12403 ) | ( n12402 & ~n12508 ) | ( n12403 & ~n12508 ) ;
  assign n12510 = ( ~n12403 & n12508 ) | ( ~n12403 & n12509 ) | ( n12508 & n12509 ) ;
  assign n12511 = ( ~n12402 & n12509 ) | ( ~n12402 & n12510 ) | ( n12509 & n12510 ) ;
  assign n12512 = n12391 & n12511 ;
  assign n12513 = n12391 | n12511 ;
  assign n12514 = ~n12512 & n12513 ;
  assign n12515 = n12105 | n12111 ;
  assign n12516 = n12514 | n12515 ;
  assign n12517 = n12514 & n12515 ;
  assign n12518 = n12516 & ~n12517 ;
  assign n12519 = x90 & n4572 ;
  assign n12520 = x89 & n4567 ;
  assign n12521 = x88 & ~n4566 ;
  assign n12522 = n4828 & n12521 ;
  assign n12523 = n12520 | n12522 ;
  assign n12524 = n12519 | n12523 ;
  assign n12525 = n4575 | n12524 ;
  assign n12526 = ( n2410 & n12524 ) | ( n2410 & n12525 ) | ( n12524 & n12525 ) ;
  assign n12527 = x38 & n12526 ;
  assign n12528 = x38 & ~n12527 ;
  assign n12529 = ( n12526 & ~n12527 ) | ( n12526 & n12528 ) | ( ~n12527 & n12528 ) ;
  assign n12530 = n12518 & n12529 ;
  assign n12531 = n12518 & ~n12530 ;
  assign n12532 = ~n12518 & n12529 ;
  assign n12533 = n12531 | n12532 ;
  assign n12534 = n12124 | n12130 ;
  assign n12535 = n12533 | n12534 ;
  assign n12536 = n12533 & n12534 ;
  assign n12537 = n12535 & ~n12536 ;
  assign n12538 = x93 & n3913 ;
  assign n12539 = x92 & n3908 ;
  assign n12540 = x91 & ~n3907 ;
  assign n12541 = n4152 & n12540 ;
  assign n12542 = n12539 | n12541 ;
  assign n12543 = n12538 | n12542 ;
  assign n12544 = n3916 | n12543 ;
  assign n12545 = ( n2931 & n12543 ) | ( n2931 & n12544 ) | ( n12543 & n12544 ) ;
  assign n12546 = x35 & n12545 ;
  assign n12547 = x35 & ~n12546 ;
  assign n12548 = ( n12545 & ~n12546 ) | ( n12545 & n12547 ) | ( ~n12546 & n12547 ) ;
  assign n12549 = n12537 & n12548 ;
  assign n12550 = n12537 & ~n12549 ;
  assign n12551 = ~n12537 & n12548 ;
  assign n12552 = n12550 | n12551 ;
  assign n12553 = n12143 | n12149 ;
  assign n12554 = n12552 | n12553 ;
  assign n12555 = n12552 & n12553 ;
  assign n12556 = n12554 & ~n12555 ;
  assign n12557 = x96 & n3314 ;
  assign n12558 = x95 & n3309 ;
  assign n12559 = x94 & ~n3308 ;
  assign n12560 = n3570 & n12559 ;
  assign n12561 = n12558 | n12560 ;
  assign n12562 = n12557 | n12561 ;
  assign n12563 = n3317 | n12562 ;
  assign n12564 = ( n3509 & n12562 ) | ( n3509 & n12563 ) | ( n12562 & n12563 ) ;
  assign n12565 = x32 & n12564 ;
  assign n12566 = x32 & ~n12565 ;
  assign n12567 = ( n12564 & ~n12565 ) | ( n12564 & n12566 ) | ( ~n12565 & n12566 ) ;
  assign n12568 = n12556 & n12567 ;
  assign n12569 = n12556 | n12567 ;
  assign n12570 = ~n12568 & n12569 ;
  assign n12571 = n12152 & n12570 ;
  assign n12572 = n12152 & ~n12571 ;
  assign n12573 = ( n12570 & ~n12571 ) | ( n12570 & n12572 ) | ( ~n12571 & n12572 ) ;
  assign n12574 = x99 & n2775 ;
  assign n12575 = x98 & n2770 ;
  assign n12576 = x97 & ~n2769 ;
  assign n12577 = n2978 & n12576 ;
  assign n12578 = n12575 | n12577 ;
  assign n12579 = n12574 | n12578 ;
  assign n12580 = n2778 | n12579 ;
  assign n12581 = ( n4325 & n12579 ) | ( n4325 & n12580 ) | ( n12579 & n12580 ) ;
  assign n12582 = x29 & n12581 ;
  assign n12583 = x29 & ~n12582 ;
  assign n12584 = ( n12581 & ~n12582 ) | ( n12581 & n12583 ) | ( ~n12582 & n12583 ) ;
  assign n12585 = n12573 & n12584 ;
  assign n12586 = n12573 & ~n12585 ;
  assign n12587 = ~n12573 & n12584 ;
  assign n12588 = n12586 | n12587 ;
  assign n12589 = n12155 | n12160 ;
  assign n12590 = n12588 | n12589 ;
  assign n12591 = n12588 & n12589 ;
  assign n12592 = n12590 & ~n12591 ;
  assign n12593 = x102 & n2280 ;
  assign n12594 = x101 & n2275 ;
  assign n12595 = x100 & ~n2274 ;
  assign n12596 = n2481 & n12595 ;
  assign n12597 = n12594 | n12596 ;
  assign n12598 = n12593 | n12597 ;
  assign n12599 = n2283 | n12598 ;
  assign n12600 = ( n5025 & n12598 ) | ( n5025 & n12599 ) | ( n12598 & n12599 ) ;
  assign n12601 = x26 & n12600 ;
  assign n12602 = x26 & ~n12601 ;
  assign n12603 = ( n12600 & ~n12601 ) | ( n12600 & n12602 ) | ( ~n12601 & n12602 ) ;
  assign n12604 = n12592 & n12603 ;
  assign n12605 = n12592 & ~n12604 ;
  assign n12606 = ~n12592 & n12603 ;
  assign n12607 = n12605 | n12606 ;
  assign n12608 = n12173 | n12179 ;
  assign n12609 = n12607 | n12608 ;
  assign n12610 = n12607 & n12608 ;
  assign n12611 = n12609 & ~n12610 ;
  assign n12612 = ( n12379 & n12380 ) | ( n12379 & ~n12611 ) | ( n12380 & ~n12611 ) ;
  assign n12613 = ( ~n12380 & n12611 ) | ( ~n12380 & n12612 ) | ( n12611 & n12612 ) ;
  assign n12614 = ( ~n12379 & n12612 ) | ( ~n12379 & n12613 ) | ( n12612 & n12613 ) ;
  assign n12615 = n12368 & n12614 ;
  assign n12616 = n12368 | n12614 ;
  assign n12617 = ~n12615 & n12616 ;
  assign n12618 = n12357 & ~n12617 ;
  assign n12619 = ~n12357 & n12617 ;
  assign n12620 = n12618 | n12619 ;
  assign n12621 = x111 & n1071 ;
  assign n12622 = x110 & n1066 ;
  assign n12623 = x109 & ~n1065 ;
  assign n12624 = n1189 & n12623 ;
  assign n12625 = n12622 | n12624 ;
  assign n12626 = n12621 | n12625 ;
  assign n12627 = n1074 | n12626 ;
  assign n12628 = ( n7492 & n12626 ) | ( n7492 & n12627 ) | ( n12626 & n12627 ) ;
  assign n12629 = x17 & n12628 ;
  assign n12630 = x17 & ~n12629 ;
  assign n12631 = ( n12628 & ~n12629 ) | ( n12628 & n12630 ) | ( ~n12629 & n12630 ) ;
  assign n12632 = n12620 & n12631 ;
  assign n12633 = n12620 | n12631 ;
  assign n12634 = ~n12632 & n12633 ;
  assign n12635 = n12230 | n12232 ;
  assign n12636 = n12634 & n12635 ;
  assign n12637 = n12634 | n12635 ;
  assign n12638 = ~n12636 & n12637 ;
  assign n12639 = n12247 | n12249 ;
  assign n12640 = ( n12356 & n12638 ) | ( n12356 & n12639 ) | ( n12638 & n12639 ) ;
  assign n12641 = ( n12638 & n12639 ) | ( n12638 & ~n12640 ) | ( n12639 & ~n12640 ) ;
  assign n12642 = ( n12356 & ~n12640 ) | ( n12356 & n12641 ) | ( ~n12640 & n12641 ) ;
  assign n12643 = n12345 & n12642 ;
  assign n12644 = n12345 | n12642 ;
  assign n12645 = ~n12643 & n12644 ;
  assign n12646 = n12264 | n12266 ;
  assign n12647 = n12645 & n12646 ;
  assign n12648 = n12645 | n12646 ;
  assign n12649 = ~n12647 & n12648 ;
  assign n12650 = x120 & n337 ;
  assign n12651 = x119 & n332 ;
  assign n12652 = x118 & ~n331 ;
  assign n12653 = n396 & n12652 ;
  assign n12654 = n12651 | n12653 ;
  assign n12655 = n12650 | n12654 ;
  assign n12656 = n340 | n12655 ;
  assign n12657 = ( n10460 & n12655 ) | ( n10460 & n12656 ) | ( n12655 & n12656 ) ;
  assign n12658 = x8 & n12657 ;
  assign n12659 = x8 & ~n12658 ;
  assign n12660 = ( n12657 & ~n12658 ) | ( n12657 & n12659 ) | ( ~n12658 & n12659 ) ;
  assign n12661 = n12649 | n12660 ;
  assign n12662 = x123 & n206 ;
  assign n12663 = x122 & n201 ;
  assign n12664 = x121 & ~n200 ;
  assign n12665 = n243 & n12664 ;
  assign n12666 = n12663 | n12665 ;
  assign n12667 = n12662 | n12666 ;
  assign n12668 = n209 | n12667 ;
  assign n12669 = ( n11219 & n12667 ) | ( n11219 & n12668 ) | ( n12667 & n12668 ) ;
  assign n12670 = x5 & n12669 ;
  assign n12671 = x5 & ~n12670 ;
  assign n12672 = ( n12669 & ~n12670 ) | ( n12669 & n12671 ) | ( ~n12670 & n12671 ) ;
  assign n12673 = ( n12660 & ~n12661 ) | ( n12660 & n12672 ) | ( ~n12661 & n12672 ) ;
  assign n12674 = ( n12649 & ~n12661 ) | ( n12649 & n12673 ) | ( ~n12661 & n12673 ) ;
  assign n12675 = n12334 | n12674 ;
  assign n12676 = ( n12649 & n12660 ) | ( n12649 & n12672 ) | ( n12660 & n12672 ) ;
  assign n12677 = n12661 & ~n12676 ;
  assign n12678 = n12675 | n12677 ;
  assign n12679 = ( n12334 & n12674 ) | ( n12334 & n12677 ) | ( n12674 & n12677 ) ;
  assign n12680 = n12678 & ~n12679 ;
  assign n12681 = x125 | x126 ;
  assign n12682 = x125 & x126 ;
  assign n12683 = n12681 & ~n12682 ;
  assign n12684 = n12301 | n12307 ;
  assign n12685 = n12683 & n12684 ;
  assign n12686 = n12683 | n12684 ;
  assign n12687 = ~n12685 & n12686 ;
  assign n12688 = x125 & n131 ;
  assign n12689 = x124 & ~n156 ;
  assign n12690 = ( n135 & n12688 ) | ( n135 & n12689 ) | ( n12688 & n12689 ) ;
  assign n12691 = x0 & x126 ;
  assign n12692 = ( ~n135 & n12688 ) | ( ~n135 & n12691 ) | ( n12688 & n12691 ) ;
  assign n12693 = n12690 | n12692 ;
  assign n12694 = n139 | n12693 ;
  assign n12695 = ( n12687 & n12693 ) | ( n12687 & n12694 ) | ( n12693 & n12694 ) ;
  assign n12696 = x2 & n12695 ;
  assign n12697 = x2 & ~n12696 ;
  assign n12698 = ( n12695 & ~n12696 ) | ( n12695 & n12697 ) | ( ~n12696 & n12697 ) ;
  assign n12699 = n12680 | n12698 ;
  assign n12700 = n12680 & n12698 ;
  assign n12701 = n12699 & ~n12700 ;
  assign n12702 = n12325 & n12701 ;
  assign n12703 = n12325 | n12701 ;
  assign n12704 = ~n12702 & n12703 ;
  assign n12705 = n12328 | n12331 ;
  assign n12706 = n12704 & n12705 ;
  assign n12707 = n12704 | n12705 ;
  assign n12708 = ~n12706 & n12707 ;
  assign n12709 = n12679 | n12700 ;
  assign n12710 = x126 & n131 ;
  assign n12711 = x125 & ~n156 ;
  assign n12712 = ( n135 & n12710 ) | ( n135 & n12711 ) | ( n12710 & n12711 ) ;
  assign n12713 = x0 & x127 ;
  assign n12714 = ( ~n135 & n12710 ) | ( ~n135 & n12713 ) | ( n12710 & n12713 ) ;
  assign n12715 = n12712 | n12714 ;
  assign n12716 = n139 | n12715 ;
  assign n12717 = ( x125 & x126 ) | ( x125 & n12684 ) | ( x126 & n12684 ) ;
  assign n12718 = ( x126 & ~x127 ) | ( x126 & n12717 ) | ( ~x127 & n12717 ) ;
  assign n12719 = ( x127 & ~n12717 ) | ( x127 & n12718 ) | ( ~n12717 & n12718 ) ;
  assign n12720 = ( ~x126 & n12718 ) | ( ~x126 & n12719 ) | ( n12718 & n12719 ) ;
  assign n12721 = ( n12715 & n12716 ) | ( n12715 & n12720 ) | ( n12716 & n12720 ) ;
  assign n12722 = x2 & n12721 ;
  assign n12723 = x2 & ~n12722 ;
  assign n12724 = ( n12721 & ~n12722 ) | ( n12721 & n12723 ) | ( ~n12722 & n12723 ) ;
  assign n12725 = x124 & n206 ;
  assign n12726 = x123 & n201 ;
  assign n12727 = x122 & ~n200 ;
  assign n12728 = n243 & n12727 ;
  assign n12729 = n12726 | n12728 ;
  assign n12730 = n12725 | n12729 ;
  assign n12731 = n209 | n12730 ;
  assign n12732 = ( n11916 & n12730 ) | ( n11916 & n12731 ) | ( n12730 & n12731 ) ;
  assign n12733 = x5 & n12732 ;
  assign n12734 = x5 & ~n12733 ;
  assign n12735 = ( n12732 & ~n12733 ) | ( n12732 & n12734 ) | ( ~n12733 & n12734 ) ;
  assign n12736 = n12632 | n12636 ;
  assign n12737 = x100 & n2775 ;
  assign n12738 = x99 & n2770 ;
  assign n12739 = x98 & ~n2769 ;
  assign n12740 = n2978 & n12739 ;
  assign n12741 = n12738 | n12740 ;
  assign n12742 = n12737 | n12741 ;
  assign n12743 = n2778 | n12742 ;
  assign n12744 = ( n4532 & n12742 ) | ( n4532 & n12743 ) | ( n12742 & n12743 ) ;
  assign n12745 = x29 & n12744 ;
  assign n12746 = x29 & ~n12745 ;
  assign n12747 = ( n12744 & ~n12745 ) | ( n12744 & n12746 ) | ( ~n12745 & n12746 ) ;
  assign n12748 = x97 & n3314 ;
  assign n12749 = x96 & n3309 ;
  assign n12750 = x95 & ~n3308 ;
  assign n12751 = n3570 & n12750 ;
  assign n12752 = n12749 | n12751 ;
  assign n12753 = n12748 | n12752 ;
  assign n12754 = n3317 | n12753 ;
  assign n12755 = ( n3707 & n12753 ) | ( n3707 & n12754 ) | ( n12753 & n12754 ) ;
  assign n12756 = x32 & n12755 ;
  assign n12757 = x32 & ~n12756 ;
  assign n12758 = ( n12755 & ~n12756 ) | ( n12755 & n12757 ) | ( ~n12756 & n12757 ) ;
  assign n12759 = n12568 | n12571 ;
  assign n12760 = n12501 | n12505 ;
  assign n12761 = x76 & n8834 ;
  assign n12762 = x75 & n8829 ;
  assign n12763 = x74 & ~n8828 ;
  assign n12764 = n9159 & n12763 ;
  assign n12765 = n12762 | n12764 ;
  assign n12766 = n12761 | n12765 ;
  assign n12767 = n8837 | n12766 ;
  assign n12768 = ( n740 & n12766 ) | ( n740 & n12767 ) | ( n12766 & n12767 ) ;
  assign n12769 = x53 & n12768 ;
  assign n12770 = x53 & ~n12769 ;
  assign n12771 = ( n12768 & ~n12769 ) | ( n12768 & n12770 ) | ( ~n12769 & n12770 ) ;
  assign n12772 = x73 & n9853 ;
  assign n12773 = x72 & n9848 ;
  assign n12774 = x71 & ~n9847 ;
  assign n12775 = n10165 & n12774 ;
  assign n12776 = n12773 | n12775 ;
  assign n12777 = n12772 | n12776 ;
  assign n12778 = ( n499 & n9856 ) | ( n499 & n12777 ) | ( n9856 & n12777 ) ;
  assign n12779 = ( x56 & ~n12777 ) | ( x56 & n12778 ) | ( ~n12777 & n12778 ) ;
  assign n12780 = ~n12778 & n12779 ;
  assign n12781 = n12777 | n12779 ;
  assign n12782 = ( ~x56 & n12780 ) | ( ~x56 & n12781 ) | ( n12780 & n12781 ) ;
  assign n12783 = n12448 | n12451 ;
  assign n12784 = x70 & n10876 ;
  assign n12785 = x69 & n10871 ;
  assign n12786 = x68 & ~n10870 ;
  assign n12787 = n11305 & n12786 ;
  assign n12788 = n12785 | n12787 ;
  assign n12789 = n12784 | n12788 ;
  assign n12790 = n10879 | n12789 ;
  assign n12791 = ( n310 & n12789 ) | ( n310 & n12790 ) | ( n12789 & n12790 ) ;
  assign n12792 = x59 & ~n12791 ;
  assign n12793 = ~x59 & n12791 ;
  assign n12794 = n12792 | n12793 ;
  assign n12795 = x67 & n11984 ;
  assign n12796 = x66 & n11979 ;
  assign n12797 = x65 & ~n11978 ;
  assign n12798 = n12430 & n12797 ;
  assign n12799 = n12796 | n12798 ;
  assign n12800 = n12795 | n12799 ;
  assign n12801 = n180 & n11987 ;
  assign n12802 = n12800 | n12801 ;
  assign n12803 = x62 & ~n12802 ;
  assign n12804 = ~x62 & n12802 ;
  assign n12805 = n12803 | n12804 ;
  assign n12806 = x62 & ~x63 ;
  assign n12807 = ~x62 & x63 ;
  assign n12808 = n12806 | n12807 ;
  assign n12809 = x64 & n12808 ;
  assign n12810 = n12441 & n12809 ;
  assign n12811 = n12441 & ~n12810 ;
  assign n12812 = ( n12809 & ~n12810 ) | ( n12809 & n12811 ) | ( ~n12810 & n12811 ) ;
  assign n12813 = n12805 & n12812 ;
  assign n12814 = n12805 | n12812 ;
  assign n12815 = ~n12813 & n12814 ;
  assign n12816 = n12794 | n12815 ;
  assign n12817 = n12794 & n12815 ;
  assign n12818 = n12816 & ~n12817 ;
  assign n12819 = n12444 & n12818 ;
  assign n12820 = n12444 | n12818 ;
  assign n12821 = ~n12819 & n12820 ;
  assign n12822 = ( n12782 & n12783 ) | ( n12782 & ~n12821 ) | ( n12783 & ~n12821 ) ;
  assign n12823 = ( ~n12783 & n12821 ) | ( ~n12783 & n12822 ) | ( n12821 & n12822 ) ;
  assign n12824 = ( ~n12782 & n12822 ) | ( ~n12782 & n12823 ) | ( n12822 & n12823 ) ;
  assign n12825 = n12771 | n12824 ;
  assign n12826 = n12771 & n12824 ;
  assign n12827 = n12825 & ~n12826 ;
  assign n12828 = n12466 | n12469 ;
  assign n12829 = n12827 & n12828 ;
  assign n12830 = n12827 | n12828 ;
  assign n12831 = ~n12829 & n12830 ;
  assign n12832 = x79 & n7812 ;
  assign n12833 = x78 & n7807 ;
  assign n12834 = x77 & ~n7806 ;
  assign n12835 = n8136 & n12834 ;
  assign n12836 = n12833 | n12835 ;
  assign n12837 = n12832 | n12836 ;
  assign n12838 = n7815 | n12837 ;
  assign n12839 = ( n961 & n12837 ) | ( n961 & n12838 ) | ( n12837 & n12838 ) ;
  assign n12840 = x50 & n12839 ;
  assign n12841 = x50 & ~n12840 ;
  assign n12842 = ( n12839 & ~n12840 ) | ( n12839 & n12841 ) | ( ~n12840 & n12841 ) ;
  assign n12843 = n12831 & n12842 ;
  assign n12844 = n12831 & ~n12843 ;
  assign n12845 = ~n12831 & n12842 ;
  assign n12846 = n12844 | n12845 ;
  assign n12847 = n12483 | n12487 ;
  assign n12848 = n12846 | n12847 ;
  assign n12849 = n12846 & n12847 ;
  assign n12850 = n12848 & ~n12849 ;
  assign n12851 = x82 & n6937 ;
  assign n12852 = x81 & n6932 ;
  assign n12853 = x80 & ~n6931 ;
  assign n12854 = n7216 & n12853 ;
  assign n12855 = n12852 | n12854 ;
  assign n12856 = n12851 | n12855 ;
  assign n12857 = n6940 | n12856 ;
  assign n12858 = ( n1371 & n12856 ) | ( n1371 & n12857 ) | ( n12856 & n12857 ) ;
  assign n12859 = x47 & n12858 ;
  assign n12860 = x47 & ~n12859 ;
  assign n12861 = ( n12858 & ~n12859 ) | ( n12858 & n12860 ) | ( ~n12859 & n12860 ) ;
  assign n12862 = n12850 | n12861 ;
  assign n12863 = n12850 & n12861 ;
  assign n12864 = n12862 & ~n12863 ;
  assign n12865 = n12760 & n12864 ;
  assign n12866 = n12760 | n12864 ;
  assign n12867 = ~n12865 & n12866 ;
  assign n12868 = x85 & n6068 ;
  assign n12869 = x84 & n6063 ;
  assign n12870 = x83 & ~n6062 ;
  assign n12871 = n6398 & n12870 ;
  assign n12872 = n12869 | n12871 ;
  assign n12873 = n12868 | n12872 ;
  assign n12874 = n6071 | n12873 ;
  assign n12875 = ( n1765 & n12873 ) | ( n1765 & n12874 ) | ( n12873 & n12874 ) ;
  assign n12876 = x44 & n12875 ;
  assign n12877 = x44 & ~n12876 ;
  assign n12878 = ( n12875 & ~n12876 ) | ( n12875 & n12877 ) | ( ~n12876 & n12877 ) ;
  assign n12879 = n12867 & n12878 ;
  assign n12880 = n12867 | n12878 ;
  assign n12881 = ~n12879 & n12880 ;
  assign n12882 = ( n12402 & n12403 ) | ( n12402 & n12508 ) | ( n12403 & n12508 ) ;
  assign n12883 = n12881 | n12882 ;
  assign n12884 = n12881 & n12882 ;
  assign n12885 = n12883 & ~n12884 ;
  assign n12886 = x88 & n5340 ;
  assign n12887 = x87 & n5335 ;
  assign n12888 = x86 & ~n5334 ;
  assign n12889 = n5580 & n12888 ;
  assign n12890 = n12887 | n12889 ;
  assign n12891 = n12886 | n12890 ;
  assign n12892 = n5343 | n12891 ;
  assign n12893 = ( n2095 & n12891 ) | ( n2095 & n12892 ) | ( n12891 & n12892 ) ;
  assign n12894 = x41 & n12893 ;
  assign n12895 = x41 & ~n12894 ;
  assign n12896 = ( n12893 & ~n12894 ) | ( n12893 & n12895 ) | ( ~n12894 & n12895 ) ;
  assign n12897 = n12885 & n12896 ;
  assign n12898 = n12885 & ~n12897 ;
  assign n12899 = ~n12885 & n12896 ;
  assign n12900 = n12898 | n12899 ;
  assign n12901 = n12512 | n12517 ;
  assign n12902 = n12900 | n12901 ;
  assign n12903 = n12900 & n12901 ;
  assign n12904 = n12902 & ~n12903 ;
  assign n12905 = x91 & n4572 ;
  assign n12906 = x90 & n4567 ;
  assign n12907 = x89 & ~n4566 ;
  assign n12908 = n4828 & n12907 ;
  assign n12909 = n12906 | n12908 ;
  assign n12910 = n12905 | n12909 ;
  assign n12911 = n4575 | n12910 ;
  assign n12912 = ( n2714 & n12910 ) | ( n2714 & n12911 ) | ( n12910 & n12911 ) ;
  assign n12913 = x38 & n12912 ;
  assign n12914 = x38 & ~n12913 ;
  assign n12915 = ( n12912 & ~n12913 ) | ( n12912 & n12914 ) | ( ~n12913 & n12914 ) ;
  assign n12916 = n12904 & n12915 ;
  assign n12917 = n12904 & ~n12916 ;
  assign n12918 = ~n12904 & n12915 ;
  assign n12919 = n12917 | n12918 ;
  assign n12920 = n12530 | n12536 ;
  assign n12921 = n12919 | n12920 ;
  assign n12922 = n12919 & n12920 ;
  assign n12923 = n12921 & ~n12922 ;
  assign n12924 = x94 & n3913 ;
  assign n12925 = x93 & n3908 ;
  assign n12926 = x92 & ~n3907 ;
  assign n12927 = n4152 & n12926 ;
  assign n12928 = n12925 | n12927 ;
  assign n12929 = n12924 | n12928 ;
  assign n12930 = n3916 | n12929 ;
  assign n12931 = ( n3271 & n12929 ) | ( n3271 & n12930 ) | ( n12929 & n12930 ) ;
  assign n12932 = x35 & n12931 ;
  assign n12933 = x35 & ~n12932 ;
  assign n12934 = ( n12931 & ~n12932 ) | ( n12931 & n12933 ) | ( ~n12932 & n12933 ) ;
  assign n12935 = n12923 | n12934 ;
  assign n12936 = n12923 & n12934 ;
  assign n12937 = n12935 & ~n12936 ;
  assign n12938 = n12549 | n12937 ;
  assign n12939 = n12555 | n12938 ;
  assign n12940 = ( n12549 & n12555 ) | ( n12549 & n12937 ) | ( n12555 & n12937 ) ;
  assign n12941 = n12939 & ~n12940 ;
  assign n12942 = ( n12758 & n12759 ) | ( n12758 & ~n12941 ) | ( n12759 & ~n12941 ) ;
  assign n12943 = ( ~n12759 & n12941 ) | ( ~n12759 & n12942 ) | ( n12941 & n12942 ) ;
  assign n12944 = ( ~n12758 & n12942 ) | ( ~n12758 & n12943 ) | ( n12942 & n12943 ) ;
  assign n12945 = n12747 & n12944 ;
  assign n12946 = n12747 | n12944 ;
  assign n12947 = ~n12945 & n12946 ;
  assign n12948 = n12585 | n12591 ;
  assign n12949 = n12947 | n12948 ;
  assign n12950 = n12947 & n12948 ;
  assign n12951 = n12949 & ~n12950 ;
  assign n12952 = x103 & n2280 ;
  assign n12953 = x102 & n2275 ;
  assign n12954 = x101 & ~n2274 ;
  assign n12955 = n2481 & n12954 ;
  assign n12956 = n12953 | n12955 ;
  assign n12957 = n12952 | n12956 ;
  assign n12958 = n2283 | n12957 ;
  assign n12959 = ( n5264 & n12957 ) | ( n5264 & n12958 ) | ( n12957 & n12958 ) ;
  assign n12960 = x26 & n12959 ;
  assign n12961 = x26 & ~n12960 ;
  assign n12962 = ( n12959 & ~n12960 ) | ( n12959 & n12961 ) | ( ~n12960 & n12961 ) ;
  assign n12963 = n12951 | n12962 ;
  assign n12964 = n12951 & n12962 ;
  assign n12965 = n12963 & ~n12964 ;
  assign n12966 = n12604 | n12610 ;
  assign n12967 = n12965 & n12966 ;
  assign n12968 = n12965 | n12966 ;
  assign n12969 = ~n12967 & n12968 ;
  assign n12970 = x106 & n1817 ;
  assign n12971 = x105 & n1812 ;
  assign n12972 = x104 & ~n1811 ;
  assign n12973 = n1977 & n12972 ;
  assign n12974 = n12971 | n12973 ;
  assign n12975 = n12970 | n12974 ;
  assign n12976 = n1820 | n12975 ;
  assign n12977 = ( n5814 & n12975 ) | ( n5814 & n12976 ) | ( n12975 & n12976 ) ;
  assign n12978 = x23 & n12977 ;
  assign n12979 = x23 & ~n12978 ;
  assign n12980 = ( n12977 & ~n12978 ) | ( n12977 & n12979 ) | ( ~n12978 & n12979 ) ;
  assign n12981 = n12969 & n12980 ;
  assign n12982 = n12969 & ~n12981 ;
  assign n12983 = ~n12969 & n12980 ;
  assign n12984 = n12982 | n12983 ;
  assign n12985 = ( n12379 & n12380 ) | ( n12379 & n12611 ) | ( n12380 & n12611 ) ;
  assign n12986 = n12984 & n12985 ;
  assign n12987 = n12984 | n12985 ;
  assign n12988 = ~n12986 & n12987 ;
  assign n12989 = x109 & n1421 ;
  assign n12990 = x108 & n1416 ;
  assign n12991 = x107 & ~n1415 ;
  assign n12992 = n1584 & n12991 ;
  assign n12993 = n12990 | n12992 ;
  assign n12994 = n12989 | n12993 ;
  assign n12995 = n1424 | n12994 ;
  assign n12996 = ( n6884 & n12994 ) | ( n6884 & n12995 ) | ( n12994 & n12995 ) ;
  assign n12997 = x20 & n12996 ;
  assign n12998 = x20 & ~n12997 ;
  assign n12999 = ( n12996 & ~n12997 ) | ( n12996 & n12998 ) | ( ~n12997 & n12998 ) ;
  assign n13000 = n12988 & n12999 ;
  assign n13001 = n12988 & ~n13000 ;
  assign n13002 = ~n12988 & n12999 ;
  assign n13003 = n13001 | n13002 ;
  assign n13004 = ( n12615 & n12617 ) | ( n12615 & ~n12619 ) | ( n12617 & ~n12619 ) ;
  assign n13005 = n13003 & n13004 ;
  assign n13006 = n13003 | n13004 ;
  assign n13007 = ~n13005 & n13006 ;
  assign n13008 = x112 & n1071 ;
  assign n13009 = x111 & n1066 ;
  assign n13010 = x110 & ~n1065 ;
  assign n13011 = n1189 & n13010 ;
  assign n13012 = n13009 | n13011 ;
  assign n13013 = n13008 | n13012 ;
  assign n13014 = n1074 | n13013 ;
  assign n13015 = ( n7789 & n13013 ) | ( n7789 & n13014 ) | ( n13013 & n13014 ) ;
  assign n13016 = x17 & n13015 ;
  assign n13017 = x17 & ~n13016 ;
  assign n13018 = ( n13015 & ~n13016 ) | ( n13015 & n13017 ) | ( ~n13016 & n13017 ) ;
  assign n13019 = n13007 & n13018 ;
  assign n13020 = n13007 & ~n13019 ;
  assign n13021 = ~n13007 & n13018 ;
  assign n13022 = n13020 | n13021 ;
  assign n13023 = n12736 & n13022 ;
  assign n13024 = n12736 | n13022 ;
  assign n13025 = ~n13023 & n13024 ;
  assign n13026 = x115 & n771 ;
  assign n13027 = x114 & n766 ;
  assign n13028 = x113 & ~n765 ;
  assign n13029 = n905 & n13028 ;
  assign n13030 = n13027 | n13029 ;
  assign n13031 = n13026 | n13030 ;
  assign n13032 = n774 | n13031 ;
  assign n13033 = ( n8749 & n13031 ) | ( n8749 & n13032 ) | ( n13031 & n13032 ) ;
  assign n13034 = x14 & n13033 ;
  assign n13035 = x14 & ~n13034 ;
  assign n13036 = ( n13033 & ~n13034 ) | ( n13033 & n13035 ) | ( ~n13034 & n13035 ) ;
  assign n13037 = n13025 & n13036 ;
  assign n13038 = n13025 | n13036 ;
  assign n13039 = ~n13037 & n13038 ;
  assign n13040 = n12640 | n13039 ;
  assign n13041 = n12640 & n13039 ;
  assign n13042 = n13040 & ~n13041 ;
  assign n13043 = x118 & n528 ;
  assign n13044 = x117 & n523 ;
  assign n13045 = x116 & ~n522 ;
  assign n13046 = n635 & n13045 ;
  assign n13047 = n13044 | n13046 ;
  assign n13048 = n13043 | n13047 ;
  assign n13049 = n531 | n13048 ;
  assign n13050 = ( n9760 & n13048 ) | ( n9760 & n13049 ) | ( n13048 & n13049 ) ;
  assign n13051 = x11 & n13050 ;
  assign n13052 = x11 & ~n13051 ;
  assign n13053 = ( n13050 & ~n13051 ) | ( n13050 & n13052 ) | ( ~n13051 & n13052 ) ;
  assign n13054 = n13042 & n13053 ;
  assign n13055 = n13042 & ~n13054 ;
  assign n13056 = ~n13042 & n13053 ;
  assign n13057 = n13055 | n13056 ;
  assign n13058 = n12643 | n12647 ;
  assign n13059 = n13057 | n13058 ;
  assign n13060 = n13057 & n13058 ;
  assign n13061 = n13059 & ~n13060 ;
  assign n13062 = x121 & n337 ;
  assign n13063 = x120 & n332 ;
  assign n13064 = x119 & ~n331 ;
  assign n13065 = n396 & n13064 ;
  assign n13066 = n13063 | n13065 ;
  assign n13067 = n13062 | n13066 ;
  assign n13068 = n340 | n13067 ;
  assign n13069 = ( n10811 & n13067 ) | ( n10811 & n13068 ) | ( n13067 & n13068 ) ;
  assign n13070 = x8 & n13069 ;
  assign n13071 = x8 & ~n13070 ;
  assign n13072 = ( n13069 & ~n13070 ) | ( n13069 & n13071 ) | ( ~n13070 & n13071 ) ;
  assign n13073 = ( n12735 & n13061 ) | ( n12735 & ~n13072 ) | ( n13061 & ~n13072 ) ;
  assign n13074 = ( ~n13061 & n13072 ) | ( ~n13061 & n13073 ) | ( n13072 & n13073 ) ;
  assign n13075 = ( ~n12735 & n13073 ) | ( ~n12735 & n13074 ) | ( n13073 & n13074 ) ;
  assign n13076 = ( n12676 & n12724 ) | ( n12676 & ~n13075 ) | ( n12724 & ~n13075 ) ;
  assign n13077 = ( ~n12676 & n13075 ) | ( ~n12676 & n13076 ) | ( n13075 & n13076 ) ;
  assign n13078 = ( ~n12724 & n13076 ) | ( ~n12724 & n13077 ) | ( n13076 & n13077 ) ;
  assign n13079 = n12709 & n13078 ;
  assign n13080 = n12709 | n13078 ;
  assign n13081 = ~n13079 & n13080 ;
  assign n13082 = n12702 | n12706 ;
  assign n13083 = n13081 & n13082 ;
  assign n13084 = n13081 | n13082 ;
  assign n13085 = ~n13083 & n13084 ;
  assign n13086 = n13079 | n13083 ;
  assign n13087 = ( n12676 & n12724 ) | ( n12676 & n13075 ) | ( n12724 & n13075 ) ;
  assign n13088 = x125 & n206 ;
  assign n13089 = x124 & n201 ;
  assign n13090 = x123 & ~n200 ;
  assign n13091 = n243 & n13090 ;
  assign n13092 = n13089 | n13091 ;
  assign n13093 = n13088 | n13092 ;
  assign n13094 = n209 | n13093 ;
  assign n13095 = ( n12310 & n13093 ) | ( n12310 & n13094 ) | ( n13093 & n13094 ) ;
  assign n13096 = x5 & n13095 ;
  assign n13097 = x5 & ~n13096 ;
  assign n13098 = ( n13095 & ~n13096 ) | ( n13095 & n13097 ) | ( ~n13096 & n13097 ) ;
  assign n13099 = n13019 | n13023 ;
  assign n13100 = n13000 | n13005 ;
  assign n13101 = n12981 | n12986 ;
  assign n13102 = x107 & n1817 ;
  assign n13103 = x106 & n1812 ;
  assign n13104 = x105 & ~n1811 ;
  assign n13105 = n1977 & n13104 ;
  assign n13106 = n13103 | n13105 ;
  assign n13107 = n13102 | n13106 ;
  assign n13108 = n1820 | n13107 ;
  assign n13109 = ( n6328 & n13107 ) | ( n6328 & n13108 ) | ( n13107 & n13108 ) ;
  assign n13110 = x23 & n13109 ;
  assign n13111 = x23 & ~n13110 ;
  assign n13112 = ( n13109 & ~n13110 ) | ( n13109 & n13111 ) | ( ~n13110 & n13111 ) ;
  assign n13113 = n229 & n11987 ;
  assign n13114 = x68 & n11984 ;
  assign n13115 = x67 & n11979 ;
  assign n13116 = x66 & ~n11978 ;
  assign n13117 = n12430 & n13116 ;
  assign n13118 = n13115 | n13117 ;
  assign n13119 = n13114 | n13118 ;
  assign n13120 = n13113 | n13119 ;
  assign n13121 = x62 | n13120 ;
  assign n13122 = ~x62 & n13121 ;
  assign n13123 = ( ~n13120 & n13121 ) | ( ~n13120 & n13122 ) | ( n13121 & n13122 ) ;
  assign n13124 = x65 & n12808 ;
  assign n13125 = x63 & x64 ;
  assign n13126 = ~n12808 & n13125 ;
  assign n13127 = n13124 | n13126 ;
  assign n13128 = n13123 & n13127 ;
  assign n13129 = n13123 & ~n13128 ;
  assign n13130 = ~n13123 & n13127 ;
  assign n13131 = n13129 | n13130 ;
  assign n13132 = n12810 | n12813 ;
  assign n13133 = n13131 | n13132 ;
  assign n13134 = n13131 & n13132 ;
  assign n13135 = n13133 & ~n13134 ;
  assign n13136 = x71 & n10876 ;
  assign n13137 = x70 & n10871 ;
  assign n13138 = x69 & ~n10870 ;
  assign n13139 = n11305 & n13138 ;
  assign n13140 = n13137 | n13139 ;
  assign n13141 = n13136 | n13140 ;
  assign n13142 = n10879 | n13141 ;
  assign n13143 = ( n376 & n13141 ) | ( n376 & n13142 ) | ( n13141 & n13142 ) ;
  assign n13144 = x59 & ~n13143 ;
  assign n13145 = ~x59 & n13143 ;
  assign n13146 = n13144 | n13145 ;
  assign n13147 = n13135 | n13146 ;
  assign n13148 = n13135 & n13146 ;
  assign n13149 = n13147 & ~n13148 ;
  assign n13150 = n12817 | n12819 ;
  assign n13151 = n13149 & n13150 ;
  assign n13152 = n13149 | n13150 ;
  assign n13153 = ~n13151 & n13152 ;
  assign n13154 = x74 & n9853 ;
  assign n13155 = x73 & n9848 ;
  assign n13156 = x72 & ~n9847 ;
  assign n13157 = n10165 & n13156 ;
  assign n13158 = n13155 | n13157 ;
  assign n13159 = n13154 | n13158 ;
  assign n13160 = n9856 | n13159 ;
  assign n13161 = ( n587 & n13159 ) | ( n587 & n13160 ) | ( n13159 & n13160 ) ;
  assign n13162 = x56 & n13161 ;
  assign n13163 = x56 & ~n13162 ;
  assign n13164 = ( n13161 & ~n13162 ) | ( n13161 & n13163 ) | ( ~n13162 & n13163 ) ;
  assign n13165 = n13153 & n13164 ;
  assign n13166 = n13153 & ~n13165 ;
  assign n13167 = ~n13153 & n13164 ;
  assign n13168 = n13166 | n13167 ;
  assign n13169 = ( n12782 & n12783 ) | ( n12782 & n12821 ) | ( n12783 & n12821 ) ;
  assign n13170 = n13168 | n13169 ;
  assign n13171 = n13168 & n13169 ;
  assign n13172 = n13170 & ~n13171 ;
  assign n13173 = x77 & n8834 ;
  assign n13174 = x76 & n8829 ;
  assign n13175 = x75 & ~n8828 ;
  assign n13176 = n9159 & n13175 ;
  assign n13177 = n13174 | n13176 ;
  assign n13178 = n13173 | n13177 ;
  assign n13179 = n8837 | n13178 ;
  assign n13180 = ( n846 & n13178 ) | ( n846 & n13179 ) | ( n13178 & n13179 ) ;
  assign n13181 = x53 & n13180 ;
  assign n13182 = x53 & ~n13181 ;
  assign n13183 = ( n13180 & ~n13181 ) | ( n13180 & n13182 ) | ( ~n13181 & n13182 ) ;
  assign n13184 = n13172 | n13183 ;
  assign n13185 = n13172 & n13183 ;
  assign n13186 = n13184 & ~n13185 ;
  assign n13187 = n12826 | n12829 ;
  assign n13188 = n13186 & n13187 ;
  assign n13189 = n13186 | n13187 ;
  assign n13190 = ~n13188 & n13189 ;
  assign n13191 = x80 & n7812 ;
  assign n13192 = x79 & n7807 ;
  assign n13193 = x78 & ~n7806 ;
  assign n13194 = n8136 & n13193 ;
  assign n13195 = n13192 | n13194 ;
  assign n13196 = n13191 | n13195 ;
  assign n13197 = n7815 | n13196 ;
  assign n13198 = ( n1147 & n13196 ) | ( n1147 & n13197 ) | ( n13196 & n13197 ) ;
  assign n13199 = x50 & n13198 ;
  assign n13200 = x50 & ~n13199 ;
  assign n13201 = ( n13198 & ~n13199 ) | ( n13198 & n13200 ) | ( ~n13199 & n13200 ) ;
  assign n13202 = n13190 & n13201 ;
  assign n13203 = n13190 & ~n13202 ;
  assign n13204 = ~n13190 & n13201 ;
  assign n13205 = n13203 | n13204 ;
  assign n13206 = n12843 | n12849 ;
  assign n13207 = n13205 | n13206 ;
  assign n13208 = n13205 & n13206 ;
  assign n13209 = n13207 & ~n13208 ;
  assign n13210 = x83 & n6937 ;
  assign n13211 = x82 & n6932 ;
  assign n13212 = x81 & ~n6931 ;
  assign n13213 = n7216 & n13212 ;
  assign n13214 = n13211 | n13213 ;
  assign n13215 = n13210 | n13214 ;
  assign n13216 = n6940 | n13215 ;
  assign n13217 = ( n1510 & n13215 ) | ( n1510 & n13216 ) | ( n13215 & n13216 ) ;
  assign n13218 = x47 & n13217 ;
  assign n13219 = x47 & ~n13218 ;
  assign n13220 = ( n13217 & ~n13218 ) | ( n13217 & n13219 ) | ( ~n13218 & n13219 ) ;
  assign n13221 = n13209 | n13220 ;
  assign n13222 = n13209 & n13220 ;
  assign n13223 = n13221 & ~n13222 ;
  assign n13224 = n12863 | n12865 ;
  assign n13225 = n13223 & n13224 ;
  assign n13226 = n13223 | n13224 ;
  assign n13227 = ~n13225 & n13226 ;
  assign n13228 = x86 & n6068 ;
  assign n13229 = x85 & n6063 ;
  assign n13230 = x84 & ~n6062 ;
  assign n13231 = n6398 & n13230 ;
  assign n13232 = n13229 | n13231 ;
  assign n13233 = n13228 | n13232 ;
  assign n13234 = n6071 | n13233 ;
  assign n13235 = ( n1921 & n13233 ) | ( n1921 & n13234 ) | ( n13233 & n13234 ) ;
  assign n13236 = x44 & n13235 ;
  assign n13237 = x44 & ~n13236 ;
  assign n13238 = ( n13235 & ~n13236 ) | ( n13235 & n13237 ) | ( ~n13236 & n13237 ) ;
  assign n13239 = n13227 & n13238 ;
  assign n13240 = n13227 & ~n13239 ;
  assign n13241 = ~n13227 & n13238 ;
  assign n13242 = n13240 | n13241 ;
  assign n13243 = n12879 | n12884 ;
  assign n13244 = n13242 | n13243 ;
  assign n13245 = n13242 & n13243 ;
  assign n13246 = n13244 & ~n13245 ;
  assign n13247 = x89 & n5340 ;
  assign n13248 = x88 & n5335 ;
  assign n13249 = x87 & ~n5334 ;
  assign n13250 = n5580 & n13249 ;
  assign n13251 = n13248 | n13250 ;
  assign n13252 = n13247 | n13251 ;
  assign n13253 = n5343 | n13252 ;
  assign n13254 = ( n2244 & n13252 ) | ( n2244 & n13253 ) | ( n13252 & n13253 ) ;
  assign n13255 = x41 & n13254 ;
  assign n13256 = x41 & ~n13255 ;
  assign n13257 = ( n13254 & ~n13255 ) | ( n13254 & n13256 ) | ( ~n13255 & n13256 ) ;
  assign n13258 = n13246 & n13257 ;
  assign n13259 = n13246 & ~n13258 ;
  assign n13260 = ~n13246 & n13257 ;
  assign n13261 = n13259 | n13260 ;
  assign n13262 = n12897 | n12903 ;
  assign n13263 = n13261 | n13262 ;
  assign n13264 = n13261 & n13262 ;
  assign n13265 = n13263 & ~n13264 ;
  assign n13266 = x92 & n4572 ;
  assign n13267 = x91 & n4567 ;
  assign n13268 = x90 & ~n4566 ;
  assign n13269 = n4828 & n13268 ;
  assign n13270 = n13267 | n13269 ;
  assign n13271 = n13266 | n13270 ;
  assign n13272 = n4575 | n13271 ;
  assign n13273 = ( n2904 & n13271 ) | ( n2904 & n13272 ) | ( n13271 & n13272 ) ;
  assign n13274 = x38 & n13273 ;
  assign n13275 = x38 & ~n13274 ;
  assign n13276 = ( n13273 & ~n13274 ) | ( n13273 & n13275 ) | ( ~n13274 & n13275 ) ;
  assign n13277 = n13265 & n13276 ;
  assign n13278 = n13265 & ~n13277 ;
  assign n13279 = ~n13265 & n13276 ;
  assign n13280 = n13278 | n13279 ;
  assign n13281 = n12916 | n12922 ;
  assign n13282 = n13280 | n13281 ;
  assign n13283 = n13280 & n13281 ;
  assign n13284 = n13282 & ~n13283 ;
  assign n13285 = x95 & n3913 ;
  assign n13286 = x94 & n3908 ;
  assign n13287 = x93 & ~n3907 ;
  assign n13288 = n4152 & n13287 ;
  assign n13289 = n13286 | n13288 ;
  assign n13290 = n13285 | n13289 ;
  assign n13291 = n3916 | n13290 ;
  assign n13292 = ( n3479 & n13290 ) | ( n3479 & n13291 ) | ( n13290 & n13291 ) ;
  assign n13293 = x35 & n13292 ;
  assign n13294 = x35 & ~n13293 ;
  assign n13295 = ( n13292 & ~n13293 ) | ( n13292 & n13294 ) | ( ~n13293 & n13294 ) ;
  assign n13296 = n13284 | n13295 ;
  assign n13297 = n13284 & n13295 ;
  assign n13298 = n13296 & ~n13297 ;
  assign n13299 = n12936 | n12940 ;
  assign n13300 = n13298 & n13299 ;
  assign n13301 = n13298 | n13299 ;
  assign n13302 = ~n13300 & n13301 ;
  assign n13303 = x98 & n3314 ;
  assign n13304 = x97 & n3309 ;
  assign n13305 = x96 & ~n3308 ;
  assign n13306 = n3570 & n13305 ;
  assign n13307 = n13304 | n13306 ;
  assign n13308 = n13303 | n13307 ;
  assign n13309 = n3317 | n13308 ;
  assign n13310 = ( n4105 & n13308 ) | ( n4105 & n13309 ) | ( n13308 & n13309 ) ;
  assign n13311 = x32 & n13310 ;
  assign n13312 = x32 & ~n13311 ;
  assign n13313 = ( n13310 & ~n13311 ) | ( n13310 & n13312 ) | ( ~n13311 & n13312 ) ;
  assign n13314 = n13302 & n13313 ;
  assign n13315 = n13302 & ~n13314 ;
  assign n13316 = ~n13302 & n13313 ;
  assign n13317 = n13315 | n13316 ;
  assign n13318 = ( n12758 & n12759 ) | ( n12758 & n12941 ) | ( n12759 & n12941 ) ;
  assign n13319 = n13317 | n13318 ;
  assign n13320 = n13317 & n13318 ;
  assign n13321 = n13319 & ~n13320 ;
  assign n13322 = x101 & n2775 ;
  assign n13323 = x100 & n2770 ;
  assign n13324 = x99 & ~n2769 ;
  assign n13325 = n2978 & n13324 ;
  assign n13326 = n13323 | n13325 ;
  assign n13327 = n13322 | n13326 ;
  assign n13328 = n2778 | n13327 ;
  assign n13329 = ( n4783 & n13327 ) | ( n4783 & n13328 ) | ( n13327 & n13328 ) ;
  assign n13330 = x29 & n13329 ;
  assign n13331 = x29 & ~n13330 ;
  assign n13332 = ( n13329 & ~n13330 ) | ( n13329 & n13331 ) | ( ~n13330 & n13331 ) ;
  assign n13333 = n13321 & n13332 ;
  assign n13334 = n13321 & ~n13333 ;
  assign n13335 = ~n13321 & n13332 ;
  assign n13336 = n13334 | n13335 ;
  assign n13337 = n12945 | n12950 ;
  assign n13338 = n13336 | n13337 ;
  assign n13339 = n13336 & n13337 ;
  assign n13340 = n13338 & ~n13339 ;
  assign n13341 = x104 & n2280 ;
  assign n13342 = x103 & n2275 ;
  assign n13343 = x102 & ~n2274 ;
  assign n13344 = n2481 & n13343 ;
  assign n13345 = n13342 | n13344 ;
  assign n13346 = n13341 | n13345 ;
  assign n13347 = n2283 | n13346 ;
  assign n13348 = ( n5295 & n13346 ) | ( n5295 & n13347 ) | ( n13346 & n13347 ) ;
  assign n13349 = x26 & n13348 ;
  assign n13350 = x26 & ~n13349 ;
  assign n13351 = ( n13348 & ~n13349 ) | ( n13348 & n13350 ) | ( ~n13349 & n13350 ) ;
  assign n13352 = ~n13340 & n13351 ;
  assign n13353 = n13340 & ~n13351 ;
  assign n13354 = n13352 | n13353 ;
  assign n13355 = n12964 | n12967 ;
  assign n13356 = ( n13112 & n13354 ) | ( n13112 & ~n13355 ) | ( n13354 & ~n13355 ) ;
  assign n13357 = ( ~n13354 & n13355 ) | ( ~n13354 & n13356 ) | ( n13355 & n13356 ) ;
  assign n13358 = ( ~n13112 & n13356 ) | ( ~n13112 & n13357 ) | ( n13356 & n13357 ) ;
  assign n13359 = n13101 & n13358 ;
  assign n13360 = n13101 | n13358 ;
  assign n13361 = ~n13359 & n13360 ;
  assign n13362 = x110 & n1421 ;
  assign n13363 = x109 & n1416 ;
  assign n13364 = x108 & ~n1415 ;
  assign n13365 = n1584 & n13364 ;
  assign n13366 = n13363 | n13365 ;
  assign n13367 = n13362 | n13366 ;
  assign n13368 = n1424 | n13367 ;
  assign n13369 = ( n7189 & n13367 ) | ( n7189 & n13368 ) | ( n13367 & n13368 ) ;
  assign n13370 = x20 & n13369 ;
  assign n13371 = x20 & ~n13370 ;
  assign n13372 = ( n13369 & ~n13370 ) | ( n13369 & n13371 ) | ( ~n13370 & n13371 ) ;
  assign n13373 = n13361 & n13372 ;
  assign n13374 = n13361 & ~n13373 ;
  assign n13375 = ~n13361 & n13372 ;
  assign n13376 = n13374 | n13375 ;
  assign n13377 = n13100 & n13376 ;
  assign n13378 = n13100 | n13376 ;
  assign n13379 = ~n13377 & n13378 ;
  assign n13380 = x113 & n1071 ;
  assign n13381 = x112 & n1066 ;
  assign n13382 = x111 & ~n1065 ;
  assign n13383 = n1189 & n13382 ;
  assign n13384 = n13381 | n13383 ;
  assign n13385 = n13380 | n13384 ;
  assign n13386 = n1074 | n13385 ;
  assign n13387 = ( n8113 & n13385 ) | ( n8113 & n13386 ) | ( n13385 & n13386 ) ;
  assign n13388 = x17 & n13387 ;
  assign n13389 = x17 & ~n13388 ;
  assign n13390 = ( n13387 & ~n13388 ) | ( n13387 & n13389 ) | ( ~n13388 & n13389 ) ;
  assign n13391 = n13379 & n13390 ;
  assign n13392 = n13379 & ~n13391 ;
  assign n13393 = ~n13379 & n13390 ;
  assign n13394 = n13392 | n13393 ;
  assign n13395 = n13099 & n13394 ;
  assign n13396 = n13099 | n13394 ;
  assign n13397 = ~n13395 & n13396 ;
  assign n13398 = x116 & n771 ;
  assign n13399 = x115 & n766 ;
  assign n13400 = x114 & ~n765 ;
  assign n13401 = n905 & n13400 ;
  assign n13402 = n13399 | n13401 ;
  assign n13403 = n13398 | n13402 ;
  assign n13404 = n774 | n13403 ;
  assign n13405 = ( n8778 & n13403 ) | ( n8778 & n13404 ) | ( n13403 & n13404 ) ;
  assign n13406 = x14 & n13405 ;
  assign n13407 = x14 & ~n13406 ;
  assign n13408 = ( n13405 & ~n13406 ) | ( n13405 & n13407 ) | ( ~n13406 & n13407 ) ;
  assign n13409 = n13397 & n13408 ;
  assign n13410 = n13397 | n13408 ;
  assign n13411 = ~n13409 & n13410 ;
  assign n13412 = n13037 | n13041 ;
  assign n13413 = n13411 & n13412 ;
  assign n13414 = n13411 | n13412 ;
  assign n13415 = ~n13413 & n13414 ;
  assign n13416 = x119 & n528 ;
  assign n13417 = x118 & n523 ;
  assign n13418 = x117 & ~n522 ;
  assign n13419 = n635 & n13418 ;
  assign n13420 = n13417 | n13419 ;
  assign n13421 = n13416 | n13420 ;
  assign n13422 = n531 | n13421 ;
  assign n13423 = ( n9789 & n13421 ) | ( n9789 & n13422 ) | ( n13421 & n13422 ) ;
  assign n13424 = x11 & n13423 ;
  assign n13425 = x11 & ~n13424 ;
  assign n13426 = ( n13423 & ~n13424 ) | ( n13423 & n13425 ) | ( ~n13424 & n13425 ) ;
  assign n13427 = n13415 & n13426 ;
  assign n13428 = n13415 | n13426 ;
  assign n13429 = ~n13427 & n13428 ;
  assign n13430 = n13054 | n13060 ;
  assign n13431 = n13429 & n13430 ;
  assign n13432 = n13429 | n13430 ;
  assign n13433 = ~n13431 & n13432 ;
  assign n13434 = x122 & n337 ;
  assign n13435 = x121 & n332 ;
  assign n13436 = x120 & ~n331 ;
  assign n13437 = n396 & n13436 ;
  assign n13438 = n13435 | n13437 ;
  assign n13439 = n13434 | n13438 ;
  assign n13440 = n340 | n13439 ;
  assign n13441 = ( n11188 & n13439 ) | ( n11188 & n13440 ) | ( n13439 & n13440 ) ;
  assign n13442 = x8 & n13441 ;
  assign n13443 = x8 & ~n13442 ;
  assign n13444 = ( n13441 & ~n13442 ) | ( n13441 & n13443 ) | ( ~n13442 & n13443 ) ;
  assign n13445 = ( n13098 & n13433 ) | ( n13098 & ~n13444 ) | ( n13433 & ~n13444 ) ;
  assign n13446 = ( ~n13433 & n13444 ) | ( ~n13433 & n13445 ) | ( n13444 & n13445 ) ;
  assign n13447 = ( ~n13098 & n13445 ) | ( ~n13098 & n13446 ) | ( n13445 & n13446 ) ;
  assign n13448 = ( n12735 & n13061 ) | ( n12735 & n13072 ) | ( n13061 & n13072 ) ;
  assign n13449 = n13447 | n13448 ;
  assign n13450 = n13447 & n13448 ;
  assign n13451 = n13449 & ~n13450 ;
  assign n13452 = x127 & n131 ;
  assign n13453 = x126 & ~n156 ;
  assign n13454 = n135 & n13453 ;
  assign n13455 = n13452 | n13454 ;
  assign n13456 = n139 | n13455 ;
  assign n13457 = ~x126 & x127 ;
  assign n13458 = x126 & ~x127 ;
  assign n13459 = ( n12682 & n12685 ) | ( n12682 & n13458 ) | ( n12685 & n13458 ) ;
  assign n13460 = n12685 & ~n13459 ;
  assign n13461 = ( n13457 & n13459 ) | ( n13457 & ~n13460 ) | ( n13459 & ~n13460 ) ;
  assign n13462 = ( n13455 & n13456 ) | ( n13455 & n13461 ) | ( n13456 & n13461 ) ;
  assign n13463 = x2 & n13462 ;
  assign n13464 = x2 & ~n13463 ;
  assign n13465 = ( n13462 & ~n13463 ) | ( n13462 & n13464 ) | ( ~n13463 & n13464 ) ;
  assign n13466 = n13451 & n13465 ;
  assign n13467 = n13451 | n13465 ;
  assign n13468 = ~n13466 & n13467 ;
  assign n13469 = n13087 & n13468 ;
  assign n13470 = n13087 | n13468 ;
  assign n13471 = ~n13469 & n13470 ;
  assign n13472 = n13086 | n13471 ;
  assign n13473 = n13086 & n13471 ;
  assign n13474 = n13472 & ~n13473 ;
  assign n13475 = n13391 | n13395 ;
  assign n13476 = n13373 | n13377 ;
  assign n13477 = n13239 | n13245 ;
  assign n13478 = x87 & n6068 ;
  assign n13479 = x86 & n6063 ;
  assign n13480 = x85 & ~n6062 ;
  assign n13481 = n6398 & n13480 ;
  assign n13482 = n13479 | n13481 ;
  assign n13483 = n13478 | n13482 ;
  assign n13484 = n6071 | n13483 ;
  assign n13485 = ( n2067 & n13483 ) | ( n2067 & n13484 ) | ( n13483 & n13484 ) ;
  assign n13486 = x44 & n13485 ;
  assign n13487 = x44 & ~n13486 ;
  assign n13488 = ( n13485 & ~n13486 ) | ( n13485 & n13487 ) | ( ~n13486 & n13487 ) ;
  assign n13489 = x84 & n6937 ;
  assign n13490 = x83 & n6932 ;
  assign n13491 = x82 & ~n6931 ;
  assign n13492 = n7216 & n13491 ;
  assign n13493 = n13490 | n13492 ;
  assign n13494 = n13489 | n13493 ;
  assign n13495 = n6940 | n13494 ;
  assign n13496 = ( n1537 & n13494 ) | ( n1537 & n13495 ) | ( n13494 & n13495 ) ;
  assign n13497 = x47 & n13496 ;
  assign n13498 = x47 & ~n13497 ;
  assign n13499 = ( n13496 & ~n13497 ) | ( n13496 & n13498 ) | ( ~n13497 & n13498 ) ;
  assign n13500 = n13222 | n13225 ;
  assign n13501 = x81 & n7812 ;
  assign n13502 = x80 & n7807 ;
  assign n13503 = x79 & ~n7806 ;
  assign n13504 = n8136 & n13503 ;
  assign n13505 = n13502 | n13504 ;
  assign n13506 = n13501 | n13505 ;
  assign n13507 = n7815 | n13506 ;
  assign n13508 = ( n1256 & n13506 ) | ( n1256 & n13507 ) | ( n13506 & n13507 ) ;
  assign n13509 = x50 & n13508 ;
  assign n13510 = x50 & ~n13509 ;
  assign n13511 = ( n13508 & ~n13509 ) | ( n13508 & n13510 ) | ( ~n13509 & n13510 ) ;
  assign n13512 = x78 & n8834 ;
  assign n13513 = x77 & n8829 ;
  assign n13514 = x76 & ~n8828 ;
  assign n13515 = n9159 & n13514 ;
  assign n13516 = n13513 | n13515 ;
  assign n13517 = n13512 | n13516 ;
  assign n13518 = n8837 | n13517 ;
  assign n13519 = ( n868 & n13517 ) | ( n868 & n13518 ) | ( n13517 & n13518 ) ;
  assign n13520 = x53 & n13519 ;
  assign n13521 = x53 & ~n13520 ;
  assign n13522 = ( n13519 & ~n13520 ) | ( n13519 & n13521 ) | ( ~n13520 & n13521 ) ;
  assign n13523 = n13185 | n13188 ;
  assign n13524 = n13165 | n13171 ;
  assign n13525 = n13148 | n13151 ;
  assign n13526 = x72 & n10876 ;
  assign n13527 = x71 & n10871 ;
  assign n13528 = x70 & ~n10870 ;
  assign n13529 = n11305 & n13528 ;
  assign n13530 = n13527 | n13529 ;
  assign n13531 = n13526 | n13530 ;
  assign n13532 = ( n435 & n10879 ) | ( n435 & n13531 ) | ( n10879 & n13531 ) ;
  assign n13533 = ( x59 & ~n13531 ) | ( x59 & n13532 ) | ( ~n13531 & n13532 ) ;
  assign n13534 = ~n13532 & n13533 ;
  assign n13535 = n13531 | n13533 ;
  assign n13536 = ( ~x59 & n13534 ) | ( ~x59 & n13535 ) | ( n13534 & n13535 ) ;
  assign n13537 = n13128 | n13134 ;
  assign n13538 = n264 & n11987 ;
  assign n13539 = x69 & n11984 ;
  assign n13540 = x68 & n11979 ;
  assign n13541 = x67 & ~n11978 ;
  assign n13542 = n12430 & n13541 ;
  assign n13543 = n13540 | n13542 ;
  assign n13544 = n13539 | n13543 ;
  assign n13545 = n13538 | n13544 ;
  assign n13546 = x62 | n13545 ;
  assign n13547 = ~x62 & n13546 ;
  assign n13548 = ( ~n13545 & n13546 ) | ( ~n13545 & n13547 ) | ( n13546 & n13547 ) ;
  assign n13549 = x66 & n12808 ;
  assign n13550 = x63 & x65 ;
  assign n13551 = ~n12808 & n13550 ;
  assign n13552 = n13549 | n13551 ;
  assign n13553 = ( n13537 & n13548 ) | ( n13537 & ~n13552 ) | ( n13548 & ~n13552 ) ;
  assign n13554 = ( ~n13548 & n13552 ) | ( ~n13548 & n13553 ) | ( n13552 & n13553 ) ;
  assign n13555 = ( ~n13537 & n13553 ) | ( ~n13537 & n13554 ) | ( n13553 & n13554 ) ;
  assign n13556 = n13536 | n13555 ;
  assign n13557 = n13525 & n13556 ;
  assign n13558 = n13536 & n13555 ;
  assign n13559 = n13556 & ~n13558 ;
  assign n13560 = ~n13557 & n13559 ;
  assign n13561 = x75 & n9853 ;
  assign n13562 = x74 & n9848 ;
  assign n13563 = x73 & ~n9847 ;
  assign n13564 = n10165 & n13563 ;
  assign n13565 = n13562 | n13564 ;
  assign n13566 = n13561 | n13565 ;
  assign n13567 = n9856 | n13566 ;
  assign n13568 = ( n609 & n13566 ) | ( n609 & n13567 ) | ( n13566 & n13567 ) ;
  assign n13569 = x56 & n13568 ;
  assign n13570 = x56 & ~n13569 ;
  assign n13571 = ( n13568 & ~n13569 ) | ( n13568 & n13570 ) | ( ~n13569 & n13570 ) ;
  assign n13572 = n13560 | n13571 ;
  assign n13573 = n13525 & ~n13559 ;
  assign n13574 = n13572 | n13573 ;
  assign n13575 = ( n13560 & n13571 ) | ( n13560 & n13573 ) | ( n13571 & n13573 ) ;
  assign n13576 = n13574 & ~n13575 ;
  assign n13577 = n13524 & n13576 ;
  assign n13578 = n13524 | n13576 ;
  assign n13579 = ~n13577 & n13578 ;
  assign n13580 = ( n13522 & n13523 ) | ( n13522 & ~n13579 ) | ( n13523 & ~n13579 ) ;
  assign n13581 = ( ~n13523 & n13579 ) | ( ~n13523 & n13580 ) | ( n13579 & n13580 ) ;
  assign n13582 = ( ~n13522 & n13580 ) | ( ~n13522 & n13581 ) | ( n13580 & n13581 ) ;
  assign n13583 = n13511 & n13582 ;
  assign n13584 = n13511 | n13582 ;
  assign n13585 = ~n13583 & n13584 ;
  assign n13586 = n13202 | n13208 ;
  assign n13587 = n13585 | n13586 ;
  assign n13588 = n13585 & n13586 ;
  assign n13589 = n13587 & ~n13588 ;
  assign n13590 = ( n13499 & n13500 ) | ( n13499 & ~n13589 ) | ( n13500 & ~n13589 ) ;
  assign n13591 = ( ~n13500 & n13589 ) | ( ~n13500 & n13590 ) | ( n13589 & n13590 ) ;
  assign n13592 = ( ~n13499 & n13590 ) | ( ~n13499 & n13591 ) | ( n13590 & n13591 ) ;
  assign n13593 = n13488 & n13592 ;
  assign n13594 = n13488 | n13592 ;
  assign n13595 = ~n13593 & n13594 ;
  assign n13596 = n13477 | n13595 ;
  assign n13597 = n13477 & n13595 ;
  assign n13598 = n13596 & ~n13597 ;
  assign n13599 = x90 & n5340 ;
  assign n13600 = x89 & n5335 ;
  assign n13601 = x88 & ~n5334 ;
  assign n13602 = n5580 & n13601 ;
  assign n13603 = n13600 | n13602 ;
  assign n13604 = n13599 | n13603 ;
  assign n13605 = n5343 | n13604 ;
  assign n13606 = ( n2410 & n13604 ) | ( n2410 & n13605 ) | ( n13604 & n13605 ) ;
  assign n13607 = x41 & n13606 ;
  assign n13608 = x41 & ~n13607 ;
  assign n13609 = ( n13606 & ~n13607 ) | ( n13606 & n13608 ) | ( ~n13607 & n13608 ) ;
  assign n13610 = n13598 & n13609 ;
  assign n13611 = n13598 & ~n13610 ;
  assign n13612 = ~n13598 & n13609 ;
  assign n13613 = n13611 | n13612 ;
  assign n13614 = n13258 | n13264 ;
  assign n13615 = n13613 | n13614 ;
  assign n13616 = n13613 & n13614 ;
  assign n13617 = n13615 & ~n13616 ;
  assign n13618 = x93 & n4572 ;
  assign n13619 = x92 & n4567 ;
  assign n13620 = x91 & ~n4566 ;
  assign n13621 = n4828 & n13620 ;
  assign n13622 = n13619 | n13621 ;
  assign n13623 = n13618 | n13622 ;
  assign n13624 = n4575 | n13623 ;
  assign n13625 = ( n2931 & n13623 ) | ( n2931 & n13624 ) | ( n13623 & n13624 ) ;
  assign n13626 = x38 & n13625 ;
  assign n13627 = x38 & ~n13626 ;
  assign n13628 = ( n13625 & ~n13626 ) | ( n13625 & n13627 ) | ( ~n13626 & n13627 ) ;
  assign n13629 = n13617 & n13628 ;
  assign n13630 = n13617 & ~n13629 ;
  assign n13631 = ~n13617 & n13628 ;
  assign n13632 = n13630 | n13631 ;
  assign n13633 = n13277 | n13283 ;
  assign n13634 = n13632 | n13633 ;
  assign n13635 = n13632 & n13633 ;
  assign n13636 = n13634 & ~n13635 ;
  assign n13637 = x96 & n3913 ;
  assign n13638 = x95 & n3908 ;
  assign n13639 = x94 & ~n3907 ;
  assign n13640 = n4152 & n13639 ;
  assign n13641 = n13638 | n13640 ;
  assign n13642 = n13637 | n13641 ;
  assign n13643 = n3916 | n13642 ;
  assign n13644 = ( n3509 & n13642 ) | ( n3509 & n13643 ) | ( n13642 & n13643 ) ;
  assign n13645 = x35 & n13644 ;
  assign n13646 = x35 & ~n13645 ;
  assign n13647 = ( n13644 & ~n13645 ) | ( n13644 & n13646 ) | ( ~n13645 & n13646 ) ;
  assign n13648 = n13636 & n13647 ;
  assign n13649 = n13636 | n13647 ;
  assign n13650 = ~n13648 & n13649 ;
  assign n13651 = n13297 | n13300 ;
  assign n13652 = n13650 & n13651 ;
  assign n13653 = n13651 & ~n13652 ;
  assign n13654 = ( n13650 & ~n13652 ) | ( n13650 & n13653 ) | ( ~n13652 & n13653 ) ;
  assign n13655 = x99 & n3314 ;
  assign n13656 = x98 & n3309 ;
  assign n13657 = x97 & ~n3308 ;
  assign n13658 = n3570 & n13657 ;
  assign n13659 = n13656 | n13658 ;
  assign n13660 = n13655 | n13659 ;
  assign n13661 = n3317 | n13660 ;
  assign n13662 = ( n4325 & n13660 ) | ( n4325 & n13661 ) | ( n13660 & n13661 ) ;
  assign n13663 = x32 & n13662 ;
  assign n13664 = x32 & ~n13663 ;
  assign n13665 = ( n13662 & ~n13663 ) | ( n13662 & n13664 ) | ( ~n13663 & n13664 ) ;
  assign n13666 = n13654 & n13665 ;
  assign n13667 = n13654 & ~n13666 ;
  assign n13668 = ~n13654 & n13665 ;
  assign n13669 = n13667 | n13668 ;
  assign n13670 = n13314 | n13320 ;
  assign n13671 = n13669 | n13670 ;
  assign n13672 = n13669 & n13670 ;
  assign n13673 = n13671 & ~n13672 ;
  assign n13674 = x102 & n2775 ;
  assign n13675 = x101 & n2770 ;
  assign n13676 = x100 & ~n2769 ;
  assign n13677 = n2978 & n13676 ;
  assign n13678 = n13675 | n13677 ;
  assign n13679 = n13674 | n13678 ;
  assign n13680 = n2778 | n13679 ;
  assign n13681 = ( n5025 & n13679 ) | ( n5025 & n13680 ) | ( n13679 & n13680 ) ;
  assign n13682 = x29 & n13681 ;
  assign n13683 = x29 & ~n13682 ;
  assign n13684 = ( n13681 & ~n13682 ) | ( n13681 & n13683 ) | ( ~n13682 & n13683 ) ;
  assign n13685 = n13673 & n13684 ;
  assign n13686 = n13673 & ~n13685 ;
  assign n13687 = ~n13673 & n13684 ;
  assign n13688 = n13686 | n13687 ;
  assign n13689 = n13333 | n13339 ;
  assign n13690 = n13688 | n13689 ;
  assign n13691 = n13688 & n13689 ;
  assign n13692 = n13690 & ~n13691 ;
  assign n13693 = x105 & n2280 ;
  assign n13694 = x104 & n2275 ;
  assign n13695 = x103 & ~n2274 ;
  assign n13696 = n2481 & n13695 ;
  assign n13697 = n13694 | n13696 ;
  assign n13698 = n13693 | n13697 ;
  assign n13699 = n2283 | n13698 ;
  assign n13700 = ( n5788 & n13698 ) | ( n5788 & n13699 ) | ( n13698 & n13699 ) ;
  assign n13701 = x26 & n13700 ;
  assign n13702 = x26 & ~n13701 ;
  assign n13703 = ( n13700 & ~n13701 ) | ( n13700 & n13702 ) | ( ~n13701 & n13702 ) ;
  assign n13704 = n13692 & n13703 ;
  assign n13705 = n13692 | n13703 ;
  assign n13706 = ~n13704 & n13705 ;
  assign n13707 = ( n13340 & n13351 ) | ( n13340 & n13355 ) | ( n13351 & n13355 ) ;
  assign n13708 = n13706 & n13707 ;
  assign n13709 = n13707 & ~n13708 ;
  assign n13710 = ( n13706 & ~n13708 ) | ( n13706 & n13709 ) | ( ~n13708 & n13709 ) ;
  assign n13711 = x108 & n1817 ;
  assign n13712 = x107 & n1812 ;
  assign n13713 = x106 & ~n1811 ;
  assign n13714 = n1977 & n13713 ;
  assign n13715 = n13712 | n13714 ;
  assign n13716 = n13711 | n13715 ;
  assign n13717 = n1820 | n13716 ;
  assign n13718 = ( n6358 & n13716 ) | ( n6358 & n13717 ) | ( n13716 & n13717 ) ;
  assign n13719 = x23 & n13718 ;
  assign n13720 = x23 & ~n13719 ;
  assign n13721 = ( n13718 & ~n13719 ) | ( n13718 & n13720 ) | ( ~n13719 & n13720 ) ;
  assign n13722 = n13710 & n13721 ;
  assign n13723 = n13710 & ~n13722 ;
  assign n13724 = ~n13710 & n13721 ;
  assign n13725 = n13723 | n13724 ;
  assign n13726 = n13354 & ~n13355 ;
  assign n13727 = ~n13354 & n13355 ;
  assign n13728 = n13726 | n13727 ;
  assign n13729 = ( n13101 & n13112 ) | ( n13101 & n13728 ) | ( n13112 & n13728 ) ;
  assign n13730 = n13725 & n13729 ;
  assign n13731 = n13725 | n13729 ;
  assign n13732 = ~n13730 & n13731 ;
  assign n13733 = x111 & n1421 ;
  assign n13734 = x110 & n1416 ;
  assign n13735 = x109 & ~n1415 ;
  assign n13736 = n1584 & n13735 ;
  assign n13737 = n13734 | n13736 ;
  assign n13738 = n13733 | n13737 ;
  assign n13739 = n1424 | n13738 ;
  assign n13740 = ( n7492 & n13738 ) | ( n7492 & n13739 ) | ( n13738 & n13739 ) ;
  assign n13741 = x20 & n13740 ;
  assign n13742 = x20 & ~n13741 ;
  assign n13743 = ( n13740 & ~n13741 ) | ( n13740 & n13742 ) | ( ~n13741 & n13742 ) ;
  assign n13744 = n13732 & n13743 ;
  assign n13745 = n13732 & ~n13744 ;
  assign n13746 = ~n13732 & n13743 ;
  assign n13747 = n13745 | n13746 ;
  assign n13748 = n13476 & n13747 ;
  assign n13749 = n13476 & ~n13748 ;
  assign n13750 = n13747 & ~n13748 ;
  assign n13751 = n13749 | n13750 ;
  assign n13752 = x114 & n1071 ;
  assign n13753 = x113 & n1066 ;
  assign n13754 = x112 & ~n1065 ;
  assign n13755 = n1189 & n13754 ;
  assign n13756 = n13753 | n13755 ;
  assign n13757 = n13752 | n13756 ;
  assign n13758 = n1074 | n13757 ;
  assign n13759 = ( n8437 & n13757 ) | ( n8437 & n13758 ) | ( n13757 & n13758 ) ;
  assign n13760 = x17 & n13759 ;
  assign n13761 = x17 & ~n13760 ;
  assign n13762 = ( n13759 & ~n13760 ) | ( n13759 & n13761 ) | ( ~n13760 & n13761 ) ;
  assign n13763 = n13751 | n13762 ;
  assign n13764 = n13751 & n13762 ;
  assign n13765 = n13763 & ~n13764 ;
  assign n13766 = n13475 & n13765 ;
  assign n13767 = n13475 | n13765 ;
  assign n13768 = ~n13766 & n13767 ;
  assign n13769 = x117 & n771 ;
  assign n13770 = x116 & n766 ;
  assign n13771 = x115 & ~n765 ;
  assign n13772 = n905 & n13771 ;
  assign n13773 = n13770 | n13772 ;
  assign n13774 = n13769 | n13773 ;
  assign n13775 = n774 | n13774 ;
  assign n13776 = ( n9118 & n13774 ) | ( n9118 & n13775 ) | ( n13774 & n13775 ) ;
  assign n13777 = x14 & n13776 ;
  assign n13778 = x14 & ~n13777 ;
  assign n13779 = ( n13776 & ~n13777 ) | ( n13776 & n13778 ) | ( ~n13777 & n13778 ) ;
  assign n13780 = n13768 & n13779 ;
  assign n13781 = n13768 & ~n13780 ;
  assign n13782 = ~n13768 & n13779 ;
  assign n13783 = n13781 | n13782 ;
  assign n13784 = n13409 | n13413 ;
  assign n13785 = n13783 | n13784 ;
  assign n13786 = n13783 & n13784 ;
  assign n13787 = n13785 & ~n13786 ;
  assign n13788 = x120 & n528 ;
  assign n13789 = x119 & n523 ;
  assign n13790 = x118 & ~n522 ;
  assign n13791 = n635 & n13790 ;
  assign n13792 = n13789 | n13791 ;
  assign n13793 = n13788 | n13792 ;
  assign n13794 = n531 | n13793 ;
  assign n13795 = ( n10460 & n13793 ) | ( n10460 & n13794 ) | ( n13793 & n13794 ) ;
  assign n13796 = x11 & n13795 ;
  assign n13797 = x11 & ~n13796 ;
  assign n13798 = ( n13795 & ~n13796 ) | ( n13795 & n13797 ) | ( ~n13796 & n13797 ) ;
  assign n13799 = n13787 | n13798 ;
  assign n13800 = x123 & n337 ;
  assign n13801 = x122 & n332 ;
  assign n13802 = x121 & ~n331 ;
  assign n13803 = n396 & n13802 ;
  assign n13804 = n13801 | n13803 ;
  assign n13805 = n13800 | n13804 ;
  assign n13806 = n340 | n13805 ;
  assign n13807 = ( n11219 & n13805 ) | ( n11219 & n13806 ) | ( n13805 & n13806 ) ;
  assign n13808 = x8 & n13807 ;
  assign n13809 = x8 & ~n13808 ;
  assign n13810 = ( n13807 & ~n13808 ) | ( n13807 & n13809 ) | ( ~n13808 & n13809 ) ;
  assign n13811 = ( n13787 & n13798 ) | ( n13787 & n13810 ) | ( n13798 & n13810 ) ;
  assign n13812 = n13799 & ~n13811 ;
  assign n13813 = n13427 | n13431 ;
  assign n13814 = ( n13798 & ~n13799 ) | ( n13798 & n13810 ) | ( ~n13799 & n13810 ) ;
  assign n13815 = ( n13787 & ~n13799 ) | ( n13787 & n13814 ) | ( ~n13799 & n13814 ) ;
  assign n13816 = n13813 | n13815 ;
  assign n13817 = n13812 | n13816 ;
  assign n13818 = ( n13812 & n13813 ) | ( n13812 & n13815 ) | ( n13813 & n13815 ) ;
  assign n13819 = n13817 & ~n13818 ;
  assign n13820 = x126 & n206 ;
  assign n13821 = x125 & n201 ;
  assign n13822 = x124 & ~n200 ;
  assign n13823 = n243 & n13822 ;
  assign n13824 = n13821 | n13823 ;
  assign n13825 = n13820 | n13824 ;
  assign n13826 = n209 | n13825 ;
  assign n13827 = ( n12687 & n13825 ) | ( n12687 & n13826 ) | ( n13825 & n13826 ) ;
  assign n13828 = x5 & n13827 ;
  assign n13829 = x5 & ~n13828 ;
  assign n13830 = ( n13827 & ~n13828 ) | ( n13827 & n13829 ) | ( ~n13828 & n13829 ) ;
  assign n13831 = n13819 & n13830 ;
  assign n13832 = n13819 & ~n13831 ;
  assign n13833 = ~n13819 & n13830 ;
  assign n13834 = n13832 | n13833 ;
  assign n13835 = x127 & n139 ;
  assign n13836 = x126 & n13835 ;
  assign n13837 = ( n12685 & n13835 ) | ( n12685 & n13836 ) | ( n13835 & n13836 ) ;
  assign n13838 = x2 | n13837 ;
  assign n13839 = x127 & ~n156 ;
  assign n13840 = n135 & n13839 ;
  assign n13841 = n13837 | n13840 ;
  assign n13842 = x2 & n13841 ;
  assign n13843 = n13838 & ~n13842 ;
  assign n13844 = n13433 & n13444 ;
  assign n13845 = n13843 | n13844 ;
  assign n13846 = n13433 & ~n13844 ;
  assign n13847 = ( n13098 & ~n13445 ) | ( n13098 & n13846 ) | ( ~n13445 & n13846 ) ;
  assign n13848 = n13845 | n13847 ;
  assign n13849 = ( n13843 & n13844 ) | ( n13843 & n13847 ) | ( n13844 & n13847 ) ;
  assign n13850 = n13848 & ~n13849 ;
  assign n13851 = n13834 & n13850 ;
  assign n13852 = n13834 | n13850 ;
  assign n13853 = ~n13851 & n13852 ;
  assign n13854 = n13450 | n13466 ;
  assign n13855 = n13853 | n13854 ;
  assign n13856 = n13853 & n13854 ;
  assign n13857 = n13855 & ~n13856 ;
  assign n13858 = n13469 | n13473 ;
  assign n13859 = n13857 | n13858 ;
  assign n13860 = n13857 & n13858 ;
  assign n13861 = n13859 & ~n13860 ;
  assign n13862 = n13849 | n13851 ;
  assign n13863 = n13818 | n13831 ;
  assign n13864 = x127 & n206 ;
  assign n13865 = x126 & n201 ;
  assign n13866 = x125 & ~n200 ;
  assign n13867 = n243 & n13866 ;
  assign n13868 = n13865 | n13867 ;
  assign n13869 = n13864 | n13868 ;
  assign n13870 = n209 | n13869 ;
  assign n13871 = ( n12720 & n13869 ) | ( n12720 & n13870 ) | ( n13869 & n13870 ) ;
  assign n13872 = x5 & n13871 ;
  assign n13873 = x5 & ~n13872 ;
  assign n13874 = ( n13871 & ~n13872 ) | ( n13871 & n13873 ) | ( ~n13872 & n13873 ) ;
  assign n13875 = n13863 & n13874 ;
  assign n13876 = n13863 & ~n13875 ;
  assign n13877 = ~n13863 & n13874 ;
  assign n13878 = n13876 | n13877 ;
  assign n13879 = x118 & n771 ;
  assign n13880 = x117 & n766 ;
  assign n13881 = x116 & ~n765 ;
  assign n13882 = n905 & n13881 ;
  assign n13883 = n13880 | n13882 ;
  assign n13884 = n13879 | n13883 ;
  assign n13885 = n774 | n13884 ;
  assign n13886 = ( n9760 & n13884 ) | ( n9760 & n13885 ) | ( n13884 & n13885 ) ;
  assign n13887 = x14 & n13886 ;
  assign n13888 = x14 & ~n13887 ;
  assign n13889 = ( n13886 & ~n13887 ) | ( n13886 & n13888 ) | ( ~n13887 & n13888 ) ;
  assign n13890 = n13764 & n13889 ;
  assign n13891 = n13889 & ~n13890 ;
  assign n13892 = ~n13766 & n13891 ;
  assign n13893 = ( n13766 & n13889 ) | ( n13766 & n13890 ) | ( n13889 & n13890 ) ;
  assign n13894 = ( n13764 & n13766 ) | ( n13764 & ~n13893 ) | ( n13766 & ~n13893 ) ;
  assign n13895 = n13892 | n13894 ;
  assign n13896 = x103 & n2775 ;
  assign n13897 = x102 & n2770 ;
  assign n13898 = x101 & ~n2769 ;
  assign n13899 = n2978 & n13898 ;
  assign n13900 = n13897 | n13899 ;
  assign n13901 = n13896 | n13900 ;
  assign n13902 = n2778 | n13901 ;
  assign n13903 = ( n5264 & n13901 ) | ( n5264 & n13902 ) | ( n13901 & n13902 ) ;
  assign n13904 = x29 & n13903 ;
  assign n13905 = x29 & ~n13904 ;
  assign n13906 = ( n13903 & ~n13904 ) | ( n13903 & n13905 ) | ( ~n13904 & n13905 ) ;
  assign n13907 = n13666 | n13906 ;
  assign n13908 = n13672 | n13907 ;
  assign n13909 = ( n13666 & n13672 ) | ( n13666 & n13906 ) | ( n13672 & n13906 ) ;
  assign n13910 = n13908 & ~n13909 ;
  assign n13911 = x100 & n3314 ;
  assign n13912 = x99 & n3309 ;
  assign n13913 = x98 & ~n3308 ;
  assign n13914 = n3570 & n13913 ;
  assign n13915 = n13912 | n13914 ;
  assign n13916 = n13911 | n13915 ;
  assign n13917 = n3317 | n13916 ;
  assign n13918 = ( n4532 & n13916 ) | ( n4532 & n13917 ) | ( n13916 & n13917 ) ;
  assign n13919 = x32 & n13918 ;
  assign n13920 = x32 & ~n13919 ;
  assign n13921 = ( n13918 & ~n13919 ) | ( n13918 & n13920 ) | ( ~n13919 & n13920 ) ;
  assign n13922 = n13648 & n13921 ;
  assign n13923 = n13921 & ~n13922 ;
  assign n13924 = ~n13652 & n13923 ;
  assign n13925 = ( n13648 & n13652 ) | ( n13648 & ~n13921 ) | ( n13652 & ~n13921 ) ;
  assign n13926 = n13924 | n13925 ;
  assign n13927 = n13629 | n13635 ;
  assign n13928 = n13610 | n13616 ;
  assign n13929 = x91 & n5340 ;
  assign n13930 = x90 & n5335 ;
  assign n13931 = x89 & ~n5334 ;
  assign n13932 = n5580 & n13931 ;
  assign n13933 = n13930 | n13932 ;
  assign n13934 = n13929 | n13933 ;
  assign n13935 = n5343 | n13934 ;
  assign n13936 = ( n2714 & n13934 ) | ( n2714 & n13935 ) | ( n13934 & n13935 ) ;
  assign n13937 = x41 & n13936 ;
  assign n13938 = x41 & ~n13937 ;
  assign n13939 = ( n13936 & ~n13937 ) | ( n13936 & n13938 ) | ( ~n13937 & n13938 ) ;
  assign n13940 = n13593 | n13597 ;
  assign n13941 = ( n13499 & n13500 ) | ( n13499 & n13589 ) | ( n13500 & n13589 ) ;
  assign n13942 = n13583 | n13588 ;
  assign n13943 = x82 & n7812 ;
  assign n13944 = x81 & n7807 ;
  assign n13945 = x80 & ~n7806 ;
  assign n13946 = n8136 & n13945 ;
  assign n13947 = n13944 | n13946 ;
  assign n13948 = n13943 | n13947 ;
  assign n13949 = n7815 | n13948 ;
  assign n13950 = ( n1371 & n13948 ) | ( n1371 & n13949 ) | ( n13948 & n13949 ) ;
  assign n13951 = x50 & n13950 ;
  assign n13952 = x50 & ~n13951 ;
  assign n13953 = ( n13950 & ~n13951 ) | ( n13950 & n13952 ) | ( ~n13951 & n13952 ) ;
  assign n13954 = ( n13522 & n13523 ) | ( n13522 & n13579 ) | ( n13523 & n13579 ) ;
  assign n13955 = x79 & n8834 ;
  assign n13956 = x78 & n8829 ;
  assign n13957 = x77 & ~n8828 ;
  assign n13958 = n9159 & n13957 ;
  assign n13959 = n13956 | n13958 ;
  assign n13960 = n13955 | n13959 ;
  assign n13961 = n8837 | n13960 ;
  assign n13962 = ( n961 & n13960 ) | ( n961 & n13961 ) | ( n13960 & n13961 ) ;
  assign n13963 = x53 & n13962 ;
  assign n13964 = x53 & ~n13963 ;
  assign n13965 = ( n13962 & ~n13963 ) | ( n13962 & n13964 ) | ( ~n13963 & n13964 ) ;
  assign n13966 = n13575 | n13577 ;
  assign n13967 = x76 & n9853 ;
  assign n13968 = x75 & n9848 ;
  assign n13969 = x74 & ~n9847 ;
  assign n13970 = n10165 & n13969 ;
  assign n13971 = n13968 | n13970 ;
  assign n13972 = n13967 | n13971 ;
  assign n13973 = n9856 | n13972 ;
  assign n13974 = ( n740 & n13972 ) | ( n740 & n13973 ) | ( n13972 & n13973 ) ;
  assign n13975 = x56 & n13974 ;
  assign n13976 = x56 & ~n13975 ;
  assign n13977 = ( n13974 & ~n13975 ) | ( n13974 & n13976 ) | ( ~n13975 & n13976 ) ;
  assign n13978 = n13557 | n13558 ;
  assign n14011 = ( n13537 & n13548 ) | ( n13537 & ~n13555 ) | ( n13548 & ~n13555 ) ;
  assign n13979 = x67 & n12808 ;
  assign n13980 = x63 & x66 ;
  assign n13981 = ~n12808 & n13980 ;
  assign n13982 = n13979 | n13981 ;
  assign n13983 = x2 & n13982 ;
  assign n13984 = x2 | n13982 ;
  assign n13985 = ~n13983 & n13984 ;
  assign n13986 = x69 & n11979 ;
  assign n13987 = x68 & ~n11978 ;
  assign n13988 = n12430 & n13987 ;
  assign n13989 = n13986 | n13988 ;
  assign n13990 = x70 & n11984 ;
  assign n13991 = n13989 | n13990 ;
  assign n13992 = ( n310 & n11987 ) | ( n310 & n13991 ) | ( n11987 & n13991 ) ;
  assign n13993 = n13991 | n13992 ;
  assign n13994 = x62 & ~n13993 ;
  assign n13995 = ~x62 & n13993 ;
  assign n13996 = n13994 | n13995 ;
  assign n13997 = n13985 & n13996 ;
  assign n13998 = n13985 | n13996 ;
  assign n13999 = ~n13997 & n13998 ;
  assign n14000 = x73 & n10876 ;
  assign n14001 = x72 & n10871 ;
  assign n14002 = x71 & ~n10870 ;
  assign n14003 = n11305 & n14002 ;
  assign n14004 = n14001 | n14003 ;
  assign n14005 = n14000 | n14004 ;
  assign n14006 = ( n499 & n10879 ) | ( n499 & n14005 ) | ( n10879 & n14005 ) ;
  assign n14007 = ( x59 & ~n14005 ) | ( x59 & n14006 ) | ( ~n14005 & n14006 ) ;
  assign n14008 = ~n14006 & n14007 ;
  assign n14009 = n14005 | n14007 ;
  assign n14010 = ( ~x59 & n14008 ) | ( ~x59 & n14009 ) | ( n14008 & n14009 ) ;
  assign n14012 = ( n13999 & n14010 ) | ( n13999 & n14011 ) | ( n14010 & n14011 ) ;
  assign n14013 = ( n13999 & n14010 ) | ( n13999 & ~n14012 ) | ( n14010 & ~n14012 ) ;
  assign n14014 = ( n14011 & ~n14012 ) | ( n14011 & n14013 ) | ( ~n14012 & n14013 ) ;
  assign n14015 = ( n13977 & n13978 ) | ( n13977 & ~n14014 ) | ( n13978 & ~n14014 ) ;
  assign n14016 = ( ~n13978 & n14014 ) | ( ~n13978 & n14015 ) | ( n14014 & n14015 ) ;
  assign n14017 = ( ~n13977 & n14015 ) | ( ~n13977 & n14016 ) | ( n14015 & n14016 ) ;
  assign n14018 = ( n13965 & ~n13966 ) | ( n13965 & n14017 ) | ( ~n13966 & n14017 ) ;
  assign n14019 = ( n13966 & ~n14017 ) | ( n13966 & n14018 ) | ( ~n14017 & n14018 ) ;
  assign n14020 = ( ~n13965 & n14018 ) | ( ~n13965 & n14019 ) | ( n14018 & n14019 ) ;
  assign n14021 = ( n13953 & ~n13954 ) | ( n13953 & n14020 ) | ( ~n13954 & n14020 ) ;
  assign n14022 = ( n13954 & ~n14020 ) | ( n13954 & n14021 ) | ( ~n14020 & n14021 ) ;
  assign n14023 = ( ~n13953 & n14021 ) | ( ~n13953 & n14022 ) | ( n14021 & n14022 ) ;
  assign n14024 = n13942 | n14023 ;
  assign n14025 = n13942 & n14023 ;
  assign n14026 = n14024 & ~n14025 ;
  assign n14027 = x85 & n6937 ;
  assign n14028 = x84 & n6932 ;
  assign n14029 = x83 & ~n6931 ;
  assign n14030 = n7216 & n14029 ;
  assign n14031 = n14028 | n14030 ;
  assign n14032 = n14027 | n14031 ;
  assign n14033 = n6940 | n14032 ;
  assign n14034 = ( n1765 & n14032 ) | ( n1765 & n14033 ) | ( n14032 & n14033 ) ;
  assign n14035 = x47 & n14034 ;
  assign n14036 = x47 & ~n14035 ;
  assign n14037 = ( n14034 & ~n14035 ) | ( n14034 & n14036 ) | ( ~n14035 & n14036 ) ;
  assign n14038 = n14026 | n14037 ;
  assign n14039 = n14026 & n14037 ;
  assign n14040 = n14038 & ~n14039 ;
  assign n14041 = x88 & n6068 ;
  assign n14042 = x87 & n6063 ;
  assign n14043 = x86 & ~n6062 ;
  assign n14044 = n6398 & n14043 ;
  assign n14045 = n14042 | n14044 ;
  assign n14046 = n14041 | n14045 ;
  assign n14047 = n6071 | n14046 ;
  assign n14048 = ( n2095 & n14046 ) | ( n2095 & n14047 ) | ( n14046 & n14047 ) ;
  assign n14049 = x44 & n14048 ;
  assign n14050 = x44 & ~n14049 ;
  assign n14051 = ( n14048 & ~n14049 ) | ( n14048 & n14050 ) | ( ~n14049 & n14050 ) ;
  assign n14052 = ( n13941 & n14040 ) | ( n13941 & n14051 ) | ( n14040 & n14051 ) ;
  assign n14053 = ( n14040 & n14051 ) | ( n14040 & ~n14052 ) | ( n14051 & ~n14052 ) ;
  assign n14054 = ( n13941 & ~n14052 ) | ( n13941 & n14053 ) | ( ~n14052 & n14053 ) ;
  assign n14055 = ( n13939 & ~n13940 ) | ( n13939 & n14054 ) | ( ~n13940 & n14054 ) ;
  assign n14056 = ( n13940 & ~n14054 ) | ( n13940 & n14055 ) | ( ~n14054 & n14055 ) ;
  assign n14057 = ( ~n13939 & n14055 ) | ( ~n13939 & n14056 ) | ( n14055 & n14056 ) ;
  assign n14058 = n13928 | n14057 ;
  assign n14059 = n13928 & n14057 ;
  assign n14060 = n14058 & ~n14059 ;
  assign n14061 = x94 & n4572 ;
  assign n14062 = x93 & n4567 ;
  assign n14063 = x92 & ~n4566 ;
  assign n14064 = n4828 & n14063 ;
  assign n14065 = n14062 | n14064 ;
  assign n14066 = n14061 | n14065 ;
  assign n14067 = n4575 | n14066 ;
  assign n14068 = ( n3271 & n14066 ) | ( n3271 & n14067 ) | ( n14066 & n14067 ) ;
  assign n14069 = x38 & n14068 ;
  assign n14070 = x38 & ~n14069 ;
  assign n14071 = ( n14068 & ~n14069 ) | ( n14068 & n14070 ) | ( ~n14069 & n14070 ) ;
  assign n14072 = n14060 | n14071 ;
  assign n14073 = n14060 & n14071 ;
  assign n14074 = n14072 & ~n14073 ;
  assign n14075 = x97 & n3913 ;
  assign n14076 = x96 & n3908 ;
  assign n14077 = x95 & ~n3907 ;
  assign n14078 = n4152 & n14077 ;
  assign n14079 = n14076 | n14078 ;
  assign n14080 = n14075 | n14079 ;
  assign n14081 = n3916 | n14080 ;
  assign n14082 = ( n3707 & n14080 ) | ( n3707 & n14081 ) | ( n14080 & n14081 ) ;
  assign n14083 = x35 & n14082 ;
  assign n14084 = x35 & ~n14083 ;
  assign n14085 = ( n14082 & ~n14083 ) | ( n14082 & n14084 ) | ( ~n14083 & n14084 ) ;
  assign n14086 = ( n13927 & n14074 ) | ( n13927 & n14085 ) | ( n14074 & n14085 ) ;
  assign n14087 = ( n14074 & n14085 ) | ( n14074 & ~n14086 ) | ( n14085 & ~n14086 ) ;
  assign n14088 = ( n13927 & ~n14086 ) | ( n13927 & n14087 ) | ( ~n14086 & n14087 ) ;
  assign n14089 = n13926 & n14088 ;
  assign n14090 = n13926 | n14088 ;
  assign n14091 = ~n14089 & n14090 ;
  assign n14092 = n13910 & ~n14091 ;
  assign n14093 = n14091 | n14092 ;
  assign n14094 = ( ~n13910 & n14092 ) | ( ~n13910 & n14093 ) | ( n14092 & n14093 ) ;
  assign n14095 = x106 & n2280 ;
  assign n14096 = x105 & n2275 ;
  assign n14097 = x104 & ~n2274 ;
  assign n14098 = n2481 & n14097 ;
  assign n14099 = n14096 | n14098 ;
  assign n14100 = n14095 | n14099 ;
  assign n14101 = n2283 | n14100 ;
  assign n14102 = ( n5814 & n14100 ) | ( n5814 & n14101 ) | ( n14100 & n14101 ) ;
  assign n14103 = x26 & n14102 ;
  assign n14104 = x26 & ~n14103 ;
  assign n14105 = ( n14102 & ~n14103 ) | ( n14102 & n14104 ) | ( ~n14103 & n14104 ) ;
  assign n14106 = n13685 | n13691 ;
  assign n14107 = n14105 | n14106 ;
  assign n14108 = n14105 & n14106 ;
  assign n14109 = n14107 & ~n14108 ;
  assign n14110 = n13704 | n13708 ;
  assign n14111 = x109 & n1817 ;
  assign n14112 = x108 & n1812 ;
  assign n14113 = x107 & ~n1811 ;
  assign n14114 = n1977 & n14113 ;
  assign n14115 = n14112 | n14114 ;
  assign n14116 = n14111 | n14115 ;
  assign n14117 = n1820 | n14116 ;
  assign n14118 = ( n6884 & n14116 ) | ( n6884 & n14117 ) | ( n14116 & n14117 ) ;
  assign n14119 = x23 & n14118 ;
  assign n14120 = x23 & ~n14119 ;
  assign n14121 = ( n14118 & ~n14119 ) | ( n14118 & n14120 ) | ( ~n14119 & n14120 ) ;
  assign n14122 = n14110 | n14121 ;
  assign n14123 = ~n14121 & n14122 ;
  assign n14124 = ( ~n14110 & n14122 ) | ( ~n14110 & n14123 ) | ( n14122 & n14123 ) ;
  assign n14125 = ( n14094 & ~n14109 ) | ( n14094 & n14124 ) | ( ~n14109 & n14124 ) ;
  assign n14126 = ( n14109 & ~n14124 ) | ( n14109 & n14125 ) | ( ~n14124 & n14125 ) ;
  assign n14127 = ( ~n14094 & n14125 ) | ( ~n14094 & n14126 ) | ( n14125 & n14126 ) ;
  assign n14128 = x115 & n1071 ;
  assign n14129 = x114 & n1066 ;
  assign n14130 = x113 & ~n1065 ;
  assign n14131 = n1189 & n14130 ;
  assign n14132 = n14129 | n14131 ;
  assign n14133 = n14128 | n14132 ;
  assign n14134 = n1074 | n14133 ;
  assign n14135 = ( n8749 & n14133 ) | ( n8749 & n14134 ) | ( n14133 & n14134 ) ;
  assign n14136 = x17 & n14135 ;
  assign n14137 = x17 & ~n14136 ;
  assign n14138 = ( n14135 & ~n14136 ) | ( n14135 & n14137 ) | ( ~n14136 & n14137 ) ;
  assign n14139 = n13744 | n14138 ;
  assign n14140 = n13748 | n14139 ;
  assign n14141 = ( n13744 & n13748 ) | ( n13744 & n14138 ) | ( n13748 & n14138 ) ;
  assign n14142 = n14140 & ~n14141 ;
  assign n14143 = x112 & n1421 ;
  assign n14144 = x111 & n1416 ;
  assign n14145 = x110 & ~n1415 ;
  assign n14146 = n1584 & n14145 ;
  assign n14147 = n14144 | n14146 ;
  assign n14148 = n14143 | n14147 ;
  assign n14149 = n1424 | n14148 ;
  assign n14150 = ( n7789 & n14148 ) | ( n7789 & n14149 ) | ( n14148 & n14149 ) ;
  assign n14151 = x20 & n14150 ;
  assign n14152 = x20 & ~n14151 ;
  assign n14153 = ( n14150 & ~n14151 ) | ( n14150 & n14152 ) | ( ~n14151 & n14152 ) ;
  assign n14154 = n13722 | n13730 ;
  assign n14155 = n14153 | n14154 ;
  assign n14156 = n14153 & n14154 ;
  assign n14157 = n14155 & ~n14156 ;
  assign n14158 = ( n14127 & n14142 ) | ( n14127 & ~n14157 ) | ( n14142 & ~n14157 ) ;
  assign n14159 = ( ~n14142 & n14157 ) | ( ~n14142 & n14158 ) | ( n14157 & n14158 ) ;
  assign n14160 = ( ~n14127 & n14158 ) | ( ~n14127 & n14159 ) | ( n14158 & n14159 ) ;
  assign n14161 = n13895 & n14160 ;
  assign n14162 = n13895 | n14160 ;
  assign n14163 = ~n14161 & n14162 ;
  assign n14164 = x121 & n528 ;
  assign n14165 = x120 & n523 ;
  assign n14166 = x119 & ~n522 ;
  assign n14167 = n635 & n14166 ;
  assign n14168 = n14165 | n14167 ;
  assign n14169 = n14164 | n14168 ;
  assign n14170 = n531 | n14169 ;
  assign n14171 = ( n10811 & n14169 ) | ( n10811 & n14170 ) | ( n14169 & n14170 ) ;
  assign n14172 = x11 & n14171 ;
  assign n14173 = x11 & ~n14172 ;
  assign n14174 = ( n14171 & ~n14172 ) | ( n14171 & n14173 ) | ( ~n14172 & n14173 ) ;
  assign n14175 = n13780 | n13786 ;
  assign n14176 = ( n14163 & n14174 ) | ( n14163 & ~n14175 ) | ( n14174 & ~n14175 ) ;
  assign n14177 = ( ~n14174 & n14175 ) | ( ~n14174 & n14176 ) | ( n14175 & n14176 ) ;
  assign n14178 = ( ~n14163 & n14176 ) | ( ~n14163 & n14177 ) | ( n14176 & n14177 ) ;
  assign n14179 = x124 & n337 ;
  assign n14180 = x123 & n332 ;
  assign n14181 = x122 & ~n331 ;
  assign n14182 = n396 & n14181 ;
  assign n14183 = n14180 | n14182 ;
  assign n14184 = n14179 | n14183 ;
  assign n14185 = n340 | n14184 ;
  assign n14186 = ( n11916 & n14184 ) | ( n11916 & n14185 ) | ( n14184 & n14185 ) ;
  assign n14187 = x8 & n14186 ;
  assign n14188 = x8 & ~n14187 ;
  assign n14189 = ( n14186 & ~n14187 ) | ( n14186 & n14188 ) | ( ~n14187 & n14188 ) ;
  assign n14190 = n13811 & n14189 ;
  assign n14191 = n14189 & ~n14190 ;
  assign n14192 = ( n13811 & ~n14190 ) | ( n13811 & n14191 ) | ( ~n14190 & n14191 ) ;
  assign n14193 = n14178 & n14192 ;
  assign n14194 = n14178 | n14192 ;
  assign n14195 = ~n14193 & n14194 ;
  assign n14196 = n13878 & n14195 ;
  assign n14197 = n13878 | n14195 ;
  assign n14198 = ~n14196 & n14197 ;
  assign n14199 = n13862 | n14198 ;
  assign n14200 = n13862 & n14198 ;
  assign n14201 = n14199 & ~n14200 ;
  assign n14202 = n13856 | n13860 ;
  assign n14203 = n14201 | n14202 ;
  assign n14204 = n14201 & n14202 ;
  assign n14205 = n14203 & ~n14204 ;
  assign n14206 = n13875 | n14196 ;
  assign n14207 = x127 & n201 ;
  assign n14208 = x126 & ~n200 ;
  assign n14209 = n243 & n14208 ;
  assign n14210 = n14207 | n14209 ;
  assign n14211 = n209 | n14210 ;
  assign n14212 = ( n13461 & n14210 ) | ( n13461 & n14211 ) | ( n14210 & n14211 ) ;
  assign n14213 = x5 & n14212 ;
  assign n14214 = x5 & ~n14213 ;
  assign n14215 = ( n14212 & ~n14213 ) | ( n14212 & n14214 ) | ( ~n14213 & n14214 ) ;
  assign n14216 = n14190 & n14215 ;
  assign n14217 = n14215 & ~n14216 ;
  assign n14218 = ~n14193 & n14217 ;
  assign n14219 = ( n14163 & n14174 ) | ( n14163 & n14175 ) | ( n14174 & n14175 ) ;
  assign n14220 = x125 & n337 ;
  assign n14221 = x124 & n332 ;
  assign n14222 = x123 & ~n331 ;
  assign n14223 = n396 & n14222 ;
  assign n14224 = n14221 | n14223 ;
  assign n14225 = n14220 | n14224 ;
  assign n14226 = n340 | n14225 ;
  assign n14227 = ( n12310 & n14225 ) | ( n12310 & n14226 ) | ( n14225 & n14226 ) ;
  assign n14228 = x8 & n14227 ;
  assign n14229 = x8 & ~n14228 ;
  assign n14230 = ( n14227 & ~n14228 ) | ( n14227 & n14229 ) | ( ~n14228 & n14229 ) ;
  assign n14231 = n14219 & n14230 ;
  assign n14232 = n14219 & ~n14231 ;
  assign n14233 = ~n14219 & n14230 ;
  assign n14234 = n14232 | n14233 ;
  assign n14235 = x101 & n3314 ;
  assign n14236 = x100 & n3309 ;
  assign n14237 = x99 & ~n3308 ;
  assign n14238 = n3570 & n14237 ;
  assign n14239 = n14236 | n14238 ;
  assign n14240 = n14235 | n14239 ;
  assign n14241 = n3317 | n14240 ;
  assign n14242 = ( n4783 & n14240 ) | ( n4783 & n14241 ) | ( n14240 & n14241 ) ;
  assign n14243 = x32 & n14242 ;
  assign n14244 = x32 & ~n14243 ;
  assign n14245 = ( n14242 & ~n14243 ) | ( n14242 & n14244 ) | ( ~n14243 & n14244 ) ;
  assign n14246 = n14086 & n14245 ;
  assign n14247 = n14086 | n14245 ;
  assign n14248 = ~n14246 & n14247 ;
  assign n14249 = x98 & n3913 ;
  assign n14250 = x97 & n3908 ;
  assign n14251 = x96 & ~n3907 ;
  assign n14252 = n4152 & n14251 ;
  assign n14253 = n14250 | n14252 ;
  assign n14254 = n14249 | n14253 ;
  assign n14255 = n3916 | n14254 ;
  assign n14256 = ( n4105 & n14254 ) | ( n4105 & n14255 ) | ( n14254 & n14255 ) ;
  assign n14257 = x35 & n14256 ;
  assign n14258 = x35 & ~n14257 ;
  assign n14259 = ( n14256 & ~n14257 ) | ( n14256 & n14258 ) | ( ~n14257 & n14258 ) ;
  assign n14260 = ( n13939 & n13940 ) | ( n13939 & n14054 ) | ( n13940 & n14054 ) ;
  assign n14261 = x92 & n5340 ;
  assign n14262 = x91 & n5335 ;
  assign n14263 = x90 & ~n5334 ;
  assign n14264 = n5580 & n14263 ;
  assign n14265 = n14262 | n14264 ;
  assign n14266 = n14261 | n14265 ;
  assign n14267 = n5343 | n14266 ;
  assign n14268 = ( n2904 & n14266 ) | ( n2904 & n14267 ) | ( n14266 & n14267 ) ;
  assign n14269 = x41 & n14268 ;
  assign n14270 = x41 & ~n14269 ;
  assign n14271 = ( n14268 & ~n14269 ) | ( n14268 & n14270 ) | ( ~n14269 & n14270 ) ;
  assign n14272 = x89 & n6068 ;
  assign n14273 = x88 & n6063 ;
  assign n14274 = x87 & ~n6062 ;
  assign n14275 = n6398 & n14274 ;
  assign n14276 = n14273 | n14275 ;
  assign n14277 = n14272 | n14276 ;
  assign n14278 = n6071 | n14277 ;
  assign n14279 = ( n2244 & n14277 ) | ( n2244 & n14278 ) | ( n14277 & n14278 ) ;
  assign n14280 = x44 & n14279 ;
  assign n14281 = x44 & ~n14280 ;
  assign n14282 = ( n14279 & ~n14280 ) | ( n14279 & n14281 ) | ( ~n14280 & n14281 ) ;
  assign n14283 = n14025 | n14039 ;
  assign n14284 = x86 & n6937 ;
  assign n14285 = x85 & n6932 ;
  assign n14286 = x84 & ~n6931 ;
  assign n14287 = n7216 & n14286 ;
  assign n14288 = n14285 | n14287 ;
  assign n14289 = n14284 | n14288 ;
  assign n14290 = n6940 | n14289 ;
  assign n14291 = ( n1921 & n14289 ) | ( n1921 & n14290 ) | ( n14289 & n14290 ) ;
  assign n14292 = x47 & n14291 ;
  assign n14293 = x47 & ~n14292 ;
  assign n14294 = ( n14291 & ~n14292 ) | ( n14291 & n14293 ) | ( ~n14292 & n14293 ) ;
  assign n14295 = ( n13953 & n13954 ) | ( n13953 & n14020 ) | ( n13954 & n14020 ) ;
  assign n14296 = x83 & n7812 ;
  assign n14297 = x82 & n7807 ;
  assign n14298 = x81 & ~n7806 ;
  assign n14299 = n8136 & n14298 ;
  assign n14300 = n14297 | n14299 ;
  assign n14301 = n14296 | n14300 ;
  assign n14302 = n7815 | n14301 ;
  assign n14303 = ( n1510 & n14301 ) | ( n1510 & n14302 ) | ( n14301 & n14302 ) ;
  assign n14304 = x50 & n14303 ;
  assign n14305 = x50 & ~n14304 ;
  assign n14306 = ( n14303 & ~n14304 ) | ( n14303 & n14305 ) | ( ~n14304 & n14305 ) ;
  assign n14307 = ( n13965 & n13966 ) | ( n13965 & n14017 ) | ( n13966 & n14017 ) ;
  assign n14308 = ( n13977 & n13978 ) | ( n13977 & n14014 ) | ( n13978 & n14014 ) ;
  assign n14309 = n13983 | n13997 ;
  assign n14310 = x71 & n11984 ;
  assign n14311 = x70 & n11979 ;
  assign n14312 = x69 & ~n11978 ;
  assign n14313 = n12430 & n14312 ;
  assign n14314 = n14311 | n14313 ;
  assign n14315 = n14310 | n14314 ;
  assign n14316 = n11987 | n14315 ;
  assign n14317 = ( n376 & n14315 ) | ( n376 & n14316 ) | ( n14315 & n14316 ) ;
  assign n14318 = x62 & ~n14317 ;
  assign n14319 = ~x62 & n14317 ;
  assign n14320 = n14318 | n14319 ;
  assign n14321 = x68 & n12808 ;
  assign n14322 = x63 & x67 ;
  assign n14323 = ~n12808 & n14322 ;
  assign n14324 = n14321 | n14323 ;
  assign n14325 = x2 & n14324 ;
  assign n14326 = n14324 & ~n14325 ;
  assign n14327 = x2 & ~n14324 ;
  assign n14328 = n14326 | n14327 ;
  assign n14329 = n14320 & n14328 ;
  assign n14330 = n14320 | n14328 ;
  assign n14331 = ~n14329 & n14330 ;
  assign n14332 = x74 & n10876 ;
  assign n14333 = x73 & n10871 ;
  assign n14334 = x72 & ~n10870 ;
  assign n14335 = n11305 & n14334 ;
  assign n14336 = n14333 | n14335 ;
  assign n14337 = n14332 | n14336 ;
  assign n14338 = n10879 | n14337 ;
  assign n14339 = ( n587 & n14337 ) | ( n587 & n14338 ) | ( n14337 & n14338 ) ;
  assign n14340 = x59 & n14339 ;
  assign n14341 = x59 & ~n14340 ;
  assign n14342 = ( n14339 & ~n14340 ) | ( n14339 & n14341 ) | ( ~n14340 & n14341 ) ;
  assign n14343 = ( n14309 & n14331 ) | ( n14309 & n14342 ) | ( n14331 & n14342 ) ;
  assign n14344 = ( n14331 & n14342 ) | ( n14331 & ~n14343 ) | ( n14342 & ~n14343 ) ;
  assign n14345 = ( n14309 & ~n14343 ) | ( n14309 & n14344 ) | ( ~n14343 & n14344 ) ;
  assign n14346 = n14012 | n14345 ;
  assign n14347 = n14012 & n14345 ;
  assign n14348 = n14346 & ~n14347 ;
  assign n14349 = x77 & n9853 ;
  assign n14350 = x76 & n9848 ;
  assign n14351 = x75 & ~n9847 ;
  assign n14352 = n10165 & n14351 ;
  assign n14353 = n14350 | n14352 ;
  assign n14354 = n14349 | n14353 ;
  assign n14355 = n9856 | n14354 ;
  assign n14356 = ( n846 & n14354 ) | ( n846 & n14355 ) | ( n14354 & n14355 ) ;
  assign n14357 = x56 & n14356 ;
  assign n14358 = x56 & ~n14357 ;
  assign n14359 = ( n14356 & ~n14357 ) | ( n14356 & n14358 ) | ( ~n14357 & n14358 ) ;
  assign n14360 = n14348 | n14359 ;
  assign n14361 = n14348 & n14359 ;
  assign n14362 = n14360 & ~n14361 ;
  assign n14363 = x80 & n8834 ;
  assign n14364 = x79 & n8829 ;
  assign n14365 = x78 & ~n8828 ;
  assign n14366 = n9159 & n14365 ;
  assign n14367 = n14364 | n14366 ;
  assign n14368 = n14363 | n14367 ;
  assign n14369 = n8837 | n14368 ;
  assign n14370 = ( n1147 & n14368 ) | ( n1147 & n14369 ) | ( n14368 & n14369 ) ;
  assign n14371 = x53 & n14370 ;
  assign n14372 = x53 & ~n14371 ;
  assign n14373 = ( n14370 & ~n14371 ) | ( n14370 & n14372 ) | ( ~n14371 & n14372 ) ;
  assign n14374 = ( n14308 & n14362 ) | ( n14308 & n14373 ) | ( n14362 & n14373 ) ;
  assign n14375 = ( n14362 & n14373 ) | ( n14362 & ~n14374 ) | ( n14373 & ~n14374 ) ;
  assign n14376 = ( n14308 & ~n14374 ) | ( n14308 & n14375 ) | ( ~n14374 & n14375 ) ;
  assign n14377 = ( n14306 & ~n14307 ) | ( n14306 & n14376 ) | ( ~n14307 & n14376 ) ;
  assign n14378 = ( n14307 & ~n14376 ) | ( n14307 & n14377 ) | ( ~n14376 & n14377 ) ;
  assign n14379 = ( ~n14306 & n14377 ) | ( ~n14306 & n14378 ) | ( n14377 & n14378 ) ;
  assign n14380 = ( n14294 & n14295 ) | ( n14294 & ~n14379 ) | ( n14295 & ~n14379 ) ;
  assign n14381 = ( ~n14295 & n14379 ) | ( ~n14295 & n14380 ) | ( n14379 & n14380 ) ;
  assign n14382 = ( ~n14294 & n14380 ) | ( ~n14294 & n14381 ) | ( n14380 & n14381 ) ;
  assign n14383 = ( n14282 & ~n14283 ) | ( n14282 & n14382 ) | ( ~n14283 & n14382 ) ;
  assign n14384 = ( n14283 & ~n14382 ) | ( n14283 & n14383 ) | ( ~n14382 & n14383 ) ;
  assign n14385 = ( ~n14282 & n14383 ) | ( ~n14282 & n14384 ) | ( n14383 & n14384 ) ;
  assign n14386 = ( ~n14052 & n14271 ) | ( ~n14052 & n14385 ) | ( n14271 & n14385 ) ;
  assign n14387 = ( n14052 & ~n14385 ) | ( n14052 & n14386 ) | ( ~n14385 & n14386 ) ;
  assign n14388 = ( ~n14271 & n14386 ) | ( ~n14271 & n14387 ) | ( n14386 & n14387 ) ;
  assign n14389 = n14260 | n14388 ;
  assign n14390 = n14260 & n14388 ;
  assign n14391 = n14389 & ~n14390 ;
  assign n14392 = x95 & n4572 ;
  assign n14393 = x94 & n4567 ;
  assign n14394 = x93 & ~n4566 ;
  assign n14395 = n4828 & n14394 ;
  assign n14396 = n14393 | n14395 ;
  assign n14397 = n14392 | n14396 ;
  assign n14398 = n4575 | n14397 ;
  assign n14399 = ( n3479 & n14397 ) | ( n3479 & n14398 ) | ( n14397 & n14398 ) ;
  assign n14400 = x38 & n14399 ;
  assign n14401 = x38 & ~n14400 ;
  assign n14402 = ( n14399 & ~n14400 ) | ( n14399 & n14401 ) | ( ~n14400 & n14401 ) ;
  assign n14403 = n14391 | n14402 ;
  assign n14404 = n14391 & n14402 ;
  assign n14405 = n14403 & ~n14404 ;
  assign n14406 = n14059 | n14073 ;
  assign n14407 = n14405 & n14406 ;
  assign n14408 = n14406 & ~n14407 ;
  assign n14409 = ( n14405 & ~n14407 ) | ( n14405 & n14408 ) | ( ~n14407 & n14408 ) ;
  assign n14410 = n14259 & ~n14409 ;
  assign n14411 = ~n14259 & n14409 ;
  assign n14412 = n14410 | n14411 ;
  assign n14413 = n14248 | n14412 ;
  assign n14414 = n14248 & n14412 ;
  assign n14415 = n14413 & ~n14414 ;
  assign n14416 = x104 & n2775 ;
  assign n14417 = x103 & n2770 ;
  assign n14418 = x102 & ~n2769 ;
  assign n14419 = n2978 & n14418 ;
  assign n14420 = n14417 | n14419 ;
  assign n14421 = n14416 | n14420 ;
  assign n14422 = n2778 | n14421 ;
  assign n14423 = ( n5295 & n14421 ) | ( n5295 & n14422 ) | ( n14421 & n14422 ) ;
  assign n14424 = x29 & n14423 ;
  assign n14425 = x29 & ~n14424 ;
  assign n14426 = ( n14423 & ~n14424 ) | ( n14423 & n14425 ) | ( ~n14424 & n14425 ) ;
  assign n14427 = ( n13652 & n13921 ) | ( n13652 & n13922 ) | ( n13921 & n13922 ) ;
  assign n14428 = n14426 & n14427 ;
  assign n14429 = n14426 & ~n14428 ;
  assign n14430 = ~n14089 & n14429 ;
  assign n14431 = ( n14089 & ~n14426 ) | ( n14089 & n14427 ) | ( ~n14426 & n14427 ) ;
  assign n14432 = n14430 | n14431 ;
  assign n14433 = n14415 & n14432 ;
  assign n14434 = n14415 | n14432 ;
  assign n14435 = ~n14433 & n14434 ;
  assign n14436 = x107 & n2280 ;
  assign n14437 = x106 & n2275 ;
  assign n14438 = x105 & ~n2274 ;
  assign n14439 = n2481 & n14438 ;
  assign n14440 = n14437 | n14439 ;
  assign n14441 = n14436 | n14440 ;
  assign n14442 = n2283 | n14441 ;
  assign n14443 = ( n6328 & n14441 ) | ( n6328 & n14442 ) | ( n14441 & n14442 ) ;
  assign n14444 = x26 & n14443 ;
  assign n14445 = x26 & ~n14444 ;
  assign n14446 = ( n14443 & ~n14444 ) | ( n14443 & n14445 ) | ( ~n14444 & n14445 ) ;
  assign n14447 = ( n13908 & n13909 ) | ( n13908 & n14091 ) | ( n13909 & n14091 ) ;
  assign n14448 = ( n14435 & n14446 ) | ( n14435 & ~n14447 ) | ( n14446 & ~n14447 ) ;
  assign n14449 = ( ~n14446 & n14447 ) | ( ~n14446 & n14448 ) | ( n14447 & n14448 ) ;
  assign n14450 = ( ~n14435 & n14448 ) | ( ~n14435 & n14449 ) | ( n14448 & n14449 ) ;
  assign n14451 = x110 & n1817 ;
  assign n14452 = x109 & n1812 ;
  assign n14453 = x108 & ~n1811 ;
  assign n14454 = n1977 & n14453 ;
  assign n14455 = n14452 | n14454 ;
  assign n14456 = n14451 | n14455 ;
  assign n14457 = n1820 | n14456 ;
  assign n14458 = ( n7189 & n14456 ) | ( n7189 & n14457 ) | ( n14456 & n14457 ) ;
  assign n14459 = x23 & n14458 ;
  assign n14460 = x23 & ~n14459 ;
  assign n14461 = ( n14458 & ~n14459 ) | ( n14458 & n14460 ) | ( ~n14459 & n14460 ) ;
  assign n14462 = ( n14094 & n14105 ) | ( n14094 & n14106 ) | ( n14105 & n14106 ) ;
  assign n14463 = ( n14450 & n14461 ) | ( n14450 & ~n14462 ) | ( n14461 & ~n14462 ) ;
  assign n14464 = ( ~n14461 & n14462 ) | ( ~n14461 & n14463 ) | ( n14462 & n14463 ) ;
  assign n14465 = ( ~n14450 & n14463 ) | ( ~n14450 & n14464 ) | ( n14463 & n14464 ) ;
  assign n14466 = x113 & n1421 ;
  assign n14467 = x112 & n1416 ;
  assign n14468 = x111 & ~n1415 ;
  assign n14469 = n1584 & n14468 ;
  assign n14470 = n14467 | n14469 ;
  assign n14471 = n14466 | n14470 ;
  assign n14472 = n1424 | n14471 ;
  assign n14473 = ( n8113 & n14471 ) | ( n8113 & n14472 ) | ( n14471 & n14472 ) ;
  assign n14474 = x20 & n14473 ;
  assign n14475 = x20 & ~n14474 ;
  assign n14476 = ( n14473 & ~n14474 ) | ( n14473 & n14475 ) | ( ~n14474 & n14475 ) ;
  assign n14477 = n14124 & ~n14127 ;
  assign n14478 = ( n13704 & n13708 ) | ( n13704 & n14121 ) | ( n13708 & n14121 ) ;
  assign n14479 = n14477 | n14478 ;
  assign n14480 = ( n14465 & n14476 ) | ( n14465 & ~n14479 ) | ( n14476 & ~n14479 ) ;
  assign n14481 = ( ~n14476 & n14479 ) | ( ~n14476 & n14480 ) | ( n14479 & n14480 ) ;
  assign n14482 = ( ~n14465 & n14480 ) | ( ~n14465 & n14481 ) | ( n14480 & n14481 ) ;
  assign n14483 = x116 & n1071 ;
  assign n14484 = x115 & n1066 ;
  assign n14485 = x114 & ~n1065 ;
  assign n14486 = n1189 & n14485 ;
  assign n14487 = n14484 | n14486 ;
  assign n14488 = n14483 | n14487 ;
  assign n14489 = n1074 | n14488 ;
  assign n14490 = ( n8778 & n14488 ) | ( n8778 & n14489 ) | ( n14488 & n14489 ) ;
  assign n14491 = x17 & n14490 ;
  assign n14492 = x17 & ~n14491 ;
  assign n14493 = ( n14490 & ~n14491 ) | ( n14490 & n14492 ) | ( ~n14491 & n14492 ) ;
  assign n14494 = ( n14127 & n14153 ) | ( n14127 & n14154 ) | ( n14153 & n14154 ) ;
  assign n14495 = ( n14482 & n14493 ) | ( n14482 & ~n14494 ) | ( n14493 & ~n14494 ) ;
  assign n14496 = ( ~n14493 & n14494 ) | ( ~n14493 & n14495 ) | ( n14494 & n14495 ) ;
  assign n14497 = ( ~n14482 & n14495 ) | ( ~n14482 & n14496 ) | ( n14495 & n14496 ) ;
  assign n14498 = x119 & n771 ;
  assign n14499 = x118 & n766 ;
  assign n14500 = x117 & ~n765 ;
  assign n14501 = n905 & n14500 ;
  assign n14502 = n14499 | n14501 ;
  assign n14503 = n14498 | n14502 ;
  assign n14504 = n774 | n14503 ;
  assign n14505 = ( n9789 & n14503 ) | ( n9789 & n14504 ) | ( n14503 & n14504 ) ;
  assign n14506 = x14 & n14505 ;
  assign n14507 = x14 & ~n14506 ;
  assign n14508 = ( n14505 & ~n14506 ) | ( n14505 & n14507 ) | ( ~n14506 & n14507 ) ;
  assign n14509 = n14142 & ~n14160 ;
  assign n14510 = n14141 | n14509 ;
  assign n14511 = ( n14497 & n14508 ) | ( n14497 & ~n14510 ) | ( n14508 & ~n14510 ) ;
  assign n14512 = ( ~n14508 & n14510 ) | ( ~n14508 & n14511 ) | ( n14510 & n14511 ) ;
  assign n14513 = ( ~n14497 & n14511 ) | ( ~n14497 & n14512 ) | ( n14511 & n14512 ) ;
  assign n14514 = x122 & n528 ;
  assign n14515 = x121 & n523 ;
  assign n14516 = x120 & ~n522 ;
  assign n14517 = n635 & n14516 ;
  assign n14518 = n14515 | n14517 ;
  assign n14519 = n14514 | n14518 ;
  assign n14520 = n531 | n14519 ;
  assign n14521 = ( n11188 & n14519 ) | ( n11188 & n14520 ) | ( n14519 & n14520 ) ;
  assign n14522 = x11 & n14521 ;
  assign n14523 = x11 & ~n14522 ;
  assign n14524 = ( n14521 & ~n14522 ) | ( n14521 & n14523 ) | ( ~n14522 & n14523 ) ;
  assign n14525 = ( n13893 & n14161 ) | ( n13893 & n14524 ) | ( n14161 & n14524 ) ;
  assign n14526 = ( n13893 & n14161 ) | ( n13893 & ~n14524 ) | ( n14161 & ~n14524 ) ;
  assign n14527 = ( n14524 & ~n14525 ) | ( n14524 & n14526 ) | ( ~n14525 & n14526 ) ;
  assign n14528 = n14513 & n14527 ;
  assign n14529 = n14513 | n14527 ;
  assign n14530 = ~n14528 & n14529 ;
  assign n14531 = n14234 & n14530 ;
  assign n14532 = n14234 | n14530 ;
  assign n14533 = ~n14531 & n14532 ;
  assign n14534 = n14218 | n14533 ;
  assign n14535 = ( n14190 & n14193 ) | ( n14190 & ~n14215 ) | ( n14193 & ~n14215 ) ;
  assign n14536 = n14534 | n14535 ;
  assign n14537 = ( n14218 & n14533 ) | ( n14218 & n14535 ) | ( n14533 & n14535 ) ;
  assign n14538 = n14536 & ~n14537 ;
  assign n14539 = ~n14206 & n14538 ;
  assign n14540 = n14200 | n14204 ;
  assign n14541 = ( n14206 & ~n14538 ) | ( n14206 & n14540 ) | ( ~n14538 & n14540 ) ;
  assign n14542 = n14206 & n14538 ;
  assign n14543 = n14206 & ~n14542 ;
  assign n14544 = n14539 | n14543 ;
  assign n14545 = ( n14200 & n14204 ) | ( n14200 & n14544 ) | ( n14204 & n14544 ) ;
  assign n14546 = ( n14539 & n14541 ) | ( n14539 & ~n14545 ) | ( n14541 & ~n14545 ) ;
  assign n14547 = x126 & n337 ;
  assign n14548 = x125 & n332 ;
  assign n14549 = x124 & ~n331 ;
  assign n14550 = n396 & n14549 ;
  assign n14551 = n14548 | n14550 ;
  assign n14552 = n14547 | n14551 ;
  assign n14553 = n340 | n14552 ;
  assign n14554 = ( n12687 & n14552 ) | ( n12687 & n14553 ) | ( n14552 & n14553 ) ;
  assign n14555 = x8 & n14554 ;
  assign n14556 = x8 & ~n14555 ;
  assign n14557 = ( n14554 & ~n14555 ) | ( n14554 & n14556 ) | ( ~n14555 & n14556 ) ;
  assign n14558 = n14525 & n14557 ;
  assign n14559 = n14557 & ~n14558 ;
  assign n14560 = ~n14528 & n14559 ;
  assign n14561 = x120 & n771 ;
  assign n14562 = x119 & n766 ;
  assign n14563 = x118 & ~n765 ;
  assign n14564 = n905 & n14563 ;
  assign n14565 = n14562 | n14564 ;
  assign n14566 = n14561 | n14565 ;
  assign n14567 = n774 | n14566 ;
  assign n14568 = ( n10460 & n14566 ) | ( n10460 & n14567 ) | ( n14566 & n14567 ) ;
  assign n14569 = x14 & n14568 ;
  assign n14570 = x14 & ~n14569 ;
  assign n14571 = ( n14568 & ~n14569 ) | ( n14568 & n14570 ) | ( ~n14569 & n14570 ) ;
  assign n14572 = n14493 & n14494 ;
  assign n14573 = n14482 & ~n14496 ;
  assign n14574 = ( n14482 & ~n14495 ) | ( n14482 & n14573 ) | ( ~n14495 & n14573 ) ;
  assign n14575 = n14572 | n14574 ;
  assign n14576 = x114 & n1421 ;
  assign n14577 = x113 & n1416 ;
  assign n14578 = x112 & ~n1415 ;
  assign n14579 = n1584 & n14578 ;
  assign n14580 = n14577 | n14579 ;
  assign n14581 = n14576 | n14580 ;
  assign n14582 = n1424 | n14581 ;
  assign n14583 = ( n8437 & n14581 ) | ( n8437 & n14582 ) | ( n14581 & n14582 ) ;
  assign n14584 = x20 & n14583 ;
  assign n14585 = x20 & ~n14584 ;
  assign n14586 = ( n14583 & ~n14584 ) | ( n14583 & n14585 ) | ( ~n14584 & n14585 ) ;
  assign n14587 = n14461 & n14462 ;
  assign n14588 = n14450 & ~n14464 ;
  assign n14589 = ( n14450 & ~n14463 ) | ( n14450 & n14588 ) | ( ~n14463 & n14588 ) ;
  assign n14590 = n14587 | n14589 ;
  assign n14591 = n14390 | n14404 ;
  assign n14592 = ( n14052 & n14271 ) | ( n14052 & n14385 ) | ( n14271 & n14385 ) ;
  assign n14593 = x93 & n5340 ;
  assign n14594 = x92 & n5335 ;
  assign n14595 = x91 & ~n5334 ;
  assign n14596 = n5580 & n14595 ;
  assign n14597 = n14594 | n14596 ;
  assign n14598 = n14593 | n14597 ;
  assign n14599 = n5343 | n14598 ;
  assign n14600 = ( n2931 & n14598 ) | ( n2931 & n14599 ) | ( n14598 & n14599 ) ;
  assign n14601 = x41 & n14600 ;
  assign n14602 = x41 & ~n14601 ;
  assign n14603 = ( n14600 & ~n14601 ) | ( n14600 & n14602 ) | ( ~n14601 & n14602 ) ;
  assign n14604 = ( n14282 & n14283 ) | ( n14282 & n14382 ) | ( n14283 & n14382 ) ;
  assign n14605 = x90 & n6068 ;
  assign n14606 = x89 & n6063 ;
  assign n14607 = x88 & ~n6062 ;
  assign n14608 = n6398 & n14607 ;
  assign n14609 = n14606 | n14608 ;
  assign n14610 = n14605 | n14609 ;
  assign n14611 = n6071 | n14610 ;
  assign n14612 = ( n2410 & n14610 ) | ( n2410 & n14611 ) | ( n14610 & n14611 ) ;
  assign n14613 = x44 & n14612 ;
  assign n14614 = x44 & ~n14613 ;
  assign n14615 = ( n14612 & ~n14613 ) | ( n14612 & n14614 ) | ( ~n14613 & n14614 ) ;
  assign n14616 = ( n14294 & n14295 ) | ( n14294 & n14379 ) | ( n14295 & n14379 ) ;
  assign n14617 = x87 & n6937 ;
  assign n14618 = x86 & n6932 ;
  assign n14619 = x85 & ~n6931 ;
  assign n14620 = n7216 & n14619 ;
  assign n14621 = n14618 | n14620 ;
  assign n14622 = n14617 | n14621 ;
  assign n14623 = n6940 | n14622 ;
  assign n14624 = ( n2067 & n14622 ) | ( n2067 & n14623 ) | ( n14622 & n14623 ) ;
  assign n14625 = x47 & n14624 ;
  assign n14626 = x47 & ~n14625 ;
  assign n14627 = ( n14624 & ~n14625 ) | ( n14624 & n14626 ) | ( ~n14625 & n14626 ) ;
  assign n14628 = ( n14306 & n14307 ) | ( n14306 & n14376 ) | ( n14307 & n14376 ) ;
  assign n14629 = x78 & n9853 ;
  assign n14630 = x77 & n9848 ;
  assign n14631 = x76 & ~n9847 ;
  assign n14632 = n10165 & n14631 ;
  assign n14633 = n14630 | n14632 ;
  assign n14634 = n14629 | n14633 ;
  assign n14635 = n9856 | n14634 ;
  assign n14636 = ( n868 & n14634 ) | ( n868 & n14635 ) | ( n14634 & n14635 ) ;
  assign n14637 = x56 & n14636 ;
  assign n14638 = x56 & ~n14637 ;
  assign n14639 = ( n14636 & ~n14637 ) | ( n14636 & n14638 ) | ( ~n14637 & n14638 ) ;
  assign n14640 = x69 & n12808 ;
  assign n14641 = x63 & x68 ;
  assign n14642 = ~n12808 & n14641 ;
  assign n14643 = n14640 | n14642 ;
  assign n14644 = x2 & n14643 ;
  assign n14645 = n14643 & ~n14644 ;
  assign n14646 = x2 & ~n14643 ;
  assign n14647 = n14645 | n14646 ;
  assign n14648 = x72 & n11984 ;
  assign n14649 = x71 & n11979 ;
  assign n14650 = x70 & ~n11978 ;
  assign n14651 = n12430 & n14650 ;
  assign n14652 = n14649 | n14651 ;
  assign n14653 = n14648 | n14652 ;
  assign n14654 = ( n435 & n11987 ) | ( n435 & n14653 ) | ( n11987 & n14653 ) ;
  assign n14655 = ( x62 & ~n14653 ) | ( x62 & n14654 ) | ( ~n14653 & n14654 ) ;
  assign n14656 = ~n14654 & n14655 ;
  assign n14657 = n14653 | n14655 ;
  assign n14658 = ( ~x62 & n14656 ) | ( ~x62 & n14657 ) | ( n14656 & n14657 ) ;
  assign n14659 = ~n14647 & n14658 ;
  assign n14660 = n14325 | n14329 ;
  assign n14661 = n14647 & ~n14658 ;
  assign n14662 = n14660 | n14661 ;
  assign n14663 = n14659 | n14662 ;
  assign n14664 = ( n14659 & n14660 ) | ( n14659 & n14661 ) | ( n14660 & n14661 ) ;
  assign n14665 = n14663 & ~n14664 ;
  assign n14666 = x75 & n10876 ;
  assign n14667 = x74 & n10871 ;
  assign n14668 = x73 & ~n10870 ;
  assign n14669 = n11305 & n14668 ;
  assign n14670 = n14667 | n14669 ;
  assign n14671 = n14666 | n14670 ;
  assign n14672 = n10879 | n14671 ;
  assign n14673 = ( n609 & n14671 ) | ( n609 & n14672 ) | ( n14671 & n14672 ) ;
  assign n14674 = x59 & n14673 ;
  assign n14675 = x59 & ~n14674 ;
  assign n14676 = ( n14673 & ~n14674 ) | ( n14673 & n14675 ) | ( ~n14674 & n14675 ) ;
  assign n14677 = n14665 | n14676 ;
  assign n14678 = n14665 & n14676 ;
  assign n14679 = n14677 & ~n14678 ;
  assign n14680 = ( n14343 & n14639 ) | ( n14343 & ~n14679 ) | ( n14639 & ~n14679 ) ;
  assign n14681 = ( ~n14343 & n14679 ) | ( ~n14343 & n14680 ) | ( n14679 & n14680 ) ;
  assign n14682 = ( ~n14639 & n14680 ) | ( ~n14639 & n14681 ) | ( n14680 & n14681 ) ;
  assign n14683 = n14347 | n14361 ;
  assign n14684 = n14682 & n14683 ;
  assign n14685 = n14682 & ~n14684 ;
  assign n14686 = ~n14682 & n14683 ;
  assign n14687 = n14685 | n14686 ;
  assign n14688 = x81 & n8834 ;
  assign n14689 = x80 & n8829 ;
  assign n14690 = x79 & ~n8828 ;
  assign n14691 = n9159 & n14690 ;
  assign n14692 = n14689 | n14691 ;
  assign n14693 = n14688 | n14692 ;
  assign n14694 = n8837 | n14693 ;
  assign n14695 = ( n1256 & n14693 ) | ( n1256 & n14694 ) | ( n14693 & n14694 ) ;
  assign n14696 = x53 & n14695 ;
  assign n14697 = x53 & ~n14696 ;
  assign n14698 = ( n14695 & ~n14696 ) | ( n14695 & n14697 ) | ( ~n14696 & n14697 ) ;
  assign n14699 = n14687 & n14698 ;
  assign n14700 = n14687 | n14698 ;
  assign n14701 = ~n14699 & n14700 ;
  assign n14702 = n14374 | n14701 ;
  assign n14703 = n14374 & n14701 ;
  assign n14704 = n14702 & ~n14703 ;
  assign n14705 = x84 & n7812 ;
  assign n14706 = x83 & n7807 ;
  assign n14707 = x82 & ~n7806 ;
  assign n14708 = n8136 & n14707 ;
  assign n14709 = n14706 | n14708 ;
  assign n14710 = n14705 | n14709 ;
  assign n14711 = n7815 | n14710 ;
  assign n14712 = ( n1537 & n14710 ) | ( n1537 & n14711 ) | ( n14710 & n14711 ) ;
  assign n14713 = x50 & n14712 ;
  assign n14714 = x50 & ~n14713 ;
  assign n14715 = ( n14712 & ~n14713 ) | ( n14712 & n14714 ) | ( ~n14713 & n14714 ) ;
  assign n14716 = n14704 | n14715 ;
  assign n14717 = n14704 & n14715 ;
  assign n14718 = n14716 & ~n14717 ;
  assign n14719 = ( n14627 & n14628 ) | ( n14627 & ~n14718 ) | ( n14628 & ~n14718 ) ;
  assign n14720 = ( ~n14628 & n14718 ) | ( ~n14628 & n14719 ) | ( n14718 & n14719 ) ;
  assign n14721 = ( ~n14627 & n14719 ) | ( ~n14627 & n14720 ) | ( n14719 & n14720 ) ;
  assign n14722 = ( n14615 & n14616 ) | ( n14615 & ~n14721 ) | ( n14616 & ~n14721 ) ;
  assign n14723 = ( ~n14616 & n14721 ) | ( ~n14616 & n14722 ) | ( n14721 & n14722 ) ;
  assign n14724 = ( ~n14615 & n14722 ) | ( ~n14615 & n14723 ) | ( n14722 & n14723 ) ;
  assign n14725 = ( n14603 & ~n14604 ) | ( n14603 & n14724 ) | ( ~n14604 & n14724 ) ;
  assign n14726 = ( n14604 & ~n14724 ) | ( n14604 & n14725 ) | ( ~n14724 & n14725 ) ;
  assign n14727 = ( ~n14603 & n14725 ) | ( ~n14603 & n14726 ) | ( n14725 & n14726 ) ;
  assign n14728 = n14592 | n14727 ;
  assign n14729 = n14592 & n14727 ;
  assign n14730 = n14728 & ~n14729 ;
  assign n14731 = x96 & n4572 ;
  assign n14732 = x95 & n4567 ;
  assign n14733 = x94 & ~n4566 ;
  assign n14734 = n4828 & n14733 ;
  assign n14735 = n14732 | n14734 ;
  assign n14736 = n14731 | n14735 ;
  assign n14737 = n4575 | n14736 ;
  assign n14738 = ( n3509 & n14736 ) | ( n3509 & n14737 ) | ( n14736 & n14737 ) ;
  assign n14739 = x38 & n14738 ;
  assign n14740 = x38 & ~n14739 ;
  assign n14741 = ( n14738 & ~n14739 ) | ( n14738 & n14740 ) | ( ~n14739 & n14740 ) ;
  assign n14742 = n14730 | n14741 ;
  assign n14743 = n14730 & n14741 ;
  assign n14744 = n14742 & ~n14743 ;
  assign n14745 = x99 & n3913 ;
  assign n14746 = x98 & n3908 ;
  assign n14747 = x97 & ~n3907 ;
  assign n14748 = n4152 & n14747 ;
  assign n14749 = n14746 | n14748 ;
  assign n14750 = n14745 | n14749 ;
  assign n14751 = n3916 | n14750 ;
  assign n14752 = ( n4325 & n14750 ) | ( n4325 & n14751 ) | ( n14750 & n14751 ) ;
  assign n14753 = x35 & n14752 ;
  assign n14754 = x35 & ~n14753 ;
  assign n14755 = ( n14752 & ~n14753 ) | ( n14752 & n14754 ) | ( ~n14753 & n14754 ) ;
  assign n14756 = ( n14591 & n14744 ) | ( n14591 & n14755 ) | ( n14744 & n14755 ) ;
  assign n14757 = ( n14744 & n14755 ) | ( n14744 & ~n14756 ) | ( n14755 & ~n14756 ) ;
  assign n14758 = ( n14591 & ~n14756 ) | ( n14591 & n14757 ) | ( ~n14756 & n14757 ) ;
  assign n14759 = x102 & n3314 ;
  assign n14760 = x101 & n3309 ;
  assign n14761 = x100 & ~n3308 ;
  assign n14762 = n3570 & n14761 ;
  assign n14763 = n14760 | n14762 ;
  assign n14764 = n14759 | n14763 ;
  assign n14765 = n3317 | n14764 ;
  assign n14766 = ( n5025 & n14764 ) | ( n5025 & n14765 ) | ( n14764 & n14765 ) ;
  assign n14767 = x32 & n14766 ;
  assign n14768 = x32 & ~n14767 ;
  assign n14769 = ( n14766 & ~n14767 ) | ( n14766 & n14768 ) | ( ~n14767 & n14768 ) ;
  assign n14770 = ( n14407 & n14409 ) | ( n14407 & ~n14411 ) | ( n14409 & ~n14411 ) ;
  assign n14771 = ( n14758 & n14769 ) | ( n14758 & ~n14770 ) | ( n14769 & ~n14770 ) ;
  assign n14772 = ( ~n14769 & n14770 ) | ( ~n14769 & n14771 ) | ( n14770 & n14771 ) ;
  assign n14773 = ( ~n14758 & n14771 ) | ( ~n14758 & n14772 ) | ( n14771 & n14772 ) ;
  assign n14774 = x105 & n2775 ;
  assign n14775 = x104 & n2770 ;
  assign n14776 = x103 & ~n2769 ;
  assign n14777 = n2978 & n14776 ;
  assign n14778 = n14775 | n14777 ;
  assign n14779 = n14774 | n14778 ;
  assign n14780 = n2778 | n14779 ;
  assign n14781 = ( n5788 & n14779 ) | ( n5788 & n14780 ) | ( n14779 & n14780 ) ;
  assign n14782 = x29 & n14781 ;
  assign n14783 = x29 & ~n14782 ;
  assign n14784 = ( n14781 & ~n14782 ) | ( n14781 & n14783 ) | ( ~n14782 & n14783 ) ;
  assign n14785 = n14246 | n14414 ;
  assign n14786 = ( n14773 & n14784 ) | ( n14773 & ~n14785 ) | ( n14784 & ~n14785 ) ;
  assign n14787 = ( ~n14784 & n14785 ) | ( ~n14784 & n14786 ) | ( n14785 & n14786 ) ;
  assign n14788 = ( ~n14773 & n14786 ) | ( ~n14773 & n14787 ) | ( n14786 & n14787 ) ;
  assign n14789 = x108 & n2280 ;
  assign n14790 = x107 & n2275 ;
  assign n14791 = x106 & ~n2274 ;
  assign n14792 = n2481 & n14791 ;
  assign n14793 = n14790 | n14792 ;
  assign n14794 = n14789 | n14793 ;
  assign n14795 = n2283 | n14794 ;
  assign n14796 = ( n6358 & n14794 ) | ( n6358 & n14795 ) | ( n14794 & n14795 ) ;
  assign n14797 = x26 & n14796 ;
  assign n14798 = x26 & ~n14797 ;
  assign n14799 = ( n14796 & ~n14797 ) | ( n14796 & n14798 ) | ( ~n14797 & n14798 ) ;
  assign n14800 = ( n14089 & n14426 ) | ( n14089 & n14428 ) | ( n14426 & n14428 ) ;
  assign n14801 = n14799 & n14800 ;
  assign n14802 = ( n14433 & n14799 ) | ( n14433 & n14801 ) | ( n14799 & n14801 ) ;
  assign n14803 = n14433 | n14800 ;
  assign n14804 = ~n14799 & n14803 ;
  assign n14805 = ( n14799 & ~n14802 ) | ( n14799 & n14804 ) | ( ~n14802 & n14804 ) ;
  assign n14806 = n14788 & n14805 ;
  assign n14807 = n14788 | n14805 ;
  assign n14808 = ~n14806 & n14807 ;
  assign n14809 = ( n14435 & n14446 ) | ( n14435 & n14447 ) | ( n14446 & n14447 ) ;
  assign n14810 = x111 & n1817 ;
  assign n14811 = x110 & n1812 ;
  assign n14812 = x109 & ~n1811 ;
  assign n14813 = n1977 & n14812 ;
  assign n14814 = n14811 | n14813 ;
  assign n14815 = n14810 | n14814 ;
  assign n14816 = n1820 | n14815 ;
  assign n14817 = ( n7492 & n14815 ) | ( n7492 & n14816 ) | ( n14815 & n14816 ) ;
  assign n14818 = x23 & n14817 ;
  assign n14819 = x23 & ~n14818 ;
  assign n14820 = ( n14817 & ~n14818 ) | ( n14817 & n14819 ) | ( ~n14818 & n14819 ) ;
  assign n14821 = ( n14808 & n14809 ) | ( n14808 & ~n14820 ) | ( n14809 & ~n14820 ) ;
  assign n14822 = ( ~n14809 & n14820 ) | ( ~n14809 & n14821 ) | ( n14820 & n14821 ) ;
  assign n14823 = ( ~n14808 & n14821 ) | ( ~n14808 & n14822 ) | ( n14821 & n14822 ) ;
  assign n14824 = ( n14586 & ~n14590 ) | ( n14586 & n14823 ) | ( ~n14590 & n14823 ) ;
  assign n14825 = ( n14590 & ~n14823 ) | ( n14590 & n14824 ) | ( ~n14823 & n14824 ) ;
  assign n14826 = ( ~n14586 & n14824 ) | ( ~n14586 & n14825 ) | ( n14824 & n14825 ) ;
  assign n14827 = ( n14465 & n14476 ) | ( n14465 & n14479 ) | ( n14476 & n14479 ) ;
  assign n14828 = x117 & n1071 ;
  assign n14829 = x116 & n1066 ;
  assign n14830 = x115 & ~n1065 ;
  assign n14831 = n1189 & n14830 ;
  assign n14832 = n14829 | n14831 ;
  assign n14833 = n14828 | n14832 ;
  assign n14834 = n1074 | n14833 ;
  assign n14835 = ( n9118 & n14833 ) | ( n9118 & n14834 ) | ( n14833 & n14834 ) ;
  assign n14836 = x17 & n14835 ;
  assign n14837 = x17 & ~n14836 ;
  assign n14838 = ( n14835 & ~n14836 ) | ( n14835 & n14837 ) | ( ~n14836 & n14837 ) ;
  assign n14839 = ( n14826 & n14827 ) | ( n14826 & ~n14838 ) | ( n14827 & ~n14838 ) ;
  assign n14840 = ( ~n14827 & n14838 ) | ( ~n14827 & n14839 ) | ( n14838 & n14839 ) ;
  assign n14841 = ( ~n14826 & n14839 ) | ( ~n14826 & n14840 ) | ( n14839 & n14840 ) ;
  assign n14842 = ( n14571 & ~n14575 ) | ( n14571 & n14841 ) | ( ~n14575 & n14841 ) ;
  assign n14843 = ( n14575 & ~n14841 ) | ( n14575 & n14842 ) | ( ~n14841 & n14842 ) ;
  assign n14844 = ( ~n14571 & n14842 ) | ( ~n14571 & n14843 ) | ( n14842 & n14843 ) ;
  assign n14845 = ( n14497 & n14508 ) | ( n14497 & n14510 ) | ( n14508 & n14510 ) ;
  assign n14846 = x123 & n528 ;
  assign n14847 = x122 & n523 ;
  assign n14848 = x121 & ~n522 ;
  assign n14849 = n635 & n14848 ;
  assign n14850 = n14847 | n14849 ;
  assign n14851 = n14846 | n14850 ;
  assign n14852 = n531 | n14851 ;
  assign n14853 = ( n11219 & n14851 ) | ( n11219 & n14852 ) | ( n14851 & n14852 ) ;
  assign n14854 = x11 & n14853 ;
  assign n14855 = x11 & ~n14854 ;
  assign n14856 = ( n14853 & ~n14854 ) | ( n14853 & n14855 ) | ( ~n14854 & n14855 ) ;
  assign n14857 = ( n14844 & n14845 ) | ( n14844 & ~n14856 ) | ( n14845 & ~n14856 ) ;
  assign n14858 = ( ~n14845 & n14856 ) | ( ~n14845 & n14857 ) | ( n14856 & n14857 ) ;
  assign n14859 = ( ~n14844 & n14857 ) | ( ~n14844 & n14858 ) | ( n14857 & n14858 ) ;
  assign n14860 = n14560 | n14859 ;
  assign n14861 = ( n14525 & n14528 ) | ( n14525 & ~n14557 ) | ( n14528 & ~n14557 ) ;
  assign n14862 = n14860 | n14861 ;
  assign n14863 = ( n14560 & n14859 ) | ( n14560 & n14861 ) | ( n14859 & n14861 ) ;
  assign n14864 = n14862 & ~n14863 ;
  assign n14865 = x127 & ~n200 ;
  assign n14866 = n243 & n14865 ;
  assign n14867 = ( x127 & n209 ) | ( x127 & n14866 ) | ( n209 & n14866 ) ;
  assign n14868 = ( x126 & n14866 ) | ( x126 & n14867 ) | ( n14866 & n14867 ) ;
  assign n14869 = ( n12685 & n14867 ) | ( n12685 & n14868 ) | ( n14867 & n14868 ) ;
  assign n14870 = x5 & n14869 ;
  assign n14871 = x5 & ~n14870 ;
  assign n14872 = ( n14869 & ~n14870 ) | ( n14869 & n14871 ) | ( ~n14870 & n14871 ) ;
  assign n14873 = n14231 & n14872 ;
  assign n14874 = n14872 & ~n14873 ;
  assign n14875 = ~n14531 & n14874 ;
  assign n14876 = n14864 | n14875 ;
  assign n14877 = ( n14231 & n14531 ) | ( n14231 & ~n14872 ) | ( n14531 & ~n14872 ) ;
  assign n14878 = n14876 | n14877 ;
  assign n14879 = ( n14864 & n14875 ) | ( n14864 & n14877 ) | ( n14875 & n14877 ) ;
  assign n14880 = n14878 & ~n14879 ;
  assign n14881 = ( n14193 & n14215 ) | ( n14193 & n14216 ) | ( n14215 & n14216 ) ;
  assign n14882 = n14537 | n14881 ;
  assign n14883 = n14880 & n14882 ;
  assign n14884 = n14882 & ~n14883 ;
  assign n14885 = ( n14880 & ~n14883 ) | ( n14880 & n14884 ) | ( ~n14883 & n14884 ) ;
  assign n14886 = n14542 | n14545 ;
  assign n14887 = n14885 | n14886 ;
  assign n14888 = ~n14886 & n14887 ;
  assign n14889 = ( ~n14885 & n14887 ) | ( ~n14885 & n14888 ) | ( n14887 & n14888 ) ;
  assign n14890 = x127 & n337 ;
  assign n14891 = x126 & n332 ;
  assign n14892 = x125 & ~n331 ;
  assign n14893 = n396 & n14892 ;
  assign n14894 = n14891 | n14893 ;
  assign n14895 = n14890 | n14894 ;
  assign n14896 = n340 | n14895 ;
  assign n14897 = ( n12720 & n14895 ) | ( n12720 & n14896 ) | ( n14895 & n14896 ) ;
  assign n14898 = x8 & n14897 ;
  assign n14899 = x8 & ~n14898 ;
  assign n14900 = ( n14897 & ~n14898 ) | ( n14897 & n14899 ) | ( ~n14898 & n14899 ) ;
  assign n14901 = ( n14528 & n14557 ) | ( n14528 & n14558 ) | ( n14557 & n14558 ) ;
  assign n14902 = n14863 | n14901 ;
  assign n14903 = x121 & n771 ;
  assign n14904 = x120 & n766 ;
  assign n14905 = x119 & ~n765 ;
  assign n14906 = n905 & n14905 ;
  assign n14907 = n14904 | n14906 ;
  assign n14908 = n14903 | n14907 ;
  assign n14909 = n774 | n14908 ;
  assign n14910 = ( n10811 & n14908 ) | ( n10811 & n14909 ) | ( n14908 & n14909 ) ;
  assign n14911 = x14 & n14910 ;
  assign n14912 = x14 & ~n14911 ;
  assign n14913 = ( n14910 & ~n14911 ) | ( n14910 & n14912 ) | ( ~n14911 & n14912 ) ;
  assign n14914 = ( n14571 & n14572 ) | ( n14571 & n14574 ) | ( n14572 & n14574 ) ;
  assign n14915 = n14913 | n14914 ;
  assign n14916 = n14571 & ~n14575 ;
  assign n14917 = ( n14841 & ~n14842 ) | ( n14841 & n14916 ) | ( ~n14842 & n14916 ) ;
  assign n14918 = n14915 | n14917 ;
  assign n14919 = ( n14913 & n14914 ) | ( n14913 & n14917 ) | ( n14914 & n14917 ) ;
  assign n14920 = n14918 & ~n14919 ;
  assign n14921 = x115 & n1421 ;
  assign n14922 = x114 & n1416 ;
  assign n14923 = x113 & ~n1415 ;
  assign n14924 = n1584 & n14923 ;
  assign n14925 = n14922 | n14924 ;
  assign n14926 = n14921 | n14925 ;
  assign n14927 = n1424 | n14926 ;
  assign n14928 = ( n8749 & n14926 ) | ( n8749 & n14927 ) | ( n14926 & n14927 ) ;
  assign n14929 = x20 & n14928 ;
  assign n14930 = x20 & ~n14929 ;
  assign n14931 = ( n14928 & ~n14929 ) | ( n14928 & n14930 ) | ( ~n14929 & n14930 ) ;
  assign n14932 = ( n14586 & n14587 ) | ( n14586 & n14589 ) | ( n14587 & n14589 ) ;
  assign n14933 = n14931 | n14932 ;
  assign n14934 = n14586 & ~n14590 ;
  assign n14935 = ( n14823 & ~n14824 ) | ( n14823 & n14934 ) | ( ~n14824 & n14934 ) ;
  assign n14936 = n14933 | n14935 ;
  assign n14937 = ( n14931 & n14932 ) | ( n14931 & n14935 ) | ( n14932 & n14935 ) ;
  assign n14938 = n14936 & ~n14937 ;
  assign n14939 = x109 & n2280 ;
  assign n14940 = x108 & n2275 ;
  assign n14941 = x107 & ~n2274 ;
  assign n14942 = n2481 & n14941 ;
  assign n14943 = n14940 | n14942 ;
  assign n14944 = n14939 | n14943 ;
  assign n14945 = n2283 | n14944 ;
  assign n14946 = ( n6884 & n14944 ) | ( n6884 & n14945 ) | ( n14944 & n14945 ) ;
  assign n14947 = x26 & n14946 ;
  assign n14948 = x26 & ~n14947 ;
  assign n14949 = ( n14946 & ~n14947 ) | ( n14946 & n14948 ) | ( ~n14947 & n14948 ) ;
  assign n14950 = n14802 | n14806 ;
  assign n14951 = ( n14773 & n14784 ) | ( n14773 & n14785 ) | ( n14784 & n14785 ) ;
  assign n14952 = x106 & n2775 ;
  assign n14953 = x105 & n2770 ;
  assign n14954 = x104 & ~n2769 ;
  assign n14955 = n2978 & n14954 ;
  assign n14956 = n14953 | n14955 ;
  assign n14957 = n14952 | n14956 ;
  assign n14958 = n2778 | n14957 ;
  assign n14959 = ( n5814 & n14957 ) | ( n5814 & n14958 ) | ( n14957 & n14958 ) ;
  assign n14960 = x29 & n14959 ;
  assign n14961 = x29 & ~n14960 ;
  assign n14962 = ( n14959 & ~n14960 ) | ( n14959 & n14961 ) | ( ~n14960 & n14961 ) ;
  assign n14963 = n14951 | n14962 ;
  assign n14964 = n14951 & n14962 ;
  assign n14965 = n14963 & ~n14964 ;
  assign n14966 = x97 & n4572 ;
  assign n14967 = x96 & n4567 ;
  assign n14968 = x95 & ~n4566 ;
  assign n14969 = n4828 & n14968 ;
  assign n14970 = n14967 | n14969 ;
  assign n14971 = n14966 | n14970 ;
  assign n14972 = n4575 | n14971 ;
  assign n14973 = ( n3707 & n14971 ) | ( n3707 & n14972 ) | ( n14971 & n14972 ) ;
  assign n14974 = x38 & n14973 ;
  assign n14975 = x38 & ~n14974 ;
  assign n14976 = ( n14973 & ~n14974 ) | ( n14973 & n14975 ) | ( ~n14974 & n14975 ) ;
  assign n14977 = x94 & n5340 ;
  assign n14978 = x93 & n5335 ;
  assign n14979 = x92 & ~n5334 ;
  assign n14980 = n5580 & n14979 ;
  assign n14981 = n14978 | n14980 ;
  assign n14982 = n14977 | n14981 ;
  assign n14983 = n5343 | n14982 ;
  assign n14984 = ( n3271 & n14982 ) | ( n3271 & n14983 ) | ( n14982 & n14983 ) ;
  assign n14985 = x41 & n14984 ;
  assign n14986 = x41 & ~n14985 ;
  assign n14987 = ( n14984 & ~n14985 ) | ( n14984 & n14986 ) | ( ~n14985 & n14986 ) ;
  assign n14988 = ( n14603 & n14604 ) | ( n14603 & n14724 ) | ( n14604 & n14724 ) ;
  assign n14989 = ( n14615 & n14616 ) | ( n14615 & n14721 ) | ( n14616 & n14721 ) ;
  assign n14990 = n14703 | n14717 ;
  assign n14991 = ( n14644 & n14658 ) | ( n14644 & ~n14659 ) | ( n14658 & ~n14659 ) ;
  assign n14992 = x70 & n12808 ;
  assign n14993 = x63 & x69 ;
  assign n14994 = ~n12808 & n14993 ;
  assign n14995 = n14992 | n14994 ;
  assign n14996 = ( x2 & x5 ) | ( x2 & ~n14995 ) | ( x5 & ~n14995 ) ;
  assign n14997 = ( ~x5 & n14995 ) | ( ~x5 & n14996 ) | ( n14995 & n14996 ) ;
  assign n14998 = ( ~x2 & n14996 ) | ( ~x2 & n14997 ) | ( n14996 & n14997 ) ;
  assign n14999 = n14991 & n14998 ;
  assign n15000 = n14991 | n14998 ;
  assign n15001 = ~n14999 & n15000 ;
  assign n15002 = x73 & n11984 ;
  assign n15003 = x72 & n11979 ;
  assign n15004 = x71 & ~n11978 ;
  assign n15005 = n12430 & n15004 ;
  assign n15006 = n15003 | n15005 ;
  assign n15007 = n15002 | n15006 ;
  assign n15008 = ( n499 & n11987 ) | ( n499 & n15007 ) | ( n11987 & n15007 ) ;
  assign n15009 = ( x62 & ~n15007 ) | ( x62 & n15008 ) | ( ~n15007 & n15008 ) ;
  assign n15010 = ~n15008 & n15009 ;
  assign n15011 = n15007 | n15009 ;
  assign n15012 = ( ~x62 & n15010 ) | ( ~x62 & n15011 ) | ( n15010 & n15011 ) ;
  assign n15013 = n15001 | n15012 ;
  assign n15014 = n15001 & n15012 ;
  assign n15015 = n15013 & ~n15014 ;
  assign n15016 = x76 & n10876 ;
  assign n15017 = x75 & n10871 ;
  assign n15018 = x74 & ~n10870 ;
  assign n15019 = n11305 & n15018 ;
  assign n15020 = n15017 | n15019 ;
  assign n15021 = n15016 | n15020 ;
  assign n15022 = n10879 | n15021 ;
  assign n15023 = ( n740 & n15021 ) | ( n740 & n15022 ) | ( n15021 & n15022 ) ;
  assign n15024 = x59 & n15023 ;
  assign n15025 = x59 & ~n15024 ;
  assign n15026 = ( n15023 & ~n15024 ) | ( n15023 & n15025 ) | ( ~n15024 & n15025 ) ;
  assign n15027 = n15015 & n15026 ;
  assign n15028 = n15015 & ~n15027 ;
  assign n15029 = ~n15015 & n15026 ;
  assign n15030 = n15028 | n15029 ;
  assign n15031 = n14664 | n14678 ;
  assign n15032 = n15030 & n15031 ;
  assign n15033 = n15030 | n15031 ;
  assign n15034 = ~n15032 & n15033 ;
  assign n15035 = x79 & n9853 ;
  assign n15036 = x78 & n9848 ;
  assign n15037 = x77 & ~n9847 ;
  assign n15038 = n10165 & n15037 ;
  assign n15039 = n15036 | n15038 ;
  assign n15040 = n15035 | n15039 ;
  assign n15041 = n9856 | n15040 ;
  assign n15042 = ( n961 & n15040 ) | ( n961 & n15041 ) | ( n15040 & n15041 ) ;
  assign n15043 = x56 & n15042 ;
  assign n15044 = x56 & ~n15043 ;
  assign n15045 = ( n15042 & ~n15043 ) | ( n15042 & n15044 ) | ( ~n15043 & n15044 ) ;
  assign n15046 = n15034 & n15045 ;
  assign n15047 = n15034 & ~n15046 ;
  assign n15048 = ~n15034 & n15045 ;
  assign n15049 = ( n14343 & n14639 ) | ( n14343 & n14679 ) | ( n14639 & n14679 ) ;
  assign n15050 = n15048 | n15049 ;
  assign n15051 = n15047 | n15050 ;
  assign n15052 = ( n15047 & n15048 ) | ( n15047 & n15049 ) | ( n15048 & n15049 ) ;
  assign n15053 = n15051 & ~n15052 ;
  assign n15054 = x82 & n8834 ;
  assign n15055 = x81 & n8829 ;
  assign n15056 = x80 & ~n8828 ;
  assign n15057 = n9159 & n15056 ;
  assign n15058 = n15055 | n15057 ;
  assign n15059 = n15054 | n15058 ;
  assign n15060 = n8837 | n15059 ;
  assign n15061 = ( n1371 & n15059 ) | ( n1371 & n15060 ) | ( n15059 & n15060 ) ;
  assign n15062 = x53 & n15061 ;
  assign n15063 = x53 & ~n15062 ;
  assign n15064 = ( n15061 & ~n15062 ) | ( n15061 & n15063 ) | ( ~n15062 & n15063 ) ;
  assign n15065 = n15053 & n15064 ;
  assign n15066 = n15053 & ~n15065 ;
  assign n15067 = ~n15053 & n15064 ;
  assign n15068 = n15066 | n15067 ;
  assign n15069 = n14684 | n14699 ;
  assign n15070 = n15068 | n15069 ;
  assign n15071 = n15068 & n15069 ;
  assign n15072 = n15070 & ~n15071 ;
  assign n15073 = x85 & n7812 ;
  assign n15074 = x84 & n7807 ;
  assign n15075 = x83 & ~n7806 ;
  assign n15076 = n8136 & n15075 ;
  assign n15077 = n15074 | n15076 ;
  assign n15078 = n15073 | n15077 ;
  assign n15079 = n7815 | n15078 ;
  assign n15080 = ( n1765 & n15078 ) | ( n1765 & n15079 ) | ( n15078 & n15079 ) ;
  assign n15081 = x50 & n15080 ;
  assign n15082 = x50 & ~n15081 ;
  assign n15083 = ( n15080 & ~n15081 ) | ( n15080 & n15082 ) | ( ~n15081 & n15082 ) ;
  assign n15084 = ( n14990 & n15072 ) | ( n14990 & ~n15083 ) | ( n15072 & ~n15083 ) ;
  assign n15085 = ( ~n15072 & n15083 ) | ( ~n15072 & n15084 ) | ( n15083 & n15084 ) ;
  assign n15086 = ( ~n14990 & n15084 ) | ( ~n14990 & n15085 ) | ( n15084 & n15085 ) ;
  assign n15087 = x88 & n6937 ;
  assign n15088 = x87 & n6932 ;
  assign n15089 = x86 & ~n6931 ;
  assign n15090 = n7216 & n15089 ;
  assign n15091 = n15088 | n15090 ;
  assign n15092 = n15087 | n15091 ;
  assign n15093 = n6940 | n15092 ;
  assign n15094 = ( n2095 & n15092 ) | ( n2095 & n15093 ) | ( n15092 & n15093 ) ;
  assign n15095 = x47 & n15094 ;
  assign n15096 = x47 & ~n15095 ;
  assign n15097 = ( n15094 & ~n15095 ) | ( n15094 & n15096 ) | ( ~n15095 & n15096 ) ;
  assign n15098 = n15086 & n15097 ;
  assign n15099 = n15086 | n15097 ;
  assign n15100 = ~n15098 & n15099 ;
  assign n15101 = ( n14627 & n14628 ) | ( n14627 & n14718 ) | ( n14628 & n14718 ) ;
  assign n15102 = n15100 | n15101 ;
  assign n15103 = n15100 & n15101 ;
  assign n15104 = n15102 & ~n15103 ;
  assign n15105 = x91 & n6068 ;
  assign n15106 = x90 & n6063 ;
  assign n15107 = x89 & ~n6062 ;
  assign n15108 = n6398 & n15107 ;
  assign n15109 = n15106 | n15108 ;
  assign n15110 = n15105 | n15109 ;
  assign n15111 = n6071 | n15110 ;
  assign n15112 = ( n2714 & n15110 ) | ( n2714 & n15111 ) | ( n15110 & n15111 ) ;
  assign n15113 = x44 & n15112 ;
  assign n15114 = x44 & ~n15113 ;
  assign n15115 = ( n15112 & ~n15113 ) | ( n15112 & n15114 ) | ( ~n15113 & n15114 ) ;
  assign n15116 = n15104 & n15115 ;
  assign n15117 = n15104 & ~n15116 ;
  assign n15118 = ~n15104 & n15115 ;
  assign n15119 = n15117 | n15118 ;
  assign n15120 = n14989 | n15119 ;
  assign n15121 = n14989 & n15119 ;
  assign n15122 = n15120 & ~n15121 ;
  assign n15123 = ( n14987 & n14988 ) | ( n14987 & ~n15122 ) | ( n14988 & ~n15122 ) ;
  assign n15124 = ( ~n14988 & n15122 ) | ( ~n14988 & n15123 ) | ( n15122 & n15123 ) ;
  assign n15125 = ( ~n14987 & n15123 ) | ( ~n14987 & n15124 ) | ( n15123 & n15124 ) ;
  assign n15126 = n14976 & n15125 ;
  assign n15127 = n14976 | n15125 ;
  assign n15128 = ~n15126 & n15127 ;
  assign n15129 = n14729 | n14743 ;
  assign n15130 = ~n15128 & n15129 ;
  assign n15131 = n15128 & ~n15129 ;
  assign n15132 = n15130 | n15131 ;
  assign n15133 = x100 & n3913 ;
  assign n15134 = x99 & n3908 ;
  assign n15135 = x98 & ~n3907 ;
  assign n15136 = n4152 & n15135 ;
  assign n15137 = n15134 | n15136 ;
  assign n15138 = n15133 | n15137 ;
  assign n15139 = n3916 | n15138 ;
  assign n15140 = ( n4532 & n15138 ) | ( n4532 & n15139 ) | ( n15138 & n15139 ) ;
  assign n15141 = x35 & n15140 ;
  assign n15142 = x35 & ~n15141 ;
  assign n15143 = ( n15140 & ~n15141 ) | ( n15140 & n15142 ) | ( ~n15141 & n15142 ) ;
  assign n15144 = n15132 & n15143 ;
  assign n15145 = n15132 | n15143 ;
  assign n15146 = ~n15144 & n15145 ;
  assign n15147 = n14756 | n15146 ;
  assign n15148 = n14756 & n15146 ;
  assign n15149 = n15147 & ~n15148 ;
  assign n15150 = x103 & n3314 ;
  assign n15151 = x102 & n3309 ;
  assign n15152 = x101 & ~n3308 ;
  assign n15153 = n3570 & n15152 ;
  assign n15154 = n15151 | n15153 ;
  assign n15155 = n15150 | n15154 ;
  assign n15156 = n3317 | n15155 ;
  assign n15157 = ( n5264 & n15155 ) | ( n5264 & n15156 ) | ( n15155 & n15156 ) ;
  assign n15158 = x32 & n15157 ;
  assign n15159 = x32 & ~n15158 ;
  assign n15160 = ( n15157 & ~n15158 ) | ( n15157 & n15159 ) | ( ~n15158 & n15159 ) ;
  assign n15161 = ( n14758 & n14769 ) | ( n14758 & n14770 ) | ( n14769 & n14770 ) ;
  assign n15162 = n15160 | n15161 ;
  assign n15163 = n15160 & n15161 ;
  assign n15164 = n15162 & ~n15163 ;
  assign n15165 = n15149 & n15164 ;
  assign n15166 = n15149 | n15164 ;
  assign n15167 = ~n15165 & n15166 ;
  assign n15168 = n14965 & n15167 ;
  assign n15169 = n14965 | n15167 ;
  assign n15170 = ~n15168 & n15169 ;
  assign n15171 = ( n14949 & ~n14950 ) | ( n14949 & n15170 ) | ( ~n14950 & n15170 ) ;
  assign n15172 = ( n14950 & ~n15170 ) | ( n14950 & n15171 ) | ( ~n15170 & n15171 ) ;
  assign n15173 = ( ~n14949 & n15171 ) | ( ~n14949 & n15172 ) | ( n15171 & n15172 ) ;
  assign n15174 = ( n14808 & n14809 ) | ( n14808 & n14820 ) | ( n14809 & n14820 ) ;
  assign n15175 = x112 & n1817 ;
  assign n15176 = x111 & n1812 ;
  assign n15177 = x110 & ~n1811 ;
  assign n15178 = n1977 & n15177 ;
  assign n15179 = n15176 | n15178 ;
  assign n15180 = n15175 | n15179 ;
  assign n15181 = n1820 | n15180 ;
  assign n15182 = ( n7789 & n15180 ) | ( n7789 & n15181 ) | ( n15180 & n15181 ) ;
  assign n15183 = x23 & n15182 ;
  assign n15184 = x23 & ~n15183 ;
  assign n15185 = ( n15182 & ~n15183 ) | ( n15182 & n15184 ) | ( ~n15183 & n15184 ) ;
  assign n15186 = ( n15173 & n15174 ) | ( n15173 & ~n15185 ) | ( n15174 & ~n15185 ) ;
  assign n15187 = ( ~n15174 & n15185 ) | ( ~n15174 & n15186 ) | ( n15185 & n15186 ) ;
  assign n15188 = ( ~n15173 & n15186 ) | ( ~n15173 & n15187 ) | ( n15186 & n15187 ) ;
  assign n15189 = n14938 & ~n15188 ;
  assign n15190 = n15188 | n15189 ;
  assign n15191 = ( ~n14938 & n15189 ) | ( ~n14938 & n15190 ) | ( n15189 & n15190 ) ;
  assign n15192 = ( n14826 & n14827 ) | ( n14826 & n14838 ) | ( n14827 & n14838 ) ;
  assign n15193 = x118 & n1071 ;
  assign n15194 = x117 & n1066 ;
  assign n15195 = x116 & ~n1065 ;
  assign n15196 = n1189 & n15195 ;
  assign n15197 = n15194 | n15196 ;
  assign n15198 = n15193 | n15197 ;
  assign n15199 = n1074 | n15198 ;
  assign n15200 = ( n9760 & n15198 ) | ( n9760 & n15199 ) | ( n15198 & n15199 ) ;
  assign n15201 = x17 & n15200 ;
  assign n15202 = x17 & ~n15201 ;
  assign n15203 = ( n15200 & ~n15201 ) | ( n15200 & n15202 ) | ( ~n15201 & n15202 ) ;
  assign n15204 = n15192 & n15203 ;
  assign n15205 = n15203 & ~n15204 ;
  assign n15206 = ( n15192 & ~n15204 ) | ( n15192 & n15205 ) | ( ~n15204 & n15205 ) ;
  assign n15207 = n15191 & n15206 ;
  assign n15208 = n15191 | n15206 ;
  assign n15209 = ~n15207 & n15208 ;
  assign n15210 = n14920 & ~n15209 ;
  assign n15211 = n15209 | n15210 ;
  assign n15212 = ( ~n14920 & n15210 ) | ( ~n14920 & n15211 ) | ( n15210 & n15211 ) ;
  assign n15213 = ( n14844 & n14845 ) | ( n14844 & n14856 ) | ( n14845 & n14856 ) ;
  assign n15214 = x124 & n528 ;
  assign n15215 = x123 & n523 ;
  assign n15216 = x122 & ~n522 ;
  assign n15217 = n635 & n15216 ;
  assign n15218 = n15215 | n15217 ;
  assign n15219 = n15214 | n15218 ;
  assign n15220 = n531 | n15219 ;
  assign n15221 = ( n11916 & n15219 ) | ( n11916 & n15220 ) | ( n15219 & n15220 ) ;
  assign n15222 = x11 & n15221 ;
  assign n15223 = x11 & ~n15222 ;
  assign n15224 = ( n15221 & ~n15222 ) | ( n15221 & n15223 ) | ( ~n15222 & n15223 ) ;
  assign n15225 = ( n15212 & n15213 ) | ( n15212 & ~n15224 ) | ( n15213 & ~n15224 ) ;
  assign n15226 = ( ~n15213 & n15224 ) | ( ~n15213 & n15225 ) | ( n15224 & n15225 ) ;
  assign n15227 = ( ~n15212 & n15225 ) | ( ~n15212 & n15226 ) | ( n15225 & n15226 ) ;
  assign n15228 = ( n14900 & ~n14902 ) | ( n14900 & n15227 ) | ( ~n14902 & n15227 ) ;
  assign n15229 = ( n14902 & ~n15227 ) | ( n14902 & n15228 ) | ( ~n15227 & n15228 ) ;
  assign n15230 = ( ~n14900 & n15228 ) | ( ~n14900 & n15229 ) | ( n15228 & n15229 ) ;
  assign n15231 = ( n14531 & n14872 ) | ( n14531 & n14873 ) | ( n14872 & n14873 ) ;
  assign n15232 = n15230 & n15231 ;
  assign n15233 = ( n14879 & n15230 ) | ( n14879 & n15232 ) | ( n15230 & n15232 ) ;
  assign n15234 = n15230 | n15231 ;
  assign n15235 = n14879 | n15234 ;
  assign n15236 = ~n15233 & n15235 ;
  assign n15237 = n14883 | n14885 ;
  assign n15238 = ( n14883 & n14886 ) | ( n14883 & n15237 ) | ( n14886 & n15237 ) ;
  assign n15239 = n15236 | n15238 ;
  assign n15240 = n15236 & n15237 ;
  assign n15241 = n14883 & n15236 ;
  assign n15242 = ( n14886 & n15240 ) | ( n14886 & n15241 ) | ( n15240 & n15241 ) ;
  assign n15243 = n15239 & ~n15242 ;
  assign n15244 = x113 & n1817 ;
  assign n15245 = x112 & n1812 ;
  assign n15246 = x111 & ~n1811 ;
  assign n15247 = n1977 & n15246 ;
  assign n15248 = n15245 | n15247 ;
  assign n15249 = n15244 | n15248 ;
  assign n15250 = n1820 | n15249 ;
  assign n15251 = ( n8113 & n15249 ) | ( n8113 & n15250 ) | ( n15249 & n15250 ) ;
  assign n15252 = x23 & n15251 ;
  assign n15253 = x23 & ~n15252 ;
  assign n15254 = ( n15251 & ~n15252 ) | ( n15251 & n15253 ) | ( ~n15252 & n15253 ) ;
  assign n15255 = ( n14949 & n14950 ) | ( n14949 & n15170 ) | ( n14950 & n15170 ) ;
  assign n15256 = n15128 & n15129 ;
  assign n15257 = n15116 | n15121 ;
  assign n15258 = n15098 | n15103 ;
  assign n15259 = x86 & n7812 ;
  assign n15260 = x85 & n7807 ;
  assign n15261 = x84 & ~n7806 ;
  assign n15262 = n8136 & n15261 ;
  assign n15263 = n15260 | n15262 ;
  assign n15264 = n15259 | n15263 ;
  assign n15265 = n7815 | n15264 ;
  assign n15266 = ( n1921 & n15264 ) | ( n1921 & n15265 ) | ( n15264 & n15265 ) ;
  assign n15267 = x50 & n15266 ;
  assign n15268 = x50 & ~n15267 ;
  assign n15269 = ( n15266 & ~n15267 ) | ( n15266 & n15268 ) | ( ~n15267 & n15268 ) ;
  assign n15270 = n15065 | n15071 ;
  assign n15271 = x83 & n8834 ;
  assign n15272 = x82 & n8829 ;
  assign n15273 = x81 & ~n8828 ;
  assign n15274 = n9159 & n15273 ;
  assign n15275 = n15272 | n15274 ;
  assign n15276 = n15271 | n15275 ;
  assign n15277 = n8837 | n15276 ;
  assign n15278 = ( n1510 & n15276 ) | ( n1510 & n15277 ) | ( n15276 & n15277 ) ;
  assign n15279 = x53 & n15278 ;
  assign n15280 = x53 & ~n15279 ;
  assign n15281 = ( n15278 & ~n15279 ) | ( n15278 & n15280 ) | ( ~n15279 & n15280 ) ;
  assign n15282 = n15046 | n15052 ;
  assign n15283 = x80 & n9853 ;
  assign n15284 = x79 & n9848 ;
  assign n15285 = x78 & ~n9847 ;
  assign n15286 = n10165 & n15285 ;
  assign n15287 = n15284 | n15286 ;
  assign n15288 = n15283 | n15287 ;
  assign n15289 = n9856 | n15288 ;
  assign n15290 = ( n1147 & n15288 ) | ( n1147 & n15289 ) | ( n15288 & n15289 ) ;
  assign n15291 = x56 & n15290 ;
  assign n15292 = x56 & ~n15291 ;
  assign n15293 = ( n15290 & ~n15291 ) | ( n15290 & n15292 ) | ( ~n15291 & n15292 ) ;
  assign n15294 = n15027 | n15032 ;
  assign n15295 = n14999 | n15014 ;
  assign n15296 = x71 & n12808 ;
  assign n15297 = x63 & x70 ;
  assign n15298 = ~n12808 & n15297 ;
  assign n15299 = n15296 | n15298 ;
  assign n15300 = n14996 | n15299 ;
  assign n15301 = n14996 & n15299 ;
  assign n15302 = n15300 & ~n15301 ;
  assign n15303 = x74 & n11984 ;
  assign n15304 = x73 & n11979 ;
  assign n15305 = x72 & ~n11978 ;
  assign n15306 = n12430 & n15305 ;
  assign n15307 = n15304 | n15306 ;
  assign n15308 = n15303 | n15307 ;
  assign n15309 = n11987 | n15308 ;
  assign n15310 = ( n587 & n15308 ) | ( n587 & n15309 ) | ( n15308 & n15309 ) ;
  assign n15311 = x62 & n15310 ;
  assign n15312 = x62 & ~n15311 ;
  assign n15313 = ( n15310 & ~n15311 ) | ( n15310 & n15312 ) | ( ~n15311 & n15312 ) ;
  assign n15314 = n15302 & n15313 ;
  assign n15315 = n15302 | n15313 ;
  assign n15316 = ~n15314 & n15315 ;
  assign n15317 = x77 & n10876 ;
  assign n15318 = x76 & n10871 ;
  assign n15319 = x75 & ~n10870 ;
  assign n15320 = n11305 & n15319 ;
  assign n15321 = n15318 | n15320 ;
  assign n15322 = n15317 | n15321 ;
  assign n15323 = n10879 | n15322 ;
  assign n15324 = ( n846 & n15322 ) | ( n846 & n15323 ) | ( n15322 & n15323 ) ;
  assign n15325 = x59 & n15324 ;
  assign n15326 = x59 & ~n15325 ;
  assign n15327 = ( n15324 & ~n15325 ) | ( n15324 & n15326 ) | ( ~n15325 & n15326 ) ;
  assign n15328 = ( n15295 & n15316 ) | ( n15295 & n15327 ) | ( n15316 & n15327 ) ;
  assign n15329 = ( n15316 & n15327 ) | ( n15316 & ~n15328 ) | ( n15327 & ~n15328 ) ;
  assign n15330 = ( n15295 & ~n15328 ) | ( n15295 & n15329 ) | ( ~n15328 & n15329 ) ;
  assign n15331 = ( n15293 & n15294 ) | ( n15293 & ~n15330 ) | ( n15294 & ~n15330 ) ;
  assign n15332 = ( ~n15294 & n15330 ) | ( ~n15294 & n15331 ) | ( n15330 & n15331 ) ;
  assign n15333 = ( ~n15293 & n15331 ) | ( ~n15293 & n15332 ) | ( n15331 & n15332 ) ;
  assign n15334 = ( n15281 & ~n15282 ) | ( n15281 & n15333 ) | ( ~n15282 & n15333 ) ;
  assign n15335 = ( n15282 & ~n15333 ) | ( n15282 & n15334 ) | ( ~n15333 & n15334 ) ;
  assign n15336 = ( ~n15281 & n15334 ) | ( ~n15281 & n15335 ) | ( n15334 & n15335 ) ;
  assign n15337 = ( n15269 & ~n15270 ) | ( n15269 & n15336 ) | ( ~n15270 & n15336 ) ;
  assign n15338 = ( n15270 & ~n15336 ) | ( n15270 & n15337 ) | ( ~n15336 & n15337 ) ;
  assign n15339 = ( ~n15269 & n15337 ) | ( ~n15269 & n15338 ) | ( n15337 & n15338 ) ;
  assign n15340 = ( n14990 & n15072 ) | ( n14990 & n15083 ) | ( n15072 & n15083 ) ;
  assign n15341 = n15339 | n15340 ;
  assign n15342 = x89 & n6937 ;
  assign n15343 = x88 & n6932 ;
  assign n15344 = x87 & ~n6931 ;
  assign n15345 = n7216 & n15344 ;
  assign n15346 = n15343 | n15345 ;
  assign n15347 = n15342 | n15346 ;
  assign n15348 = n6940 | n15347 ;
  assign n15349 = ( n2244 & n15347 ) | ( n2244 & n15348 ) | ( n15347 & n15348 ) ;
  assign n15350 = x47 & n15349 ;
  assign n15351 = x47 & ~n15350 ;
  assign n15352 = ( n15349 & ~n15350 ) | ( n15349 & n15351 ) | ( ~n15350 & n15351 ) ;
  assign n15353 = ( n15340 & ~n15341 ) | ( n15340 & n15352 ) | ( ~n15341 & n15352 ) ;
  assign n15354 = ( n15339 & ~n15341 ) | ( n15339 & n15353 ) | ( ~n15341 & n15353 ) ;
  assign n15355 = n15258 | n15354 ;
  assign n15356 = ( n15339 & n15340 ) | ( n15339 & n15352 ) | ( n15340 & n15352 ) ;
  assign n15357 = n15341 & ~n15356 ;
  assign n15358 = n15355 | n15357 ;
  assign n15359 = ( n15258 & n15354 ) | ( n15258 & n15357 ) | ( n15354 & n15357 ) ;
  assign n15360 = n15358 & ~n15359 ;
  assign n15361 = x92 & n6068 ;
  assign n15362 = x91 & n6063 ;
  assign n15363 = x90 & ~n6062 ;
  assign n15364 = n6398 & n15363 ;
  assign n15365 = n15362 | n15364 ;
  assign n15366 = n15361 | n15365 ;
  assign n15367 = n6071 | n15366 ;
  assign n15368 = ( n2904 & n15366 ) | ( n2904 & n15367 ) | ( n15366 & n15367 ) ;
  assign n15369 = x44 & n15368 ;
  assign n15370 = x44 & ~n15369 ;
  assign n15371 = ( n15368 & ~n15369 ) | ( n15368 & n15370 ) | ( ~n15369 & n15370 ) ;
  assign n15372 = n15360 & ~n15371 ;
  assign n15373 = n15371 | n15372 ;
  assign n15374 = ( ~n15360 & n15372 ) | ( ~n15360 & n15373 ) | ( n15372 & n15373 ) ;
  assign n15375 = n15257 | n15374 ;
  assign n15376 = n15257 & n15374 ;
  assign n15377 = n15375 & ~n15376 ;
  assign n15378 = x95 & n5340 ;
  assign n15379 = x94 & n5335 ;
  assign n15380 = x93 & ~n5334 ;
  assign n15381 = n5580 & n15380 ;
  assign n15382 = n15379 | n15381 ;
  assign n15383 = n15378 | n15382 ;
  assign n15384 = n5343 | n15383 ;
  assign n15385 = ( n3479 & n15383 ) | ( n3479 & n15384 ) | ( n15383 & n15384 ) ;
  assign n15386 = x41 & n15385 ;
  assign n15387 = x41 & ~n15386 ;
  assign n15388 = ( n15385 & ~n15386 ) | ( n15385 & n15387 ) | ( ~n15386 & n15387 ) ;
  assign n15389 = n15377 | n15388 ;
  assign n15390 = n15377 & n15388 ;
  assign n15391 = n15389 & ~n15390 ;
  assign n15392 = n14987 | n15122 ;
  assign n15393 = ( n14988 & ~n15125 ) | ( n14988 & n15392 ) | ( ~n15125 & n15392 ) ;
  assign n15394 = n15391 & n15393 ;
  assign n15395 = n15391 | n15393 ;
  assign n15396 = ~n15394 & n15395 ;
  assign n15397 = x98 & n4572 ;
  assign n15398 = x97 & n4567 ;
  assign n15399 = x96 & ~n4566 ;
  assign n15400 = n4828 & n15399 ;
  assign n15401 = n15398 | n15400 ;
  assign n15402 = n15397 | n15401 ;
  assign n15403 = n4575 | n15402 ;
  assign n15404 = ( n4105 & n15402 ) | ( n4105 & n15403 ) | ( n15402 & n15403 ) ;
  assign n15405 = x38 & n15404 ;
  assign n15406 = x38 & ~n15405 ;
  assign n15407 = ( n15404 & ~n15405 ) | ( n15404 & n15406 ) | ( ~n15405 & n15406 ) ;
  assign n15408 = n15396 & n15407 ;
  assign n15409 = n15396 | n15407 ;
  assign n15410 = ~n15408 & n15409 ;
  assign n15411 = n15126 | n15410 ;
  assign n15412 = n15256 | n15411 ;
  assign n15413 = ( n15126 & n15256 ) | ( n15126 & n15410 ) | ( n15256 & n15410 ) ;
  assign n15414 = n15412 & ~n15413 ;
  assign n15415 = x101 & n3913 ;
  assign n15416 = x100 & n3908 ;
  assign n15417 = x99 & ~n3907 ;
  assign n15418 = n4152 & n15417 ;
  assign n15419 = n15416 | n15418 ;
  assign n15420 = n15415 | n15419 ;
  assign n15421 = n3916 | n15420 ;
  assign n15422 = ( n4783 & n15420 ) | ( n4783 & n15421 ) | ( n15420 & n15421 ) ;
  assign n15423 = x35 & n15422 ;
  assign n15424 = x35 & ~n15423 ;
  assign n15425 = ( n15422 & ~n15423 ) | ( n15422 & n15424 ) | ( ~n15423 & n15424 ) ;
  assign n15426 = n15414 & ~n15425 ;
  assign n15427 = n15425 | n15426 ;
  assign n15428 = ( ~n15414 & n15426 ) | ( ~n15414 & n15427 ) | ( n15426 & n15427 ) ;
  assign n15429 = x104 & n3314 ;
  assign n15430 = x103 & n3309 ;
  assign n15431 = x102 & ~n3308 ;
  assign n15432 = n3570 & n15431 ;
  assign n15433 = n15430 | n15432 ;
  assign n15434 = n15429 | n15433 ;
  assign n15435 = n3317 | n15434 ;
  assign n15436 = ( n5295 & n15434 ) | ( n5295 & n15435 ) | ( n15434 & n15435 ) ;
  assign n15437 = x32 & n15436 ;
  assign n15438 = x32 & ~n15437 ;
  assign n15439 = ( n15436 & ~n15437 ) | ( n15436 & n15438 ) | ( ~n15437 & n15438 ) ;
  assign n15440 = n15144 | n15148 ;
  assign n15441 = ( n15428 & n15439 ) | ( n15428 & ~n15440 ) | ( n15439 & ~n15440 ) ;
  assign n15442 = ( ~n15439 & n15440 ) | ( ~n15439 & n15441 ) | ( n15440 & n15441 ) ;
  assign n15443 = ( ~n15428 & n15441 ) | ( ~n15428 & n15442 ) | ( n15441 & n15442 ) ;
  assign n15444 = x107 & n2775 ;
  assign n15445 = x106 & n2770 ;
  assign n15446 = x105 & ~n2769 ;
  assign n15447 = n2978 & n15446 ;
  assign n15448 = n15445 | n15447 ;
  assign n15449 = n15444 | n15448 ;
  assign n15450 = n2778 | n15449 ;
  assign n15451 = ( n6328 & n15449 ) | ( n6328 & n15450 ) | ( n15449 & n15450 ) ;
  assign n15452 = x29 & n15451 ;
  assign n15453 = x29 & ~n15452 ;
  assign n15454 = ( n15451 & ~n15452 ) | ( n15451 & n15453 ) | ( ~n15452 & n15453 ) ;
  assign n15455 = n15163 | n15165 ;
  assign n15456 = ( n15443 & n15454 ) | ( n15443 & ~n15455 ) | ( n15454 & ~n15455 ) ;
  assign n15457 = ( ~n15454 & n15455 ) | ( ~n15454 & n15456 ) | ( n15455 & n15456 ) ;
  assign n15458 = ( ~n15443 & n15456 ) | ( ~n15443 & n15457 ) | ( n15456 & n15457 ) ;
  assign n15459 = x110 & n2280 ;
  assign n15460 = x109 & n2275 ;
  assign n15461 = x108 & ~n2274 ;
  assign n15462 = n2481 & n15461 ;
  assign n15463 = n15460 | n15462 ;
  assign n15464 = n15459 | n15463 ;
  assign n15465 = n2283 | n15464 ;
  assign n15466 = ( n7189 & n15464 ) | ( n7189 & n15465 ) | ( n15464 & n15465 ) ;
  assign n15467 = x26 & n15466 ;
  assign n15468 = x26 & ~n15467 ;
  assign n15469 = ( n15466 & ~n15467 ) | ( n15466 & n15468 ) | ( ~n15467 & n15468 ) ;
  assign n15470 = n14964 | n15168 ;
  assign n15471 = ( n15458 & n15469 ) | ( n15458 & ~n15470 ) | ( n15469 & ~n15470 ) ;
  assign n15472 = ( ~n15469 & n15470 ) | ( ~n15469 & n15471 ) | ( n15470 & n15471 ) ;
  assign n15473 = ( ~n15458 & n15471 ) | ( ~n15458 & n15472 ) | ( n15471 & n15472 ) ;
  assign n15474 = ( n15254 & ~n15255 ) | ( n15254 & n15473 ) | ( ~n15255 & n15473 ) ;
  assign n15475 = ( n15255 & ~n15473 ) | ( n15255 & n15474 ) | ( ~n15473 & n15474 ) ;
  assign n15476 = ( ~n15254 & n15474 ) | ( ~n15254 & n15475 ) | ( n15474 & n15475 ) ;
  assign n15477 = ( n15173 & n15174 ) | ( n15173 & n15185 ) | ( n15174 & n15185 ) ;
  assign n15478 = x116 & n1421 ;
  assign n15479 = x115 & n1416 ;
  assign n15480 = x114 & ~n1415 ;
  assign n15481 = n1584 & n15480 ;
  assign n15482 = n15479 | n15481 ;
  assign n15483 = n15478 | n15482 ;
  assign n15484 = n1424 | n15483 ;
  assign n15485 = ( n8778 & n15483 ) | ( n8778 & n15484 ) | ( n15483 & n15484 ) ;
  assign n15486 = x20 & n15485 ;
  assign n15487 = x20 & ~n15486 ;
  assign n15488 = ( n15485 & ~n15486 ) | ( n15485 & n15487 ) | ( ~n15486 & n15487 ) ;
  assign n15489 = ( n15476 & n15477 ) | ( n15476 & ~n15488 ) | ( n15477 & ~n15488 ) ;
  assign n15490 = ( ~n15477 & n15488 ) | ( ~n15477 & n15489 ) | ( n15488 & n15489 ) ;
  assign n15491 = ( ~n15476 & n15489 ) | ( ~n15476 & n15490 ) | ( n15489 & n15490 ) ;
  assign n15492 = x122 & n771 ;
  assign n15493 = x121 & n766 ;
  assign n15494 = x120 & ~n765 ;
  assign n15495 = n905 & n15494 ;
  assign n15496 = n15493 | n15495 ;
  assign n15497 = n15492 | n15496 ;
  assign n15498 = n774 | n15497 ;
  assign n15499 = ( n11188 & n15497 ) | ( n11188 & n15498 ) | ( n15497 & n15498 ) ;
  assign n15500 = x14 & n15499 ;
  assign n15501 = x14 & ~n15500 ;
  assign n15502 = ( n15499 & ~n15500 ) | ( n15499 & n15501 ) | ( ~n15500 & n15501 ) ;
  assign n15503 = n15204 | n15502 ;
  assign n15504 = n15207 | n15503 ;
  assign n15505 = ( n15204 & n15207 ) | ( n15204 & n15502 ) | ( n15207 & n15502 ) ;
  assign n15506 = n15504 & ~n15505 ;
  assign n15507 = x119 & n1071 ;
  assign n15508 = x118 & n1066 ;
  assign n15509 = x117 & ~n1065 ;
  assign n15510 = n1189 & n15509 ;
  assign n15511 = n15508 | n15510 ;
  assign n15512 = n15507 | n15511 ;
  assign n15513 = n1074 | n15512 ;
  assign n15514 = ( n9789 & n15512 ) | ( n9789 & n15513 ) | ( n15512 & n15513 ) ;
  assign n15515 = x17 & n15514 ;
  assign n15516 = x17 & ~n15515 ;
  assign n15517 = ( n15514 & ~n15515 ) | ( n15514 & n15516 ) | ( ~n15515 & n15516 ) ;
  assign n15518 = ( n14936 & n14937 ) | ( n14936 & n15188 ) | ( n14937 & n15188 ) ;
  assign n15519 = n15517 | n15518 ;
  assign n15520 = n15517 & n15518 ;
  assign n15521 = n15519 & ~n15520 ;
  assign n15522 = ( n15491 & n15506 ) | ( n15491 & ~n15521 ) | ( n15506 & ~n15521 ) ;
  assign n15523 = ( ~n15506 & n15521 ) | ( ~n15506 & n15522 ) | ( n15521 & n15522 ) ;
  assign n15524 = ( ~n15491 & n15522 ) | ( ~n15491 & n15523 ) | ( n15522 & n15523 ) ;
  assign n15525 = ( n15212 & n15213 ) | ( n15212 & n15224 ) | ( n15213 & n15224 ) ;
  assign n15526 = x127 & n332 ;
  assign n15527 = x126 & ~n331 ;
  assign n15528 = n396 & n15527 ;
  assign n15529 = n15526 | n15528 ;
  assign n15530 = n340 | n15529 ;
  assign n15531 = ( n13461 & n15529 ) | ( n13461 & n15530 ) | ( n15529 & n15530 ) ;
  assign n15532 = x8 & n15531 ;
  assign n15533 = x8 & ~n15532 ;
  assign n15534 = ( n15531 & ~n15532 ) | ( n15531 & n15533 ) | ( ~n15532 & n15533 ) ;
  assign n15535 = n15525 & n15534 ;
  assign n15536 = n15525 | n15534 ;
  assign n15537 = ~n15535 & n15536 ;
  assign n15538 = x125 & n528 ;
  assign n15539 = x124 & n523 ;
  assign n15540 = x123 & ~n522 ;
  assign n15541 = n635 & n15540 ;
  assign n15542 = n15539 | n15541 ;
  assign n15543 = n15538 | n15542 ;
  assign n15544 = n531 | n15543 ;
  assign n15545 = ( n12310 & n15543 ) | ( n12310 & n15544 ) | ( n15543 & n15544 ) ;
  assign n15546 = x11 & n15545 ;
  assign n15547 = x11 & ~n15546 ;
  assign n15548 = ( n15545 & ~n15546 ) | ( n15545 & n15547 ) | ( ~n15546 & n15547 ) ;
  assign n15549 = ( n14918 & n14919 ) | ( n14918 & n15209 ) | ( n14919 & n15209 ) ;
  assign n15550 = n15548 | n15549 ;
  assign n15551 = n15548 & n15549 ;
  assign n15552 = n15550 & ~n15551 ;
  assign n15553 = ( n15524 & n15537 ) | ( n15524 & ~n15552 ) | ( n15537 & ~n15552 ) ;
  assign n15554 = ( ~n15537 & n15552 ) | ( ~n15537 & n15553 ) | ( n15552 & n15553 ) ;
  assign n15555 = ( ~n15524 & n15553 ) | ( ~n15524 & n15554 ) | ( n15553 & n15554 ) ;
  assign n15556 = ( n14900 & n14902 ) | ( n14900 & n15227 ) | ( n14902 & n15227 ) ;
  assign n15557 = n15555 & n15556 ;
  assign n15558 = n15556 & ~n15557 ;
  assign n15559 = ( n15555 & ~n15557 ) | ( n15555 & n15558 ) | ( ~n15557 & n15558 ) ;
  assign n15560 = n15233 | n15242 ;
  assign n15561 = n15559 | n15560 ;
  assign n15562 = n15559 & n15560 ;
  assign n15563 = n15561 & ~n15562 ;
  assign n15564 = ( n15524 & n15548 ) | ( n15524 & n15549 ) | ( n15548 & n15549 ) ;
  assign n15565 = x127 & ~n331 ;
  assign n15566 = n396 & n15565 ;
  assign n15567 = ( x127 & n340 ) | ( x127 & n15566 ) | ( n340 & n15566 ) ;
  assign n15568 = ( x126 & n15566 ) | ( x126 & n15567 ) | ( n15566 & n15567 ) ;
  assign n15569 = ( n12685 & n15567 ) | ( n12685 & n15568 ) | ( n15567 & n15568 ) ;
  assign n15570 = x8 & n15569 ;
  assign n15571 = x8 & ~n15570 ;
  assign n15572 = ( n15569 & ~n15570 ) | ( n15569 & n15571 ) | ( ~n15570 & n15571 ) ;
  assign n15573 = n15564 & n15572 ;
  assign n15574 = n15564 & ~n15573 ;
  assign n15575 = n15506 & ~n15524 ;
  assign n15576 = n15505 | n15575 ;
  assign n15577 = x126 & n528 ;
  assign n15578 = x125 & n523 ;
  assign n15579 = x124 & ~n522 ;
  assign n15580 = n635 & n15579 ;
  assign n15581 = n15578 | n15580 ;
  assign n15582 = n15577 | n15581 ;
  assign n15583 = n531 | n15582 ;
  assign n15584 = ( n12687 & n15582 ) | ( n12687 & n15583 ) | ( n15582 & n15583 ) ;
  assign n15585 = x11 & n15584 ;
  assign n15586 = x11 & ~n15585 ;
  assign n15587 = ( n15584 & ~n15585 ) | ( n15584 & n15586 ) | ( ~n15585 & n15586 ) ;
  assign n15588 = n15576 & n15587 ;
  assign n15589 = n15576 & ~n15588 ;
  assign n15590 = ~n15576 & n15587 ;
  assign n15591 = x114 & n1817 ;
  assign n15592 = x113 & n1812 ;
  assign n15593 = x112 & ~n1811 ;
  assign n15594 = n1977 & n15593 ;
  assign n15595 = n15592 | n15594 ;
  assign n15596 = n15591 | n15595 ;
  assign n15597 = n1820 | n15596 ;
  assign n15598 = ( n8437 & n15596 ) | ( n8437 & n15597 ) | ( n15596 & n15597 ) ;
  assign n15599 = x23 & n15598 ;
  assign n15600 = x23 & ~n15599 ;
  assign n15601 = ( n15598 & ~n15599 ) | ( n15598 & n15600 ) | ( ~n15599 & n15600 ) ;
  assign n15602 = ( n15458 & n15469 ) | ( n15458 & n15470 ) | ( n15469 & n15470 ) ;
  assign n15603 = n15601 | n15602 ;
  assign n15604 = n15601 & n15602 ;
  assign n15605 = n15603 & ~n15604 ;
  assign n15606 = x111 & n2280 ;
  assign n15607 = x110 & n2275 ;
  assign n15608 = x109 & ~n2274 ;
  assign n15609 = n2481 & n15608 ;
  assign n15610 = n15607 | n15609 ;
  assign n15611 = n15606 | n15610 ;
  assign n15612 = n2283 | n15611 ;
  assign n15613 = ( n7492 & n15611 ) | ( n7492 & n15612 ) | ( n15611 & n15612 ) ;
  assign n15614 = x26 & n15613 ;
  assign n15615 = x26 & ~n15614 ;
  assign n15616 = ( n15613 & ~n15614 ) | ( n15613 & n15615 ) | ( ~n15614 & n15615 ) ;
  assign n15617 = n15454 & n15455 ;
  assign n15618 = n15616 & n15617 ;
  assign n15619 = n15616 & ~n15618 ;
  assign n15620 = n15443 & ~n15457 ;
  assign n15621 = ( n15443 & ~n15456 ) | ( n15443 & n15620 ) | ( ~n15456 & n15620 ) ;
  assign n15622 = n15619 & ~n15621 ;
  assign n15623 = ( ~n15616 & n15617 ) | ( ~n15616 & n15621 ) | ( n15617 & n15621 ) ;
  assign n15624 = n15622 | n15623 ;
  assign n15625 = ( n15428 & n15439 ) | ( n15428 & n15440 ) | ( n15439 & n15440 ) ;
  assign n15626 = x108 & n2775 ;
  assign n15627 = x107 & n2770 ;
  assign n15628 = x106 & ~n2769 ;
  assign n15629 = n2978 & n15628 ;
  assign n15630 = n15627 | n15629 ;
  assign n15631 = n15626 | n15630 ;
  assign n15632 = n2778 | n15631 ;
  assign n15633 = ( n6358 & n15631 ) | ( n6358 & n15632 ) | ( n15631 & n15632 ) ;
  assign n15634 = x29 & n15633 ;
  assign n15635 = x29 & ~n15634 ;
  assign n15636 = ( n15633 & ~n15634 ) | ( n15633 & n15635 ) | ( ~n15634 & n15635 ) ;
  assign n15637 = n15625 & n15636 ;
  assign n15638 = n15625 & ~n15637 ;
  assign n15639 = ~n15625 & n15636 ;
  assign n15640 = n15638 | n15639 ;
  assign n15641 = x102 & n3913 ;
  assign n15642 = x101 & n3908 ;
  assign n15643 = x100 & ~n3907 ;
  assign n15644 = n4152 & n15643 ;
  assign n15645 = n15642 | n15644 ;
  assign n15646 = n15641 | n15645 ;
  assign n15647 = n3916 | n15646 ;
  assign n15648 = ( n5025 & n15646 ) | ( n5025 & n15647 ) | ( n15646 & n15647 ) ;
  assign n15649 = x35 & n15648 ;
  assign n15650 = x35 & ~n15649 ;
  assign n15651 = ( n15648 & ~n15649 ) | ( n15648 & n15650 ) | ( ~n15649 & n15650 ) ;
  assign n15652 = x105 & n3314 ;
  assign n15653 = x104 & n3309 ;
  assign n15654 = x103 & ~n3308 ;
  assign n15655 = n3570 & n15654 ;
  assign n15656 = n15653 | n15655 ;
  assign n15657 = n15652 | n15656 ;
  assign n15658 = n3317 | n15657 ;
  assign n15659 = ( n5788 & n15657 ) | ( n5788 & n15658 ) | ( n15657 & n15658 ) ;
  assign n15660 = x32 & n15659 ;
  assign n15661 = x32 & ~n15660 ;
  assign n15662 = ( n15659 & ~n15660 ) | ( n15659 & n15661 ) | ( ~n15660 & n15661 ) ;
  assign n15663 = ( n15412 & n15413 ) | ( n15412 & n15425 ) | ( n15413 & n15425 ) ;
  assign n15664 = n15662 | n15663 ;
  assign n15665 = n15662 & n15663 ;
  assign n15666 = n15664 & ~n15665 ;
  assign n15667 = n15394 | n15408 ;
  assign n15668 = n15376 | n15390 ;
  assign n15669 = ( n15358 & n15359 ) | ( n15358 & n15371 ) | ( n15359 & n15371 ) ;
  assign n15670 = x93 & n6068 ;
  assign n15671 = x92 & n6063 ;
  assign n15672 = x91 & ~n6062 ;
  assign n15673 = n6398 & n15672 ;
  assign n15674 = n15671 | n15673 ;
  assign n15675 = n15670 | n15674 ;
  assign n15676 = n6071 | n15675 ;
  assign n15677 = ( n2931 & n15675 ) | ( n2931 & n15676 ) | ( n15675 & n15676 ) ;
  assign n15678 = x44 & n15677 ;
  assign n15679 = x44 & ~n15678 ;
  assign n15680 = ( n15677 & ~n15678 ) | ( n15677 & n15679 ) | ( ~n15678 & n15679 ) ;
  assign n15681 = x90 & n6937 ;
  assign n15682 = x89 & n6932 ;
  assign n15683 = x88 & ~n6931 ;
  assign n15684 = n7216 & n15683 ;
  assign n15685 = n15682 | n15684 ;
  assign n15686 = n15681 | n15685 ;
  assign n15687 = n6940 | n15686 ;
  assign n15688 = ( n2410 & n15686 ) | ( n2410 & n15687 ) | ( n15686 & n15687 ) ;
  assign n15689 = x47 & n15688 ;
  assign n15690 = x47 & ~n15689 ;
  assign n15691 = ( n15688 & ~n15689 ) | ( n15688 & n15690 ) | ( ~n15689 & n15690 ) ;
  assign n15692 = ( n15269 & n15270 ) | ( n15269 & n15336 ) | ( n15270 & n15336 ) ;
  assign n15693 = ( n15281 & n15282 ) | ( n15281 & n15333 ) | ( n15282 & n15333 ) ;
  assign n15694 = ( n15293 & n15294 ) | ( n15293 & n15330 ) | ( n15294 & n15330 ) ;
  assign n15695 = x81 & n9853 ;
  assign n15696 = x80 & n9848 ;
  assign n15697 = x79 & ~n9847 ;
  assign n15698 = n10165 & n15697 ;
  assign n15699 = n15696 | n15698 ;
  assign n15700 = n15695 | n15699 ;
  assign n15701 = n9856 | n15700 ;
  assign n15702 = ( n1256 & n15700 ) | ( n1256 & n15701 ) | ( n15700 & n15701 ) ;
  assign n15703 = x56 & n15702 ;
  assign n15704 = x56 & ~n15703 ;
  assign n15705 = ( n15702 & ~n15703 ) | ( n15702 & n15704 ) | ( ~n15703 & n15704 ) ;
  assign n15706 = x78 & n10876 ;
  assign n15707 = x77 & n10871 ;
  assign n15708 = x76 & ~n10870 ;
  assign n15709 = n11305 & n15708 ;
  assign n15710 = n15707 | n15709 ;
  assign n15711 = n15706 | n15710 ;
  assign n15712 = n10879 | n15711 ;
  assign n15713 = ( n868 & n15711 ) | ( n868 & n15712 ) | ( n15711 & n15712 ) ;
  assign n15714 = x59 & n15713 ;
  assign n15715 = x59 & ~n15714 ;
  assign n15716 = ( n15713 & ~n15714 ) | ( n15713 & n15715 ) | ( ~n15714 & n15715 ) ;
  assign n15717 = x72 & n12808 ;
  assign n15718 = x63 & x71 ;
  assign n15719 = ~n12808 & n15718 ;
  assign n15720 = n15717 | n15719 ;
  assign n15721 = ~n15299 & n15720 ;
  assign n15722 = n15299 & ~n15720 ;
  assign n15723 = n15301 | n15722 ;
  assign n15724 = ( n15300 & ~n15313 ) | ( n15300 & n15723 ) | ( ~n15313 & n15723 ) ;
  assign n15725 = n15721 | n15724 ;
  assign n15726 = ~n15722 & n15725 ;
  assign n15727 = ~n15721 & n15726 ;
  assign n15728 = ( ~n15300 & n15314 ) | ( ~n15300 & n15725 ) | ( n15314 & n15725 ) ;
  assign n15729 = n15727 | n15728 ;
  assign n15730 = x75 & n11984 ;
  assign n15731 = x74 & n11979 ;
  assign n15732 = x73 & ~n11978 ;
  assign n15733 = n12430 & n15732 ;
  assign n15734 = n15731 | n15733 ;
  assign n15735 = n15730 | n15734 ;
  assign n15736 = n11987 | n15735 ;
  assign n15737 = ( n609 & n15735 ) | ( n609 & n15736 ) | ( n15735 & n15736 ) ;
  assign n15738 = x62 & n15737 ;
  assign n15739 = x62 & ~n15738 ;
  assign n15740 = ( n15737 & ~n15738 ) | ( n15737 & n15739 ) | ( ~n15738 & n15739 ) ;
  assign n15741 = ( n15716 & n15729 ) | ( n15716 & ~n15740 ) | ( n15729 & ~n15740 ) ;
  assign n15742 = ( ~n15729 & n15740 ) | ( ~n15729 & n15741 ) | ( n15740 & n15741 ) ;
  assign n15743 = ( ~n15716 & n15741 ) | ( ~n15716 & n15742 ) | ( n15741 & n15742 ) ;
  assign n15744 = ( ~n15328 & n15705 ) | ( ~n15328 & n15743 ) | ( n15705 & n15743 ) ;
  assign n15745 = ( n15328 & ~n15743 ) | ( n15328 & n15744 ) | ( ~n15743 & n15744 ) ;
  assign n15746 = ( ~n15705 & n15744 ) | ( ~n15705 & n15745 ) | ( n15744 & n15745 ) ;
  assign n15747 = n15694 | n15746 ;
  assign n15748 = n15694 & n15746 ;
  assign n15749 = n15747 & ~n15748 ;
  assign n15750 = x84 & n8834 ;
  assign n15751 = x83 & n8829 ;
  assign n15752 = x82 & ~n8828 ;
  assign n15753 = n9159 & n15752 ;
  assign n15754 = n15751 | n15753 ;
  assign n15755 = n15750 | n15754 ;
  assign n15756 = n8837 | n15755 ;
  assign n15757 = ( n1537 & n15755 ) | ( n1537 & n15756 ) | ( n15755 & n15756 ) ;
  assign n15758 = x53 & n15757 ;
  assign n15759 = x53 & ~n15758 ;
  assign n15760 = ( n15757 & ~n15758 ) | ( n15757 & n15759 ) | ( ~n15758 & n15759 ) ;
  assign n15761 = n15749 | n15760 ;
  assign n15762 = n15749 & n15760 ;
  assign n15763 = n15761 & ~n15762 ;
  assign n15764 = x87 & n7812 ;
  assign n15765 = x86 & n7807 ;
  assign n15766 = x85 & ~n7806 ;
  assign n15767 = n8136 & n15766 ;
  assign n15768 = n15765 | n15767 ;
  assign n15769 = n15764 | n15768 ;
  assign n15770 = n7815 | n15769 ;
  assign n15771 = ( n2067 & n15769 ) | ( n2067 & n15770 ) | ( n15769 & n15770 ) ;
  assign n15772 = x50 & n15771 ;
  assign n15773 = x50 & ~n15772 ;
  assign n15774 = ( n15771 & ~n15772 ) | ( n15771 & n15773 ) | ( ~n15772 & n15773 ) ;
  assign n15775 = ( n15693 & ~n15763 ) | ( n15693 & n15774 ) | ( ~n15763 & n15774 ) ;
  assign n15776 = ( n15763 & ~n15774 ) | ( n15763 & n15775 ) | ( ~n15774 & n15775 ) ;
  assign n15777 = ( ~n15693 & n15775 ) | ( ~n15693 & n15776 ) | ( n15775 & n15776 ) ;
  assign n15778 = ( n15691 & n15692 ) | ( n15691 & ~n15777 ) | ( n15692 & ~n15777 ) ;
  assign n15779 = ( ~n15692 & n15777 ) | ( ~n15692 & n15778 ) | ( n15777 & n15778 ) ;
  assign n15780 = ( ~n15691 & n15778 ) | ( ~n15691 & n15779 ) | ( n15778 & n15779 ) ;
  assign n15781 = ( n15356 & n15680 ) | ( n15356 & ~n15780 ) | ( n15680 & ~n15780 ) ;
  assign n15782 = ( ~n15356 & n15780 ) | ( ~n15356 & n15781 ) | ( n15780 & n15781 ) ;
  assign n15783 = ( ~n15680 & n15781 ) | ( ~n15680 & n15782 ) | ( n15781 & n15782 ) ;
  assign n15784 = n15669 | n15783 ;
  assign n15785 = n15669 & n15783 ;
  assign n15786 = n15784 & ~n15785 ;
  assign n15787 = x96 & n5340 ;
  assign n15788 = x95 & n5335 ;
  assign n15789 = x94 & ~n5334 ;
  assign n15790 = n5580 & n15789 ;
  assign n15791 = n15788 | n15790 ;
  assign n15792 = n15787 | n15791 ;
  assign n15793 = n5343 | n15792 ;
  assign n15794 = ( n3509 & n15792 ) | ( n3509 & n15793 ) | ( n15792 & n15793 ) ;
  assign n15795 = x41 & n15794 ;
  assign n15796 = x41 & ~n15795 ;
  assign n15797 = ( n15794 & ~n15795 ) | ( n15794 & n15796 ) | ( ~n15795 & n15796 ) ;
  assign n15798 = n15786 | n15797 ;
  assign n15799 = n15786 & n15797 ;
  assign n15800 = n15798 & ~n15799 ;
  assign n15801 = x99 & n4572 ;
  assign n15802 = x98 & n4567 ;
  assign n15803 = x97 & ~n4566 ;
  assign n15804 = n4828 & n15803 ;
  assign n15805 = n15802 | n15804 ;
  assign n15806 = n15801 | n15805 ;
  assign n15807 = n4575 | n15806 ;
  assign n15808 = ( n4325 & n15806 ) | ( n4325 & n15807 ) | ( n15806 & n15807 ) ;
  assign n15809 = x38 & n15808 ;
  assign n15810 = x38 & ~n15809 ;
  assign n15811 = ( n15808 & ~n15809 ) | ( n15808 & n15810 ) | ( ~n15809 & n15810 ) ;
  assign n15812 = ( n15668 & n15800 ) | ( n15668 & n15811 ) | ( n15800 & n15811 ) ;
  assign n15813 = ( n15800 & n15811 ) | ( n15800 & ~n15812 ) | ( n15811 & ~n15812 ) ;
  assign n15814 = ( n15668 & ~n15812 ) | ( n15668 & n15813 ) | ( ~n15812 & n15813 ) ;
  assign n15815 = n15667 | n15814 ;
  assign n15816 = n15667 & n15814 ;
  assign n15817 = n15815 & ~n15816 ;
  assign n15818 = ( n15651 & n15666 ) | ( n15651 & ~n15817 ) | ( n15666 & ~n15817 ) ;
  assign n15819 = ( ~n15666 & n15817 ) | ( ~n15666 & n15818 ) | ( n15817 & n15818 ) ;
  assign n15820 = ( ~n15651 & n15818 ) | ( ~n15651 & n15819 ) | ( n15818 & n15819 ) ;
  assign n15821 = n15640 & n15820 ;
  assign n15822 = n15640 | n15820 ;
  assign n15823 = ~n15821 & n15822 ;
  assign n15824 = n15624 & n15823 ;
  assign n15825 = n15624 | n15823 ;
  assign n15826 = ~n15824 & n15825 ;
  assign n15827 = n15605 | n15826 ;
  assign n15828 = n15605 & n15826 ;
  assign n15829 = n15827 & ~n15828 ;
  assign n15830 = x117 & n1421 ;
  assign n15831 = x116 & n1416 ;
  assign n15832 = x115 & ~n1415 ;
  assign n15833 = n1584 & n15832 ;
  assign n15834 = n15831 | n15833 ;
  assign n15835 = n15830 | n15834 ;
  assign n15836 = n1424 | n15835 ;
  assign n15837 = ( n9118 & n15835 ) | ( n9118 & n15836 ) | ( n15835 & n15836 ) ;
  assign n15838 = x20 & n15837 ;
  assign n15839 = x20 & ~n15838 ;
  assign n15840 = ( n15837 & ~n15838 ) | ( n15837 & n15839 ) | ( ~n15838 & n15839 ) ;
  assign n15841 = ( n14802 & n14806 ) | ( n14802 & n14949 ) | ( n14806 & n14949 ) ;
  assign n15842 = n15254 & n15841 ;
  assign n15843 = ( n15254 & n15255 ) | ( n15254 & n15842 ) | ( n15255 & n15842 ) ;
  assign n15844 = n15840 & n15843 ;
  assign n15845 = n15840 & ~n15844 ;
  assign n15846 = n15254 & ~n15255 ;
  assign n15847 = ( n15473 & ~n15474 ) | ( n15473 & n15846 ) | ( ~n15474 & n15846 ) ;
  assign n15848 = n15845 & ~n15847 ;
  assign n15849 = ( ~n15840 & n15843 ) | ( ~n15840 & n15847 ) | ( n15843 & n15847 ) ;
  assign n15850 = n15848 | n15849 ;
  assign n15851 = n15829 & n15850 ;
  assign n15852 = n15829 | n15850 ;
  assign n15853 = ~n15851 & n15852 ;
  assign n15854 = ( n15476 & n15477 ) | ( n15476 & n15488 ) | ( n15477 & n15488 ) ;
  assign n15855 = x120 & n1071 ;
  assign n15856 = x119 & n1066 ;
  assign n15857 = x118 & ~n1065 ;
  assign n15858 = n1189 & n15857 ;
  assign n15859 = n15856 | n15858 ;
  assign n15860 = n15855 | n15859 ;
  assign n15861 = n1074 | n15860 ;
  assign n15862 = ( n10460 & n15860 ) | ( n10460 & n15861 ) | ( n15860 & n15861 ) ;
  assign n15863 = x17 & n15862 ;
  assign n15864 = x17 & ~n15863 ;
  assign n15865 = ( n15862 & ~n15863 ) | ( n15862 & n15864 ) | ( ~n15863 & n15864 ) ;
  assign n15866 = ( n15853 & n15854 ) | ( n15853 & ~n15865 ) | ( n15854 & ~n15865 ) ;
  assign n15867 = ( ~n15854 & n15865 ) | ( ~n15854 & n15866 ) | ( n15865 & n15866 ) ;
  assign n15868 = ( ~n15853 & n15866 ) | ( ~n15853 & n15867 ) | ( n15866 & n15867 ) ;
  assign n15869 = x123 & n771 ;
  assign n15870 = x122 & n766 ;
  assign n15871 = x121 & ~n765 ;
  assign n15872 = n905 & n15871 ;
  assign n15873 = n15870 | n15872 ;
  assign n15874 = n15869 | n15873 ;
  assign n15875 = n774 | n15874 ;
  assign n15876 = ( n11219 & n15874 ) | ( n11219 & n15875 ) | ( n15874 & n15875 ) ;
  assign n15877 = x14 & n15876 ;
  assign n15878 = x14 & ~n15877 ;
  assign n15879 = ( n15876 & ~n15877 ) | ( n15876 & n15878 ) | ( ~n15877 & n15878 ) ;
  assign n15880 = ( n15491 & n15517 ) | ( n15491 & n15518 ) | ( n15517 & n15518 ) ;
  assign n15881 = ( n15868 & n15879 ) | ( n15868 & ~n15880 ) | ( n15879 & ~n15880 ) ;
  assign n15882 = ( ~n15879 & n15880 ) | ( ~n15879 & n15881 ) | ( n15880 & n15881 ) ;
  assign n15883 = ( ~n15868 & n15881 ) | ( ~n15868 & n15882 ) | ( n15881 & n15882 ) ;
  assign n15884 = n15590 | n15883 ;
  assign n15885 = n15589 | n15884 ;
  assign n15886 = ( n15589 & n15590 ) | ( n15589 & n15883 ) | ( n15590 & n15883 ) ;
  assign n15887 = n15885 & ~n15886 ;
  assign n15888 = ~n15564 & n15572 ;
  assign n15889 = n15887 | n15888 ;
  assign n15890 = n15574 | n15889 ;
  assign n15891 = ( n15574 & n15887 ) | ( n15574 & n15888 ) | ( n15887 & n15888 ) ;
  assign n15892 = n15890 & ~n15891 ;
  assign n15893 = n15557 | n15562 ;
  assign n15894 = ( n15525 & n15534 ) | ( n15525 & ~n15555 ) | ( n15534 & ~n15555 ) ;
  assign n15895 = ( n15892 & ~n15893 ) | ( n15892 & n15894 ) | ( ~n15893 & n15894 ) ;
  assign n15896 = ( n15893 & ~n15894 ) | ( n15893 & n15895 ) | ( ~n15894 & n15895 ) ;
  assign n15897 = ( ~n15892 & n15895 ) | ( ~n15892 & n15896 ) | ( n15895 & n15896 ) ;
  assign n15898 = n15573 | n15891 ;
  assign n15899 = x127 & n528 ;
  assign n15900 = x126 & n523 ;
  assign n15901 = x125 & ~n522 ;
  assign n15902 = n635 & n15901 ;
  assign n15903 = n15900 | n15902 ;
  assign n15904 = n15899 | n15903 ;
  assign n15905 = n531 | n15904 ;
  assign n15906 = ( n12720 & n15904 ) | ( n12720 & n15905 ) | ( n15904 & n15905 ) ;
  assign n15907 = x11 & n15906 ;
  assign n15908 = x11 & ~n15907 ;
  assign n15909 = ( n15906 & ~n15907 ) | ( n15906 & n15908 ) | ( ~n15907 & n15908 ) ;
  assign n15910 = n15588 | n15886 ;
  assign n15911 = x118 & n1421 ;
  assign n15912 = x117 & n1416 ;
  assign n15913 = x116 & ~n1415 ;
  assign n15914 = n1584 & n15913 ;
  assign n15915 = n15912 | n15914 ;
  assign n15916 = n15911 | n15915 ;
  assign n15917 = n1424 | n15916 ;
  assign n15918 = ( n9760 & n15916 ) | ( n9760 & n15917 ) | ( n15916 & n15917 ) ;
  assign n15919 = x20 & n15918 ;
  assign n15920 = x20 & ~n15919 ;
  assign n15921 = ( n15918 & ~n15919 ) | ( n15918 & n15920 ) | ( ~n15919 & n15920 ) ;
  assign n15922 = ( n15840 & n15844 ) | ( n15840 & n15847 ) | ( n15844 & n15847 ) ;
  assign n15923 = n15921 & n15922 ;
  assign n15924 = ( n15851 & n15921 ) | ( n15851 & n15923 ) | ( n15921 & n15923 ) ;
  assign n15925 = n15851 | n15922 ;
  assign n15926 = ~n15921 & n15925 ;
  assign n15927 = ( n15921 & ~n15924 ) | ( n15921 & n15926 ) | ( ~n15924 & n15926 ) ;
  assign n15928 = ( n15616 & n15618 ) | ( n15616 & n15621 ) | ( n15618 & n15621 ) ;
  assign n15929 = x112 & n2280 ;
  assign n15930 = x111 & n2275 ;
  assign n15931 = x110 & ~n2274 ;
  assign n15932 = n2481 & n15931 ;
  assign n15933 = n15930 | n15932 ;
  assign n15934 = n15929 | n15933 ;
  assign n15935 = n2283 | n15934 ;
  assign n15936 = ( n7789 & n15934 ) | ( n7789 & n15935 ) | ( n15934 & n15935 ) ;
  assign n15937 = x26 & n15936 ;
  assign n15938 = x26 & ~n15937 ;
  assign n15939 = ( n15936 & ~n15937 ) | ( n15936 & n15938 ) | ( ~n15937 & n15938 ) ;
  assign n15940 = n15928 | n15939 ;
  assign n15941 = n15824 | n15940 ;
  assign n15942 = ( n15824 & n15928 ) | ( n15824 & n15939 ) | ( n15928 & n15939 ) ;
  assign n15943 = n15941 & ~n15942 ;
  assign n15944 = x109 & n2775 ;
  assign n15945 = x108 & n2770 ;
  assign n15946 = x107 & ~n2769 ;
  assign n15947 = n2978 & n15946 ;
  assign n15948 = n15945 | n15947 ;
  assign n15949 = n15944 | n15948 ;
  assign n15950 = n2778 | n15949 ;
  assign n15951 = ( n6884 & n15949 ) | ( n6884 & n15950 ) | ( n15949 & n15950 ) ;
  assign n15952 = x29 & n15951 ;
  assign n15953 = x29 & ~n15952 ;
  assign n15954 = ( n15951 & ~n15952 ) | ( n15951 & n15953 ) | ( ~n15952 & n15953 ) ;
  assign n15955 = n15637 | n15821 ;
  assign n15956 = ( n15662 & n15663 ) | ( n15662 & ~n15820 ) | ( n15663 & ~n15820 ) ;
  assign n15957 = x106 & n3314 ;
  assign n15958 = x105 & n3309 ;
  assign n15959 = x104 & ~n3308 ;
  assign n15960 = n3570 & n15959 ;
  assign n15961 = n15958 | n15960 ;
  assign n15962 = n15957 | n15961 ;
  assign n15963 = n3317 | n15962 ;
  assign n15964 = ( n5814 & n15962 ) | ( n5814 & n15963 ) | ( n15962 & n15963 ) ;
  assign n15965 = x32 & n15964 ;
  assign n15966 = x32 & ~n15965 ;
  assign n15967 = ( n15964 & ~n15965 ) | ( n15964 & n15966 ) | ( ~n15965 & n15966 ) ;
  assign n15968 = n15956 & n15967 ;
  assign n15969 = n15956 & ~n15968 ;
  assign n15970 = ~n15956 & n15967 ;
  assign n15971 = n15969 | n15970 ;
  assign n15972 = x103 & n3913 ;
  assign n15973 = x102 & n3908 ;
  assign n15974 = x101 & ~n3907 ;
  assign n15975 = n4152 & n15974 ;
  assign n15976 = n15973 | n15975 ;
  assign n15977 = n15972 | n15976 ;
  assign n15978 = n3916 | n15977 ;
  assign n15979 = ( n5264 & n15977 ) | ( n5264 & n15978 ) | ( n15977 & n15978 ) ;
  assign n15980 = x35 & n15979 ;
  assign n15981 = x35 & ~n15980 ;
  assign n15982 = ( n15979 & ~n15980 ) | ( n15979 & n15981 ) | ( ~n15980 & n15981 ) ;
  assign n15983 = x100 & n4572 ;
  assign n15984 = x99 & n4567 ;
  assign n15985 = x98 & ~n4566 ;
  assign n15986 = n4828 & n15985 ;
  assign n15987 = n15984 | n15986 ;
  assign n15988 = n15983 | n15987 ;
  assign n15989 = n4575 | n15988 ;
  assign n15990 = ( n4532 & n15988 ) | ( n4532 & n15989 ) | ( n15988 & n15989 ) ;
  assign n15991 = x38 & n15990 ;
  assign n15992 = x38 & ~n15991 ;
  assign n15993 = ( n15990 & ~n15991 ) | ( n15990 & n15992 ) | ( ~n15991 & n15992 ) ;
  assign n15994 = n15785 | n15799 ;
  assign n15995 = ( n15356 & n15680 ) | ( n15356 & n15780 ) | ( n15680 & n15780 ) ;
  assign n15996 = x91 & n6937 ;
  assign n15997 = x90 & n6932 ;
  assign n15998 = x89 & ~n6931 ;
  assign n15999 = n7216 & n15998 ;
  assign n16000 = n15997 | n15999 ;
  assign n16001 = n15996 | n16000 ;
  assign n16002 = n6940 | n16001 ;
  assign n16003 = ( n2714 & n16001 ) | ( n2714 & n16002 ) | ( n16001 & n16002 ) ;
  assign n16004 = x47 & n16003 ;
  assign n16005 = x47 & ~n16004 ;
  assign n16006 = ( n16003 & ~n16004 ) | ( n16003 & n16005 ) | ( ~n16004 & n16005 ) ;
  assign n16007 = x88 & n7812 ;
  assign n16008 = x87 & n7807 ;
  assign n16009 = x86 & ~n7806 ;
  assign n16010 = n8136 & n16009 ;
  assign n16011 = n16008 | n16010 ;
  assign n16012 = n16007 | n16011 ;
  assign n16013 = n7815 | n16012 ;
  assign n16014 = ( n2095 & n16012 ) | ( n2095 & n16013 ) | ( n16012 & n16013 ) ;
  assign n16015 = x50 & n16014 ;
  assign n16016 = x50 & ~n16015 ;
  assign n16017 = ( n16014 & ~n16015 ) | ( n16014 & n16016 ) | ( ~n16015 & n16016 ) ;
  assign n16018 = x79 & n10876 ;
  assign n16019 = x78 & n10871 ;
  assign n16020 = x77 & ~n10870 ;
  assign n16021 = n11305 & n16020 ;
  assign n16022 = n16019 | n16021 ;
  assign n16023 = n16018 | n16022 ;
  assign n16024 = n10879 | n16023 ;
  assign n16025 = ( n961 & n16023 ) | ( n961 & n16024 ) | ( n16023 & n16024 ) ;
  assign n16026 = x59 & n16025 ;
  assign n16027 = x59 & ~n16026 ;
  assign n16028 = ( n16025 & ~n16026 ) | ( n16025 & n16027 ) | ( ~n16026 & n16027 ) ;
  assign n16029 = x76 & n11984 ;
  assign n16030 = x75 & n11979 ;
  assign n16031 = x74 & ~n11978 ;
  assign n16032 = n12430 & n16031 ;
  assign n16033 = n16030 | n16032 ;
  assign n16034 = n16029 | n16033 ;
  assign n16035 = n11987 | n16034 ;
  assign n16036 = ( n740 & n16034 ) | ( n740 & n16035 ) | ( n16034 & n16035 ) ;
  assign n16037 = x62 & n16036 ;
  assign n16038 = x62 & ~n16037 ;
  assign n16039 = ( n16036 & ~n16037 ) | ( n16036 & n16038 ) | ( ~n16037 & n16038 ) ;
  assign n16040 = x73 & n12808 ;
  assign n16041 = x63 & x72 ;
  assign n16042 = ~n12808 & n16041 ;
  assign n16043 = n16040 | n16042 ;
  assign n16044 = ( x8 & ~n15720 ) | ( x8 & n16043 ) | ( ~n15720 & n16043 ) ;
  assign n16045 = ( ~x8 & n15720 ) | ( ~x8 & n16043 ) | ( n15720 & n16043 ) ;
  assign n16046 = ( ~n16043 & n16044 ) | ( ~n16043 & n16045 ) | ( n16044 & n16045 ) ;
  assign n16047 = ( n15726 & n16039 ) | ( n15726 & ~n16046 ) | ( n16039 & ~n16046 ) ;
  assign n16048 = ( ~n15726 & n16046 ) | ( ~n15726 & n16047 ) | ( n16046 & n16047 ) ;
  assign n16049 = ( ~n16039 & n16047 ) | ( ~n16039 & n16048 ) | ( n16047 & n16048 ) ;
  assign n16050 = n16028 & n16049 ;
  assign n16051 = n16028 | n16049 ;
  assign n16052 = ~n16050 & n16051 ;
  assign n16053 = ( n15716 & n15729 ) | ( n15716 & n15740 ) | ( n15729 & n15740 ) ;
  assign n16054 = n16052 | n16053 ;
  assign n16055 = n16052 & n16053 ;
  assign n16056 = n16054 & ~n16055 ;
  assign n16057 = x82 & n9853 ;
  assign n16058 = x81 & n9848 ;
  assign n16059 = x80 & ~n9847 ;
  assign n16060 = n10165 & n16059 ;
  assign n16061 = n16058 | n16060 ;
  assign n16062 = n16057 | n16061 ;
  assign n16063 = n9856 | n16062 ;
  assign n16064 = ( n1371 & n16062 ) | ( n1371 & n16063 ) | ( n16062 & n16063 ) ;
  assign n16065 = x56 & n16064 ;
  assign n16066 = x56 & ~n16065 ;
  assign n16067 = ( n16064 & ~n16065 ) | ( n16064 & n16066 ) | ( ~n16065 & n16066 ) ;
  assign n16068 = n16056 & n16067 ;
  assign n16069 = n16056 & ~n16068 ;
  assign n16070 = ( n15328 & n15705 ) | ( n15328 & n15743 ) | ( n15705 & n15743 ) ;
  assign n16071 = ~n16056 & n16067 ;
  assign n16072 = n16070 | n16071 ;
  assign n16073 = n16069 | n16072 ;
  assign n16074 = ( n16069 & n16070 ) | ( n16069 & n16071 ) | ( n16070 & n16071 ) ;
  assign n16075 = n16073 & ~n16074 ;
  assign n16076 = x85 & n8834 ;
  assign n16077 = x84 & n8829 ;
  assign n16078 = x83 & ~n8828 ;
  assign n16079 = n9159 & n16078 ;
  assign n16080 = n16077 | n16079 ;
  assign n16081 = n16076 | n16080 ;
  assign n16082 = n8837 | n16081 ;
  assign n16083 = ( n1765 & n16081 ) | ( n1765 & n16082 ) | ( n16081 & n16082 ) ;
  assign n16084 = x53 & n16083 ;
  assign n16085 = x53 & ~n16084 ;
  assign n16086 = ( n16083 & ~n16084 ) | ( n16083 & n16085 ) | ( ~n16084 & n16085 ) ;
  assign n16087 = n16075 & n16086 ;
  assign n16088 = n16075 & ~n16087 ;
  assign n16089 = ~n16075 & n16086 ;
  assign n16090 = n16088 | n16089 ;
  assign n16091 = n15748 | n15762 ;
  assign n16092 = n16090 & n16091 ;
  assign n16093 = n16090 | n16091 ;
  assign n16094 = ~n16092 & n16093 ;
  assign n16095 = ( n15693 & n15763 ) | ( n15693 & n15774 ) | ( n15763 & n15774 ) ;
  assign n16096 = ( n16017 & n16094 ) | ( n16017 & n16095 ) | ( n16094 & n16095 ) ;
  assign n16097 = ( n16094 & n16095 ) | ( n16094 & ~n16096 ) | ( n16095 & ~n16096 ) ;
  assign n16098 = ( n16017 & ~n16096 ) | ( n16017 & n16097 ) | ( ~n16096 & n16097 ) ;
  assign n16099 = n16006 & n16098 ;
  assign n16100 = n16006 | n16098 ;
  assign n16101 = ~n16099 & n16100 ;
  assign n16102 = ( n15691 & n15692 ) | ( n15691 & n15777 ) | ( n15692 & n15777 ) ;
  assign n16103 = n16101 | n16102 ;
  assign n16104 = n16101 & n16102 ;
  assign n16105 = n16103 & ~n16104 ;
  assign n16106 = x94 & n6068 ;
  assign n16107 = x93 & n6063 ;
  assign n16108 = x92 & ~n6062 ;
  assign n16109 = n6398 & n16108 ;
  assign n16110 = n16107 | n16109 ;
  assign n16111 = n16106 | n16110 ;
  assign n16112 = n6071 | n16111 ;
  assign n16113 = ( n3271 & n16111 ) | ( n3271 & n16112 ) | ( n16111 & n16112 ) ;
  assign n16114 = x44 & n16113 ;
  assign n16115 = x44 & ~n16114 ;
  assign n16116 = ( n16113 & ~n16114 ) | ( n16113 & n16115 ) | ( ~n16114 & n16115 ) ;
  assign n16117 = ( n15995 & n16105 ) | ( n15995 & ~n16116 ) | ( n16105 & ~n16116 ) ;
  assign n16118 = ( ~n16105 & n16116 ) | ( ~n16105 & n16117 ) | ( n16116 & n16117 ) ;
  assign n16119 = ( ~n15995 & n16117 ) | ( ~n15995 & n16118 ) | ( n16117 & n16118 ) ;
  assign n16120 = x97 & n5340 ;
  assign n16121 = x96 & n5335 ;
  assign n16122 = x95 & ~n5334 ;
  assign n16123 = n5580 & n16122 ;
  assign n16124 = n16121 | n16123 ;
  assign n16125 = n16120 | n16124 ;
  assign n16126 = n5343 | n16125 ;
  assign n16127 = ( n3707 & n16125 ) | ( n3707 & n16126 ) | ( n16125 & n16126 ) ;
  assign n16128 = x41 & n16127 ;
  assign n16129 = x41 & ~n16128 ;
  assign n16130 = ( n16127 & ~n16128 ) | ( n16127 & n16129 ) | ( ~n16128 & n16129 ) ;
  assign n16131 = ( n15994 & n16119 ) | ( n15994 & ~n16130 ) | ( n16119 & ~n16130 ) ;
  assign n16132 = ( ~n16119 & n16130 ) | ( ~n16119 & n16131 ) | ( n16130 & n16131 ) ;
  assign n16133 = ( ~n15994 & n16131 ) | ( ~n15994 & n16132 ) | ( n16131 & n16132 ) ;
  assign n16134 = n15993 & n16133 ;
  assign n16135 = n15993 | n16133 ;
  assign n16136 = ~n16134 & n16135 ;
  assign n16137 = n15812 | n16136 ;
  assign n16138 = n15812 & n16136 ;
  assign n16139 = n16137 & ~n16138 ;
  assign n16140 = ( n15651 & n15667 ) | ( n15651 & n15814 ) | ( n15667 & n15814 ) ;
  assign n16141 = ( n15982 & n16139 ) | ( n15982 & n16140 ) | ( n16139 & n16140 ) ;
  assign n16142 = ( n16139 & n16140 ) | ( n16139 & ~n16141 ) | ( n16140 & ~n16141 ) ;
  assign n16143 = ( n15982 & ~n16141 ) | ( n15982 & n16142 ) | ( ~n16141 & n16142 ) ;
  assign n16144 = n15971 & n16143 ;
  assign n16145 = n15971 | n16143 ;
  assign n16146 = ~n16144 & n16145 ;
  assign n16147 = ( n15954 & ~n15955 ) | ( n15954 & n16146 ) | ( ~n15955 & n16146 ) ;
  assign n16148 = ( n15955 & ~n16146 ) | ( n15955 & n16147 ) | ( ~n16146 & n16147 ) ;
  assign n16149 = ( ~n15954 & n16147 ) | ( ~n15954 & n16148 ) | ( n16147 & n16148 ) ;
  assign n16150 = n15943 & ~n16149 ;
  assign n16151 = n16149 | n16150 ;
  assign n16152 = ( ~n15943 & n16150 ) | ( ~n15943 & n16151 ) | ( n16150 & n16151 ) ;
  assign n16153 = x115 & n1817 ;
  assign n16154 = x114 & n1812 ;
  assign n16155 = x113 & ~n1811 ;
  assign n16156 = n1977 & n16155 ;
  assign n16157 = n16154 | n16156 ;
  assign n16158 = n16153 | n16157 ;
  assign n16159 = n1820 | n16158 ;
  assign n16160 = ( n8749 & n16158 ) | ( n8749 & n16159 ) | ( n16158 & n16159 ) ;
  assign n16161 = x23 & n16160 ;
  assign n16162 = x23 & ~n16161 ;
  assign n16163 = ( n16160 & ~n16161 ) | ( n16160 & n16162 ) | ( ~n16161 & n16162 ) ;
  assign n16164 = n15604 | n15828 ;
  assign n16165 = ( n16152 & n16163 ) | ( n16152 & ~n16164 ) | ( n16163 & ~n16164 ) ;
  assign n16166 = ( ~n16163 & n16164 ) | ( ~n16163 & n16165 ) | ( n16164 & n16165 ) ;
  assign n16167 = ( ~n16152 & n16165 ) | ( ~n16152 & n16166 ) | ( n16165 & n16166 ) ;
  assign n16168 = n15927 & n16167 ;
  assign n16169 = n15927 | n16167 ;
  assign n16170 = ~n16168 & n16169 ;
  assign n16171 = ( n15853 & n15854 ) | ( n15853 & n15865 ) | ( n15854 & n15865 ) ;
  assign n16172 = x121 & n1071 ;
  assign n16173 = x120 & n1066 ;
  assign n16174 = x119 & ~n1065 ;
  assign n16175 = n1189 & n16174 ;
  assign n16176 = n16173 | n16175 ;
  assign n16177 = n16172 | n16176 ;
  assign n16178 = n1074 | n16177 ;
  assign n16179 = ( n10811 & n16177 ) | ( n10811 & n16178 ) | ( n16177 & n16178 ) ;
  assign n16180 = x17 & n16179 ;
  assign n16181 = x17 & ~n16180 ;
  assign n16182 = ( n16179 & ~n16180 ) | ( n16179 & n16181 ) | ( ~n16180 & n16181 ) ;
  assign n16183 = n16171 | n16182 ;
  assign n16184 = n16171 & n16182 ;
  assign n16185 = n16183 & ~n16184 ;
  assign n16186 = n15879 & n15880 ;
  assign n16187 = n15868 & ~n15882 ;
  assign n16188 = ( n15868 & ~n15881 ) | ( n15868 & n16187 ) | ( ~n15881 & n16187 ) ;
  assign n16189 = n16186 | n16188 ;
  assign n16190 = x124 & n771 ;
  assign n16191 = x123 & n766 ;
  assign n16192 = x122 & ~n765 ;
  assign n16193 = n905 & n16192 ;
  assign n16194 = n16191 | n16193 ;
  assign n16195 = n16190 | n16194 ;
  assign n16196 = n774 | n16195 ;
  assign n16197 = ( n11916 & n16195 ) | ( n11916 & n16196 ) | ( n16195 & n16196 ) ;
  assign n16198 = x14 & n16197 ;
  assign n16199 = x14 & ~n16198 ;
  assign n16200 = ( n16197 & ~n16198 ) | ( n16197 & n16199 ) | ( ~n16198 & n16199 ) ;
  assign n16201 = n16189 | n16200 ;
  assign n16202 = ~n16200 & n16201 ;
  assign n16203 = ( ~n16189 & n16201 ) | ( ~n16189 & n16202 ) | ( n16201 & n16202 ) ;
  assign n16204 = ( n16170 & ~n16185 ) | ( n16170 & n16203 ) | ( ~n16185 & n16203 ) ;
  assign n16205 = ( n16185 & ~n16203 ) | ( n16185 & n16204 ) | ( ~n16203 & n16204 ) ;
  assign n16206 = ( ~n16170 & n16204 ) | ( ~n16170 & n16205 ) | ( n16204 & n16205 ) ;
  assign n16207 = ( n15909 & ~n15910 ) | ( n15909 & n16206 ) | ( ~n15910 & n16206 ) ;
  assign n16208 = ( n15910 & ~n16206 ) | ( n15910 & n16207 ) | ( ~n16206 & n16207 ) ;
  assign n16209 = ( ~n15909 & n16207 ) | ( ~n15909 & n16208 ) | ( n16207 & n16208 ) ;
  assign n16210 = n15573 & n16209 ;
  assign n16211 = ( n15891 & n16209 ) | ( n15891 & n16210 ) | ( n16209 & n16210 ) ;
  assign n16212 = n15898 & ~n16211 ;
  assign n16213 = ( n15557 & n15892 ) | ( n15557 & n15894 ) | ( n15892 & n15894 ) ;
  assign n16214 = n15892 | n15894 ;
  assign n16215 = ( n15562 & n16213 ) | ( n15562 & n16214 ) | ( n16213 & n16214 ) ;
  assign n16216 = n16209 & ~n16210 ;
  assign n16217 = ~n15891 & n16216 ;
  assign n16218 = n16215 | n16217 ;
  assign n16219 = n16212 | n16218 ;
  assign n16220 = n16212 | n16217 ;
  assign n16221 = n16213 & n16220 ;
  assign n16222 = n16214 & n16220 ;
  assign n16223 = ( n15562 & n16221 ) | ( n15562 & n16222 ) | ( n16221 & n16222 ) ;
  assign n16224 = n16219 & ~n16223 ;
  assign n16225 = n16203 & ~n16206 ;
  assign n16226 = ( n16186 & n16188 ) | ( n16186 & n16200 ) | ( n16188 & n16200 ) ;
  assign n16227 = n16225 | n16226 ;
  assign n16228 = x127 & n523 ;
  assign n16229 = x126 & ~n522 ;
  assign n16230 = n635 & n16229 ;
  assign n16231 = n16228 | n16230 ;
  assign n16232 = n531 | n16231 ;
  assign n16233 = ( n13461 & n16231 ) | ( n13461 & n16232 ) | ( n16231 & n16232 ) ;
  assign n16234 = x11 & n16233 ;
  assign n16235 = x11 & ~n16234 ;
  assign n16236 = ( n16233 & ~n16234 ) | ( n16233 & n16235 ) | ( ~n16234 & n16235 ) ;
  assign n16237 = n16227 & n16236 ;
  assign n16238 = n16227 & ~n16237 ;
  assign n16239 = ~n16227 & n16236 ;
  assign n16240 = x113 & n2280 ;
  assign n16241 = x112 & n2275 ;
  assign n16242 = x111 & ~n2274 ;
  assign n16243 = n2481 & n16242 ;
  assign n16244 = n16241 | n16243 ;
  assign n16245 = n16240 | n16244 ;
  assign n16246 = n2283 | n16245 ;
  assign n16247 = ( n8113 & n16245 ) | ( n8113 & n16246 ) | ( n16245 & n16246 ) ;
  assign n16248 = x26 & n16247 ;
  assign n16249 = x26 & ~n16248 ;
  assign n16250 = ( n16247 & ~n16248 ) | ( n16247 & n16249 ) | ( ~n16248 & n16249 ) ;
  assign n16251 = ( n15637 & n15821 ) | ( n15637 & n15954 ) | ( n15821 & n15954 ) ;
  assign n16252 = n16250 & n16251 ;
  assign n16253 = n16250 & ~n16252 ;
  assign n16254 = ( n15954 & n15955 ) | ( n15954 & n16146 ) | ( n15955 & n16146 ) ;
  assign n16255 = ~n15955 & n16254 ;
  assign n16256 = ( n16146 & ~n16147 ) | ( n16146 & n16255 ) | ( ~n16147 & n16255 ) ;
  assign n16257 = n16253 & ~n16256 ;
  assign n16258 = ( ~n16250 & n16251 ) | ( ~n16250 & n16256 ) | ( n16251 & n16256 ) ;
  assign n16259 = n16257 | n16258 ;
  assign n16260 = x110 & n2775 ;
  assign n16261 = x109 & n2770 ;
  assign n16262 = x108 & ~n2769 ;
  assign n16263 = n2978 & n16262 ;
  assign n16264 = n16261 | n16263 ;
  assign n16265 = n16260 | n16264 ;
  assign n16266 = n2778 | n16265 ;
  assign n16267 = ( n7189 & n16265 ) | ( n7189 & n16266 ) | ( n16265 & n16266 ) ;
  assign n16268 = x29 & n16267 ;
  assign n16269 = x29 & ~n16268 ;
  assign n16270 = ( n16267 & ~n16268 ) | ( n16267 & n16269 ) | ( ~n16268 & n16269 ) ;
  assign n16271 = n15968 & n16270 ;
  assign n16272 = n16270 & ~n16271 ;
  assign n16273 = ~n16144 & n16272 ;
  assign n16274 = ( n15968 & n16144 ) | ( n15968 & ~n16270 ) | ( n16144 & ~n16270 ) ;
  assign n16275 = n16273 | n16274 ;
  assign n16276 = x104 & n3913 ;
  assign n16277 = x103 & n3908 ;
  assign n16278 = x102 & ~n3907 ;
  assign n16279 = n4152 & n16278 ;
  assign n16280 = n16277 | n16279 ;
  assign n16281 = n16276 | n16280 ;
  assign n16282 = n3916 | n16281 ;
  assign n16283 = ( n5295 & n16281 ) | ( n5295 & n16282 ) | ( n16281 & n16282 ) ;
  assign n16284 = x35 & n16283 ;
  assign n16285 = x35 & ~n16284 ;
  assign n16286 = ( n16283 & ~n16284 ) | ( n16283 & n16285 ) | ( ~n16284 & n16285 ) ;
  assign n16287 = ( n15994 & n16119 ) | ( n15994 & n16130 ) | ( n16119 & n16130 ) ;
  assign n16288 = n16099 | n16104 ;
  assign n16289 = x92 & n6937 ;
  assign n16290 = x91 & n6932 ;
  assign n16291 = x90 & ~n6931 ;
  assign n16292 = n7216 & n16291 ;
  assign n16293 = n16290 | n16292 ;
  assign n16294 = n16289 | n16293 ;
  assign n16295 = n6940 | n16294 ;
  assign n16296 = ( n2904 & n16294 ) | ( n2904 & n16295 ) | ( n16294 & n16295 ) ;
  assign n16297 = x47 & n16296 ;
  assign n16298 = x47 & ~n16297 ;
  assign n16299 = ( n16296 & ~n16297 ) | ( n16296 & n16298 ) | ( ~n16297 & n16298 ) ;
  assign n16300 = n16087 | n16092 ;
  assign n16301 = n16068 | n16074 ;
  assign n16302 = x80 & n10876 ;
  assign n16303 = x79 & n10871 ;
  assign n16304 = x78 & ~n10870 ;
  assign n16305 = n11305 & n16304 ;
  assign n16306 = n16303 | n16305 ;
  assign n16307 = n16302 | n16306 ;
  assign n16308 = n10879 | n16307 ;
  assign n16309 = ( n1147 & n16307 ) | ( n1147 & n16308 ) | ( n16307 & n16308 ) ;
  assign n16310 = x59 & n16309 ;
  assign n16311 = x59 & ~n16310 ;
  assign n16312 = ( n16309 & ~n16310 ) | ( n16309 & n16311 ) | ( ~n16310 & n16311 ) ;
  assign n16313 = x77 & n11984 ;
  assign n16314 = x76 & n11979 ;
  assign n16315 = x75 & ~n11978 ;
  assign n16316 = n12430 & n16315 ;
  assign n16317 = n16314 | n16316 ;
  assign n16318 = n16313 | n16317 ;
  assign n16319 = n11987 | n16318 ;
  assign n16320 = ( n846 & n16318 ) | ( n846 & n16319 ) | ( n16318 & n16319 ) ;
  assign n16321 = ~x62 & n16320 ;
  assign n16322 = x62 & ~n16320 ;
  assign n16323 = n16321 | n16322 ;
  assign n16324 = x74 & n12808 ;
  assign n16325 = x63 & x73 ;
  assign n16326 = ~n12808 & n16325 ;
  assign n16327 = n16324 | n16326 ;
  assign n16328 = n16045 & ~n16327 ;
  assign n16329 = n16045 & ~n16328 ;
  assign n16330 = n16045 | n16327 ;
  assign n16331 = ~n16329 & n16330 ;
  assign n16332 = n16323 & ~n16331 ;
  assign n16333 = ~n16323 & n16331 ;
  assign n16334 = n16332 | n16333 ;
  assign n16335 = ( n15726 & ~n16039 ) | ( n15726 & n16046 ) | ( ~n16039 & n16046 ) ;
  assign n16336 = n16334 | n16335 ;
  assign n16337 = ~n16335 & n16336 ;
  assign n16338 = ( ~n16334 & n16336 ) | ( ~n16334 & n16337 ) | ( n16336 & n16337 ) ;
  assign n16339 = ~n16312 & n16338 ;
  assign n16340 = n16312 & ~n16338 ;
  assign n16341 = n16050 | n16055 ;
  assign n16342 = n16340 | n16341 ;
  assign n16343 = n16339 | n16342 ;
  assign n16344 = ( n16339 & n16340 ) | ( n16339 & n16341 ) | ( n16340 & n16341 ) ;
  assign n16345 = n16343 & ~n16344 ;
  assign n16346 = x83 & n9853 ;
  assign n16347 = x82 & n9848 ;
  assign n16348 = x81 & ~n9847 ;
  assign n16349 = n10165 & n16348 ;
  assign n16350 = n16347 | n16349 ;
  assign n16351 = n16346 | n16350 ;
  assign n16352 = n9856 | n16351 ;
  assign n16353 = ( n1510 & n16351 ) | ( n1510 & n16352 ) | ( n16351 & n16352 ) ;
  assign n16354 = x56 & n16353 ;
  assign n16355 = x56 & ~n16354 ;
  assign n16356 = ( n16353 & ~n16354 ) | ( n16353 & n16355 ) | ( ~n16354 & n16355 ) ;
  assign n16357 = n16345 & ~n16356 ;
  assign n16358 = n16356 | n16357 ;
  assign n16359 = ( ~n16345 & n16357 ) | ( ~n16345 & n16358 ) | ( n16357 & n16358 ) ;
  assign n16360 = n16301 | n16359 ;
  assign n16361 = x86 & n8834 ;
  assign n16362 = x85 & n8829 ;
  assign n16363 = x84 & ~n8828 ;
  assign n16364 = n9159 & n16363 ;
  assign n16365 = n16362 | n16364 ;
  assign n16366 = n16361 | n16365 ;
  assign n16367 = n8837 | n16366 ;
  assign n16368 = ( n1921 & n16366 ) | ( n1921 & n16367 ) | ( n16366 & n16367 ) ;
  assign n16369 = x53 & n16368 ;
  assign n16370 = x53 & ~n16369 ;
  assign n16371 = ( n16368 & ~n16369 ) | ( n16368 & n16370 ) | ( ~n16369 & n16370 ) ;
  assign n16372 = ( n16359 & ~n16360 ) | ( n16359 & n16371 ) | ( ~n16360 & n16371 ) ;
  assign n16373 = ( n16301 & ~n16360 ) | ( n16301 & n16372 ) | ( ~n16360 & n16372 ) ;
  assign n16374 = n16300 | n16373 ;
  assign n16375 = ( n16301 & n16359 ) | ( n16301 & n16371 ) | ( n16359 & n16371 ) ;
  assign n16376 = n16360 & ~n16375 ;
  assign n16377 = n16374 | n16376 ;
  assign n16378 = ( n16300 & n16373 ) | ( n16300 & n16376 ) | ( n16373 & n16376 ) ;
  assign n16379 = n16377 & ~n16378 ;
  assign n16380 = x89 & n7812 ;
  assign n16381 = x88 & n7807 ;
  assign n16382 = x87 & ~n7806 ;
  assign n16383 = n8136 & n16382 ;
  assign n16384 = n16381 | n16383 ;
  assign n16385 = n16380 | n16384 ;
  assign n16386 = n7815 | n16385 ;
  assign n16387 = ( n2244 & n16385 ) | ( n2244 & n16386 ) | ( n16385 & n16386 ) ;
  assign n16388 = x50 & n16387 ;
  assign n16389 = x50 & ~n16388 ;
  assign n16390 = ( n16387 & ~n16388 ) | ( n16387 & n16389 ) | ( ~n16388 & n16389 ) ;
  assign n16391 = n16379 & ~n16390 ;
  assign n16392 = n16390 | n16391 ;
  assign n16393 = ( ~n16379 & n16391 ) | ( ~n16379 & n16392 ) | ( n16391 & n16392 ) ;
  assign n16394 = ( ~n16096 & n16299 ) | ( ~n16096 & n16393 ) | ( n16299 & n16393 ) ;
  assign n16395 = ( n16096 & ~n16393 ) | ( n16096 & n16394 ) | ( ~n16393 & n16394 ) ;
  assign n16396 = ( ~n16299 & n16394 ) | ( ~n16299 & n16395 ) | ( n16394 & n16395 ) ;
  assign n16397 = n16288 | n16396 ;
  assign n16398 = n16288 & n16396 ;
  assign n16399 = n16397 & ~n16398 ;
  assign n16400 = x95 & n6068 ;
  assign n16401 = x94 & n6063 ;
  assign n16402 = x93 & ~n6062 ;
  assign n16403 = n6398 & n16402 ;
  assign n16404 = n16401 | n16403 ;
  assign n16405 = n16400 | n16404 ;
  assign n16406 = n6071 | n16405 ;
  assign n16407 = ( n3479 & n16405 ) | ( n3479 & n16406 ) | ( n16405 & n16406 ) ;
  assign n16408 = x44 & n16407 ;
  assign n16409 = x44 & ~n16408 ;
  assign n16410 = ( n16407 & ~n16408 ) | ( n16407 & n16409 ) | ( ~n16408 & n16409 ) ;
  assign n16411 = n16399 | n16410 ;
  assign n16412 = n16399 & n16410 ;
  assign n16413 = n16411 & ~n16412 ;
  assign n16414 = ( n15995 & n16105 ) | ( n15995 & n16116 ) | ( n16105 & n16116 ) ;
  assign n16415 = n16413 & n16414 ;
  assign n16416 = n16413 | n16414 ;
  assign n16417 = ~n16415 & n16416 ;
  assign n16418 = x98 & n5340 ;
  assign n16419 = x97 & n5335 ;
  assign n16420 = x96 & ~n5334 ;
  assign n16421 = n5580 & n16420 ;
  assign n16422 = n16419 | n16421 ;
  assign n16423 = n16418 | n16422 ;
  assign n16424 = n5343 | n16423 ;
  assign n16425 = ( n4105 & n16423 ) | ( n4105 & n16424 ) | ( n16423 & n16424 ) ;
  assign n16426 = x41 & n16425 ;
  assign n16427 = x41 & ~n16426 ;
  assign n16428 = ( n16425 & ~n16426 ) | ( n16425 & n16427 ) | ( ~n16426 & n16427 ) ;
  assign n16429 = n16417 & n16428 ;
  assign n16430 = n16417 | n16428 ;
  assign n16431 = ~n16429 & n16430 ;
  assign n16432 = x101 & n4572 ;
  assign n16433 = x100 & n4567 ;
  assign n16434 = x99 & ~n4566 ;
  assign n16435 = n4828 & n16434 ;
  assign n16436 = n16433 | n16435 ;
  assign n16437 = n16432 | n16436 ;
  assign n16438 = n4575 | n16437 ;
  assign n16439 = ( n4783 & n16437 ) | ( n4783 & n16438 ) | ( n16437 & n16438 ) ;
  assign n16440 = x38 & n16439 ;
  assign n16441 = x38 & ~n16440 ;
  assign n16442 = ( n16439 & ~n16440 ) | ( n16439 & n16441 ) | ( ~n16440 & n16441 ) ;
  assign n16443 = ( n16287 & ~n16431 ) | ( n16287 & n16442 ) | ( ~n16431 & n16442 ) ;
  assign n16444 = ( n16431 & ~n16442 ) | ( n16431 & n16443 ) | ( ~n16442 & n16443 ) ;
  assign n16445 = ( ~n16287 & n16443 ) | ( ~n16287 & n16444 ) | ( n16443 & n16444 ) ;
  assign n16446 = n16134 | n16138 ;
  assign n16447 = n16445 & n16446 ;
  assign n16448 = n16446 & ~n16447 ;
  assign n16449 = ( n16445 & ~n16447 ) | ( n16445 & n16448 ) | ( ~n16447 & n16448 ) ;
  assign n16450 = n16286 & n16449 ;
  assign n16451 = n16286 | n16449 ;
  assign n16452 = ~n16450 & n16451 ;
  assign n16453 = x107 & n3314 ;
  assign n16454 = x106 & n3309 ;
  assign n16455 = x105 & ~n3308 ;
  assign n16456 = n3570 & n16455 ;
  assign n16457 = n16454 | n16456 ;
  assign n16458 = n16453 | n16457 ;
  assign n16459 = n3317 | n16458 ;
  assign n16460 = ( n6328 & n16458 ) | ( n6328 & n16459 ) | ( n16458 & n16459 ) ;
  assign n16461 = x32 & n16460 ;
  assign n16462 = x32 & ~n16461 ;
  assign n16463 = ( n16460 & ~n16461 ) | ( n16460 & n16462 ) | ( ~n16461 & n16462 ) ;
  assign n16464 = ( ~n16141 & n16452 ) | ( ~n16141 & n16463 ) | ( n16452 & n16463 ) ;
  assign n16465 = ( n16141 & ~n16463 ) | ( n16141 & n16464 ) | ( ~n16463 & n16464 ) ;
  assign n16466 = ( ~n16452 & n16464 ) | ( ~n16452 & n16465 ) | ( n16464 & n16465 ) ;
  assign n16467 = n16275 & n16466 ;
  assign n16468 = n16275 | n16466 ;
  assign n16469 = ~n16467 & n16468 ;
  assign n16470 = n16259 & n16469 ;
  assign n16471 = n16259 | n16469 ;
  assign n16472 = ~n16470 & n16471 ;
  assign n16473 = x119 & n1421 ;
  assign n16474 = x118 & n1416 ;
  assign n16475 = x117 & ~n1415 ;
  assign n16476 = n1584 & n16475 ;
  assign n16477 = n16474 | n16476 ;
  assign n16478 = n16473 | n16477 ;
  assign n16479 = n1424 | n16478 ;
  assign n16480 = ( n9789 & n16478 ) | ( n9789 & n16479 ) | ( n16478 & n16479 ) ;
  assign n16481 = x20 & n16480 ;
  assign n16482 = x20 & ~n16481 ;
  assign n16483 = ( n16480 & ~n16481 ) | ( n16480 & n16482 ) | ( ~n16481 & n16482 ) ;
  assign n16484 = ( n16152 & n16163 ) | ( n16152 & n16164 ) | ( n16163 & n16164 ) ;
  assign n16485 = n16483 | n16484 ;
  assign n16486 = n16483 & n16484 ;
  assign n16487 = n16485 & ~n16486 ;
  assign n16488 = x116 & n1817 ;
  assign n16489 = x115 & n1812 ;
  assign n16490 = x114 & ~n1811 ;
  assign n16491 = n1977 & n16490 ;
  assign n16492 = n16489 | n16491 ;
  assign n16493 = n16488 | n16492 ;
  assign n16494 = n1820 | n16493 ;
  assign n16495 = ( n8778 & n16493 ) | ( n8778 & n16494 ) | ( n16493 & n16494 ) ;
  assign n16496 = x23 & n16495 ;
  assign n16497 = x23 & ~n16496 ;
  assign n16498 = ( n16495 & ~n16496 ) | ( n16495 & n16497 ) | ( ~n16496 & n16497 ) ;
  assign n16499 = ( n15941 & n15942 ) | ( n15941 & n16149 ) | ( n15942 & n16149 ) ;
  assign n16500 = n16498 | n16499 ;
  assign n16501 = n16498 & n16499 ;
  assign n16502 = n16500 & ~n16501 ;
  assign n16503 = ( n16472 & n16487 ) | ( n16472 & ~n16502 ) | ( n16487 & ~n16502 ) ;
  assign n16504 = ( ~n16487 & n16502 ) | ( ~n16487 & n16503 ) | ( n16502 & n16503 ) ;
  assign n16505 = ( ~n16472 & n16503 ) | ( ~n16472 & n16504 ) | ( n16503 & n16504 ) ;
  assign n16506 = x122 & n1071 ;
  assign n16507 = x121 & n1066 ;
  assign n16508 = x120 & ~n1065 ;
  assign n16509 = n1189 & n16508 ;
  assign n16510 = n16507 | n16509 ;
  assign n16511 = n16506 | n16510 ;
  assign n16512 = n1074 | n16511 ;
  assign n16513 = ( n11188 & n16511 ) | ( n11188 & n16512 ) | ( n16511 & n16512 ) ;
  assign n16514 = x17 & n16513 ;
  assign n16515 = x17 & ~n16514 ;
  assign n16516 = ( n16513 & ~n16514 ) | ( n16513 & n16515 ) | ( ~n16514 & n16515 ) ;
  assign n16517 = ( n15924 & n16168 ) | ( n15924 & n16516 ) | ( n16168 & n16516 ) ;
  assign n16518 = ( n15924 & n16168 ) | ( n15924 & ~n16516 ) | ( n16168 & ~n16516 ) ;
  assign n16519 = ( n16516 & ~n16517 ) | ( n16516 & n16518 ) | ( ~n16517 & n16518 ) ;
  assign n16520 = n16505 & n16519 ;
  assign n16521 = n16505 | n16519 ;
  assign n16522 = ~n16520 & n16521 ;
  assign n16523 = ( n16170 & n16171 ) | ( n16170 & n16182 ) | ( n16171 & n16182 ) ;
  assign n16524 = x125 & n771 ;
  assign n16525 = x124 & n766 ;
  assign n16526 = x123 & ~n765 ;
  assign n16527 = n905 & n16526 ;
  assign n16528 = n16525 | n16527 ;
  assign n16529 = n16524 | n16528 ;
  assign n16530 = n774 | n16529 ;
  assign n16531 = ( n12310 & n16529 ) | ( n12310 & n16530 ) | ( n16529 & n16530 ) ;
  assign n16532 = x14 & n16531 ;
  assign n16533 = x14 & ~n16532 ;
  assign n16534 = ( n16531 & ~n16532 ) | ( n16531 & n16533 ) | ( ~n16532 & n16533 ) ;
  assign n16535 = n16523 & n16534 ;
  assign n16536 = n16534 & ~n16535 ;
  assign n16537 = ( n16523 & ~n16535 ) | ( n16523 & n16536 ) | ( ~n16535 & n16536 ) ;
  assign n16538 = n16522 & n16537 ;
  assign n16539 = n16522 | n16537 ;
  assign n16540 = ~n16538 & n16539 ;
  assign n16541 = n16239 | n16540 ;
  assign n16542 = n16238 | n16541 ;
  assign n16543 = ( n16238 & n16239 ) | ( n16238 & n16540 ) | ( n16239 & n16540 ) ;
  assign n16544 = n16542 & ~n16543 ;
  assign n16545 = ( n15909 & n15910 ) | ( n15909 & n16206 ) | ( n15910 & n16206 ) ;
  assign n16546 = n16544 & ~n16545 ;
  assign n16547 = n16211 | n16221 ;
  assign n16548 = n16544 & n16545 ;
  assign n16549 = n16545 & ~n16548 ;
  assign n16550 = n16546 | n16549 ;
  assign n16551 = n16547 & n16550 ;
  assign n16552 = n16211 | n16222 ;
  assign n16553 = n16550 & n16552 ;
  assign n16554 = ( n15562 & n16551 ) | ( n15562 & n16553 ) | ( n16551 & n16553 ) ;
  assign n16555 = ( n15562 & n16547 ) | ( n15562 & n16552 ) | ( n16547 & n16552 ) ;
  assign n16556 = ( ~n16544 & n16545 ) | ( ~n16544 & n16555 ) | ( n16545 & n16555 ) ;
  assign n16557 = ( n16546 & ~n16554 ) | ( n16546 & n16556 ) | ( ~n16554 & n16556 ) ;
  assign n16558 = n16237 | n16543 ;
  assign n16559 = x127 & ~n522 ;
  assign n16560 = n635 & n16559 ;
  assign n16561 = ( x127 & n531 ) | ( x127 & n16560 ) | ( n531 & n16560 ) ;
  assign n16562 = ( x126 & n16560 ) | ( x126 & n16561 ) | ( n16560 & n16561 ) ;
  assign n16563 = ( n12685 & n16561 ) | ( n12685 & n16562 ) | ( n16561 & n16562 ) ;
  assign n16564 = x11 & n16563 ;
  assign n16565 = x11 & ~n16564 ;
  assign n16566 = ( n16563 & ~n16564 ) | ( n16563 & n16565 ) | ( ~n16564 & n16565 ) ;
  assign n16567 = n16535 | n16538 ;
  assign n16568 = ( n16472 & n16498 ) | ( n16472 & n16499 ) | ( n16498 & n16499 ) ;
  assign n16569 = x120 & n1421 ;
  assign n16570 = x119 & n1416 ;
  assign n16571 = x118 & ~n1415 ;
  assign n16572 = n1584 & n16571 ;
  assign n16573 = n16570 | n16572 ;
  assign n16574 = n16569 | n16573 ;
  assign n16575 = n1424 | n16574 ;
  assign n16576 = ( n10460 & n16574 ) | ( n10460 & n16575 ) | ( n16574 & n16575 ) ;
  assign n16577 = x20 & n16576 ;
  assign n16578 = x20 & ~n16577 ;
  assign n16579 = ( n16576 & ~n16577 ) | ( n16576 & n16578 ) | ( ~n16577 & n16578 ) ;
  assign n16580 = n16568 & n16579 ;
  assign n16581 = n16568 & ~n16580 ;
  assign n16582 = ~n16568 & n16579 ;
  assign n16583 = n16581 | n16582 ;
  assign n16584 = x108 & n3314 ;
  assign n16585 = x107 & n3309 ;
  assign n16586 = x106 & ~n3308 ;
  assign n16587 = n3570 & n16586 ;
  assign n16588 = n16585 | n16587 ;
  assign n16589 = n16584 | n16588 ;
  assign n16590 = n3317 | n16589 ;
  assign n16591 = ( n6358 & n16589 ) | ( n6358 & n16590 ) | ( n16589 & n16590 ) ;
  assign n16592 = x32 & n16591 ;
  assign n16593 = x32 & ~n16592 ;
  assign n16594 = ( n16591 & ~n16592 ) | ( n16591 & n16593 ) | ( ~n16592 & n16593 ) ;
  assign n16595 = n16447 | n16594 ;
  assign n16596 = n16450 | n16595 ;
  assign n16597 = ( n16447 & n16450 ) | ( n16447 & n16594 ) | ( n16450 & n16594 ) ;
  assign n16598 = n16596 & ~n16597 ;
  assign n16599 = ( n16287 & n16431 ) | ( n16287 & n16442 ) | ( n16431 & n16442 ) ;
  assign n16600 = n16415 | n16429 ;
  assign n16601 = n16398 | n16412 ;
  assign n16602 = ( n16096 & n16299 ) | ( n16096 & n16393 ) | ( n16299 & n16393 ) ;
  assign n16603 = ( n16377 & n16378 ) | ( n16377 & n16390 ) | ( n16378 & n16390 ) ;
  assign n16604 = x78 & n11984 ;
  assign n16605 = x77 & n11979 ;
  assign n16606 = x76 & ~n11978 ;
  assign n16607 = n12430 & n16606 ;
  assign n16608 = n16605 | n16607 ;
  assign n16609 = n16604 | n16608 ;
  assign n16610 = n11987 | n16609 ;
  assign n16611 = ( n868 & n16609 ) | ( n868 & n16610 ) | ( n16609 & n16610 ) ;
  assign n16612 = x62 & n16611 ;
  assign n16613 = x62 & ~n16612 ;
  assign n16614 = ( n16611 & ~n16612 ) | ( n16611 & n16613 ) | ( ~n16612 & n16613 ) ;
  assign n16615 = n16328 | n16332 ;
  assign n16616 = x75 & n12808 ;
  assign n16617 = x63 & x74 ;
  assign n16618 = ~n12808 & n16617 ;
  assign n16619 = n16616 | n16618 ;
  assign n16620 = ~n16327 & n16619 ;
  assign n16621 = n16327 | n16620 ;
  assign n16622 = n16619 & ~n16620 ;
  assign n16623 = n16621 & ~n16622 ;
  assign n16624 = n16615 | n16623 ;
  assign n16625 = n16328 & ~n16623 ;
  assign n16626 = ( n16332 & ~n16623 ) | ( n16332 & n16625 ) | ( ~n16623 & n16625 ) ;
  assign n16627 = ( ~n16615 & n16624 ) | ( ~n16615 & n16626 ) | ( n16624 & n16626 ) ;
  assign n16628 = n16614 & ~n16627 ;
  assign n16629 = ~n16614 & n16627 ;
  assign n16630 = n16628 | n16629 ;
  assign n16631 = x81 & n10876 ;
  assign n16632 = x80 & n10871 ;
  assign n16633 = x79 & ~n10870 ;
  assign n16634 = n11305 & n16633 ;
  assign n16635 = n16632 | n16634 ;
  assign n16636 = n16631 | n16635 ;
  assign n16637 = n10879 | n16636 ;
  assign n16638 = ( n1256 & n16636 ) | ( n1256 & n16637 ) | ( n16636 & n16637 ) ;
  assign n16639 = x59 & n16638 ;
  assign n16640 = x59 & ~n16639 ;
  assign n16641 = ( n16638 & ~n16639 ) | ( n16638 & n16640 ) | ( ~n16639 & n16640 ) ;
  assign n16642 = ~n16630 & n16641 ;
  assign n16643 = n16630 | n16642 ;
  assign n16644 = n16630 & n16641 ;
  assign n16645 = ( n16334 & n16335 ) | ( n16334 & n16339 ) | ( n16335 & n16339 ) ;
  assign n16646 = ~n16644 & n16645 ;
  assign n16647 = n16643 & n16646 ;
  assign n16648 = ( n16643 & ~n16644 ) | ( n16643 & n16645 ) | ( ~n16644 & n16645 ) ;
  assign n16649 = ~n16647 & n16648 ;
  assign n16650 = x84 & n9853 ;
  assign n16651 = x83 & n9848 ;
  assign n16652 = x82 & ~n9847 ;
  assign n16653 = n10165 & n16652 ;
  assign n16654 = n16651 | n16653 ;
  assign n16655 = n16650 | n16654 ;
  assign n16656 = n9856 | n16655 ;
  assign n16657 = ( n1537 & n16655 ) | ( n1537 & n16656 ) | ( n16655 & n16656 ) ;
  assign n16658 = x56 & n16657 ;
  assign n16659 = x56 & ~n16658 ;
  assign n16660 = ( n16657 & ~n16658 ) | ( n16657 & n16659 ) | ( ~n16658 & n16659 ) ;
  assign n16661 = n16649 | n16660 ;
  assign n16662 = n16649 & n16660 ;
  assign n16663 = n16661 & ~n16662 ;
  assign n16664 = ( n16343 & n16344 ) | ( n16343 & n16356 ) | ( n16344 & n16356 ) ;
  assign n16665 = ~n16663 & n16664 ;
  assign n16666 = n16663 & n16664 ;
  assign n16667 = n16663 & ~n16666 ;
  assign n16668 = x87 & n8834 ;
  assign n16669 = x86 & n8829 ;
  assign n16670 = x85 & ~n8828 ;
  assign n16671 = n9159 & n16670 ;
  assign n16672 = n16669 | n16671 ;
  assign n16673 = n16668 | n16672 ;
  assign n16674 = n8837 | n16673 ;
  assign n16675 = ( n2067 & n16673 ) | ( n2067 & n16674 ) | ( n16673 & n16674 ) ;
  assign n16676 = x53 & n16675 ;
  assign n16677 = x53 & ~n16676 ;
  assign n16678 = ( n16675 & ~n16676 ) | ( n16675 & n16677 ) | ( ~n16676 & n16677 ) ;
  assign n16679 = n16667 | n16678 ;
  assign n16680 = n16665 | n16679 ;
  assign n16681 = ( n16665 & n16667 ) | ( n16665 & n16678 ) | ( n16667 & n16678 ) ;
  assign n16682 = n16680 & ~n16681 ;
  assign n16683 = n16375 & n16682 ;
  assign n16684 = n16375 | n16682 ;
  assign n16685 = ~n16683 & n16684 ;
  assign n16686 = x90 & n7812 ;
  assign n16687 = x89 & n7807 ;
  assign n16688 = x88 & ~n7806 ;
  assign n16689 = n8136 & n16688 ;
  assign n16690 = n16687 | n16689 ;
  assign n16691 = n16686 | n16690 ;
  assign n16692 = n7815 | n16691 ;
  assign n16693 = ( n2410 & n16691 ) | ( n2410 & n16692 ) | ( n16691 & n16692 ) ;
  assign n16694 = x50 & n16693 ;
  assign n16695 = x50 & ~n16694 ;
  assign n16696 = ( n16693 & ~n16694 ) | ( n16693 & n16695 ) | ( ~n16694 & n16695 ) ;
  assign n16697 = n16685 & n16696 ;
  assign n16698 = n16685 | n16696 ;
  assign n16699 = ~n16697 & n16698 ;
  assign n16700 = x93 & n6937 ;
  assign n16701 = x92 & n6932 ;
  assign n16702 = x91 & ~n6931 ;
  assign n16703 = n7216 & n16702 ;
  assign n16704 = n16701 | n16703 ;
  assign n16705 = n16700 | n16704 ;
  assign n16706 = n6940 | n16705 ;
  assign n16707 = ( n2931 & n16705 ) | ( n2931 & n16706 ) | ( n16705 & n16706 ) ;
  assign n16708 = x47 & n16707 ;
  assign n16709 = x47 & ~n16708 ;
  assign n16710 = ( n16707 & ~n16708 ) | ( n16707 & n16709 ) | ( ~n16708 & n16709 ) ;
  assign n16711 = ( n16603 & n16699 ) | ( n16603 & n16710 ) | ( n16699 & n16710 ) ;
  assign n16712 = ( n16699 & n16710 ) | ( n16699 & ~n16711 ) | ( n16710 & ~n16711 ) ;
  assign n16713 = ( n16603 & ~n16711 ) | ( n16603 & n16712 ) | ( ~n16711 & n16712 ) ;
  assign n16714 = n16602 | n16713 ;
  assign n16715 = n16602 & n16713 ;
  assign n16716 = n16714 & ~n16715 ;
  assign n16717 = x96 & n6068 ;
  assign n16718 = x95 & n6063 ;
  assign n16719 = x94 & ~n6062 ;
  assign n16720 = n6398 & n16719 ;
  assign n16721 = n16718 | n16720 ;
  assign n16722 = n16717 | n16721 ;
  assign n16723 = n6071 | n16722 ;
  assign n16724 = ( n3509 & n16722 ) | ( n3509 & n16723 ) | ( n16722 & n16723 ) ;
  assign n16725 = x44 & n16724 ;
  assign n16726 = x44 & ~n16725 ;
  assign n16727 = ( n16724 & ~n16725 ) | ( n16724 & n16726 ) | ( ~n16725 & n16726 ) ;
  assign n16728 = n16716 | n16727 ;
  assign n16729 = n16716 & n16727 ;
  assign n16730 = n16728 & ~n16729 ;
  assign n16731 = x99 & n5340 ;
  assign n16732 = x98 & n5335 ;
  assign n16733 = x97 & ~n5334 ;
  assign n16734 = n5580 & n16733 ;
  assign n16735 = n16732 | n16734 ;
  assign n16736 = n16731 | n16735 ;
  assign n16737 = n5343 | n16736 ;
  assign n16738 = ( n4325 & n16736 ) | ( n4325 & n16737 ) | ( n16736 & n16737 ) ;
  assign n16739 = x41 & n16738 ;
  assign n16740 = x41 & ~n16739 ;
  assign n16741 = ( n16738 & ~n16739 ) | ( n16738 & n16740 ) | ( ~n16739 & n16740 ) ;
  assign n16742 = ( n16601 & n16730 ) | ( n16601 & n16741 ) | ( n16730 & n16741 ) ;
  assign n16743 = ( n16730 & n16741 ) | ( n16730 & ~n16742 ) | ( n16741 & ~n16742 ) ;
  assign n16744 = ( n16601 & ~n16742 ) | ( n16601 & n16743 ) | ( ~n16742 & n16743 ) ;
  assign n16745 = n16600 | n16744 ;
  assign n16746 = n16600 & n16744 ;
  assign n16747 = n16745 & ~n16746 ;
  assign n16748 = x102 & n4572 ;
  assign n16749 = x101 & n4567 ;
  assign n16750 = x100 & ~n4566 ;
  assign n16751 = n4828 & n16750 ;
  assign n16752 = n16749 | n16751 ;
  assign n16753 = n16748 | n16752 ;
  assign n16754 = n4575 | n16753 ;
  assign n16755 = ( n5025 & n16753 ) | ( n5025 & n16754 ) | ( n16753 & n16754 ) ;
  assign n16756 = x38 & n16755 ;
  assign n16757 = x38 & ~n16756 ;
  assign n16758 = ( n16755 & ~n16756 ) | ( n16755 & n16757 ) | ( ~n16756 & n16757 ) ;
  assign n16759 = n16747 | n16758 ;
  assign n16760 = n16747 & n16758 ;
  assign n16761 = n16759 & ~n16760 ;
  assign n16762 = x105 & n3913 ;
  assign n16763 = x104 & n3908 ;
  assign n16764 = x103 & ~n3907 ;
  assign n16765 = n4152 & n16764 ;
  assign n16766 = n16763 | n16765 ;
  assign n16767 = n16762 | n16766 ;
  assign n16768 = n3916 | n16767 ;
  assign n16769 = ( n5788 & n16767 ) | ( n5788 & n16768 ) | ( n16767 & n16768 ) ;
  assign n16770 = x35 & n16769 ;
  assign n16771 = x35 & ~n16770 ;
  assign n16772 = ( n16769 & ~n16770 ) | ( n16769 & n16771 ) | ( ~n16770 & n16771 ) ;
  assign n16773 = ( n16599 & n16761 ) | ( n16599 & n16772 ) | ( n16761 & n16772 ) ;
  assign n16774 = ( n16761 & n16772 ) | ( n16761 & ~n16773 ) | ( n16772 & ~n16773 ) ;
  assign n16775 = ( n16599 & ~n16773 ) | ( n16599 & n16774 ) | ( ~n16773 & n16774 ) ;
  assign n16776 = n16598 & ~n16775 ;
  assign n16777 = n16775 | n16776 ;
  assign n16778 = ( ~n16598 & n16776 ) | ( ~n16598 & n16777 ) | ( n16776 & n16777 ) ;
  assign n16779 = x114 & n2280 ;
  assign n16780 = x113 & n2275 ;
  assign n16781 = x112 & ~n2274 ;
  assign n16782 = n2481 & n16781 ;
  assign n16783 = n16780 | n16782 ;
  assign n16784 = n16779 | n16783 ;
  assign n16785 = n2283 | n16784 ;
  assign n16786 = ( n8437 & n16784 ) | ( n8437 & n16785 ) | ( n16784 & n16785 ) ;
  assign n16787 = x26 & n16786 ;
  assign n16788 = x26 & ~n16787 ;
  assign n16789 = ( n16786 & ~n16787 ) | ( n16786 & n16788 ) | ( ~n16787 & n16788 ) ;
  assign n16790 = ( n16144 & n16270 ) | ( n16144 & n16271 ) | ( n16270 & n16271 ) ;
  assign n16791 = n16789 | n16790 ;
  assign n16792 = n16467 | n16791 ;
  assign n16793 = ( n16467 & n16789 ) | ( n16467 & n16790 ) | ( n16789 & n16790 ) ;
  assign n16794 = n16792 & ~n16793 ;
  assign n16795 = ( n16141 & n16452 ) | ( n16141 & n16463 ) | ( n16452 & n16463 ) ;
  assign n16796 = x111 & n2775 ;
  assign n16797 = x110 & n2770 ;
  assign n16798 = x109 & ~n2769 ;
  assign n16799 = n2978 & n16798 ;
  assign n16800 = n16797 | n16799 ;
  assign n16801 = n16796 | n16800 ;
  assign n16802 = n2778 | n16801 ;
  assign n16803 = ( n7492 & n16801 ) | ( n7492 & n16802 ) | ( n16801 & n16802 ) ;
  assign n16804 = x29 & n16803 ;
  assign n16805 = x29 & ~n16804 ;
  assign n16806 = ( n16803 & ~n16804 ) | ( n16803 & n16805 ) | ( ~n16804 & n16805 ) ;
  assign n16807 = n16795 | n16806 ;
  assign n16808 = n16795 & n16806 ;
  assign n16809 = n16807 & ~n16808 ;
  assign n16810 = ( n16778 & n16794 ) | ( n16778 & ~n16809 ) | ( n16794 & ~n16809 ) ;
  assign n16811 = ( ~n16794 & n16809 ) | ( ~n16794 & n16810 ) | ( n16809 & n16810 ) ;
  assign n16812 = ( ~n16778 & n16810 ) | ( ~n16778 & n16811 ) | ( n16810 & n16811 ) ;
  assign n16813 = x117 & n1817 ;
  assign n16814 = x116 & n1812 ;
  assign n16815 = x115 & ~n1811 ;
  assign n16816 = n1977 & n16815 ;
  assign n16817 = n16814 | n16816 ;
  assign n16818 = n16813 | n16817 ;
  assign n16819 = n1820 | n16818 ;
  assign n16820 = ( n9118 & n16818 ) | ( n9118 & n16819 ) | ( n16818 & n16819 ) ;
  assign n16821 = x23 & n16820 ;
  assign n16822 = x23 & ~n16821 ;
  assign n16823 = ( n16820 & ~n16821 ) | ( n16820 & n16822 ) | ( ~n16821 & n16822 ) ;
  assign n16824 = ( n16250 & n16252 ) | ( n16250 & n16256 ) | ( n16252 & n16256 ) ;
  assign n16825 = n16823 & n16824 ;
  assign n16826 = ( n16470 & n16823 ) | ( n16470 & n16825 ) | ( n16823 & n16825 ) ;
  assign n16827 = n16470 | n16824 ;
  assign n16828 = ~n16823 & n16827 ;
  assign n16829 = ( n16823 & ~n16826 ) | ( n16823 & n16828 ) | ( ~n16826 & n16828 ) ;
  assign n16830 = n16812 & n16829 ;
  assign n16831 = n16812 | n16829 ;
  assign n16832 = ~n16830 & n16831 ;
  assign n16833 = n16583 & n16832 ;
  assign n16834 = n16583 | n16832 ;
  assign n16835 = ~n16833 & n16834 ;
  assign n16836 = x126 & n771 ;
  assign n16837 = x125 & n766 ;
  assign n16838 = x124 & ~n765 ;
  assign n16839 = n905 & n16838 ;
  assign n16840 = n16837 | n16839 ;
  assign n16841 = n16836 | n16840 ;
  assign n16842 = n774 | n16841 ;
  assign n16843 = ( n12687 & n16841 ) | ( n12687 & n16842 ) | ( n16841 & n16842 ) ;
  assign n16844 = x14 & n16843 ;
  assign n16845 = x14 & ~n16844 ;
  assign n16846 = ( n16843 & ~n16844 ) | ( n16843 & n16845 ) | ( ~n16844 & n16845 ) ;
  assign n16847 = n16517 | n16846 ;
  assign n16848 = n16520 | n16847 ;
  assign n16849 = ( n16517 & n16520 ) | ( n16517 & n16846 ) | ( n16520 & n16846 ) ;
  assign n16850 = n16848 & ~n16849 ;
  assign n16851 = x123 & n1071 ;
  assign n16852 = x122 & n1066 ;
  assign n16853 = x121 & ~n1065 ;
  assign n16854 = n1189 & n16853 ;
  assign n16855 = n16852 | n16854 ;
  assign n16856 = n16851 | n16855 ;
  assign n16857 = n1074 | n16856 ;
  assign n16858 = ( n11219 & n16856 ) | ( n11219 & n16857 ) | ( n16856 & n16857 ) ;
  assign n16859 = x17 & n16858 ;
  assign n16860 = x17 & ~n16859 ;
  assign n16861 = ( n16858 & ~n16859 ) | ( n16858 & n16860 ) | ( ~n16859 & n16860 ) ;
  assign n16862 = ( n16483 & n16484 ) | ( n16483 & ~n16505 ) | ( n16484 & ~n16505 ) ;
  assign n16863 = n16861 | n16862 ;
  assign n16864 = n16861 & n16862 ;
  assign n16865 = n16863 & ~n16864 ;
  assign n16866 = ( n16835 & n16850 ) | ( n16835 & ~n16865 ) | ( n16850 & ~n16865 ) ;
  assign n16867 = ( ~n16850 & n16865 ) | ( ~n16850 & n16866 ) | ( n16865 & n16866 ) ;
  assign n16868 = ( ~n16835 & n16866 ) | ( ~n16835 & n16867 ) | ( n16866 & n16867 ) ;
  assign n16869 = ( n16566 & ~n16567 ) | ( n16566 & n16868 ) | ( ~n16567 & n16868 ) ;
  assign n16870 = ( n16567 & ~n16868 ) | ( n16567 & n16869 ) | ( ~n16868 & n16869 ) ;
  assign n16871 = ( ~n16566 & n16869 ) | ( ~n16566 & n16870 ) | ( n16869 & n16870 ) ;
  assign n16872 = n16558 & n16871 ;
  assign n16873 = n16558 & ~n16872 ;
  assign n16874 = n16871 & ~n16872 ;
  assign n16875 = n16873 | n16874 ;
  assign n16876 = n16548 | n16551 ;
  assign n16877 = n16875 & n16876 ;
  assign n16878 = n16548 | n16553 ;
  assign n16879 = n16875 & n16878 ;
  assign n16880 = ( n15562 & n16877 ) | ( n15562 & n16879 ) | ( n16877 & n16879 ) ;
  assign n16881 = ( n15562 & n16876 ) | ( n15562 & n16878 ) | ( n16876 & n16878 ) ;
  assign n16882 = ~n16880 & n16881 ;
  assign n16883 = ( n16875 & ~n16880 ) | ( n16875 & n16882 ) | ( ~n16880 & n16882 ) ;
  assign n16884 = ( n16566 & n16567 ) | ( n16566 & n16868 ) | ( n16567 & n16868 ) ;
  assign n16885 = ~n16567 & n16884 ;
  assign n16886 = ( n16868 & ~n16869 ) | ( n16868 & n16885 ) | ( ~n16869 & n16885 ) ;
  assign n16887 = ( n16535 & n16538 ) | ( n16535 & n16566 ) | ( n16538 & n16566 ) ;
  assign n16888 = n16886 | n16887 ;
  assign n16889 = x115 & n2280 ;
  assign n16890 = x114 & n2275 ;
  assign n16891 = x113 & ~n2274 ;
  assign n16892 = n2481 & n16891 ;
  assign n16893 = n16890 | n16892 ;
  assign n16894 = n16889 | n16893 ;
  assign n16895 = n2283 | n16894 ;
  assign n16896 = ( n8749 & n16894 ) | ( n8749 & n16895 ) | ( n16894 & n16895 ) ;
  assign n16897 = x26 & n16896 ;
  assign n16898 = x26 & ~n16897 ;
  assign n16899 = ( n16896 & ~n16897 ) | ( n16896 & n16898 ) | ( ~n16897 & n16898 ) ;
  assign n16900 = n16778 & n16809 ;
  assign n16901 = ( n16778 & n16792 ) | ( n16778 & n16809 ) | ( n16792 & n16809 ) ;
  assign n16902 = ( n16793 & ~n16900 ) | ( n16793 & n16901 ) | ( ~n16900 & n16901 ) ;
  assign n16903 = n16899 | n16902 ;
  assign n16904 = n16899 & n16902 ;
  assign n16905 = n16903 & ~n16904 ;
  assign n16906 = x118 & n1817 ;
  assign n16907 = x117 & n1812 ;
  assign n16908 = x116 & ~n1811 ;
  assign n16909 = n1977 & n16908 ;
  assign n16910 = n16907 | n16909 ;
  assign n16911 = n16906 | n16910 ;
  assign n16912 = n1820 | n16911 ;
  assign n16913 = ( n9760 & n16911 ) | ( n9760 & n16912 ) | ( n16911 & n16912 ) ;
  assign n16914 = x23 & n16913 ;
  assign n16915 = x23 & ~n16914 ;
  assign n16916 = ( n16913 & ~n16914 ) | ( n16913 & n16915 ) | ( ~n16914 & n16915 ) ;
  assign n16917 = n16826 & n16916 ;
  assign n16918 = n16916 & ~n16917 ;
  assign n16919 = ~n16830 & n16918 ;
  assign n16920 = ( n16826 & n16830 ) | ( n16826 & ~n16916 ) | ( n16830 & ~n16916 ) ;
  assign n16921 = n16919 | n16920 ;
  assign n16922 = n16808 | n16900 ;
  assign n16923 = ( n16596 & n16597 ) | ( n16596 & n16775 ) | ( n16597 & n16775 ) ;
  assign n16924 = x109 & n3314 ;
  assign n16925 = x108 & n3309 ;
  assign n16926 = x107 & ~n3308 ;
  assign n16927 = n3570 & n16926 ;
  assign n16928 = n16925 | n16927 ;
  assign n16929 = n16924 | n16928 ;
  assign n16930 = n3317 | n16929 ;
  assign n16931 = ( n6884 & n16929 ) | ( n6884 & n16930 ) | ( n16929 & n16930 ) ;
  assign n16932 = x32 & n16931 ;
  assign n16933 = x32 & ~n16932 ;
  assign n16934 = ( n16931 & ~n16932 ) | ( n16931 & n16933 ) | ( ~n16932 & n16933 ) ;
  assign n16935 = n16923 & n16934 ;
  assign n16936 = n16923 & ~n16935 ;
  assign n16937 = x106 & n3913 ;
  assign n16938 = x105 & n3908 ;
  assign n16939 = x104 & ~n3907 ;
  assign n16940 = n4152 & n16939 ;
  assign n16941 = n16938 | n16940 ;
  assign n16942 = n16937 | n16941 ;
  assign n16943 = n3916 | n16942 ;
  assign n16944 = ( n5814 & n16942 ) | ( n5814 & n16943 ) | ( n16942 & n16943 ) ;
  assign n16945 = x35 & n16944 ;
  assign n16946 = x35 & ~n16945 ;
  assign n16947 = ( n16944 & ~n16945 ) | ( n16944 & n16946 ) | ( ~n16945 & n16946 ) ;
  assign n16948 = x103 & n4572 ;
  assign n16949 = x102 & n4567 ;
  assign n16950 = x101 & ~n4566 ;
  assign n16951 = n4828 & n16950 ;
  assign n16952 = n16949 | n16951 ;
  assign n16953 = n16948 | n16952 ;
  assign n16954 = n4575 | n16953 ;
  assign n16955 = ( n5264 & n16953 ) | ( n5264 & n16954 ) | ( n16953 & n16954 ) ;
  assign n16956 = x38 & n16955 ;
  assign n16957 = x38 & ~n16956 ;
  assign n16958 = ( n16955 & ~n16956 ) | ( n16955 & n16957 ) | ( ~n16956 & n16957 ) ;
  assign n16959 = n16715 | n16729 ;
  assign n16960 = x91 & n7812 ;
  assign n16961 = x90 & n7807 ;
  assign n16962 = x89 & ~n7806 ;
  assign n16963 = n8136 & n16962 ;
  assign n16964 = n16961 | n16963 ;
  assign n16965 = n16960 | n16964 ;
  assign n16966 = n7815 | n16965 ;
  assign n16967 = ( n2714 & n16965 ) | ( n2714 & n16966 ) | ( n16965 & n16966 ) ;
  assign n16968 = x50 & n16967 ;
  assign n16969 = x50 & ~n16968 ;
  assign n16970 = ( n16967 & ~n16968 ) | ( n16967 & n16969 ) | ( ~n16968 & n16969 ) ;
  assign n16971 = x88 & n8834 ;
  assign n16972 = x87 & n8829 ;
  assign n16973 = x86 & ~n8828 ;
  assign n16974 = n9159 & n16973 ;
  assign n16975 = n16972 | n16974 ;
  assign n16976 = n16971 | n16975 ;
  assign n16977 = n8837 | n16976 ;
  assign n16978 = ( n2095 & n16976 ) | ( n2095 & n16977 ) | ( n16976 & n16977 ) ;
  assign n16979 = x53 & n16978 ;
  assign n16980 = x53 & ~n16979 ;
  assign n16981 = ( n16978 & ~n16979 ) | ( n16978 & n16980 ) | ( ~n16979 & n16980 ) ;
  assign n16982 = n16628 | n16642 ;
  assign n16983 = x79 & n11984 ;
  assign n16984 = x78 & n11979 ;
  assign n16985 = x77 & ~n11978 ;
  assign n16986 = n12430 & n16985 ;
  assign n16987 = n16984 | n16986 ;
  assign n16988 = n16983 | n16987 ;
  assign n16989 = n11987 | n16988 ;
  assign n16990 = ( n961 & n16988 ) | ( n961 & n16989 ) | ( n16988 & n16989 ) ;
  assign n16991 = ~x62 & n16990 ;
  assign n16992 = x62 & ~n16990 ;
  assign n16993 = n16991 | n16992 ;
  assign n16994 = x76 & n12808 ;
  assign n16995 = x63 & x75 ;
  assign n16996 = ~n12808 & n16995 ;
  assign n16997 = n16994 | n16996 ;
  assign n16998 = ( x11 & ~n16327 ) | ( x11 & n16997 ) | ( ~n16327 & n16997 ) ;
  assign n16999 = ( ~x11 & n16327 ) | ( ~x11 & n16997 ) | ( n16327 & n16997 ) ;
  assign n17000 = ( ~n16997 & n16998 ) | ( ~n16997 & n16999 ) | ( n16998 & n16999 ) ;
  assign n17001 = n16993 & ~n17000 ;
  assign n17002 = ~n16993 & n17000 ;
  assign n17003 = n17001 | n17002 ;
  assign n17004 = n16620 | n16626 ;
  assign n17005 = ~n17003 & n17004 ;
  assign n17006 = n17003 | n17005 ;
  assign n17007 = n17003 & n17004 ;
  assign n17008 = n17006 & ~n17007 ;
  assign n17009 = x82 & n10876 ;
  assign n17010 = x81 & n10871 ;
  assign n17011 = x80 & ~n10870 ;
  assign n17012 = n11305 & n17011 ;
  assign n17013 = n17010 | n17012 ;
  assign n17014 = n17009 | n17013 ;
  assign n17015 = n10879 | n17014 ;
  assign n17016 = ( n1371 & n17014 ) | ( n1371 & n17015 ) | ( n17014 & n17015 ) ;
  assign n17017 = x59 & n17016 ;
  assign n17018 = x59 & ~n17017 ;
  assign n17019 = ( n17016 & ~n17017 ) | ( n17016 & n17018 ) | ( ~n17017 & n17018 ) ;
  assign n17020 = ~n17008 & n17019 ;
  assign n17021 = n17008 & ~n17019 ;
  assign n17022 = n17020 | n17021 ;
  assign n17023 = ~n16982 & n17022 ;
  assign n17024 = n16982 & ~n17022 ;
  assign n17025 = n17023 | n17024 ;
  assign n17026 = x85 & n9853 ;
  assign n17027 = x84 & n9848 ;
  assign n17028 = x83 & ~n9847 ;
  assign n17029 = n10165 & n17028 ;
  assign n17030 = n17027 | n17029 ;
  assign n17031 = n17026 | n17030 ;
  assign n17032 = n9856 | n17031 ;
  assign n17033 = ( n1765 & n17031 ) | ( n1765 & n17032 ) | ( n17031 & n17032 ) ;
  assign n17034 = x56 & n17033 ;
  assign n17035 = x56 & ~n17034 ;
  assign n17036 = ( n17033 & ~n17034 ) | ( n17033 & n17035 ) | ( ~n17034 & n17035 ) ;
  assign n17037 = ~n17025 & n17036 ;
  assign n17038 = n17025 | n17037 ;
  assign n17039 = n17025 & n17036 ;
  assign n17040 = n16648 & ~n16662 ;
  assign n17041 = ~n17039 & n17040 ;
  assign n17042 = n17038 & n17041 ;
  assign n17043 = ( n17038 & ~n17039 ) | ( n17038 & n17040 ) | ( ~n17039 & n17040 ) ;
  assign n17044 = ~n17042 & n17043 ;
  assign n17045 = n16666 | n16681 ;
  assign n17046 = ( n16981 & n17044 ) | ( n16981 & n17045 ) | ( n17044 & n17045 ) ;
  assign n17047 = ( n17044 & n17045 ) | ( n17044 & ~n17046 ) | ( n17045 & ~n17046 ) ;
  assign n17048 = ( n16981 & ~n17046 ) | ( n16981 & n17047 ) | ( ~n17046 & n17047 ) ;
  assign n17049 = n16970 & n17048 ;
  assign n17050 = n16970 | n17048 ;
  assign n17051 = ~n17049 & n17050 ;
  assign n17052 = n16683 | n16697 ;
  assign n17053 = n17051 | n17052 ;
  assign n17054 = n17051 & n17052 ;
  assign n17055 = n17053 & ~n17054 ;
  assign n17056 = x94 & n6937 ;
  assign n17057 = x93 & n6932 ;
  assign n17058 = x92 & ~n6931 ;
  assign n17059 = n7216 & n17058 ;
  assign n17060 = n17057 | n17059 ;
  assign n17061 = n17056 | n17060 ;
  assign n17062 = n6940 | n17061 ;
  assign n17063 = ( n3271 & n17061 ) | ( n3271 & n17062 ) | ( n17061 & n17062 ) ;
  assign n17064 = x47 & n17063 ;
  assign n17065 = x47 & ~n17064 ;
  assign n17066 = ( n17063 & ~n17064 ) | ( n17063 & n17065 ) | ( ~n17064 & n17065 ) ;
  assign n17067 = n17055 & n17066 ;
  assign n17068 = n17055 | n17066 ;
  assign n17069 = n16711 & n17068 ;
  assign n17070 = ~n17067 & n17069 ;
  assign n17071 = n16711 & ~n17070 ;
  assign n17072 = ( n17055 & n17066 ) | ( n17055 & ~n17069 ) | ( n17066 & ~n17069 ) ;
  assign n17073 = ( ~n17067 & n17071 ) | ( ~n17067 & n17072 ) | ( n17071 & n17072 ) ;
  assign n17074 = x97 & n6068 ;
  assign n17075 = x96 & n6063 ;
  assign n17076 = x95 & ~n6062 ;
  assign n17077 = n6398 & n17076 ;
  assign n17078 = n17075 | n17077 ;
  assign n17079 = n17074 | n17078 ;
  assign n17080 = n6071 | n17079 ;
  assign n17081 = ( n3707 & n17079 ) | ( n3707 & n17080 ) | ( n17079 & n17080 ) ;
  assign n17082 = x44 & n17081 ;
  assign n17083 = x44 & ~n17082 ;
  assign n17084 = ( n17081 & ~n17082 ) | ( n17081 & n17083 ) | ( ~n17082 & n17083 ) ;
  assign n17085 = ( n16959 & n17073 ) | ( n16959 & ~n17084 ) | ( n17073 & ~n17084 ) ;
  assign n17086 = ( ~n17073 & n17084 ) | ( ~n17073 & n17085 ) | ( n17084 & n17085 ) ;
  assign n17087 = ( ~n16959 & n17085 ) | ( ~n16959 & n17086 ) | ( n17085 & n17086 ) ;
  assign n17088 = x100 & n5340 ;
  assign n17089 = x99 & n5335 ;
  assign n17090 = x98 & ~n5334 ;
  assign n17091 = n5580 & n17090 ;
  assign n17092 = n17089 | n17091 ;
  assign n17093 = n17088 | n17092 ;
  assign n17094 = n5343 | n17093 ;
  assign n17095 = ( n4532 & n17093 ) | ( n4532 & n17094 ) | ( n17093 & n17094 ) ;
  assign n17096 = x41 & n17095 ;
  assign n17097 = x41 & ~n17096 ;
  assign n17098 = ( n17095 & ~n17096 ) | ( n17095 & n17097 ) | ( ~n17096 & n17097 ) ;
  assign n17099 = n17087 & n17098 ;
  assign n17100 = n17087 | n17098 ;
  assign n17101 = ~n17099 & n17100 ;
  assign n17102 = n16742 | n17101 ;
  assign n17103 = n16742 & n17101 ;
  assign n17104 = n17102 & ~n17103 ;
  assign n17105 = n16746 | n16760 ;
  assign n17106 = ( n16958 & n17104 ) | ( n16958 & n17105 ) | ( n17104 & n17105 ) ;
  assign n17107 = ( n17104 & n17105 ) | ( n17104 & ~n17106 ) | ( n17105 & ~n17106 ) ;
  assign n17108 = ( n16958 & ~n17106 ) | ( n16958 & n17107 ) | ( ~n17106 & n17107 ) ;
  assign n17109 = n16947 & n17108 ;
  assign n17110 = n16947 | n17108 ;
  assign n17111 = ~n17109 & n17110 ;
  assign n17112 = n16773 | n17111 ;
  assign n17113 = n16773 & n17111 ;
  assign n17114 = n17112 & ~n17113 ;
  assign n17115 = ~n16923 & n16934 ;
  assign n17116 = n17114 | n17115 ;
  assign n17117 = n16936 | n17116 ;
  assign n17118 = ( n16936 & n17114 ) | ( n16936 & n17115 ) | ( n17114 & n17115 ) ;
  assign n17119 = n17117 & ~n17118 ;
  assign n17120 = x112 & n2775 ;
  assign n17121 = x111 & n2770 ;
  assign n17122 = x110 & ~n2769 ;
  assign n17123 = n2978 & n17122 ;
  assign n17124 = n17121 | n17123 ;
  assign n17125 = n17120 | n17124 ;
  assign n17126 = n2778 | n17125 ;
  assign n17127 = ( n7789 & n17125 ) | ( n7789 & n17126 ) | ( n17125 & n17126 ) ;
  assign n17128 = x29 & n17127 ;
  assign n17129 = x29 & ~n17128 ;
  assign n17130 = ( n17127 & ~n17128 ) | ( n17127 & n17129 ) | ( ~n17128 & n17129 ) ;
  assign n17131 = ( n16922 & n17119 ) | ( n16922 & ~n17130 ) | ( n17119 & ~n17130 ) ;
  assign n17132 = ( ~n17119 & n17130 ) | ( ~n17119 & n17131 ) | ( n17130 & n17131 ) ;
  assign n17133 = ( ~n16922 & n17131 ) | ( ~n16922 & n17132 ) | ( n17131 & n17132 ) ;
  assign n17134 = ( n16905 & ~n16921 ) | ( n16905 & n17133 ) | ( ~n16921 & n17133 ) ;
  assign n17135 = ( n16921 & ~n17133 ) | ( n16921 & n17134 ) | ( ~n17133 & n17134 ) ;
  assign n17136 = ( ~n16905 & n17134 ) | ( ~n16905 & n17135 ) | ( n17134 & n17135 ) ;
  assign n17137 = x124 & n1071 ;
  assign n17138 = x123 & n1066 ;
  assign n17139 = x122 & ~n1065 ;
  assign n17140 = n1189 & n17139 ;
  assign n17141 = n17138 | n17140 ;
  assign n17142 = n17137 | n17141 ;
  assign n17143 = n1074 | n17142 ;
  assign n17144 = ( n11916 & n17142 ) | ( n11916 & n17143 ) | ( n17142 & n17143 ) ;
  assign n17145 = x17 & n17144 ;
  assign n17146 = x17 & ~n17145 ;
  assign n17147 = ( n17144 & ~n17145 ) | ( n17144 & n17146 ) | ( ~n17145 & n17146 ) ;
  assign n17148 = ( n16835 & n16861 ) | ( n16835 & n16862 ) | ( n16861 & n16862 ) ;
  assign n17149 = ~n17147 & n17148 ;
  assign n17150 = n17147 & ~n17148 ;
  assign n17151 = n17149 | n17150 ;
  assign n17152 = x121 & n1421 ;
  assign n17153 = x120 & n1416 ;
  assign n17154 = x119 & ~n1415 ;
  assign n17155 = n1584 & n17154 ;
  assign n17156 = n17153 | n17155 ;
  assign n17157 = n17152 | n17156 ;
  assign n17158 = n1424 | n17157 ;
  assign n17159 = ( n10811 & n17157 ) | ( n10811 & n17158 ) | ( n17157 & n17158 ) ;
  assign n17160 = x20 & n17159 ;
  assign n17161 = x20 & ~n17160 ;
  assign n17162 = ( n17159 & ~n17160 ) | ( n17159 & n17161 ) | ( ~n17160 & n17161 ) ;
  assign n17163 = n16580 | n17162 ;
  assign n17164 = n16833 | n17163 ;
  assign n17165 = ( n16580 & n16833 ) | ( n16580 & n17162 ) | ( n16833 & n17162 ) ;
  assign n17166 = n17164 & ~n17165 ;
  assign n17167 = ( n17136 & n17151 ) | ( n17136 & ~n17166 ) | ( n17151 & ~n17166 ) ;
  assign n17168 = ( ~n17151 & n17166 ) | ( ~n17151 & n17167 ) | ( n17166 & n17167 ) ;
  assign n17169 = ( ~n17136 & n17167 ) | ( ~n17136 & n17168 ) | ( n17167 & n17168 ) ;
  assign n17170 = x127 & n771 ;
  assign n17171 = x126 & n766 ;
  assign n17172 = x125 & ~n765 ;
  assign n17173 = n905 & n17172 ;
  assign n17174 = n17171 | n17173 ;
  assign n17175 = n17170 | n17174 ;
  assign n17176 = n774 | n17175 ;
  assign n17177 = ( n12720 & n17175 ) | ( n12720 & n17176 ) | ( n17175 & n17176 ) ;
  assign n17178 = x14 & n17177 ;
  assign n17179 = x14 & ~n17178 ;
  assign n17180 = ( n17177 & ~n17178 ) | ( n17177 & n17179 ) | ( ~n17178 & n17179 ) ;
  assign n17181 = n16850 & ~n16868 ;
  assign n17182 = n16849 | n17181 ;
  assign n17183 = ( n17169 & n17180 ) | ( n17169 & ~n17182 ) | ( n17180 & ~n17182 ) ;
  assign n17184 = ( ~n17180 & n17182 ) | ( ~n17180 & n17183 ) | ( n17182 & n17183 ) ;
  assign n17185 = ( ~n17169 & n17183 ) | ( ~n17169 & n17184 ) | ( n17183 & n17184 ) ;
  assign n17186 = n16887 & n17185 ;
  assign n17187 = ( n16886 & n17185 ) | ( n16886 & n17186 ) | ( n17185 & n17186 ) ;
  assign n17188 = n16888 & ~n17187 ;
  assign n17189 = n16872 | n16877 ;
  assign n17190 = n16872 | n16879 ;
  assign n17191 = ( n15562 & n17189 ) | ( n15562 & n17190 ) | ( n17189 & n17190 ) ;
  assign n17192 = n17185 & ~n17186 ;
  assign n17193 = ~n16886 & n17192 ;
  assign n17194 = n17191 | n17193 ;
  assign n17195 = n17188 | n17194 ;
  assign n17196 = n17188 | n17193 ;
  assign n17197 = n17191 & n17196 ;
  assign n17198 = n17195 & ~n17197 ;
  assign n17199 = ( n17169 & n17180 ) | ( n17169 & n17182 ) | ( n17180 & n17182 ) ;
  assign n17200 = n17136 & n17166 ;
  assign n17201 = n17136 | n17166 ;
  assign n17202 = ~n17200 & n17201 ;
  assign n17203 = ( n17147 & n17148 ) | ( n17147 & n17202 ) | ( n17148 & n17202 ) ;
  assign n17204 = x127 & n766 ;
  assign n17205 = x126 & ~n765 ;
  assign n17206 = n905 & n17205 ;
  assign n17207 = n17204 | n17206 ;
  assign n17208 = n774 | n17207 ;
  assign n17209 = ( n13461 & n17207 ) | ( n13461 & n17208 ) | ( n17207 & n17208 ) ;
  assign n17210 = x14 & n17209 ;
  assign n17211 = x14 & ~n17210 ;
  assign n17212 = ( n17209 & ~n17210 ) | ( n17209 & n17211 ) | ( ~n17210 & n17211 ) ;
  assign n17213 = n17203 & n17212 ;
  assign n17214 = n17203 & ~n17213 ;
  assign n17215 = ~n17203 & n17212 ;
  assign n17216 = n17165 | n17200 ;
  assign n17217 = x125 & n1071 ;
  assign n17218 = x124 & n1066 ;
  assign n17219 = x123 & ~n1065 ;
  assign n17220 = n1189 & n17219 ;
  assign n17221 = n17218 | n17220 ;
  assign n17222 = n17217 | n17221 ;
  assign n17223 = n1074 | n17222 ;
  assign n17224 = ( n12310 & n17222 ) | ( n12310 & n17223 ) | ( n17222 & n17223 ) ;
  assign n17225 = x17 & n17224 ;
  assign n17226 = x17 & ~n17225 ;
  assign n17227 = ( n17224 & ~n17225 ) | ( n17224 & n17226 ) | ( ~n17225 & n17226 ) ;
  assign n17228 = n17216 & n17227 ;
  assign n17229 = n17216 & ~n17228 ;
  assign n17230 = ~n17216 & n17227 ;
  assign n17231 = n17229 | n17230 ;
  assign n17232 = ( n16830 & n16916 ) | ( n16830 & n16917 ) | ( n16916 & n16917 ) ;
  assign n17233 = n16905 & n17133 ;
  assign n17234 = ~n17232 & n17233 ;
  assign n17235 = n16905 | n17133 ;
  assign n17236 = ( n16919 & n16920 ) | ( n16919 & n17235 ) | ( n16920 & n17235 ) ;
  assign n17237 = ( n17232 & ~n17234 ) | ( n17232 & n17236 ) | ( ~n17234 & n17236 ) ;
  assign n17238 = x122 & n1421 ;
  assign n17239 = x121 & n1416 ;
  assign n17240 = x120 & ~n1415 ;
  assign n17241 = n1584 & n17240 ;
  assign n17242 = n17239 | n17241 ;
  assign n17243 = n17238 | n17242 ;
  assign n17244 = n1424 | n17243 ;
  assign n17245 = ( n11188 & n17243 ) | ( n11188 & n17244 ) | ( n17243 & n17244 ) ;
  assign n17246 = x20 & n17245 ;
  assign n17247 = x20 & ~n17246 ;
  assign n17248 = ( n17245 & ~n17246 ) | ( n17245 & n17247 ) | ( ~n17246 & n17247 ) ;
  assign n17249 = n17237 & n17248 ;
  assign n17250 = n17237 | n17248 ;
  assign n17251 = ~n17249 & n17250 ;
  assign n17252 = n16904 | n17233 ;
  assign n17253 = x119 & n1817 ;
  assign n17254 = x118 & n1812 ;
  assign n17255 = x117 & ~n1811 ;
  assign n17256 = n1977 & n17255 ;
  assign n17257 = n17254 | n17256 ;
  assign n17258 = n17253 | n17257 ;
  assign n17259 = n1820 | n17258 ;
  assign n17260 = ( n9789 & n17258 ) | ( n9789 & n17259 ) | ( n17258 & n17259 ) ;
  assign n17261 = x23 & n17260 ;
  assign n17262 = x23 & ~n17261 ;
  assign n17263 = ( n17260 & ~n17261 ) | ( n17260 & n17262 ) | ( ~n17261 & n17262 ) ;
  assign n17264 = n17252 & n17263 ;
  assign n17265 = n17252 & ~n17264 ;
  assign n17266 = ~n17252 & n17263 ;
  assign n17267 = n17265 | n17266 ;
  assign n17268 = x113 & n2775 ;
  assign n17269 = x112 & n2770 ;
  assign n17270 = x111 & ~n2769 ;
  assign n17271 = n2978 & n17270 ;
  assign n17272 = n17269 | n17271 ;
  assign n17273 = n17268 | n17272 ;
  assign n17274 = n2778 | n17273 ;
  assign n17275 = ( n8113 & n17273 ) | ( n8113 & n17274 ) | ( n17273 & n17274 ) ;
  assign n17276 = x29 & n17275 ;
  assign n17277 = x29 & ~n17276 ;
  assign n17278 = ( n17275 & ~n17276 ) | ( n17275 & n17277 ) | ( ~n17276 & n17277 ) ;
  assign n17279 = n16935 & n17278 ;
  assign n17280 = n17278 & ~n17279 ;
  assign n17281 = ~n17118 & n17280 ;
  assign n17282 = ( n16935 & n17118 ) | ( n16935 & ~n17278 ) | ( n17118 & ~n17278 ) ;
  assign n17283 = n17281 | n17282 ;
  assign n17284 = x104 & n4572 ;
  assign n17285 = x103 & n4567 ;
  assign n17286 = x102 & ~n4566 ;
  assign n17287 = n4828 & n17286 ;
  assign n17288 = n17285 | n17287 ;
  assign n17289 = n17284 | n17288 ;
  assign n17290 = n4575 | n17289 ;
  assign n17291 = ( n5295 & n17289 ) | ( n5295 & n17290 ) | ( n17289 & n17290 ) ;
  assign n17292 = x38 & n17291 ;
  assign n17293 = x38 & ~n17292 ;
  assign n17294 = ( n17291 & ~n17292 ) | ( n17291 & n17293 ) | ( ~n17292 & n17293 ) ;
  assign n17295 = ( n16959 & n17073 ) | ( n16959 & n17084 ) | ( n17073 & n17084 ) ;
  assign n17296 = n17067 | n17070 ;
  assign n17297 = n17049 | n17054 ;
  assign n17298 = x89 & n8834 ;
  assign n17299 = x88 & n8829 ;
  assign n17300 = x87 & ~n8828 ;
  assign n17301 = n9159 & n17300 ;
  assign n17302 = n17299 | n17301 ;
  assign n17303 = n17298 | n17302 ;
  assign n17304 = n8837 | n17303 ;
  assign n17305 = ( n2244 & n17303 ) | ( n2244 & n17304 ) | ( n17303 & n17304 ) ;
  assign n17306 = x53 & n17305 ;
  assign n17307 = x53 & ~n17306 ;
  assign n17308 = ( n17305 & ~n17306 ) | ( n17305 & n17307 ) | ( ~n17306 & n17307 ) ;
  assign n17309 = n17001 | n17005 ;
  assign n17310 = x80 & n11984 ;
  assign n17311 = x79 & n11979 ;
  assign n17312 = x78 & ~n11978 ;
  assign n17313 = n12430 & n17312 ;
  assign n17314 = n17311 | n17313 ;
  assign n17315 = n17310 | n17314 ;
  assign n17316 = n11987 | n17315 ;
  assign n17317 = ( n1147 & n17315 ) | ( n1147 & n17316 ) | ( n17315 & n17316 ) ;
  assign n17318 = ~x62 & n17317 ;
  assign n17319 = x62 & ~n17317 ;
  assign n17320 = n17318 | n17319 ;
  assign n17321 = x77 & n12808 ;
  assign n17322 = x63 & x76 ;
  assign n17323 = ~n12808 & n17322 ;
  assign n17324 = n17321 | n17323 ;
  assign n17325 = ( n16999 & n17320 ) | ( n16999 & ~n17324 ) | ( n17320 & ~n17324 ) ;
  assign n17326 = ( ~n17320 & n17324 ) | ( ~n17320 & n17325 ) | ( n17324 & n17325 ) ;
  assign n17327 = ( ~n16999 & n17325 ) | ( ~n16999 & n17326 ) | ( n17325 & n17326 ) ;
  assign n17328 = ~n17309 & n17327 ;
  assign n17329 = n17309 & ~n17327 ;
  assign n17330 = n17328 | n17329 ;
  assign n17331 = x83 & n10876 ;
  assign n17332 = x82 & n10871 ;
  assign n17333 = x81 & ~n10870 ;
  assign n17334 = n11305 & n17333 ;
  assign n17335 = n17332 | n17334 ;
  assign n17336 = n17331 | n17335 ;
  assign n17337 = n10879 | n17336 ;
  assign n17338 = ( n1510 & n17336 ) | ( n1510 & n17337 ) | ( n17336 & n17337 ) ;
  assign n17339 = x59 & n17338 ;
  assign n17340 = x59 & ~n17339 ;
  assign n17341 = ( n17338 & ~n17339 ) | ( n17338 & n17340 ) | ( ~n17339 & n17340 ) ;
  assign n17342 = n17330 & n17341 ;
  assign n17343 = ( n17309 & ~n17327 ) | ( n17309 & n17341 ) | ( ~n17327 & n17341 ) ;
  assign n17344 = n17328 | n17343 ;
  assign n17345 = ~n17342 & n17344 ;
  assign n17346 = n17020 | n17024 ;
  assign n17347 = n17345 & ~n17346 ;
  assign n17348 = ~n17345 & n17346 ;
  assign n17349 = n17347 | n17348 ;
  assign n17350 = x86 & n9853 ;
  assign n17351 = x85 & n9848 ;
  assign n17352 = x84 & ~n9847 ;
  assign n17353 = n10165 & n17352 ;
  assign n17354 = n17351 | n17353 ;
  assign n17355 = n17350 | n17354 ;
  assign n17356 = n9856 | n17355 ;
  assign n17357 = ( n1921 & n17355 ) | ( n1921 & n17356 ) | ( n17355 & n17356 ) ;
  assign n17358 = x56 & n17357 ;
  assign n17359 = x56 & ~n17358 ;
  assign n17360 = ( n17357 & ~n17358 ) | ( n17357 & n17359 ) | ( ~n17358 & n17359 ) ;
  assign n17361 = n17349 & n17360 ;
  assign n17362 = ( ~n17345 & n17346 ) | ( ~n17345 & n17360 ) | ( n17346 & n17360 ) ;
  assign n17363 = n17347 | n17362 ;
  assign n17364 = ~n17361 & n17363 ;
  assign n17365 = ~n17037 & n17043 ;
  assign n17366 = ( n17308 & n17364 ) | ( n17308 & ~n17365 ) | ( n17364 & ~n17365 ) ;
  assign n17367 = ( ~n17364 & n17365 ) | ( ~n17364 & n17366 ) | ( n17365 & n17366 ) ;
  assign n17368 = ( ~n17308 & n17366 ) | ( ~n17308 & n17367 ) | ( n17366 & n17367 ) ;
  assign n17369 = n17046 | n17368 ;
  assign n17370 = n17046 & n17368 ;
  assign n17371 = n17369 & ~n17370 ;
  assign n17372 = x92 & n7812 ;
  assign n17373 = x91 & n7807 ;
  assign n17374 = x90 & ~n7806 ;
  assign n17375 = n8136 & n17374 ;
  assign n17376 = n17373 | n17375 ;
  assign n17377 = n17372 | n17376 ;
  assign n17378 = n7815 | n17377 ;
  assign n17379 = ( n2904 & n17377 ) | ( n2904 & n17378 ) | ( n17377 & n17378 ) ;
  assign n17380 = x50 & n17379 ;
  assign n17381 = x50 & ~n17380 ;
  assign n17382 = ( n17379 & ~n17380 ) | ( n17379 & n17381 ) | ( ~n17380 & n17381 ) ;
  assign n17383 = n17371 | n17382 ;
  assign n17384 = n17371 & n17382 ;
  assign n17385 = n17383 & ~n17384 ;
  assign n17386 = x95 & n6937 ;
  assign n17387 = x94 & n6932 ;
  assign n17388 = x93 & ~n6931 ;
  assign n17389 = n7216 & n17388 ;
  assign n17390 = n17387 | n17389 ;
  assign n17391 = n17386 | n17390 ;
  assign n17392 = n6940 | n17391 ;
  assign n17393 = ( n3479 & n17391 ) | ( n3479 & n17392 ) | ( n17391 & n17392 ) ;
  assign n17394 = x47 & n17393 ;
  assign n17395 = x47 & ~n17394 ;
  assign n17396 = ( n17393 & ~n17394 ) | ( n17393 & n17395 ) | ( ~n17394 & n17395 ) ;
  assign n17397 = ( n17297 & ~n17385 ) | ( n17297 & n17396 ) | ( ~n17385 & n17396 ) ;
  assign n17398 = ( n17385 & ~n17396 ) | ( n17385 & n17397 ) | ( ~n17396 & n17397 ) ;
  assign n17399 = ( ~n17297 & n17397 ) | ( ~n17297 & n17398 ) | ( n17397 & n17398 ) ;
  assign n17400 = n17296 & n17399 ;
  assign n17401 = n17296 | n17399 ;
  assign n17402 = ~n17400 & n17401 ;
  assign n17403 = x98 & n6068 ;
  assign n17404 = x97 & n6063 ;
  assign n17405 = x96 & ~n6062 ;
  assign n17406 = n6398 & n17405 ;
  assign n17407 = n17404 | n17406 ;
  assign n17408 = n17403 | n17407 ;
  assign n17409 = n6071 | n17408 ;
  assign n17410 = ( n4105 & n17408 ) | ( n4105 & n17409 ) | ( n17408 & n17409 ) ;
  assign n17411 = x44 & n17410 ;
  assign n17412 = x44 & ~n17411 ;
  assign n17413 = ( n17410 & ~n17411 ) | ( n17410 & n17412 ) | ( ~n17411 & n17412 ) ;
  assign n17414 = n17402 & n17413 ;
  assign n17415 = n17402 | n17413 ;
  assign n17416 = ~n17414 & n17415 ;
  assign n17417 = n17295 & n17416 ;
  assign n17418 = n17295 & ~n17417 ;
  assign n17419 = x101 & n5340 ;
  assign n17420 = x100 & n5335 ;
  assign n17421 = x99 & ~n5334 ;
  assign n17422 = n5580 & n17421 ;
  assign n17423 = n17420 | n17422 ;
  assign n17424 = n17419 | n17423 ;
  assign n17425 = n5343 | n17424 ;
  assign n17426 = ( n4783 & n17424 ) | ( n4783 & n17425 ) | ( n17424 & n17425 ) ;
  assign n17427 = x41 & n17426 ;
  assign n17428 = x41 & ~n17427 ;
  assign n17429 = ( n17426 & ~n17427 ) | ( n17426 & n17428 ) | ( ~n17427 & n17428 ) ;
  assign n17430 = n17416 & ~n17417 ;
  assign n17431 = n17429 | n17430 ;
  assign n17432 = n17418 | n17431 ;
  assign n17433 = ( n17418 & n17429 ) | ( n17418 & n17430 ) | ( n17429 & n17430 ) ;
  assign n17434 = n17432 & ~n17433 ;
  assign n17435 = n17099 | n17103 ;
  assign n17436 = n17434 & n17435 ;
  assign n17437 = n17435 & ~n17436 ;
  assign n17438 = ( n17434 & ~n17436 ) | ( n17434 & n17437 ) | ( ~n17436 & n17437 ) ;
  assign n17439 = n17294 & n17438 ;
  assign n17440 = n17294 | n17438 ;
  assign n17441 = ~n17439 & n17440 ;
  assign n17442 = x107 & n3913 ;
  assign n17443 = x106 & n3908 ;
  assign n17444 = x105 & ~n3907 ;
  assign n17445 = n4152 & n17444 ;
  assign n17446 = n17443 | n17445 ;
  assign n17447 = n17442 | n17446 ;
  assign n17448 = n3916 | n17447 ;
  assign n17449 = ( n6328 & n17447 ) | ( n6328 & n17448 ) | ( n17447 & n17448 ) ;
  assign n17450 = x35 & n17449 ;
  assign n17451 = x35 & ~n17450 ;
  assign n17452 = ( n17449 & ~n17450 ) | ( n17449 & n17451 ) | ( ~n17450 & n17451 ) ;
  assign n17453 = ( n17106 & n17441 ) | ( n17106 & n17452 ) | ( n17441 & n17452 ) ;
  assign n17454 = ( n17441 & n17452 ) | ( n17441 & ~n17453 ) | ( n17452 & ~n17453 ) ;
  assign n17455 = ( n17106 & ~n17453 ) | ( n17106 & n17454 ) | ( ~n17453 & n17454 ) ;
  assign n17456 = n17109 | n17113 ;
  assign n17457 = x110 & n3314 ;
  assign n17458 = x109 & n3309 ;
  assign n17459 = x108 & ~n3308 ;
  assign n17460 = n3570 & n17459 ;
  assign n17461 = n17458 | n17460 ;
  assign n17462 = n17457 | n17461 ;
  assign n17463 = n3317 | n17462 ;
  assign n17464 = ( n7189 & n17462 ) | ( n7189 & n17463 ) | ( n17462 & n17463 ) ;
  assign n17465 = x32 & n17464 ;
  assign n17466 = x32 & ~n17465 ;
  assign n17467 = ( n17464 & ~n17465 ) | ( n17464 & n17466 ) | ( ~n17465 & n17466 ) ;
  assign n17468 = ( n17455 & n17456 ) | ( n17455 & ~n17467 ) | ( n17456 & ~n17467 ) ;
  assign n17469 = ( ~n17456 & n17467 ) | ( ~n17456 & n17468 ) | ( n17467 & n17468 ) ;
  assign n17470 = ( ~n17455 & n17468 ) | ( ~n17455 & n17469 ) | ( n17468 & n17469 ) ;
  assign n17471 = n17283 & n17470 ;
  assign n17472 = n17283 | n17470 ;
  assign n17473 = ~n17471 & n17472 ;
  assign n17474 = x116 & n2280 ;
  assign n17475 = x115 & n2275 ;
  assign n17476 = x114 & ~n2274 ;
  assign n17477 = n2481 & n17476 ;
  assign n17478 = n17475 | n17477 ;
  assign n17479 = n17474 | n17478 ;
  assign n17480 = n2283 | n17479 ;
  assign n17481 = ( n8778 & n17479 ) | ( n8778 & n17480 ) | ( n17479 & n17480 ) ;
  assign n17482 = x26 & n17481 ;
  assign n17483 = x26 & ~n17482 ;
  assign n17484 = ( n17481 & ~n17482 ) | ( n17481 & n17483 ) | ( ~n17482 & n17483 ) ;
  assign n17485 = ( n16922 & n17119 ) | ( n16922 & n17130 ) | ( n17119 & n17130 ) ;
  assign n17486 = ( n17473 & n17484 ) | ( n17473 & ~n17485 ) | ( n17484 & ~n17485 ) ;
  assign n17487 = ( ~n17484 & n17485 ) | ( ~n17484 & n17486 ) | ( n17485 & n17486 ) ;
  assign n17488 = ( ~n17473 & n17486 ) | ( ~n17473 & n17487 ) | ( n17486 & n17487 ) ;
  assign n17489 = n17267 & n17488 ;
  assign n17490 = n17267 | n17488 ;
  assign n17491 = ~n17489 & n17490 ;
  assign n17492 = ~n17251 & n17491 ;
  assign n17493 = n17251 & ~n17491 ;
  assign n17494 = n17492 | n17493 ;
  assign n17495 = n17231 & n17494 ;
  assign n17496 = n17231 | n17494 ;
  assign n17497 = ~n17495 & n17496 ;
  assign n17498 = n17215 | n17497 ;
  assign n17499 = n17214 | n17498 ;
  assign n17500 = ( n17214 & n17215 ) | ( n17214 & n17497 ) | ( n17215 & n17497 ) ;
  assign n17501 = n17499 & ~n17500 ;
  assign n17502 = n17199 & n17501 ;
  assign n17503 = n17199 & ~n17502 ;
  assign n17504 = ~n17199 & n17501 ;
  assign n17505 = n17503 | n17504 ;
  assign n17506 = n17187 | n17197 ;
  assign n17507 = n17505 | n17506 ;
  assign n17508 = ~n17506 & n17507 ;
  assign n17509 = ( ~n17505 & n17507 ) | ( ~n17505 & n17508 ) | ( n17507 & n17508 ) ;
  assign n17510 = x127 & ~n765 ;
  assign n17511 = n905 & n17510 ;
  assign n17512 = ( x127 & n774 ) | ( x127 & n17511 ) | ( n774 & n17511 ) ;
  assign n17513 = ( x126 & n17511 ) | ( x126 & n17512 ) | ( n17511 & n17512 ) ;
  assign n17514 = ( n12685 & n17512 ) | ( n12685 & n17513 ) | ( n17512 & n17513 ) ;
  assign n17515 = x14 & n17514 ;
  assign n17516 = x14 & ~n17515 ;
  assign n17517 = ( n17514 & ~n17515 ) | ( n17514 & n17516 ) | ( ~n17515 & n17516 ) ;
  assign n17518 = n17228 & n17517 ;
  assign n17519 = n17517 & ~n17518 ;
  assign n17520 = ~n17495 & n17519 ;
  assign n17521 = x117 & n2280 ;
  assign n17522 = x116 & n2275 ;
  assign n17523 = x115 & ~n2274 ;
  assign n17524 = n2481 & n17523 ;
  assign n17525 = n17522 | n17524 ;
  assign n17526 = n17521 | n17525 ;
  assign n17527 = n2283 | n17526 ;
  assign n17528 = ( n9118 & n17526 ) | ( n9118 & n17527 ) | ( n17526 & n17527 ) ;
  assign n17529 = x26 & n17528 ;
  assign n17530 = x26 & ~n17529 ;
  assign n17531 = ( n17528 & ~n17529 ) | ( n17528 & n17530 ) | ( ~n17529 & n17530 ) ;
  assign n17532 = ( n17118 & n17278 ) | ( n17118 & n17279 ) | ( n17278 & n17279 ) ;
  assign n17533 = n17531 & n17532 ;
  assign n17534 = ( n17471 & n17531 ) | ( n17471 & n17533 ) | ( n17531 & n17533 ) ;
  assign n17535 = n17531 | n17532 ;
  assign n17536 = n17471 | n17535 ;
  assign n17537 = ~n17534 & n17536 ;
  assign n17538 = n17400 | n17414 ;
  assign n17539 = x99 & n6068 ;
  assign n17540 = x98 & n6063 ;
  assign n17541 = x97 & ~n6062 ;
  assign n17542 = n6398 & n17541 ;
  assign n17543 = n17540 | n17542 ;
  assign n17544 = n17539 | n17543 ;
  assign n17545 = n6071 | n17544 ;
  assign n17546 = ( n4325 & n17544 ) | ( n4325 & n17545 ) | ( n17544 & n17545 ) ;
  assign n17547 = x44 & n17546 ;
  assign n17548 = x44 & ~n17547 ;
  assign n17549 = ( n17546 & ~n17547 ) | ( n17546 & n17548 ) | ( ~n17547 & n17548 ) ;
  assign n17550 = ( ~n17308 & n17364 ) | ( ~n17308 & n17365 ) | ( n17364 & n17365 ) ;
  assign n17551 = x84 & n10876 ;
  assign n17552 = x83 & n10871 ;
  assign n17553 = x82 & ~n10870 ;
  assign n17554 = n11305 & n17553 ;
  assign n17555 = n17552 | n17554 ;
  assign n17556 = n17551 | n17555 ;
  assign n17557 = n10879 | n17556 ;
  assign n17558 = ( n1537 & n17556 ) | ( n1537 & n17557 ) | ( n17556 & n17557 ) ;
  assign n17559 = x59 & n17558 ;
  assign n17560 = x59 & ~n17559 ;
  assign n17561 = ( n17558 & ~n17559 ) | ( n17558 & n17560 ) | ( ~n17559 & n17560 ) ;
  assign n17562 = x78 & n12808 ;
  assign n17563 = x63 & x77 ;
  assign n17564 = ~n12808 & n17563 ;
  assign n17565 = n17562 | n17564 ;
  assign n17566 = ~n17324 & n17565 ;
  assign n17567 = n17324 & ~n17565 ;
  assign n17568 = n17566 | n17567 ;
  assign n17569 = x81 & n11984 ;
  assign n17570 = x80 & n11979 ;
  assign n17571 = x79 & ~n11978 ;
  assign n17572 = n12430 & n17571 ;
  assign n17573 = n17570 | n17572 ;
  assign n17574 = n17569 | n17573 ;
  assign n17575 = n11987 | n17574 ;
  assign n17576 = ( n1256 & n17574 ) | ( n1256 & n17575 ) | ( n17574 & n17575 ) ;
  assign n17577 = x62 & n17576 ;
  assign n17578 = x62 & ~n17577 ;
  assign n17579 = ( n17576 & ~n17577 ) | ( n17576 & n17578 ) | ( ~n17577 & n17578 ) ;
  assign n17580 = ~n17568 & n17579 ;
  assign n17581 = n17568 & ~n17579 ;
  assign n17582 = n17580 | n17581 ;
  assign n17583 = ( ~n17325 & n17561 ) | ( ~n17325 & n17582 ) | ( n17561 & n17582 ) ;
  assign n17584 = ( n17325 & ~n17582 ) | ( n17325 & n17583 ) | ( ~n17582 & n17583 ) ;
  assign n17585 = ( ~n17561 & n17583 ) | ( ~n17561 & n17584 ) | ( n17583 & n17584 ) ;
  assign n17586 = ~n17343 & n17585 ;
  assign n17587 = n17343 & ~n17585 ;
  assign n17588 = n17586 | n17587 ;
  assign n17589 = x87 & n9853 ;
  assign n17590 = x86 & n9848 ;
  assign n17591 = x85 & ~n9847 ;
  assign n17592 = n10165 & n17591 ;
  assign n17593 = n17590 | n17592 ;
  assign n17594 = n17589 | n17593 ;
  assign n17595 = n9856 | n17594 ;
  assign n17596 = ( n2067 & n17594 ) | ( n2067 & n17595 ) | ( n17594 & n17595 ) ;
  assign n17597 = x56 & n17596 ;
  assign n17598 = x56 & ~n17597 ;
  assign n17599 = ( n17596 & ~n17597 ) | ( n17596 & n17598 ) | ( ~n17597 & n17598 ) ;
  assign n17600 = n17588 & ~n17599 ;
  assign n17601 = ~n17588 & n17599 ;
  assign n17602 = n17600 | n17601 ;
  assign n17603 = n17362 & ~n17602 ;
  assign n17604 = ~n17362 & n17602 ;
  assign n17605 = n17603 | n17604 ;
  assign n17606 = x90 & n8834 ;
  assign n17607 = x89 & n8829 ;
  assign n17608 = x88 & ~n8828 ;
  assign n17609 = n9159 & n17608 ;
  assign n17610 = n17607 | n17609 ;
  assign n17611 = n17606 | n17610 ;
  assign n17612 = n8837 | n17611 ;
  assign n17613 = ( n2410 & n17611 ) | ( n2410 & n17612 ) | ( n17611 & n17612 ) ;
  assign n17614 = x53 & n17613 ;
  assign n17615 = x53 & ~n17614 ;
  assign n17616 = ( n17613 & ~n17614 ) | ( n17613 & n17615 ) | ( ~n17614 & n17615 ) ;
  assign n17617 = ~n17605 & n17616 ;
  assign n17618 = n17605 & ~n17616 ;
  assign n17619 = n17617 | n17618 ;
  assign n17620 = n17550 | n17619 ;
  assign n17621 = n17550 & n17619 ;
  assign n17622 = n17620 & ~n17621 ;
  assign n17623 = x93 & n7812 ;
  assign n17624 = x92 & n7807 ;
  assign n17625 = x91 & ~n7806 ;
  assign n17626 = n8136 & n17625 ;
  assign n17627 = n17624 | n17626 ;
  assign n17628 = n17623 | n17627 ;
  assign n17629 = n7815 | n17628 ;
  assign n17630 = ( n2931 & n17628 ) | ( n2931 & n17629 ) | ( n17628 & n17629 ) ;
  assign n17631 = x50 & n17630 ;
  assign n17632 = x50 & ~n17631 ;
  assign n17633 = ( n17630 & ~n17631 ) | ( n17630 & n17632 ) | ( ~n17631 & n17632 ) ;
  assign n17634 = n17622 & ~n17633 ;
  assign n17635 = n17633 | n17634 ;
  assign n17636 = ( ~n17622 & n17634 ) | ( ~n17622 & n17635 ) | ( n17634 & n17635 ) ;
  assign n17637 = n17370 | n17384 ;
  assign n17638 = n17636 & n17637 ;
  assign n17639 = n17636 & ~n17638 ;
  assign n17640 = n17637 & ~n17638 ;
  assign n17641 = n17639 | n17640 ;
  assign n17642 = x96 & n6937 ;
  assign n17643 = x95 & n6932 ;
  assign n17644 = x94 & ~n6931 ;
  assign n17645 = n7216 & n17644 ;
  assign n17646 = n17643 | n17645 ;
  assign n17647 = n17642 | n17646 ;
  assign n17648 = n6940 | n17647 ;
  assign n17649 = ( n3509 & n17647 ) | ( n3509 & n17648 ) | ( n17647 & n17648 ) ;
  assign n17650 = x47 & n17649 ;
  assign n17651 = x47 & ~n17650 ;
  assign n17652 = ( n17649 & ~n17650 ) | ( n17649 & n17651 ) | ( ~n17650 & n17651 ) ;
  assign n17653 = n17641 & ~n17652 ;
  assign n17654 = ~n17641 & n17652 ;
  assign n17655 = n17653 | n17654 ;
  assign n17656 = ( n17297 & n17385 ) | ( n17297 & n17396 ) | ( n17385 & n17396 ) ;
  assign n17657 = ( n17549 & n17655 ) | ( n17549 & ~n17656 ) | ( n17655 & ~n17656 ) ;
  assign n17658 = ( ~n17655 & n17656 ) | ( ~n17655 & n17657 ) | ( n17656 & n17657 ) ;
  assign n17659 = ( ~n17549 & n17657 ) | ( ~n17549 & n17658 ) | ( n17657 & n17658 ) ;
  assign n17660 = n17538 | n17659 ;
  assign n17661 = n17538 & n17659 ;
  assign n17662 = n17660 & ~n17661 ;
  assign n17663 = x102 & n5340 ;
  assign n17664 = x101 & n5335 ;
  assign n17665 = x100 & ~n5334 ;
  assign n17666 = n5580 & n17665 ;
  assign n17667 = n17664 | n17666 ;
  assign n17668 = n17663 | n17667 ;
  assign n17669 = n5343 | n17668 ;
  assign n17670 = ( n5025 & n17668 ) | ( n5025 & n17669 ) | ( n17668 & n17669 ) ;
  assign n17671 = x41 & n17670 ;
  assign n17672 = x41 & ~n17671 ;
  assign n17673 = ( n17670 & ~n17671 ) | ( n17670 & n17672 ) | ( ~n17671 & n17672 ) ;
  assign n17674 = n17662 | n17673 ;
  assign n17675 = n17662 & n17673 ;
  assign n17676 = n17674 & ~n17675 ;
  assign n17677 = n17417 | n17433 ;
  assign n17678 = n17676 & n17677 ;
  assign n17679 = n17676 | n17677 ;
  assign n17680 = ~n17678 & n17679 ;
  assign n17681 = x105 & n4572 ;
  assign n17682 = x104 & n4567 ;
  assign n17683 = x103 & ~n4566 ;
  assign n17684 = n4828 & n17683 ;
  assign n17685 = n17682 | n17684 ;
  assign n17686 = n17681 | n17685 ;
  assign n17687 = n4575 | n17686 ;
  assign n17688 = ( n5788 & n17686 ) | ( n5788 & n17687 ) | ( n17686 & n17687 ) ;
  assign n17689 = x38 & n17688 ;
  assign n17690 = x38 & ~n17689 ;
  assign n17691 = ( n17688 & ~n17689 ) | ( n17688 & n17690 ) | ( ~n17689 & n17690 ) ;
  assign n17692 = n17680 & n17691 ;
  assign n17693 = n17680 | n17691 ;
  assign n17694 = ~n17692 & n17693 ;
  assign n17695 = n17436 | n17439 ;
  assign n17696 = n17694 & n17695 ;
  assign n17697 = n17694 | n17695 ;
  assign n17698 = ~n17696 & n17697 ;
  assign n17699 = x108 & n3913 ;
  assign n17700 = x107 & n3908 ;
  assign n17701 = x106 & ~n3907 ;
  assign n17702 = n4152 & n17701 ;
  assign n17703 = n17700 | n17702 ;
  assign n17704 = n17699 | n17703 ;
  assign n17705 = n3916 | n17704 ;
  assign n17706 = ( n6358 & n17704 ) | ( n6358 & n17705 ) | ( n17704 & n17705 ) ;
  assign n17707 = x35 & n17706 ;
  assign n17708 = x35 & ~n17707 ;
  assign n17709 = ( n17706 & ~n17707 ) | ( n17706 & n17708 ) | ( ~n17707 & n17708 ) ;
  assign n17710 = n17698 & n17709 ;
  assign n17711 = n17698 & ~n17710 ;
  assign n17712 = ~n17698 & n17709 ;
  assign n17713 = n17711 | n17712 ;
  assign n17714 = x111 & n3314 ;
  assign n17715 = x110 & n3309 ;
  assign n17716 = x109 & ~n3308 ;
  assign n17717 = n3570 & n17716 ;
  assign n17718 = n17715 | n17717 ;
  assign n17719 = n17714 | n17718 ;
  assign n17720 = n3317 | n17719 ;
  assign n17721 = ( n7492 & n17719 ) | ( n7492 & n17720 ) | ( n17719 & n17720 ) ;
  assign n17722 = x32 & n17721 ;
  assign n17723 = x32 & ~n17722 ;
  assign n17724 = ( n17721 & ~n17722 ) | ( n17721 & n17723 ) | ( ~n17722 & n17723 ) ;
  assign n17725 = ( ~n17453 & n17713 ) | ( ~n17453 & n17724 ) | ( n17713 & n17724 ) ;
  assign n17726 = ( n17453 & ~n17724 ) | ( n17453 & n17725 ) | ( ~n17724 & n17725 ) ;
  assign n17727 = ( ~n17713 & n17725 ) | ( ~n17713 & n17726 ) | ( n17725 & n17726 ) ;
  assign n17728 = x114 & n2775 ;
  assign n17729 = x113 & n2770 ;
  assign n17730 = x112 & ~n2769 ;
  assign n17731 = n2978 & n17730 ;
  assign n17732 = n17729 | n17731 ;
  assign n17733 = n17728 | n17732 ;
  assign n17734 = n2778 | n17733 ;
  assign n17735 = ( n8437 & n17733 ) | ( n8437 & n17734 ) | ( n17733 & n17734 ) ;
  assign n17736 = x29 & n17735 ;
  assign n17737 = x29 & ~n17736 ;
  assign n17738 = ( n17735 & ~n17736 ) | ( n17735 & n17737 ) | ( ~n17736 & n17737 ) ;
  assign n17739 = ( n17455 & n17456 ) | ( n17455 & n17467 ) | ( n17456 & n17467 ) ;
  assign n17740 = ( n17727 & n17738 ) | ( n17727 & ~n17739 ) | ( n17738 & ~n17739 ) ;
  assign n17741 = ( ~n17738 & n17739 ) | ( ~n17738 & n17740 ) | ( n17739 & n17740 ) ;
  assign n17742 = ( ~n17727 & n17740 ) | ( ~n17727 & n17741 ) | ( n17740 & n17741 ) ;
  assign n17743 = n17537 & ~n17742 ;
  assign n17744 = n17742 | n17743 ;
  assign n17745 = ( ~n17537 & n17743 ) | ( ~n17537 & n17744 ) | ( n17743 & n17744 ) ;
  assign n17746 = x123 & n1421 ;
  assign n17747 = x122 & n1416 ;
  assign n17748 = x121 & ~n1415 ;
  assign n17749 = n1584 & n17748 ;
  assign n17750 = n17747 | n17749 ;
  assign n17751 = n17746 | n17750 ;
  assign n17752 = n1424 | n17751 ;
  assign n17753 = ( n11219 & n17751 ) | ( n11219 & n17752 ) | ( n17751 & n17752 ) ;
  assign n17754 = x20 & n17753 ;
  assign n17755 = x20 & ~n17754 ;
  assign n17756 = ( n17753 & ~n17754 ) | ( n17753 & n17755 ) | ( ~n17754 & n17755 ) ;
  assign n17757 = n17264 | n17756 ;
  assign n17758 = n17489 | n17757 ;
  assign n17759 = ( n17264 & n17489 ) | ( n17264 & n17756 ) | ( n17489 & n17756 ) ;
  assign n17760 = n17758 & ~n17759 ;
  assign n17761 = x120 & n1817 ;
  assign n17762 = x119 & n1812 ;
  assign n17763 = x118 & ~n1811 ;
  assign n17764 = n1977 & n17763 ;
  assign n17765 = n17762 | n17764 ;
  assign n17766 = n17761 | n17765 ;
  assign n17767 = n1820 | n17766 ;
  assign n17768 = ( n10460 & n17766 ) | ( n10460 & n17767 ) | ( n17766 & n17767 ) ;
  assign n17769 = x23 & n17768 ;
  assign n17770 = x23 & ~n17769 ;
  assign n17771 = ( n17768 & ~n17769 ) | ( n17768 & n17770 ) | ( ~n17769 & n17770 ) ;
  assign n17772 = ( n17473 & n17484 ) | ( n17473 & n17485 ) | ( n17484 & n17485 ) ;
  assign n17773 = n17771 | n17772 ;
  assign n17774 = n17771 & n17772 ;
  assign n17775 = n17773 & ~n17774 ;
  assign n17776 = ( n17745 & n17760 ) | ( n17745 & ~n17775 ) | ( n17760 & ~n17775 ) ;
  assign n17777 = ( ~n17760 & n17775 ) | ( ~n17760 & n17776 ) | ( n17775 & n17776 ) ;
  assign n17778 = ( ~n17745 & n17776 ) | ( ~n17745 & n17777 ) | ( n17776 & n17777 ) ;
  assign n17779 = x126 & n1071 ;
  assign n17780 = x125 & n1066 ;
  assign n17781 = x124 & ~n1065 ;
  assign n17782 = n1189 & n17781 ;
  assign n17783 = n17780 | n17782 ;
  assign n17784 = n17779 | n17783 ;
  assign n17785 = n1074 | n17784 ;
  assign n17786 = ( n12687 & n17784 ) | ( n12687 & n17785 ) | ( n17784 & n17785 ) ;
  assign n17787 = x17 & n17786 ;
  assign n17788 = x17 & ~n17787 ;
  assign n17789 = ( n17786 & ~n17787 ) | ( n17786 & n17788 ) | ( ~n17787 & n17788 ) ;
  assign n17790 = ( n17249 & n17251 ) | ( n17249 & ~n17493 ) | ( n17251 & ~n17493 ) ;
  assign n17791 = ( n17778 & n17789 ) | ( n17778 & ~n17790 ) | ( n17789 & ~n17790 ) ;
  assign n17792 = ( ~n17789 & n17790 ) | ( ~n17789 & n17791 ) | ( n17790 & n17791 ) ;
  assign n17793 = ( ~n17778 & n17791 ) | ( ~n17778 & n17792 ) | ( n17791 & n17792 ) ;
  assign n17794 = n17520 | n17793 ;
  assign n17795 = ( n17228 & n17495 ) | ( n17228 & ~n17517 ) | ( n17495 & ~n17517 ) ;
  assign n17796 = n17794 | n17795 ;
  assign n17797 = ( n17520 & n17793 ) | ( n17520 & n17795 ) | ( n17793 & n17795 ) ;
  assign n17798 = n17796 & ~n17797 ;
  assign n17799 = n17213 | n17798 ;
  assign n17800 = n17500 | n17799 ;
  assign n17801 = ( n17213 & n17500 ) | ( n17213 & n17798 ) | ( n17500 & n17798 ) ;
  assign n17802 = n17800 & ~n17801 ;
  assign n17803 = n17502 | n17505 ;
  assign n17804 = ( n17502 & n17506 ) | ( n17502 & n17803 ) | ( n17506 & n17803 ) ;
  assign n17805 = n17802 | n17804 ;
  assign n17806 = n17802 & n17803 ;
  assign n17807 = n17502 & n17802 ;
  assign n17808 = ( n17506 & n17806 ) | ( n17506 & n17807 ) | ( n17806 & n17807 ) ;
  assign n17809 = n17805 & ~n17808 ;
  assign n17810 = ( n17495 & n17517 ) | ( n17495 & n17518 ) | ( n17517 & n17518 ) ;
  assign n17811 = n17797 | n17810 ;
  assign n17812 = ( n17453 & n17713 ) | ( n17453 & n17724 ) | ( n17713 & n17724 ) ;
  assign n17813 = x112 & n3314 ;
  assign n17814 = x111 & n3309 ;
  assign n17815 = x110 & ~n3308 ;
  assign n17816 = n3570 & n17815 ;
  assign n17817 = n17814 | n17816 ;
  assign n17818 = n17813 | n17817 ;
  assign n17819 = n3317 | n17818 ;
  assign n17820 = ( n7789 & n17818 ) | ( n7789 & n17819 ) | ( n17818 & n17819 ) ;
  assign n17821 = x32 & n17820 ;
  assign n17822 = x32 & ~n17821 ;
  assign n17823 = ( n17820 & ~n17821 ) | ( n17820 & n17822 ) | ( ~n17821 & n17822 ) ;
  assign n17824 = n17812 & n17823 ;
  assign n17825 = n17812 & ~n17824 ;
  assign n17826 = x106 & n4572 ;
  assign n17827 = x105 & n4567 ;
  assign n17828 = x104 & ~n4566 ;
  assign n17829 = n4828 & n17828 ;
  assign n17830 = n17827 | n17829 ;
  assign n17831 = n17826 | n17830 ;
  assign n17832 = n4575 | n17831 ;
  assign n17833 = ( n5814 & n17831 ) | ( n5814 & n17832 ) | ( n17831 & n17832 ) ;
  assign n17834 = x38 & n17833 ;
  assign n17835 = x38 & ~n17834 ;
  assign n17836 = ( n17833 & ~n17834 ) | ( n17833 & n17835 ) | ( ~n17834 & n17835 ) ;
  assign n17837 = x103 & n5340 ;
  assign n17838 = x102 & n5335 ;
  assign n17839 = x101 & ~n5334 ;
  assign n17840 = n5580 & n17839 ;
  assign n17841 = n17838 | n17840 ;
  assign n17842 = n17837 | n17841 ;
  assign n17843 = n5343 | n17842 ;
  assign n17844 = ( n5264 & n17842 ) | ( n5264 & n17843 ) | ( n17842 & n17843 ) ;
  assign n17845 = x41 & n17844 ;
  assign n17846 = x41 & ~n17845 ;
  assign n17847 = ( n17844 & ~n17845 ) | ( n17844 & n17846 ) | ( ~n17845 & n17846 ) ;
  assign n17848 = ( n17549 & n17655 ) | ( n17549 & n17656 ) | ( n17655 & n17656 ) ;
  assign n17849 = ( n17638 & n17641 ) | ( n17638 & ~n17653 ) | ( n17641 & ~n17653 ) ;
  assign n17850 = ( n17550 & n17619 ) | ( n17550 & n17634 ) | ( n17619 & n17634 ) ;
  assign n17851 = x94 & n7812 ;
  assign n17852 = x93 & n7807 ;
  assign n17853 = x92 & ~n7806 ;
  assign n17854 = n8136 & n17853 ;
  assign n17855 = n17852 | n17854 ;
  assign n17856 = n17851 | n17855 ;
  assign n17857 = n7815 | n17856 ;
  assign n17858 = ( n3271 & n17856 ) | ( n3271 & n17857 ) | ( n17856 & n17857 ) ;
  assign n17859 = x50 & n17858 ;
  assign n17860 = x50 & ~n17859 ;
  assign n17861 = ( n17858 & ~n17859 ) | ( n17858 & n17860 ) | ( ~n17859 & n17860 ) ;
  assign n17862 = n17587 | n17601 ;
  assign n17863 = n17566 | n17580 ;
  assign n17864 = x82 & n11984 ;
  assign n17865 = x81 & n11979 ;
  assign n17866 = x80 & ~n11978 ;
  assign n17867 = n12430 & n17866 ;
  assign n17868 = n17865 | n17867 ;
  assign n17869 = n17864 | n17868 ;
  assign n17870 = n11987 | n17869 ;
  assign n17871 = ( n1371 & n17869 ) | ( n1371 & n17870 ) | ( n17869 & n17870 ) ;
  assign n17872 = ~x62 & n17871 ;
  assign n17873 = x62 & ~n17871 ;
  assign n17874 = n17872 | n17873 ;
  assign n17875 = x79 & n12808 ;
  assign n17876 = x63 & x78 ;
  assign n17877 = ~n12808 & n17876 ;
  assign n17878 = n17875 | n17877 ;
  assign n17879 = ~x14 & n17878 ;
  assign n17880 = n17878 & ~n17879 ;
  assign n17881 = x14 | n17878 ;
  assign n17882 = ~n17880 & n17881 ;
  assign n17883 = n17324 & ~n17882 ;
  assign n17884 = ~n17324 & n17882 ;
  assign n17885 = n17883 | n17884 ;
  assign n17886 = ( n17863 & n17874 ) | ( n17863 & ~n17885 ) | ( n17874 & ~n17885 ) ;
  assign n17887 = ( ~n17874 & n17885 ) | ( ~n17874 & n17886 ) | ( n17885 & n17886 ) ;
  assign n17888 = ( ~n17863 & n17886 ) | ( ~n17863 & n17887 ) | ( n17886 & n17887 ) ;
  assign n17889 = x85 & n10876 ;
  assign n17890 = x84 & n10871 ;
  assign n17891 = x83 & ~n10870 ;
  assign n17892 = n11305 & n17891 ;
  assign n17893 = n17890 | n17892 ;
  assign n17894 = n17889 | n17893 ;
  assign n17895 = n10879 | n17894 ;
  assign n17896 = ( n1765 & n17894 ) | ( n1765 & n17895 ) | ( n17894 & n17895 ) ;
  assign n17897 = x59 & n17896 ;
  assign n17898 = x59 & ~n17897 ;
  assign n17899 = ( n17896 & ~n17897 ) | ( n17896 & n17898 ) | ( ~n17897 & n17898 ) ;
  assign n17900 = ~n17888 & n17899 ;
  assign n17901 = n17888 | n17900 ;
  assign n17902 = n17888 & n17899 ;
  assign n17903 = n17584 | n17902 ;
  assign n17904 = n17901 & ~n17903 ;
  assign n17905 = ( n17584 & ~n17901 ) | ( n17584 & n17902 ) | ( ~n17901 & n17902 ) ;
  assign n17906 = n17904 | n17905 ;
  assign n17907 = x88 & n9853 ;
  assign n17908 = x87 & n9848 ;
  assign n17909 = x86 & ~n9847 ;
  assign n17910 = n10165 & n17909 ;
  assign n17911 = n17908 | n17910 ;
  assign n17912 = n17907 | n17911 ;
  assign n17913 = n9856 | n17912 ;
  assign n17914 = ( n2095 & n17912 ) | ( n2095 & n17913 ) | ( n17912 & n17913 ) ;
  assign n17915 = x56 & n17914 ;
  assign n17916 = x56 & ~n17915 ;
  assign n17917 = ( n17914 & ~n17915 ) | ( n17914 & n17916 ) | ( ~n17915 & n17916 ) ;
  assign n17918 = ( n17862 & n17906 ) | ( n17862 & ~n17917 ) | ( n17906 & ~n17917 ) ;
  assign n17919 = ( n17862 & ~n17906 ) | ( n17862 & n17917 ) | ( ~n17906 & n17917 ) ;
  assign n17920 = ( ~n17862 & n17918 ) | ( ~n17862 & n17919 ) | ( n17918 & n17919 ) ;
  assign n17921 = x91 & n8834 ;
  assign n17922 = x90 & n8829 ;
  assign n17923 = x89 & ~n8828 ;
  assign n17924 = n9159 & n17923 ;
  assign n17925 = n17922 | n17924 ;
  assign n17926 = n17921 | n17925 ;
  assign n17927 = n8837 | n17926 ;
  assign n17928 = ( n2714 & n17926 ) | ( n2714 & n17927 ) | ( n17926 & n17927 ) ;
  assign n17929 = x53 & n17928 ;
  assign n17930 = x53 & ~n17929 ;
  assign n17931 = ( n17928 & ~n17929 ) | ( n17928 & n17930 ) | ( ~n17929 & n17930 ) ;
  assign n17932 = ~n17920 & n17931 ;
  assign n17933 = n17920 | n17932 ;
  assign n17934 = n17920 & n17931 ;
  assign n17935 = n17603 | n17617 ;
  assign n17936 = n17934 | n17935 ;
  assign n17937 = n17933 & ~n17936 ;
  assign n17938 = ( ~n17933 & n17934 ) | ( ~n17933 & n17935 ) | ( n17934 & n17935 ) ;
  assign n17939 = n17937 | n17938 ;
  assign n17940 = n17861 & ~n17939 ;
  assign n17941 = n17939 | n17940 ;
  assign n17942 = ( ~n17861 & n17940 ) | ( ~n17861 & n17941 ) | ( n17940 & n17941 ) ;
  assign n17943 = n17850 & n17942 ;
  assign n17944 = n17850 | n17942 ;
  assign n17945 = ~n17943 & n17944 ;
  assign n17946 = x97 & n6937 ;
  assign n17947 = x96 & n6932 ;
  assign n17948 = x95 & ~n6931 ;
  assign n17949 = n7216 & n17948 ;
  assign n17950 = n17947 | n17949 ;
  assign n17951 = n17946 | n17950 ;
  assign n17952 = n6940 | n17951 ;
  assign n17953 = ( n3707 & n17951 ) | ( n3707 & n17952 ) | ( n17951 & n17952 ) ;
  assign n17954 = x47 & n17953 ;
  assign n17955 = x47 & ~n17954 ;
  assign n17956 = ( n17953 & ~n17954 ) | ( n17953 & n17955 ) | ( ~n17954 & n17955 ) ;
  assign n17957 = n17945 & n17956 ;
  assign n17958 = n17945 & ~n17957 ;
  assign n17959 = ~n17945 & n17956 ;
  assign n17960 = n17958 | n17959 ;
  assign n17961 = n17849 & n17960 ;
  assign n17962 = n17960 & ~n17961 ;
  assign n17963 = ( n17849 & ~n17961 ) | ( n17849 & n17962 ) | ( ~n17961 & n17962 ) ;
  assign n17964 = x100 & n6068 ;
  assign n17965 = x99 & n6063 ;
  assign n17966 = x98 & ~n6062 ;
  assign n17967 = n6398 & n17966 ;
  assign n17968 = n17965 | n17967 ;
  assign n17969 = n17964 | n17968 ;
  assign n17970 = n6071 | n17969 ;
  assign n17971 = ( n4532 & n17969 ) | ( n4532 & n17970 ) | ( n17969 & n17970 ) ;
  assign n17972 = x44 & n17971 ;
  assign n17973 = x44 & ~n17972 ;
  assign n17974 = ( n17971 & ~n17972 ) | ( n17971 & n17973 ) | ( ~n17972 & n17973 ) ;
  assign n17975 = n17963 & n17974 ;
  assign n17976 = n17963 | n17974 ;
  assign n17977 = ~n17975 & n17976 ;
  assign n17978 = n17848 | n17977 ;
  assign n17979 = n17848 & n17977 ;
  assign n17980 = n17978 & ~n17979 ;
  assign n17981 = n17661 | n17675 ;
  assign n17982 = ( n17847 & n17980 ) | ( n17847 & n17981 ) | ( n17980 & n17981 ) ;
  assign n17983 = ( n17980 & n17981 ) | ( n17980 & ~n17982 ) | ( n17981 & ~n17982 ) ;
  assign n17984 = ( n17847 & ~n17982 ) | ( n17847 & n17983 ) | ( ~n17982 & n17983 ) ;
  assign n17985 = n17836 & n17984 ;
  assign n17986 = n17836 | n17984 ;
  assign n17987 = ~n17985 & n17986 ;
  assign n17988 = n17678 | n17692 ;
  assign n17989 = n17987 | n17988 ;
  assign n17990 = n17987 & n17988 ;
  assign n17991 = n17989 & ~n17990 ;
  assign n17992 = x109 & n3913 ;
  assign n17993 = x108 & n3908 ;
  assign n17994 = x107 & ~n3907 ;
  assign n17995 = n4152 & n17994 ;
  assign n17996 = n17993 | n17995 ;
  assign n17997 = n17992 | n17996 ;
  assign n17998 = n3916 | n17997 ;
  assign n17999 = ( n6884 & n17997 ) | ( n6884 & n17998 ) | ( n17997 & n17998 ) ;
  assign n18000 = x35 & n17999 ;
  assign n18001 = x35 & ~n18000 ;
  assign n18002 = ( n17999 & ~n18000 ) | ( n17999 & n18001 ) | ( ~n18000 & n18001 ) ;
  assign n18003 = n17991 & n18002 ;
  assign n18004 = n17991 & ~n18003 ;
  assign n18005 = ~n17991 & n18002 ;
  assign n18006 = n18004 | n18005 ;
  assign n18007 = n17696 | n17710 ;
  assign n18008 = n18006 | n18007 ;
  assign n18009 = n18006 & n18007 ;
  assign n18010 = n18008 & ~n18009 ;
  assign n18011 = ~n17812 & n17823 ;
  assign n18012 = n18010 | n18011 ;
  assign n18013 = n17825 | n18012 ;
  assign n18014 = ( n17825 & n18010 ) | ( n17825 & n18011 ) | ( n18010 & n18011 ) ;
  assign n18015 = n18013 & ~n18014 ;
  assign n18016 = x115 & n2775 ;
  assign n18017 = x114 & n2770 ;
  assign n18018 = x113 & ~n2769 ;
  assign n18019 = n2978 & n18018 ;
  assign n18020 = n18017 | n18019 ;
  assign n18021 = n18016 | n18020 ;
  assign n18022 = n2778 | n18021 ;
  assign n18023 = ( n8749 & n18021 ) | ( n8749 & n18022 ) | ( n18021 & n18022 ) ;
  assign n18024 = x29 & n18023 ;
  assign n18025 = x29 & ~n18024 ;
  assign n18026 = ( n18023 & ~n18024 ) | ( n18023 & n18025 ) | ( ~n18024 & n18025 ) ;
  assign n18027 = ( n17727 & n17738 ) | ( n17727 & n17739 ) | ( n17738 & n17739 ) ;
  assign n18028 = n18026 | n18027 ;
  assign n18029 = n18026 & n18027 ;
  assign n18030 = n18028 & ~n18029 ;
  assign n18031 = n18015 & n18030 ;
  assign n18032 = n18030 & ~n18031 ;
  assign n18033 = ( n18015 & ~n18031 ) | ( n18015 & n18032 ) | ( ~n18031 & n18032 ) ;
  assign n18034 = x121 & n1817 ;
  assign n18035 = x120 & n1812 ;
  assign n18036 = x119 & ~n1811 ;
  assign n18037 = n1977 & n18036 ;
  assign n18038 = n18035 | n18037 ;
  assign n18039 = n18034 | n18038 ;
  assign n18040 = n1820 | n18039 ;
  assign n18041 = ( n10811 & n18039 ) | ( n10811 & n18040 ) | ( n18039 & n18040 ) ;
  assign n18042 = x23 & n18041 ;
  assign n18043 = x23 & ~n18042 ;
  assign n18044 = ( n18041 & ~n18042 ) | ( n18041 & n18043 ) | ( ~n18042 & n18043 ) ;
  assign n18045 = n17745 & n17775 ;
  assign n18046 = n17774 | n18045 ;
  assign n18047 = ~n18044 & n18046 ;
  assign n18048 = n18044 & ~n18046 ;
  assign n18049 = n18047 | n18048 ;
  assign n18050 = x118 & n2280 ;
  assign n18051 = x117 & n2275 ;
  assign n18052 = x116 & ~n2274 ;
  assign n18053 = n2481 & n18052 ;
  assign n18054 = n18051 | n18053 ;
  assign n18055 = n18050 | n18054 ;
  assign n18056 = n2283 | n18055 ;
  assign n18057 = ( n9760 & n18055 ) | ( n9760 & n18056 ) | ( n18055 & n18056 ) ;
  assign n18058 = x26 & n18057 ;
  assign n18059 = x26 & ~n18058 ;
  assign n18060 = ( n18057 & ~n18058 ) | ( n18057 & n18059 ) | ( ~n18058 & n18059 ) ;
  assign n18061 = ( n17534 & n17536 ) | ( n17534 & n17742 ) | ( n17536 & n17742 ) ;
  assign n18062 = n18060 | n18061 ;
  assign n18063 = n18060 & n18061 ;
  assign n18064 = n18062 & ~n18063 ;
  assign n18065 = ( n18033 & n18049 ) | ( n18033 & ~n18064 ) | ( n18049 & ~n18064 ) ;
  assign n18066 = ( ~n18049 & n18064 ) | ( ~n18049 & n18065 ) | ( n18064 & n18065 ) ;
  assign n18067 = ( ~n18033 & n18065 ) | ( ~n18033 & n18066 ) | ( n18065 & n18066 ) ;
  assign n18068 = x124 & n1421 ;
  assign n18069 = x123 & n1416 ;
  assign n18070 = x122 & ~n1415 ;
  assign n18071 = n1584 & n18070 ;
  assign n18072 = n18069 | n18071 ;
  assign n18073 = n18068 | n18072 ;
  assign n18074 = n1424 | n18073 ;
  assign n18075 = ( n11916 & n18073 ) | ( n11916 & n18074 ) | ( n18073 & n18074 ) ;
  assign n18076 = x20 & n18075 ;
  assign n18077 = x20 & ~n18076 ;
  assign n18078 = ( n18075 & ~n18076 ) | ( n18075 & n18077 ) | ( ~n18076 & n18077 ) ;
  assign n18079 = ( n17745 & n17760 ) | ( n17745 & n17775 ) | ( n17760 & n17775 ) ;
  assign n18080 = ( n17759 & ~n18045 ) | ( n17759 & n18079 ) | ( ~n18045 & n18079 ) ;
  assign n18081 = n18078 | n18080 ;
  assign n18082 = n18078 & n18080 ;
  assign n18083 = n18081 & ~n18082 ;
  assign n18084 = x127 & n1071 ;
  assign n18085 = x126 & n1066 ;
  assign n18086 = x125 & ~n1065 ;
  assign n18087 = n1189 & n18086 ;
  assign n18088 = n18085 | n18087 ;
  assign n18089 = n18084 | n18088 ;
  assign n18090 = n1074 | n18089 ;
  assign n18091 = ( n12720 & n18089 ) | ( n12720 & n18090 ) | ( n18089 & n18090 ) ;
  assign n18092 = x17 & n18091 ;
  assign n18093 = x17 & ~n18092 ;
  assign n18094 = ( n18091 & ~n18092 ) | ( n18091 & n18093 ) | ( ~n18092 & n18093 ) ;
  assign n18095 = ( n17778 & n17789 ) | ( n17778 & n17790 ) | ( n17789 & n17790 ) ;
  assign n18096 = n18094 & n18095 ;
  assign n18097 = n18094 | n18095 ;
  assign n18098 = ~n18096 & n18097 ;
  assign n18099 = ( n18067 & ~n18083 ) | ( n18067 & n18098 ) | ( ~n18083 & n18098 ) ;
  assign n18100 = ( n18083 & ~n18098 ) | ( n18083 & n18099 ) | ( ~n18098 & n18099 ) ;
  assign n18101 = ( ~n18067 & n18099 ) | ( ~n18067 & n18100 ) | ( n18099 & n18100 ) ;
  assign n18102 = n17811 | n18101 ;
  assign n18103 = n17811 & n18101 ;
  assign n18104 = n18102 & ~n18103 ;
  assign n18105 = n17801 | n17806 ;
  assign n18106 = n17801 | n17807 ;
  assign n18107 = ( n17506 & n18105 ) | ( n17506 & n18106 ) | ( n18105 & n18106 ) ;
  assign n18108 = n18104 | n18107 ;
  assign n18109 = n18104 & n18105 ;
  assign n18110 = n18104 & n18106 ;
  assign n18111 = ( n17506 & n18109 ) | ( n17506 & n18110 ) | ( n18109 & n18110 ) ;
  assign n18112 = n18108 & ~n18111 ;
  assign n18113 = x113 & n3314 ;
  assign n18114 = x112 & n3309 ;
  assign n18115 = x111 & ~n3308 ;
  assign n18116 = n3570 & n18115 ;
  assign n18117 = n18114 | n18116 ;
  assign n18118 = n18113 | n18117 ;
  assign n18119 = n3317 | n18118 ;
  assign n18120 = ( n8113 & n18118 ) | ( n8113 & n18119 ) | ( n18118 & n18119 ) ;
  assign n18121 = x32 & n18120 ;
  assign n18122 = x32 & ~n18121 ;
  assign n18123 = ( n18120 & ~n18121 ) | ( n18120 & n18122 ) | ( ~n18121 & n18122 ) ;
  assign n18124 = n18003 | n18009 ;
  assign n18125 = n18123 | n18124 ;
  assign n18126 = n18123 & n18124 ;
  assign n18127 = n18125 & ~n18126 ;
  assign n18128 = x116 & n2775 ;
  assign n18129 = x115 & n2770 ;
  assign n18130 = x114 & ~n2769 ;
  assign n18131 = n2978 & n18130 ;
  assign n18132 = n18129 | n18131 ;
  assign n18133 = n18128 | n18132 ;
  assign n18134 = n2778 | n18133 ;
  assign n18135 = ( n8778 & n18133 ) | ( n8778 & n18134 ) | ( n18133 & n18134 ) ;
  assign n18136 = x29 & n18135 ;
  assign n18137 = x29 & ~n18136 ;
  assign n18138 = ( n18135 & ~n18136 ) | ( n18135 & n18137 ) | ( ~n18136 & n18137 ) ;
  assign n18139 = n17824 & n18138 ;
  assign n18140 = n18138 & ~n18139 ;
  assign n18141 = ~n18014 & n18140 ;
  assign n18142 = ( n17824 & n18014 ) | ( n17824 & ~n18138 ) | ( n18014 & ~n18138 ) ;
  assign n18143 = n18141 | n18142 ;
  assign n18144 = x110 & n3913 ;
  assign n18145 = x109 & n3908 ;
  assign n18146 = x108 & ~n3907 ;
  assign n18147 = n4152 & n18146 ;
  assign n18148 = n18145 | n18147 ;
  assign n18149 = n18144 | n18148 ;
  assign n18150 = n3916 | n18149 ;
  assign n18151 = ( n7189 & n18149 ) | ( n7189 & n18150 ) | ( n18149 & n18150 ) ;
  assign n18152 = x35 & n18151 ;
  assign n18153 = x35 & ~n18152 ;
  assign n18154 = ( n18151 & ~n18152 ) | ( n18151 & n18153 ) | ( ~n18152 & n18153 ) ;
  assign n18155 = n17985 | n17990 ;
  assign n18156 = x107 & n4572 ;
  assign n18157 = x106 & n4567 ;
  assign n18158 = x105 & ~n4566 ;
  assign n18159 = n4828 & n18158 ;
  assign n18160 = n18157 | n18159 ;
  assign n18161 = n18156 | n18160 ;
  assign n18162 = n4575 | n18161 ;
  assign n18163 = ( n6328 & n18161 ) | ( n6328 & n18162 ) | ( n18161 & n18162 ) ;
  assign n18164 = x38 & n18163 ;
  assign n18165 = x38 & ~n18164 ;
  assign n18166 = ( n18163 & ~n18164 ) | ( n18163 & n18165 ) | ( ~n18164 & n18165 ) ;
  assign n18167 = n17975 | n17979 ;
  assign n18168 = n17957 | n17961 ;
  assign n18169 = n17932 | n17938 ;
  assign n18170 = n17900 | n17905 ;
  assign n18171 = x86 & n10876 ;
  assign n18172 = x85 & n10871 ;
  assign n18173 = x84 & ~n10870 ;
  assign n18174 = n11305 & n18173 ;
  assign n18175 = n18172 | n18174 ;
  assign n18176 = n18171 | n18175 ;
  assign n18177 = n10879 | n18176 ;
  assign n18178 = ( n1921 & n18176 ) | ( n1921 & n18177 ) | ( n18176 & n18177 ) ;
  assign n18179 = x59 & n18178 ;
  assign n18180 = x59 & ~n18179 ;
  assign n18181 = ( n18178 & ~n18179 ) | ( n18178 & n18180 ) | ( ~n18179 & n18180 ) ;
  assign n18182 = x80 & n12808 ;
  assign n18183 = x63 & x79 ;
  assign n18184 = ~n12808 & n18183 ;
  assign n18185 = n18182 | n18184 ;
  assign n18186 = ~n17879 & n18185 ;
  assign n18187 = ~n17883 & n18186 ;
  assign n18188 = ( n17879 & n17883 ) | ( n17879 & ~n18185 ) | ( n17883 & ~n18185 ) ;
  assign n18189 = n18187 | n18188 ;
  assign n18190 = x83 & n11984 ;
  assign n18191 = x82 & n11979 ;
  assign n18192 = x81 & ~n11978 ;
  assign n18193 = n12430 & n18192 ;
  assign n18194 = n18191 | n18193 ;
  assign n18195 = n18190 | n18194 ;
  assign n18196 = n11987 | n18195 ;
  assign n18197 = ( n1510 & n18195 ) | ( n1510 & n18196 ) | ( n18195 & n18196 ) ;
  assign n18198 = x62 & n18197 ;
  assign n18199 = x62 & ~n18198 ;
  assign n18200 = ( n18197 & ~n18198 ) | ( n18197 & n18199 ) | ( ~n18198 & n18199 ) ;
  assign n18201 = ~n18189 & n18200 ;
  assign n18202 = n18189 & ~n18200 ;
  assign n18203 = n18201 | n18202 ;
  assign n18204 = ( ~n17886 & n18181 ) | ( ~n17886 & n18203 ) | ( n18181 & n18203 ) ;
  assign n18205 = ( n17886 & ~n18203 ) | ( n17886 & n18204 ) | ( ~n18203 & n18204 ) ;
  assign n18206 = ( ~n18181 & n18204 ) | ( ~n18181 & n18205 ) | ( n18204 & n18205 ) ;
  assign n18207 = ~n18170 & n18206 ;
  assign n18208 = n18170 & ~n18206 ;
  assign n18209 = n18207 | n18208 ;
  assign n18210 = x89 & n9853 ;
  assign n18211 = x88 & n9848 ;
  assign n18212 = x87 & ~n9847 ;
  assign n18213 = n10165 & n18212 ;
  assign n18214 = n18211 | n18213 ;
  assign n18215 = n18210 | n18214 ;
  assign n18216 = n9856 | n18215 ;
  assign n18217 = ( n2244 & n18215 ) | ( n2244 & n18216 ) | ( n18215 & n18216 ) ;
  assign n18218 = x56 & n18217 ;
  assign n18219 = x56 & ~n18218 ;
  assign n18220 = ( n18217 & ~n18218 ) | ( n18217 & n18219 ) | ( ~n18218 & n18219 ) ;
  assign n18221 = n18209 & n18220 ;
  assign n18222 = ~n17919 & n18221 ;
  assign n18223 = ( n18170 & ~n18206 ) | ( n18170 & n18220 ) | ( ~n18206 & n18220 ) ;
  assign n18224 = n18207 | n18223 ;
  assign n18225 = ( n17919 & ~n18222 ) | ( n17919 & n18224 ) | ( ~n18222 & n18224 ) ;
  assign n18226 = ~n18221 & n18224 ;
  assign n18227 = ( n17919 & n18222 ) | ( n17919 & n18226 ) | ( n18222 & n18226 ) ;
  assign n18228 = n18225 & ~n18227 ;
  assign n18229 = x92 & n8834 ;
  assign n18230 = x91 & n8829 ;
  assign n18231 = x90 & ~n8828 ;
  assign n18232 = n9159 & n18231 ;
  assign n18233 = n18230 | n18232 ;
  assign n18234 = n18229 | n18233 ;
  assign n18235 = n8837 | n18234 ;
  assign n18236 = ( n2904 & n18234 ) | ( n2904 & n18235 ) | ( n18234 & n18235 ) ;
  assign n18237 = x53 & n18236 ;
  assign n18238 = x53 & ~n18237 ;
  assign n18239 = ( n18236 & ~n18237 ) | ( n18236 & n18238 ) | ( ~n18237 & n18238 ) ;
  assign n18240 = ( n18169 & n18228 ) | ( n18169 & ~n18239 ) | ( n18228 & ~n18239 ) ;
  assign n18241 = ( ~n18228 & n18239 ) | ( ~n18228 & n18240 ) | ( n18239 & n18240 ) ;
  assign n18242 = ( ~n18169 & n18240 ) | ( ~n18169 & n18241 ) | ( n18240 & n18241 ) ;
  assign n18243 = x95 & n7812 ;
  assign n18244 = x94 & n7807 ;
  assign n18245 = x93 & ~n7806 ;
  assign n18246 = n8136 & n18245 ;
  assign n18247 = n18244 | n18246 ;
  assign n18248 = n18243 | n18247 ;
  assign n18249 = n7815 | n18248 ;
  assign n18250 = ( n3479 & n18248 ) | ( n3479 & n18249 ) | ( n18248 & n18249 ) ;
  assign n18251 = x50 & n18250 ;
  assign n18252 = x50 & ~n18251 ;
  assign n18253 = ( n18250 & ~n18251 ) | ( n18250 & n18252 ) | ( ~n18251 & n18252 ) ;
  assign n18254 = n18242 | n18253 ;
  assign n18255 = ~n18253 & n18254 ;
  assign n18256 = ( ~n18242 & n18254 ) | ( ~n18242 & n18255 ) | ( n18254 & n18255 ) ;
  assign n18257 = ~n17940 & n17944 ;
  assign n18258 = n18256 & n18257 ;
  assign n18259 = n18256 | n18257 ;
  assign n18260 = ~n18258 & n18259 ;
  assign n18261 = x98 & n6937 ;
  assign n18262 = x97 & n6932 ;
  assign n18263 = x96 & ~n6931 ;
  assign n18264 = n7216 & n18263 ;
  assign n18265 = n18262 | n18264 ;
  assign n18266 = n18261 | n18265 ;
  assign n18267 = n6940 | n18266 ;
  assign n18268 = ( n4105 & n18266 ) | ( n4105 & n18267 ) | ( n18266 & n18267 ) ;
  assign n18269 = x47 & n18268 ;
  assign n18270 = x47 & ~n18269 ;
  assign n18271 = ( n18268 & ~n18269 ) | ( n18268 & n18270 ) | ( ~n18269 & n18270 ) ;
  assign n18272 = n18260 | n18271 ;
  assign n18273 = n18260 & n18271 ;
  assign n18274 = n18272 & ~n18273 ;
  assign n18275 = n18168 & n18274 ;
  assign n18276 = n18168 & ~n18275 ;
  assign n18277 = ~n18168 & n18274 ;
  assign n18278 = x101 & n6068 ;
  assign n18279 = x100 & n6063 ;
  assign n18280 = x99 & ~n6062 ;
  assign n18281 = n6398 & n18280 ;
  assign n18282 = n18279 | n18281 ;
  assign n18283 = n18278 | n18282 ;
  assign n18284 = n6071 | n18283 ;
  assign n18285 = ( n4783 & n18283 ) | ( n4783 & n18284 ) | ( n18283 & n18284 ) ;
  assign n18286 = x44 & n18285 ;
  assign n18287 = x44 & ~n18286 ;
  assign n18288 = ( n18285 & ~n18286 ) | ( n18285 & n18287 ) | ( ~n18286 & n18287 ) ;
  assign n18289 = n18277 | n18288 ;
  assign n18290 = n18276 | n18289 ;
  assign n18291 = ( n18276 & n18277 ) | ( n18276 & n18288 ) | ( n18277 & n18288 ) ;
  assign n18292 = n18290 & ~n18291 ;
  assign n18293 = x104 & n5340 ;
  assign n18294 = x103 & n5335 ;
  assign n18295 = x102 & ~n5334 ;
  assign n18296 = n5580 & n18295 ;
  assign n18297 = n18294 | n18296 ;
  assign n18298 = n18293 | n18297 ;
  assign n18299 = n5343 | n18298 ;
  assign n18300 = ( n5295 & n18298 ) | ( n5295 & n18299 ) | ( n18298 & n18299 ) ;
  assign n18301 = x41 & n18300 ;
  assign n18302 = x41 & ~n18301 ;
  assign n18303 = ( n18300 & ~n18301 ) | ( n18300 & n18302 ) | ( ~n18301 & n18302 ) ;
  assign n18304 = ( n18167 & n18292 ) | ( n18167 & n18303 ) | ( n18292 & n18303 ) ;
  assign n18305 = ( n18292 & n18303 ) | ( n18292 & ~n18304 ) | ( n18303 & ~n18304 ) ;
  assign n18306 = ( n18167 & ~n18304 ) | ( n18167 & n18305 ) | ( ~n18304 & n18305 ) ;
  assign n18307 = ( n17982 & n18166 ) | ( n17982 & ~n18306 ) | ( n18166 & ~n18306 ) ;
  assign n18308 = ( ~n17982 & n18306 ) | ( ~n17982 & n18307 ) | ( n18306 & n18307 ) ;
  assign n18309 = ( ~n18166 & n18307 ) | ( ~n18166 & n18308 ) | ( n18307 & n18308 ) ;
  assign n18310 = ( n18154 & n18155 ) | ( n18154 & ~n18309 ) | ( n18155 & ~n18309 ) ;
  assign n18311 = ( ~n18155 & n18309 ) | ( ~n18155 & n18310 ) | ( n18309 & n18310 ) ;
  assign n18312 = ( ~n18154 & n18310 ) | ( ~n18154 & n18311 ) | ( n18310 & n18311 ) ;
  assign n18313 = ( n18127 & ~n18143 ) | ( n18127 & n18312 ) | ( ~n18143 & n18312 ) ;
  assign n18314 = ( n18143 & ~n18312 ) | ( n18143 & n18313 ) | ( ~n18312 & n18313 ) ;
  assign n18315 = ( ~n18127 & n18313 ) | ( ~n18127 & n18314 ) | ( n18313 & n18314 ) ;
  assign n18316 = x122 & n1817 ;
  assign n18317 = x121 & n1812 ;
  assign n18318 = x120 & ~n1811 ;
  assign n18319 = n1977 & n18318 ;
  assign n18320 = n18317 | n18319 ;
  assign n18321 = n18316 | n18320 ;
  assign n18322 = n1820 | n18321 ;
  assign n18323 = ( n11188 & n18321 ) | ( n11188 & n18322 ) | ( n18321 & n18322 ) ;
  assign n18324 = x23 & n18323 ;
  assign n18325 = x23 & ~n18324 ;
  assign n18326 = ( n18323 & ~n18324 ) | ( n18323 & n18325 ) | ( ~n18324 & n18325 ) ;
  assign n18327 = ( n18033 & n18060 ) | ( n18033 & n18061 ) | ( n18060 & n18061 ) ;
  assign n18328 = n18326 | n18327 ;
  assign n18329 = n18326 & n18327 ;
  assign n18330 = n18328 & ~n18329 ;
  assign n18331 = n18029 | n18031 ;
  assign n18332 = x119 & n2280 ;
  assign n18333 = x118 & n2275 ;
  assign n18334 = x117 & ~n2274 ;
  assign n18335 = n2481 & n18334 ;
  assign n18336 = n18333 | n18335 ;
  assign n18337 = n18332 | n18336 ;
  assign n18338 = n2283 | n18337 ;
  assign n18339 = ( n9789 & n18337 ) | ( n9789 & n18338 ) | ( n18337 & n18338 ) ;
  assign n18340 = x26 & n18339 ;
  assign n18341 = x26 & ~n18340 ;
  assign n18342 = ( n18339 & ~n18340 ) | ( n18339 & n18341 ) | ( ~n18340 & n18341 ) ;
  assign n18343 = n18331 | n18342 ;
  assign n18344 = n18331 & n18342 ;
  assign n18345 = n18343 & ~n18344 ;
  assign n18346 = ( n18315 & n18330 ) | ( n18315 & ~n18345 ) | ( n18330 & ~n18345 ) ;
  assign n18347 = ( ~n18330 & n18345 ) | ( ~n18330 & n18346 ) | ( n18345 & n18346 ) ;
  assign n18348 = ( ~n18315 & n18346 ) | ( ~n18315 & n18347 ) | ( n18346 & n18347 ) ;
  assign n18349 = x127 & n1066 ;
  assign n18350 = x126 & ~n1065 ;
  assign n18351 = n1189 & n18350 ;
  assign n18352 = n18349 | n18351 ;
  assign n18353 = n1074 | n18352 ;
  assign n18354 = ( n13461 & n18352 ) | ( n13461 & n18353 ) | ( n18352 & n18353 ) ;
  assign n18355 = x17 & n18354 ;
  assign n18356 = x17 & ~n18355 ;
  assign n18357 = ( n18354 & ~n18355 ) | ( n18354 & n18356 ) | ( ~n18355 & n18356 ) ;
  assign n18358 = ( n18067 & n18078 ) | ( n18067 & n18080 ) | ( n18078 & n18080 ) ;
  assign n18359 = n18357 & n18358 ;
  assign n18360 = n18357 | n18358 ;
  assign n18361 = ~n18359 & n18360 ;
  assign n18362 = x125 & n1421 ;
  assign n18363 = x124 & n1416 ;
  assign n18364 = x123 & ~n1415 ;
  assign n18365 = n1584 & n18364 ;
  assign n18366 = n18363 | n18365 ;
  assign n18367 = n18362 | n18366 ;
  assign n18368 = n1424 | n18367 ;
  assign n18369 = ( n12310 & n18367 ) | ( n12310 & n18368 ) | ( n18367 & n18368 ) ;
  assign n18370 = x20 & n18369 ;
  assign n18371 = x20 & ~n18370 ;
  assign n18372 = ( n18369 & ~n18370 ) | ( n18369 & n18371 ) | ( ~n18370 & n18371 ) ;
  assign n18373 = ( n18044 & n18046 ) | ( n18044 & ~n18067 ) | ( n18046 & ~n18067 ) ;
  assign n18374 = n18372 | n18373 ;
  assign n18375 = n18372 & n18373 ;
  assign n18376 = n18374 & ~n18375 ;
  assign n18377 = ( n18348 & n18361 ) | ( n18348 & ~n18376 ) | ( n18361 & ~n18376 ) ;
  assign n18378 = ( ~n18361 & n18376 ) | ( ~n18361 & n18377 ) | ( n18376 & n18377 ) ;
  assign n18379 = ( ~n18348 & n18377 ) | ( ~n18348 & n18378 ) | ( n18377 & n18378 ) ;
  assign n18380 = ( n18094 & n18095 ) | ( n18094 & ~n18101 ) | ( n18095 & ~n18101 ) ;
  assign n18381 = n18379 | n18380 ;
  assign n18382 = n18379 & n18380 ;
  assign n18383 = n18381 & ~n18382 ;
  assign n18384 = n18103 | n18109 ;
  assign n18385 = n18103 | n18110 ;
  assign n18386 = ( n17506 & n18384 ) | ( n17506 & n18385 ) | ( n18384 & n18385 ) ;
  assign n18387 = n18383 | n18386 ;
  assign n18388 = n18383 & n18384 ;
  assign n18389 = n18383 & n18385 ;
  assign n18390 = ( n17506 & n18388 ) | ( n17506 & n18389 ) | ( n18388 & n18389 ) ;
  assign n18391 = n18387 & ~n18390 ;
  assign n18392 = n18348 & n18376 ;
  assign n18393 = n18348 | n18376 ;
  assign n18394 = ~n18392 & n18393 ;
  assign n18395 = ( n18357 & n18358 ) | ( n18357 & n18394 ) | ( n18358 & n18394 ) ;
  assign n18396 = n18375 | n18392 ;
  assign n18397 = x127 & ~n1065 ;
  assign n18398 = n1189 & n18397 ;
  assign n18399 = ( x127 & n1074 ) | ( x127 & n18398 ) | ( n1074 & n18398 ) ;
  assign n18400 = ( x126 & n18398 ) | ( x126 & n18399 ) | ( n18398 & n18399 ) ;
  assign n18401 = ( n12685 & n18399 ) | ( n12685 & n18400 ) | ( n18399 & n18400 ) ;
  assign n18402 = x17 & n18401 ;
  assign n18403 = x17 & ~n18402 ;
  assign n18404 = ( n18401 & ~n18402 ) | ( n18401 & n18403 ) | ( ~n18402 & n18403 ) ;
  assign n18405 = n18396 & n18404 ;
  assign n18406 = n18396 & ~n18405 ;
  assign n18407 = x126 & n1421 ;
  assign n18408 = x125 & n1416 ;
  assign n18409 = x124 & ~n1415 ;
  assign n18410 = n1584 & n18409 ;
  assign n18411 = n18408 | n18410 ;
  assign n18412 = n18407 | n18411 ;
  assign n18413 = n1424 | n18412 ;
  assign n18414 = ( n12687 & n18412 ) | ( n12687 & n18413 ) | ( n18412 & n18413 ) ;
  assign n18415 = x20 & n18414 ;
  assign n18416 = x20 & ~n18415 ;
  assign n18417 = ( n18414 & ~n18415 ) | ( n18414 & n18416 ) | ( ~n18415 & n18416 ) ;
  assign n18418 = ( n18326 & n18327 ) | ( n18326 & ~n18348 ) | ( n18327 & ~n18348 ) ;
  assign n18419 = n18417 | n18418 ;
  assign n18420 = n18417 & n18418 ;
  assign n18421 = n18419 & ~n18420 ;
  assign n18422 = x120 & n2280 ;
  assign n18423 = x119 & n2275 ;
  assign n18424 = x118 & ~n2274 ;
  assign n18425 = n2481 & n18424 ;
  assign n18426 = n18423 | n18425 ;
  assign n18427 = n18422 | n18426 ;
  assign n18428 = n2283 | n18427 ;
  assign n18429 = ( n10460 & n18427 ) | ( n10460 & n18428 ) | ( n18427 & n18428 ) ;
  assign n18430 = x26 & n18429 ;
  assign n18431 = x26 & ~n18430 ;
  assign n18432 = ( n18429 & ~n18430 ) | ( n18429 & n18431 ) | ( ~n18430 & n18431 ) ;
  assign n18433 = ( n18014 & n18138 ) | ( n18014 & n18139 ) | ( n18138 & n18139 ) ;
  assign n18434 = n18127 & n18312 ;
  assign n18435 = ~n18433 & n18434 ;
  assign n18436 = n18127 | n18312 ;
  assign n18437 = ( n18141 & n18142 ) | ( n18141 & n18436 ) | ( n18142 & n18436 ) ;
  assign n18438 = ( n18433 & ~n18435 ) | ( n18433 & n18437 ) | ( ~n18435 & n18437 ) ;
  assign n18439 = n18432 & n18438 ;
  assign n18440 = n18432 | n18438 ;
  assign n18441 = ~n18439 & n18440 ;
  assign n18442 = n18315 & n18345 ;
  assign n18443 = x123 & n1817 ;
  assign n18444 = x122 & n1812 ;
  assign n18445 = x121 & ~n1811 ;
  assign n18446 = n1977 & n18445 ;
  assign n18447 = n18444 | n18446 ;
  assign n18448 = n18443 | n18447 ;
  assign n18449 = n1820 | n18448 ;
  assign n18450 = ( n11219 & n18448 ) | ( n11219 & n18449 ) | ( n18448 & n18449 ) ;
  assign n18451 = x23 & n18450 ;
  assign n18452 = x23 & ~n18451 ;
  assign n18453 = ( n18450 & ~n18451 ) | ( n18450 & n18452 ) | ( ~n18451 & n18452 ) ;
  assign n18454 = n18344 & n18453 ;
  assign n18455 = n18453 & ~n18454 ;
  assign n18456 = ~n18442 & n18455 ;
  assign n18457 = ( n18344 & n18442 ) | ( n18344 & ~n18453 ) | ( n18442 & ~n18453 ) ;
  assign n18458 = n18456 | n18457 ;
  assign n18459 = ( n18154 & n18155 ) | ( n18154 & n18309 ) | ( n18155 & n18309 ) ;
  assign n18460 = x114 & n3314 ;
  assign n18461 = x113 & n3309 ;
  assign n18462 = x112 & ~n3308 ;
  assign n18463 = n3570 & n18462 ;
  assign n18464 = n18461 | n18463 ;
  assign n18465 = n18460 | n18464 ;
  assign n18466 = n3317 | n18465 ;
  assign n18467 = ( n8437 & n18465 ) | ( n8437 & n18466 ) | ( n18465 & n18466 ) ;
  assign n18468 = x32 & n18467 ;
  assign n18469 = x32 & ~n18468 ;
  assign n18470 = ( n18467 & ~n18468 ) | ( n18467 & n18469 ) | ( ~n18468 & n18469 ) ;
  assign n18471 = n18459 | n18470 ;
  assign n18472 = n18459 & n18470 ;
  assign n18473 = n18471 & ~n18472 ;
  assign n18474 = x117 & n2775 ;
  assign n18475 = x116 & n2770 ;
  assign n18476 = x115 & ~n2769 ;
  assign n18477 = n2978 & n18476 ;
  assign n18478 = n18475 | n18477 ;
  assign n18479 = n18474 | n18478 ;
  assign n18480 = n2778 | n18479 ;
  assign n18481 = ( n9118 & n18479 ) | ( n9118 & n18480 ) | ( n18479 & n18480 ) ;
  assign n18482 = x29 & n18481 ;
  assign n18483 = x29 & ~n18482 ;
  assign n18484 = ( n18481 & ~n18482 ) | ( n18481 & n18483 ) | ( ~n18482 & n18483 ) ;
  assign n18485 = n18126 & n18484 ;
  assign n18486 = n18484 & ~n18485 ;
  assign n18487 = ~n18434 & n18486 ;
  assign n18488 = ( n18126 & n18434 ) | ( n18126 & ~n18484 ) | ( n18434 & ~n18484 ) ;
  assign n18489 = n18487 | n18488 ;
  assign n18490 = ( n17982 & n18166 ) | ( n17982 & n18306 ) | ( n18166 & n18306 ) ;
  assign n18491 = n18275 | n18291 ;
  assign n18492 = x102 & n6068 ;
  assign n18493 = x101 & n6063 ;
  assign n18494 = x100 & ~n6062 ;
  assign n18495 = n6398 & n18494 ;
  assign n18496 = n18493 | n18495 ;
  assign n18497 = n18492 | n18496 ;
  assign n18498 = n6071 | n18497 ;
  assign n18499 = ( n5025 & n18497 ) | ( n5025 & n18498 ) | ( n18497 & n18498 ) ;
  assign n18500 = x44 & n18499 ;
  assign n18501 = x44 & ~n18500 ;
  assign n18502 = ( n18499 & ~n18500 ) | ( n18499 & n18501 ) | ( ~n18500 & n18501 ) ;
  assign n18503 = x96 & n7812 ;
  assign n18504 = x95 & n7807 ;
  assign n18505 = x94 & ~n7806 ;
  assign n18506 = n8136 & n18505 ;
  assign n18507 = n18504 | n18506 ;
  assign n18508 = n18503 | n18507 ;
  assign n18509 = n7815 | n18508 ;
  assign n18510 = ( n3509 & n18508 ) | ( n3509 & n18509 ) | ( n18508 & n18509 ) ;
  assign n18511 = x50 & n18510 ;
  assign n18512 = x50 & ~n18511 ;
  assign n18513 = ( n18510 & ~n18511 ) | ( n18510 & n18512 ) | ( ~n18511 & n18512 ) ;
  assign n18514 = ( n17919 & ~n18226 ) | ( n17919 & n18239 ) | ( ~n18226 & n18239 ) ;
  assign n18515 = x93 & n8834 ;
  assign n18516 = x92 & n8829 ;
  assign n18517 = x91 & ~n8828 ;
  assign n18518 = n9159 & n18517 ;
  assign n18519 = n18516 | n18518 ;
  assign n18520 = n18515 | n18519 ;
  assign n18521 = n8837 | n18520 ;
  assign n18522 = ( n2931 & n18520 ) | ( n2931 & n18521 ) | ( n18520 & n18521 ) ;
  assign n18523 = x53 & n18522 ;
  assign n18524 = x53 & ~n18523 ;
  assign n18525 = ( n18522 & ~n18523 ) | ( n18522 & n18524 ) | ( ~n18523 & n18524 ) ;
  assign n18526 = n18188 | n18201 ;
  assign n18527 = x81 & n12808 ;
  assign n18528 = x63 & x80 ;
  assign n18529 = ~n12808 & n18528 ;
  assign n18530 = n18527 | n18529 ;
  assign n18531 = ~n18185 & n18530 ;
  assign n18532 = x84 & n11984 ;
  assign n18533 = x83 & n11979 ;
  assign n18534 = x82 & ~n11978 ;
  assign n18535 = n12430 & n18534 ;
  assign n18536 = n18533 | n18535 ;
  assign n18537 = n18532 | n18536 ;
  assign n18538 = n11987 | n18537 ;
  assign n18539 = ( n1537 & n18537 ) | ( n1537 & n18538 ) | ( n18537 & n18538 ) ;
  assign n18540 = ~x62 & n18539 ;
  assign n18541 = x62 & ~n18539 ;
  assign n18542 = n18540 | n18541 ;
  assign n18543 = ( n18185 & ~n18530 ) | ( n18185 & n18542 ) | ( ~n18530 & n18542 ) ;
  assign n18544 = n18531 | n18543 ;
  assign n18545 = ~n18526 & n18544 ;
  assign n18546 = n18185 & ~n18530 ;
  assign n18547 = ( n18531 & n18542 ) | ( n18531 & n18546 ) | ( n18542 & n18546 ) ;
  assign n18548 = n18545 & ~n18547 ;
  assign n18549 = ( n18526 & ~n18544 ) | ( n18526 & n18547 ) | ( ~n18544 & n18547 ) ;
  assign n18550 = n18548 | n18549 ;
  assign n18551 = x87 & n10876 ;
  assign n18552 = x86 & n10871 ;
  assign n18553 = x85 & ~n10870 ;
  assign n18554 = n11305 & n18553 ;
  assign n18555 = n18552 | n18554 ;
  assign n18556 = n18551 | n18555 ;
  assign n18557 = n10879 | n18556 ;
  assign n18558 = ( n2067 & n18556 ) | ( n2067 & n18557 ) | ( n18556 & n18557 ) ;
  assign n18559 = x59 & n18558 ;
  assign n18560 = x59 & ~n18559 ;
  assign n18561 = ( n18558 & ~n18559 ) | ( n18558 & n18560 ) | ( ~n18559 & n18560 ) ;
  assign n18562 = n18550 & ~n18561 ;
  assign n18563 = ~n18550 & n18561 ;
  assign n18564 = n18562 | n18563 ;
  assign n18565 = n18205 & ~n18564 ;
  assign n18566 = ~n18205 & n18564 ;
  assign n18567 = n18565 | n18566 ;
  assign n18568 = x90 & n9853 ;
  assign n18569 = x89 & n9848 ;
  assign n18570 = x88 & ~n9847 ;
  assign n18571 = n10165 & n18570 ;
  assign n18572 = n18569 | n18571 ;
  assign n18573 = n18568 | n18572 ;
  assign n18574 = n9856 | n18573 ;
  assign n18575 = ( n2410 & n18573 ) | ( n2410 & n18574 ) | ( n18573 & n18574 ) ;
  assign n18576 = x56 & n18575 ;
  assign n18577 = x56 & ~n18576 ;
  assign n18578 = ( n18575 & ~n18576 ) | ( n18575 & n18577 ) | ( ~n18576 & n18577 ) ;
  assign n18579 = ~n18567 & n18578 ;
  assign n18580 = n18567 & ~n18578 ;
  assign n18581 = n18579 | n18580 ;
  assign n18582 = ( n18223 & n18525 ) | ( n18223 & ~n18581 ) | ( n18525 & ~n18581 ) ;
  assign n18583 = ( ~n18223 & n18581 ) | ( ~n18223 & n18582 ) | ( n18581 & n18582 ) ;
  assign n18584 = ( ~n18525 & n18582 ) | ( ~n18525 & n18583 ) | ( n18582 & n18583 ) ;
  assign n18585 = ( n18513 & ~n18514 ) | ( n18513 & n18584 ) | ( ~n18514 & n18584 ) ;
  assign n18586 = ( n18514 & ~n18584 ) | ( n18514 & n18585 ) | ( ~n18584 & n18585 ) ;
  assign n18587 = ( ~n18513 & n18585 ) | ( ~n18513 & n18586 ) | ( n18585 & n18586 ) ;
  assign n18588 = ( n18169 & n18253 ) | ( n18169 & n18256 ) | ( n18253 & n18256 ) ;
  assign n18589 = n18587 & ~n18588 ;
  assign n18590 = ~n18587 & n18588 ;
  assign n18591 = n18589 | n18590 ;
  assign n18592 = x99 & n6937 ;
  assign n18593 = x98 & n6932 ;
  assign n18594 = x97 & ~n6931 ;
  assign n18595 = n7216 & n18594 ;
  assign n18596 = n18593 | n18595 ;
  assign n18597 = n18592 | n18596 ;
  assign n18598 = n6940 | n18597 ;
  assign n18599 = ( n4325 & n18597 ) | ( n4325 & n18598 ) | ( n18597 & n18598 ) ;
  assign n18600 = x47 & n18599 ;
  assign n18601 = x47 & ~n18600 ;
  assign n18602 = ( n18599 & ~n18600 ) | ( n18599 & n18601 ) | ( ~n18600 & n18601 ) ;
  assign n18603 = n18591 & n18602 ;
  assign n18604 = ( ~n18587 & n18588 ) | ( ~n18587 & n18602 ) | ( n18588 & n18602 ) ;
  assign n18605 = n18589 | n18604 ;
  assign n18606 = ~n18603 & n18605 ;
  assign n18607 = n18259 & ~n18273 ;
  assign n18608 = ( n18502 & n18606 ) | ( n18502 & ~n18607 ) | ( n18606 & ~n18607 ) ;
  assign n18609 = ( ~n18606 & n18607 ) | ( ~n18606 & n18608 ) | ( n18607 & n18608 ) ;
  assign n18610 = ( ~n18502 & n18608 ) | ( ~n18502 & n18609 ) | ( n18608 & n18609 ) ;
  assign n18611 = n18491 & n18610 ;
  assign n18612 = n18491 | n18610 ;
  assign n18613 = ~n18611 & n18612 ;
  assign n18614 = x105 & n5340 ;
  assign n18615 = x104 & n5335 ;
  assign n18616 = x103 & ~n5334 ;
  assign n18617 = n5580 & n18616 ;
  assign n18618 = n18615 | n18617 ;
  assign n18619 = n18614 | n18618 ;
  assign n18620 = n5343 | n18619 ;
  assign n18621 = ( n5788 & n18619 ) | ( n5788 & n18620 ) | ( n18619 & n18620 ) ;
  assign n18622 = x41 & n18621 ;
  assign n18623 = x41 & ~n18622 ;
  assign n18624 = ( n18621 & ~n18622 ) | ( n18621 & n18623 ) | ( ~n18622 & n18623 ) ;
  assign n18625 = n18613 & n18624 ;
  assign n18626 = n18613 | n18624 ;
  assign n18627 = ~n18625 & n18626 ;
  assign n18628 = n18304 & n18627 ;
  assign n18629 = n18304 | n18627 ;
  assign n18630 = ~n18628 & n18629 ;
  assign n18631 = x108 & n4572 ;
  assign n18632 = x107 & n4567 ;
  assign n18633 = x106 & ~n4566 ;
  assign n18634 = n4828 & n18633 ;
  assign n18635 = n18632 | n18634 ;
  assign n18636 = n18631 | n18635 ;
  assign n18637 = n4575 | n18636 ;
  assign n18638 = ( n6358 & n18636 ) | ( n6358 & n18637 ) | ( n18636 & n18637 ) ;
  assign n18639 = x38 & n18638 ;
  assign n18640 = x38 & ~n18639 ;
  assign n18641 = ( n18638 & ~n18639 ) | ( n18638 & n18640 ) | ( ~n18639 & n18640 ) ;
  assign n18642 = n18630 & n18641 ;
  assign n18643 = n18630 | n18641 ;
  assign n18644 = ~n18642 & n18643 ;
  assign n18645 = x111 & n3913 ;
  assign n18646 = x110 & n3908 ;
  assign n18647 = x109 & ~n3907 ;
  assign n18648 = n4152 & n18647 ;
  assign n18649 = n18646 | n18648 ;
  assign n18650 = n18645 | n18649 ;
  assign n18651 = n3916 | n18650 ;
  assign n18652 = ( n7492 & n18650 ) | ( n7492 & n18651 ) | ( n18650 & n18651 ) ;
  assign n18653 = x35 & n18652 ;
  assign n18654 = x35 & ~n18653 ;
  assign n18655 = ( n18652 & ~n18653 ) | ( n18652 & n18654 ) | ( ~n18653 & n18654 ) ;
  assign n18656 = ( n18490 & n18644 ) | ( n18490 & n18655 ) | ( n18644 & n18655 ) ;
  assign n18657 = ( n18644 & n18655 ) | ( n18644 & ~n18656 ) | ( n18655 & ~n18656 ) ;
  assign n18658 = ( n18490 & ~n18656 ) | ( n18490 & n18657 ) | ( ~n18656 & n18657 ) ;
  assign n18659 = ( n18473 & ~n18489 ) | ( n18473 & n18658 ) | ( ~n18489 & n18658 ) ;
  assign n18660 = ( n18489 & ~n18658 ) | ( n18489 & n18659 ) | ( ~n18658 & n18659 ) ;
  assign n18661 = ( ~n18473 & n18659 ) | ( ~n18473 & n18660 ) | ( n18659 & n18660 ) ;
  assign n18662 = ( n18441 & ~n18458 ) | ( n18441 & n18661 ) | ( ~n18458 & n18661 ) ;
  assign n18663 = ( n18458 & ~n18661 ) | ( n18458 & n18662 ) | ( ~n18661 & n18662 ) ;
  assign n18664 = ( ~n18441 & n18662 ) | ( ~n18441 & n18663 ) | ( n18662 & n18663 ) ;
  assign n18665 = n18421 | n18664 ;
  assign n18666 = n18421 & n18664 ;
  assign n18667 = n18665 & ~n18666 ;
  assign n18668 = ~n18396 & n18404 ;
  assign n18669 = n18667 | n18668 ;
  assign n18670 = n18406 | n18669 ;
  assign n18671 = ( n18406 & n18667 ) | ( n18406 & n18668 ) | ( n18667 & n18668 ) ;
  assign n18672 = n18670 & ~n18671 ;
  assign n18673 = n18395 & n18672 ;
  assign n18674 = n18395 & ~n18673 ;
  assign n18675 = n18382 | n18388 ;
  assign n18676 = n18382 | n18389 ;
  assign n18677 = ( n17506 & n18675 ) | ( n17506 & n18676 ) | ( n18675 & n18676 ) ;
  assign n18678 = ~n18395 & n18672 ;
  assign n18679 = n18677 | n18678 ;
  assign n18680 = n18674 | n18679 ;
  assign n18681 = n18674 | n18678 ;
  assign n18682 = n18675 & n18681 ;
  assign n18683 = n18676 & n18681 ;
  assign n18684 = ( n17506 & n18682 ) | ( n17506 & n18683 ) | ( n18682 & n18683 ) ;
  assign n18685 = n18680 & ~n18684 ;
  assign n18686 = n18405 | n18671 ;
  assign n18687 = x127 & n1421 ;
  assign n18688 = x126 & n1416 ;
  assign n18689 = x125 & ~n1415 ;
  assign n18690 = n1584 & n18689 ;
  assign n18691 = n18688 | n18690 ;
  assign n18692 = n18687 | n18691 ;
  assign n18693 = n1424 | n18692 ;
  assign n18694 = ( n12720 & n18692 ) | ( n12720 & n18693 ) | ( n18692 & n18693 ) ;
  assign n18695 = x20 & n18694 ;
  assign n18696 = x20 & ~n18695 ;
  assign n18697 = ( n18694 & ~n18695 ) | ( n18694 & n18696 ) | ( ~n18695 & n18696 ) ;
  assign n18698 = n18420 | n18666 ;
  assign n18699 = x118 & n2775 ;
  assign n18700 = x117 & n2770 ;
  assign n18701 = x116 & ~n2769 ;
  assign n18702 = n2978 & n18701 ;
  assign n18703 = n18700 | n18702 ;
  assign n18704 = n18699 | n18703 ;
  assign n18705 = n2778 | n18704 ;
  assign n18706 = ( n9760 & n18704 ) | ( n9760 & n18705 ) | ( n18704 & n18705 ) ;
  assign n18707 = x29 & n18706 ;
  assign n18708 = x29 & ~n18707 ;
  assign n18709 = ( n18706 & ~n18707 ) | ( n18706 & n18708 ) | ( ~n18707 & n18708 ) ;
  assign n18710 = ( n18434 & n18484 ) | ( n18434 & n18485 ) | ( n18484 & n18485 ) ;
  assign n18711 = n18473 & n18658 ;
  assign n18712 = ~n18710 & n18711 ;
  assign n18713 = n18473 | n18658 ;
  assign n18714 = ( n18487 & n18488 ) | ( n18487 & n18713 ) | ( n18488 & n18713 ) ;
  assign n18715 = ( n18710 & ~n18712 ) | ( n18710 & n18714 ) | ( ~n18712 & n18714 ) ;
  assign n18716 = n18709 & n18715 ;
  assign n18717 = n18709 | n18715 ;
  assign n18718 = ~n18716 & n18717 ;
  assign n18719 = x106 & n5340 ;
  assign n18720 = x105 & n5335 ;
  assign n18721 = x104 & ~n5334 ;
  assign n18722 = n5580 & n18721 ;
  assign n18723 = n18720 | n18722 ;
  assign n18724 = n18719 | n18723 ;
  assign n18725 = n5343 | n18724 ;
  assign n18726 = ( n5814 & n18724 ) | ( n5814 & n18725 ) | ( n18724 & n18725 ) ;
  assign n18727 = x41 & n18726 ;
  assign n18728 = x41 & ~n18727 ;
  assign n18729 = ( n18726 & ~n18727 ) | ( n18726 & n18728 ) | ( ~n18727 & n18728 ) ;
  assign n18730 = ( ~n18502 & n18606 ) | ( ~n18502 & n18607 ) | ( n18606 & n18607 ) ;
  assign n18731 = x85 & n11984 ;
  assign n18732 = x84 & n11979 ;
  assign n18733 = x83 & ~n11978 ;
  assign n18734 = n12430 & n18733 ;
  assign n18735 = n18732 | n18734 ;
  assign n18736 = n18731 | n18735 ;
  assign n18737 = n11987 | n18736 ;
  assign n18738 = ( n1765 & n18736 ) | ( n1765 & n18737 ) | ( n18736 & n18737 ) ;
  assign n18739 = ~x62 & n18738 ;
  assign n18740 = x62 & ~n18738 ;
  assign n18741 = n18739 | n18740 ;
  assign n18742 = x82 & n12808 ;
  assign n18743 = x63 & x81 ;
  assign n18744 = ~n12808 & n18743 ;
  assign n18745 = n18742 | n18744 ;
  assign n18746 = ~x17 & n18745 ;
  assign n18747 = x17 & ~n18745 ;
  assign n18748 = n18746 | n18747 ;
  assign n18749 = n18530 & ~n18748 ;
  assign n18750 = ~n18530 & n18748 ;
  assign n18751 = n18749 | n18750 ;
  assign n18752 = n18741 & ~n18751 ;
  assign n18753 = ~n18741 & n18751 ;
  assign n18754 = n18752 | n18753 ;
  assign n18755 = n18543 | n18754 ;
  assign n18756 = n18543 & n18754 ;
  assign n18757 = x88 & n10876 ;
  assign n18758 = x87 & n10871 ;
  assign n18759 = x86 & ~n10870 ;
  assign n18760 = n11305 & n18759 ;
  assign n18761 = n18758 | n18760 ;
  assign n18762 = n18757 | n18761 ;
  assign n18763 = n10879 | n18762 ;
  assign n18764 = ( n2095 & n18762 ) | ( n2095 & n18763 ) | ( n18762 & n18763 ) ;
  assign n18765 = x59 & n18764 ;
  assign n18766 = x59 & ~n18765 ;
  assign n18767 = ( n18764 & ~n18765 ) | ( n18764 & n18766 ) | ( ~n18765 & n18766 ) ;
  assign n18768 = n18756 | n18767 ;
  assign n18769 = n18755 & ~n18768 ;
  assign n18770 = ( ~n18755 & n18756 ) | ( ~n18755 & n18767 ) | ( n18756 & n18767 ) ;
  assign n18771 = n18769 | n18770 ;
  assign n18772 = n18549 | n18563 ;
  assign n18773 = ~n18771 & n18772 ;
  assign n18774 = n18771 & ~n18772 ;
  assign n18775 = n18773 | n18774 ;
  assign n18776 = x91 & n9853 ;
  assign n18777 = x90 & n9848 ;
  assign n18778 = x89 & ~n9847 ;
  assign n18779 = n10165 & n18778 ;
  assign n18780 = n18777 | n18779 ;
  assign n18781 = n18776 | n18780 ;
  assign n18782 = n9856 | n18781 ;
  assign n18783 = ( n2714 & n18781 ) | ( n2714 & n18782 ) | ( n18781 & n18782 ) ;
  assign n18784 = x56 & n18783 ;
  assign n18785 = x56 & ~n18784 ;
  assign n18786 = ( n18783 & ~n18784 ) | ( n18783 & n18785 ) | ( ~n18784 & n18785 ) ;
  assign n18787 = ~n18775 & n18786 ;
  assign n18788 = n18775 | n18787 ;
  assign n18789 = n18775 & n18786 ;
  assign n18790 = n18565 | n18579 ;
  assign n18791 = n18789 | n18790 ;
  assign n18792 = n18788 & ~n18791 ;
  assign n18793 = ( ~n18788 & n18789 ) | ( ~n18788 & n18790 ) | ( n18789 & n18790 ) ;
  assign n18794 = n18792 | n18793 ;
  assign n18795 = x94 & n8834 ;
  assign n18796 = x93 & n8829 ;
  assign n18797 = x92 & ~n8828 ;
  assign n18798 = n9159 & n18797 ;
  assign n18799 = n18796 | n18798 ;
  assign n18800 = n18795 | n18799 ;
  assign n18801 = n8837 | n18800 ;
  assign n18802 = ( n3271 & n18800 ) | ( n3271 & n18801 ) | ( n18800 & n18801 ) ;
  assign n18803 = x53 & n18802 ;
  assign n18804 = x53 & ~n18803 ;
  assign n18805 = ( n18802 & ~n18803 ) | ( n18802 & n18804 ) | ( ~n18803 & n18804 ) ;
  assign n18806 = ~n18794 & n18805 ;
  assign n18807 = n18794 | n18806 ;
  assign n18808 = n18794 & n18805 ;
  assign n18809 = n18582 | n18808 ;
  assign n18810 = n18807 & ~n18809 ;
  assign n18811 = ( n18582 & ~n18807 ) | ( n18582 & n18808 ) | ( ~n18807 & n18808 ) ;
  assign n18812 = n18810 | n18811 ;
  assign n18813 = n18514 & ~n18584 ;
  assign n18814 = x97 & n7812 ;
  assign n18815 = x96 & n7807 ;
  assign n18816 = x95 & ~n7806 ;
  assign n18817 = n8136 & n18816 ;
  assign n18818 = n18815 | n18817 ;
  assign n18819 = n18814 | n18818 ;
  assign n18820 = n7815 | n18819 ;
  assign n18821 = ( n3707 & n18819 ) | ( n3707 & n18820 ) | ( n18819 & n18820 ) ;
  assign n18822 = x50 & n18821 ;
  assign n18823 = x50 & ~n18822 ;
  assign n18824 = ( n18821 & ~n18822 ) | ( n18821 & n18823 ) | ( ~n18822 & n18823 ) ;
  assign n18825 = n18813 | n18824 ;
  assign n18826 = n18514 & n18584 ;
  assign n18827 = ( n18513 & n18587 ) | ( n18513 & n18826 ) | ( n18587 & n18826 ) ;
  assign n18828 = n18825 | n18827 ;
  assign n18829 = ( n18813 & n18824 ) | ( n18813 & n18827 ) | ( n18824 & n18827 ) ;
  assign n18830 = n18828 & ~n18829 ;
  assign n18831 = n18812 & n18830 ;
  assign n18832 = n18812 | n18830 ;
  assign n18833 = ~n18831 & n18832 ;
  assign n18834 = x100 & n6937 ;
  assign n18835 = x99 & n6932 ;
  assign n18836 = x98 & ~n6931 ;
  assign n18837 = n7216 & n18836 ;
  assign n18838 = n18835 | n18837 ;
  assign n18839 = n18834 | n18838 ;
  assign n18840 = n6940 | n18839 ;
  assign n18841 = ( n4532 & n18839 ) | ( n4532 & n18840 ) | ( n18839 & n18840 ) ;
  assign n18842 = x47 & n18841 ;
  assign n18843 = x47 & ~n18842 ;
  assign n18844 = ( n18841 & ~n18842 ) | ( n18841 & n18843 ) | ( ~n18842 & n18843 ) ;
  assign n18845 = ~n18833 & n18844 ;
  assign n18846 = n18833 & ~n18844 ;
  assign n18847 = n18845 | n18846 ;
  assign n18848 = ~n18604 & n18847 ;
  assign n18849 = n18604 & ~n18847 ;
  assign n18850 = n18848 | n18849 ;
  assign n18851 = x103 & n6068 ;
  assign n18852 = x102 & n6063 ;
  assign n18853 = x101 & ~n6062 ;
  assign n18854 = n6398 & n18853 ;
  assign n18855 = n18852 | n18854 ;
  assign n18856 = n18851 | n18855 ;
  assign n18857 = n6071 | n18856 ;
  assign n18858 = ( n5264 & n18856 ) | ( n5264 & n18857 ) | ( n18856 & n18857 ) ;
  assign n18859 = x44 & n18858 ;
  assign n18860 = x44 & ~n18859 ;
  assign n18861 = ( n18858 & ~n18859 ) | ( n18858 & n18860 ) | ( ~n18859 & n18860 ) ;
  assign n18862 = ( n18730 & n18850 ) | ( n18730 & ~n18861 ) | ( n18850 & ~n18861 ) ;
  assign n18863 = ( ~n18850 & n18861 ) | ( ~n18850 & n18862 ) | ( n18861 & n18862 ) ;
  assign n18864 = ( ~n18730 & n18862 ) | ( ~n18730 & n18863 ) | ( n18862 & n18863 ) ;
  assign n18865 = n18729 & n18864 ;
  assign n18866 = n18729 | n18864 ;
  assign n18867 = ~n18865 & n18866 ;
  assign n18868 = n18611 | n18625 ;
  assign n18869 = n18867 | n18868 ;
  assign n18870 = n18867 & n18868 ;
  assign n18871 = n18869 & ~n18870 ;
  assign n18872 = x109 & n4572 ;
  assign n18873 = x108 & n4567 ;
  assign n18874 = x107 & ~n4566 ;
  assign n18875 = n4828 & n18874 ;
  assign n18876 = n18873 | n18875 ;
  assign n18877 = n18872 | n18876 ;
  assign n18878 = n4575 | n18877 ;
  assign n18879 = ( n6884 & n18877 ) | ( n6884 & n18878 ) | ( n18877 & n18878 ) ;
  assign n18880 = x38 & n18879 ;
  assign n18881 = x38 & ~n18880 ;
  assign n18882 = ( n18879 & ~n18880 ) | ( n18879 & n18881 ) | ( ~n18880 & n18881 ) ;
  assign n18883 = n18871 & n18882 ;
  assign n18884 = n18871 & ~n18883 ;
  assign n18885 = ~n18871 & n18882 ;
  assign n18886 = n18628 | n18642 ;
  assign n18887 = n18885 | n18886 ;
  assign n18888 = n18884 | n18887 ;
  assign n18889 = ( n18884 & n18885 ) | ( n18884 & n18886 ) | ( n18885 & n18886 ) ;
  assign n18890 = n18888 & ~n18889 ;
  assign n18891 = x112 & n3913 ;
  assign n18892 = x111 & n3908 ;
  assign n18893 = x110 & ~n3907 ;
  assign n18894 = n4152 & n18893 ;
  assign n18895 = n18892 | n18894 ;
  assign n18896 = n18891 | n18895 ;
  assign n18897 = n3916 | n18896 ;
  assign n18898 = ( n7789 & n18896 ) | ( n7789 & n18897 ) | ( n18896 & n18897 ) ;
  assign n18899 = x35 & n18898 ;
  assign n18900 = x35 & ~n18899 ;
  assign n18901 = ( n18898 & ~n18899 ) | ( n18898 & n18900 ) | ( ~n18899 & n18900 ) ;
  assign n18902 = n18890 & n18901 ;
  assign n18903 = n18890 & ~n18902 ;
  assign n18904 = ~n18890 & n18901 ;
  assign n18905 = n18656 | n18904 ;
  assign n18906 = n18903 | n18905 ;
  assign n18907 = ( n18656 & n18903 ) | ( n18656 & n18904 ) | ( n18903 & n18904 ) ;
  assign n18908 = n18906 & ~n18907 ;
  assign n18909 = x115 & n3314 ;
  assign n18910 = x114 & n3309 ;
  assign n18911 = x113 & ~n3308 ;
  assign n18912 = n3570 & n18911 ;
  assign n18913 = n18910 | n18912 ;
  assign n18914 = n18909 | n18913 ;
  assign n18915 = n3317 | n18914 ;
  assign n18916 = ( n8749 & n18914 ) | ( n8749 & n18915 ) | ( n18914 & n18915 ) ;
  assign n18917 = x32 & n18916 ;
  assign n18918 = x32 & ~n18917 ;
  assign n18919 = ( n18916 & ~n18917 ) | ( n18916 & n18918 ) | ( ~n18917 & n18918 ) ;
  assign n18920 = n18472 | n18711 ;
  assign n18921 = ( n18908 & n18919 ) | ( n18908 & ~n18920 ) | ( n18919 & ~n18920 ) ;
  assign n18922 = ( ~n18919 & n18920 ) | ( ~n18919 & n18921 ) | ( n18920 & n18921 ) ;
  assign n18923 = ( ~n18908 & n18921 ) | ( ~n18908 & n18922 ) | ( n18921 & n18922 ) ;
  assign n18924 = n18718 & n18923 ;
  assign n18925 = n18718 & ~n18924 ;
  assign n18926 = n18923 & ~n18924 ;
  assign n18927 = n18925 | n18926 ;
  assign n18928 = x121 & n2280 ;
  assign n18929 = x120 & n2275 ;
  assign n18930 = x119 & ~n2274 ;
  assign n18931 = n2481 & n18930 ;
  assign n18932 = n18929 | n18931 ;
  assign n18933 = n18928 | n18932 ;
  assign n18934 = n2283 | n18933 ;
  assign n18935 = ( n10811 & n18933 ) | ( n10811 & n18934 ) | ( n18933 & n18934 ) ;
  assign n18936 = x26 & n18935 ;
  assign n18937 = x26 & ~n18936 ;
  assign n18938 = ( n18935 & ~n18936 ) | ( n18935 & n18937 ) | ( ~n18936 & n18937 ) ;
  assign n18939 = n18441 & n18661 ;
  assign n18940 = n18439 | n18939 ;
  assign n18941 = ( n18927 & n18938 ) | ( n18927 & ~n18940 ) | ( n18938 & ~n18940 ) ;
  assign n18942 = ( ~n18938 & n18940 ) | ( ~n18938 & n18941 ) | ( n18940 & n18941 ) ;
  assign n18943 = ( ~n18927 & n18941 ) | ( ~n18927 & n18942 ) | ( n18941 & n18942 ) ;
  assign n18944 = x124 & n1817 ;
  assign n18945 = x123 & n1812 ;
  assign n18946 = x122 & ~n1811 ;
  assign n18947 = n1977 & n18946 ;
  assign n18948 = n18945 | n18947 ;
  assign n18949 = n18944 | n18948 ;
  assign n18950 = n1820 | n18949 ;
  assign n18951 = ( n11916 & n18949 ) | ( n11916 & n18950 ) | ( n18949 & n18950 ) ;
  assign n18952 = x23 & n18951 ;
  assign n18953 = x23 & ~n18952 ;
  assign n18954 = ( n18951 & ~n18952 ) | ( n18951 & n18953 ) | ( ~n18952 & n18953 ) ;
  assign n18955 = ( n18442 & n18453 ) | ( n18442 & n18454 ) | ( n18453 & n18454 ) ;
  assign n18956 = n18939 & ~n18955 ;
  assign n18957 = n18441 | n18661 ;
  assign n18958 = ( n18456 & n18457 ) | ( n18456 & n18957 ) | ( n18457 & n18957 ) ;
  assign n18959 = ( n18955 & ~n18956 ) | ( n18955 & n18958 ) | ( ~n18956 & n18958 ) ;
  assign n18960 = ( n18943 & n18954 ) | ( n18943 & ~n18959 ) | ( n18954 & ~n18959 ) ;
  assign n18961 = ( ~n18954 & n18959 ) | ( ~n18954 & n18960 ) | ( n18959 & n18960 ) ;
  assign n18962 = ( ~n18943 & n18960 ) | ( ~n18943 & n18961 ) | ( n18960 & n18961 ) ;
  assign n18963 = ( n18697 & ~n18698 ) | ( n18697 & n18962 ) | ( ~n18698 & n18962 ) ;
  assign n18964 = ( n18698 & ~n18962 ) | ( n18698 & n18963 ) | ( ~n18962 & n18963 ) ;
  assign n18965 = ( ~n18697 & n18963 ) | ( ~n18697 & n18964 ) | ( n18963 & n18964 ) ;
  assign n18966 = ~n18686 & n18965 ;
  assign n18967 = n18673 | n18682 ;
  assign n18968 = n18686 & n18965 ;
  assign n18969 = n18686 & ~n18968 ;
  assign n18970 = n18966 | n18969 ;
  assign n18971 = n18967 & n18970 ;
  assign n18972 = n18673 | n18683 ;
  assign n18973 = n18970 & n18972 ;
  assign n18974 = ( n17506 & n18971 ) | ( n17506 & n18973 ) | ( n18971 & n18973 ) ;
  assign n18975 = ( n17506 & n18967 ) | ( n17506 & n18972 ) | ( n18967 & n18972 ) ;
  assign n18976 = ( n18686 & ~n18965 ) | ( n18686 & n18975 ) | ( ~n18965 & n18975 ) ;
  assign n18977 = ( n18966 & ~n18974 ) | ( n18966 & n18976 ) | ( ~n18974 & n18976 ) ;
  assign n18978 = ( n18943 & n18954 ) | ( n18943 & n18959 ) | ( n18954 & n18959 ) ;
  assign n18979 = x127 & n1416 ;
  assign n18980 = x126 & ~n1415 ;
  assign n18981 = n1584 & n18980 ;
  assign n18982 = n18979 | n18981 ;
  assign n18983 = n1424 | n18982 ;
  assign n18984 = ( n13461 & n18982 ) | ( n13461 & n18983 ) | ( n18982 & n18983 ) ;
  assign n18985 = x20 & n18984 ;
  assign n18986 = x20 & ~n18985 ;
  assign n18987 = ( n18984 & ~n18985 ) | ( n18984 & n18986 ) | ( ~n18985 & n18986 ) ;
  assign n18988 = n18978 & n18987 ;
  assign n18989 = n18978 & ~n18988 ;
  assign n18990 = ~n18978 & n18987 ;
  assign n18991 = x122 & n2280 ;
  assign n18992 = x121 & n2275 ;
  assign n18993 = x120 & ~n2274 ;
  assign n18994 = n2481 & n18993 ;
  assign n18995 = n18992 | n18994 ;
  assign n18996 = n18991 | n18995 ;
  assign n18997 = n2283 | n18996 ;
  assign n18998 = ( n11188 & n18996 ) | ( n11188 & n18997 ) | ( n18996 & n18997 ) ;
  assign n18999 = x26 & n18998 ;
  assign n19000 = x26 & ~n18999 ;
  assign n19001 = ( n18998 & ~n18999 ) | ( n18998 & n19000 ) | ( ~n18999 & n19000 ) ;
  assign n19002 = n18716 | n19001 ;
  assign n19003 = n18924 | n19002 ;
  assign n19004 = ( n18716 & n18924 ) | ( n18716 & n19001 ) | ( n18924 & n19001 ) ;
  assign n19005 = n19003 & ~n19004 ;
  assign n19006 = x113 & n3913 ;
  assign n19007 = x112 & n3908 ;
  assign n19008 = x111 & ~n3907 ;
  assign n19009 = n4152 & n19008 ;
  assign n19010 = n19007 | n19009 ;
  assign n19011 = n19006 | n19010 ;
  assign n19012 = n3916 | n19011 ;
  assign n19013 = ( n8113 & n19011 ) | ( n8113 & n19012 ) | ( n19011 & n19012 ) ;
  assign n19014 = x35 & n19013 ;
  assign n19015 = x35 & ~n19014 ;
  assign n19016 = ( n19013 & ~n19014 ) | ( n19013 & n19015 ) | ( ~n19014 & n19015 ) ;
  assign n19017 = n18883 | n18889 ;
  assign n19018 = x110 & n4572 ;
  assign n19019 = x109 & n4567 ;
  assign n19020 = x108 & ~n4566 ;
  assign n19021 = n4828 & n19020 ;
  assign n19022 = n19019 | n19021 ;
  assign n19023 = n19018 | n19022 ;
  assign n19024 = n4575 | n19023 ;
  assign n19025 = ( n7189 & n19023 ) | ( n7189 & n19024 ) | ( n19023 & n19024 ) ;
  assign n19026 = x38 & n19025 ;
  assign n19027 = x38 & ~n19026 ;
  assign n19028 = ( n19025 & ~n19026 ) | ( n19025 & n19027 ) | ( ~n19026 & n19027 ) ;
  assign n19029 = n18806 | n18811 ;
  assign n19030 = x95 & n8834 ;
  assign n19031 = x94 & n8829 ;
  assign n19032 = x93 & ~n8828 ;
  assign n19033 = n9159 & n19032 ;
  assign n19034 = n19031 | n19033 ;
  assign n19035 = n19030 | n19034 ;
  assign n19036 = n8837 | n19035 ;
  assign n19037 = ( n3479 & n19035 ) | ( n3479 & n19036 ) | ( n19035 & n19036 ) ;
  assign n19038 = x53 & n19037 ;
  assign n19039 = x53 & ~n19038 ;
  assign n19040 = ( n19037 & ~n19038 ) | ( n19037 & n19039 ) | ( ~n19038 & n19039 ) ;
  assign n19041 = n18787 | n18793 ;
  assign n19042 = x92 & n9853 ;
  assign n19043 = x91 & n9848 ;
  assign n19044 = x90 & ~n9847 ;
  assign n19045 = n10165 & n19044 ;
  assign n19046 = n19043 | n19045 ;
  assign n19047 = n19042 | n19046 ;
  assign n19048 = n9856 | n19047 ;
  assign n19049 = ( n2904 & n19047 ) | ( n2904 & n19048 ) | ( n19047 & n19048 ) ;
  assign n19050 = x56 & n19049 ;
  assign n19051 = x56 & ~n19050 ;
  assign n19052 = ( n19049 & ~n19050 ) | ( n19049 & n19051 ) | ( ~n19050 & n19051 ) ;
  assign n19053 = n18770 | n18773 ;
  assign n19054 = x89 & n10876 ;
  assign n19055 = x88 & n10871 ;
  assign n19056 = x87 & ~n10870 ;
  assign n19057 = n11305 & n19056 ;
  assign n19058 = n19055 | n19057 ;
  assign n19059 = n19054 | n19058 ;
  assign n19060 = n10879 | n19059 ;
  assign n19061 = ( n2244 & n19059 ) | ( n2244 & n19060 ) | ( n19059 & n19060 ) ;
  assign n19062 = x59 & n19061 ;
  assign n19063 = x59 & ~n19062 ;
  assign n19064 = ( n19061 & ~n19062 ) | ( n19061 & n19063 ) | ( ~n19062 & n19063 ) ;
  assign n19065 = x86 & n11984 ;
  assign n19066 = x85 & n11979 ;
  assign n19067 = x84 & ~n11978 ;
  assign n19068 = n12430 & n19067 ;
  assign n19069 = n19066 | n19068 ;
  assign n19070 = n19065 | n19069 ;
  assign n19071 = n11987 | n19070 ;
  assign n19072 = ( n1921 & n19070 ) | ( n1921 & n19071 ) | ( n19070 & n19071 ) ;
  assign n19073 = ~x62 & n19072 ;
  assign n19074 = x83 & n12808 ;
  assign n19075 = x63 & x82 ;
  assign n19076 = ~n12808 & n19075 ;
  assign n19077 = n19074 | n19076 ;
  assign n19078 = n18746 | n18749 ;
  assign n19079 = n19077 & ~n19078 ;
  assign n19080 = ~n19077 & n19078 ;
  assign n19081 = n19079 | n19080 ;
  assign n19082 = x62 & ~n19072 ;
  assign n19083 = n19081 & ~n19082 ;
  assign n19084 = ~n19073 & n19083 ;
  assign n19085 = ( n19073 & ~n19081 ) | ( n19073 & n19082 ) | ( ~n19081 & n19082 ) ;
  assign n19086 = n19084 | n19085 ;
  assign n19087 = ( n18752 & ~n18754 ) | ( n18752 & n18755 ) | ( ~n18754 & n18755 ) ;
  assign n19088 = ( n19064 & n19086 ) | ( n19064 & ~n19087 ) | ( n19086 & ~n19087 ) ;
  assign n19089 = ( ~n19086 & n19087 ) | ( ~n19086 & n19088 ) | ( n19087 & n19088 ) ;
  assign n19090 = ( ~n19064 & n19088 ) | ( ~n19064 & n19089 ) | ( n19088 & n19089 ) ;
  assign n19091 = ( n19052 & ~n19053 ) | ( n19052 & n19090 ) | ( ~n19053 & n19090 ) ;
  assign n19092 = ( n19052 & n19053 ) | ( n19052 & ~n19090 ) | ( n19053 & ~n19090 ) ;
  assign n19093 = ( ~n19052 & n19091 ) | ( ~n19052 & n19092 ) | ( n19091 & n19092 ) ;
  assign n19094 = ( n19040 & ~n19041 ) | ( n19040 & n19093 ) | ( ~n19041 & n19093 ) ;
  assign n19095 = ( n19041 & ~n19093 ) | ( n19041 & n19094 ) | ( ~n19093 & n19094 ) ;
  assign n19096 = ( ~n19040 & n19094 ) | ( ~n19040 & n19095 ) | ( n19094 & n19095 ) ;
  assign n19097 = ~n19029 & n19096 ;
  assign n19098 = n19029 & ~n19096 ;
  assign n19099 = n19097 | n19098 ;
  assign n19100 = x98 & n7812 ;
  assign n19101 = x97 & n7807 ;
  assign n19102 = x96 & ~n7806 ;
  assign n19103 = n8136 & n19102 ;
  assign n19104 = n19101 | n19103 ;
  assign n19105 = n19100 | n19104 ;
  assign n19106 = n7815 | n19105 ;
  assign n19107 = ( n4105 & n19105 ) | ( n4105 & n19106 ) | ( n19105 & n19106 ) ;
  assign n19108 = x50 & n19107 ;
  assign n19109 = x50 & ~n19108 ;
  assign n19110 = ( n19107 & ~n19108 ) | ( n19107 & n19109 ) | ( ~n19108 & n19109 ) ;
  assign n19111 = n19099 & n19110 ;
  assign n19112 = ( n19029 & ~n19096 ) | ( n19029 & n19110 ) | ( ~n19096 & n19110 ) ;
  assign n19113 = n19097 | n19112 ;
  assign n19114 = ~n19111 & n19113 ;
  assign n19115 = ( n18829 & n18830 ) | ( n18829 & ~n18831 ) | ( n18830 & ~n18831 ) ;
  assign n19116 = n19114 & ~n19115 ;
  assign n19117 = ~n19114 & n19115 ;
  assign n19118 = n19116 | n19117 ;
  assign n19119 = x101 & n6937 ;
  assign n19120 = x100 & n6932 ;
  assign n19121 = x99 & ~n6931 ;
  assign n19122 = n7216 & n19121 ;
  assign n19123 = n19120 | n19122 ;
  assign n19124 = n19119 | n19123 ;
  assign n19125 = n6940 | n19124 ;
  assign n19126 = ( n4783 & n19124 ) | ( n4783 & n19125 ) | ( n19124 & n19125 ) ;
  assign n19127 = x47 & n19126 ;
  assign n19128 = x47 & ~n19127 ;
  assign n19129 = ( n19126 & ~n19127 ) | ( n19126 & n19128 ) | ( ~n19127 & n19128 ) ;
  assign n19130 = n19118 & ~n19129 ;
  assign n19131 = ~n19118 & n19129 ;
  assign n19132 = n19130 | n19131 ;
  assign n19133 = n18845 | n18849 ;
  assign n19134 = n19132 & n19133 ;
  assign n19135 = ~n19132 & n19133 ;
  assign n19136 = n19132 | n19135 ;
  assign n19137 = x104 & n6068 ;
  assign n19138 = x103 & n6063 ;
  assign n19139 = x102 & ~n6062 ;
  assign n19140 = n6398 & n19139 ;
  assign n19141 = n19138 | n19140 ;
  assign n19142 = n19137 | n19141 ;
  assign n19143 = n6071 | n19142 ;
  assign n19144 = ( n5295 & n19142 ) | ( n5295 & n19143 ) | ( n19142 & n19143 ) ;
  assign n19145 = x44 & n19144 ;
  assign n19146 = x44 & ~n19145 ;
  assign n19147 = ( n19144 & ~n19145 ) | ( n19144 & n19146 ) | ( ~n19145 & n19146 ) ;
  assign n19148 = n19136 & ~n19147 ;
  assign n19149 = ~n19134 & n19148 ;
  assign n19150 = ( n19134 & ~n19136 ) | ( n19134 & n19147 ) | ( ~n19136 & n19147 ) ;
  assign n19151 = n19149 | n19150 ;
  assign n19152 = n18862 | n19151 ;
  assign n19153 = n18862 & n19151 ;
  assign n19154 = n19152 & ~n19153 ;
  assign n19155 = x107 & n5340 ;
  assign n19156 = x106 & n5335 ;
  assign n19157 = x105 & ~n5334 ;
  assign n19158 = n5580 & n19157 ;
  assign n19159 = n19156 | n19158 ;
  assign n19160 = n19155 | n19159 ;
  assign n19161 = n5343 | n19160 ;
  assign n19162 = ( n6328 & n19160 ) | ( n6328 & n19161 ) | ( n19160 & n19161 ) ;
  assign n19163 = x41 & n19162 ;
  assign n19164 = x41 & ~n19163 ;
  assign n19165 = ( n19162 & ~n19163 ) | ( n19162 & n19164 ) | ( ~n19163 & n19164 ) ;
  assign n19166 = n19154 & ~n19165 ;
  assign n19167 = n19165 | n19166 ;
  assign n19168 = ( ~n19154 & n19166 ) | ( ~n19154 & n19167 ) | ( n19166 & n19167 ) ;
  assign n19169 = n18865 | n18870 ;
  assign n19170 = ( n19028 & n19168 ) | ( n19028 & ~n19169 ) | ( n19168 & ~n19169 ) ;
  assign n19171 = ( ~n19168 & n19169 ) | ( ~n19168 & n19170 ) | ( n19169 & n19170 ) ;
  assign n19172 = ( ~n19028 & n19170 ) | ( ~n19028 & n19171 ) | ( n19170 & n19171 ) ;
  assign n19173 = ( n19016 & ~n19017 ) | ( n19016 & n19172 ) | ( ~n19017 & n19172 ) ;
  assign n19174 = ( n19017 & ~n19172 ) | ( n19017 & n19173 ) | ( ~n19172 & n19173 ) ;
  assign n19175 = ( ~n19016 & n19173 ) | ( ~n19016 & n19174 ) | ( n19173 & n19174 ) ;
  assign n19176 = x119 & n2775 ;
  assign n19177 = x118 & n2770 ;
  assign n19178 = x117 & ~n2769 ;
  assign n19179 = n2978 & n19178 ;
  assign n19180 = n19177 | n19179 ;
  assign n19181 = n19176 | n19180 ;
  assign n19182 = n2778 | n19181 ;
  assign n19183 = ( n9789 & n19181 ) | ( n9789 & n19182 ) | ( n19181 & n19182 ) ;
  assign n19184 = x29 & n19183 ;
  assign n19185 = x29 & ~n19184 ;
  assign n19186 = ( n19183 & ~n19184 ) | ( n19183 & n19185 ) | ( ~n19184 & n19185 ) ;
  assign n19187 = ( n18908 & n18919 ) | ( n18908 & n18920 ) | ( n18919 & n18920 ) ;
  assign n19188 = n19186 | n19187 ;
  assign n19189 = n19186 & n19187 ;
  assign n19190 = n19188 & ~n19189 ;
  assign n19191 = x116 & n3314 ;
  assign n19192 = x115 & n3309 ;
  assign n19193 = x114 & ~n3308 ;
  assign n19194 = n3570 & n19193 ;
  assign n19195 = n19192 | n19194 ;
  assign n19196 = n19191 | n19195 ;
  assign n19197 = n3317 | n19196 ;
  assign n19198 = ( n8778 & n19196 ) | ( n8778 & n19197 ) | ( n19196 & n19197 ) ;
  assign n19199 = x32 & n19198 ;
  assign n19200 = x32 & ~n19199 ;
  assign n19201 = ( n19198 & ~n19199 ) | ( n19198 & n19200 ) | ( ~n19199 & n19200 ) ;
  assign n19202 = n18902 | n19201 ;
  assign n19203 = n18907 | n19202 ;
  assign n19204 = ( n18902 & n18907 ) | ( n18902 & n19201 ) | ( n18907 & n19201 ) ;
  assign n19205 = n19203 & ~n19204 ;
  assign n19206 = ( n19175 & n19190 ) | ( n19175 & ~n19205 ) | ( n19190 & ~n19205 ) ;
  assign n19207 = ( ~n19190 & n19205 ) | ( ~n19190 & n19206 ) | ( n19205 & n19206 ) ;
  assign n19208 = ( ~n19175 & n19206 ) | ( ~n19175 & n19207 ) | ( n19206 & n19207 ) ;
  assign n19209 = n19005 & n19208 ;
  assign n19210 = n19005 | n19208 ;
  assign n19211 = ~n19209 & n19210 ;
  assign n19212 = x125 & n1817 ;
  assign n19213 = x124 & n1812 ;
  assign n19214 = x123 & ~n1811 ;
  assign n19215 = n1977 & n19214 ;
  assign n19216 = n19213 | n19215 ;
  assign n19217 = n19212 | n19216 ;
  assign n19218 = n1820 | n19217 ;
  assign n19219 = ( n12310 & n19217 ) | ( n12310 & n19218 ) | ( n19217 & n19218 ) ;
  assign n19220 = x23 & n19219 ;
  assign n19221 = x23 & ~n19220 ;
  assign n19222 = ( n19219 & ~n19220 ) | ( n19219 & n19221 ) | ( ~n19220 & n19221 ) ;
  assign n19223 = ( n18927 & n18938 ) | ( n18927 & n18940 ) | ( n18938 & n18940 ) ;
  assign n19224 = n19222 | n19223 ;
  assign n19225 = n19222 & n19223 ;
  assign n19226 = n19224 & ~n19225 ;
  assign n19227 = n19211 & n19226 ;
  assign n19228 = n19226 & ~n19227 ;
  assign n19229 = ( n19211 & ~n19227 ) | ( n19211 & n19228 ) | ( ~n19227 & n19228 ) ;
  assign n19230 = n18990 | n19229 ;
  assign n19231 = n18989 | n19230 ;
  assign n19232 = ( n18989 & n18990 ) | ( n18989 & n19229 ) | ( n18990 & n19229 ) ;
  assign n19233 = n19231 & ~n19232 ;
  assign n19234 = ( n18697 & n18698 ) | ( n18697 & n18962 ) | ( n18698 & n18962 ) ;
  assign n19235 = n19233 & ~n19234 ;
  assign n19236 = n18968 | n18971 ;
  assign n19237 = n19233 & n19234 ;
  assign n19238 = n19234 & ~n19237 ;
  assign n19239 = n19235 | n19238 ;
  assign n19240 = n19236 & n19239 ;
  assign n19241 = n18968 | n18973 ;
  assign n19242 = n19239 & n19241 ;
  assign n19243 = ( n17506 & n19240 ) | ( n17506 & n19242 ) | ( n19240 & n19242 ) ;
  assign n19244 = ( n17506 & n19236 ) | ( n17506 & n19241 ) | ( n19236 & n19241 ) ;
  assign n19245 = ( ~n19233 & n19234 ) | ( ~n19233 & n19244 ) | ( n19234 & n19244 ) ;
  assign n19246 = ( n19235 & ~n19243 ) | ( n19235 & n19245 ) | ( ~n19243 & n19245 ) ;
  assign n19247 = n18988 | n19232 ;
  assign n19248 = n19225 | n19227 ;
  assign n19249 = x127 & ~n1415 ;
  assign n19250 = n1584 & n19249 ;
  assign n19251 = ( x127 & n1424 ) | ( x127 & n19250 ) | ( n1424 & n19250 ) ;
  assign n19252 = ( x126 & n19250 ) | ( x126 & n19251 ) | ( n19250 & n19251 ) ;
  assign n19253 = ( n12685 & n19251 ) | ( n12685 & n19252 ) | ( n19251 & n19252 ) ;
  assign n19254 = x20 & n19253 ;
  assign n19255 = x20 & ~n19254 ;
  assign n19256 = ( n19253 & ~n19254 ) | ( n19253 & n19255 ) | ( ~n19254 & n19255 ) ;
  assign n19257 = n19248 & n19256 ;
  assign n19258 = n19248 & ~n19257 ;
  assign n19259 = x126 & n1817 ;
  assign n19260 = x125 & n1812 ;
  assign n19261 = x124 & ~n1811 ;
  assign n19262 = n1977 & n19261 ;
  assign n19263 = n19260 | n19262 ;
  assign n19264 = n19259 | n19263 ;
  assign n19265 = n1820 | n19264 ;
  assign n19266 = ( n12687 & n19264 ) | ( n12687 & n19265 ) | ( n19264 & n19265 ) ;
  assign n19267 = x23 & n19266 ;
  assign n19268 = x23 & ~n19267 ;
  assign n19269 = ( n19266 & ~n19267 ) | ( n19266 & n19268 ) | ( ~n19267 & n19268 ) ;
  assign n19270 = ( n19004 & n19209 ) | ( n19004 & n19269 ) | ( n19209 & n19269 ) ;
  assign n19271 = ( n19004 & n19209 ) | ( n19004 & ~n19269 ) | ( n19209 & ~n19269 ) ;
  assign n19272 = ( n19269 & ~n19270 ) | ( n19269 & n19271 ) | ( ~n19270 & n19271 ) ;
  assign n19273 = x114 & n3913 ;
  assign n19274 = x113 & n3908 ;
  assign n19275 = x112 & ~n3907 ;
  assign n19276 = n4152 & n19275 ;
  assign n19277 = n19274 | n19276 ;
  assign n19278 = n19273 | n19277 ;
  assign n19279 = n3916 | n19278 ;
  assign n19280 = ( n8437 & n19278 ) | ( n8437 & n19279 ) | ( n19278 & n19279 ) ;
  assign n19281 = x35 & n19280 ;
  assign n19282 = x35 & ~n19281 ;
  assign n19283 = ( n19280 & ~n19281 ) | ( n19280 & n19282 ) | ( ~n19281 & n19282 ) ;
  assign n19284 = ( n19016 & n19017 ) | ( n19016 & n19172 ) | ( n19017 & n19172 ) ;
  assign n19285 = x117 & n3314 ;
  assign n19286 = x116 & n3309 ;
  assign n19287 = x115 & ~n3308 ;
  assign n19288 = n3570 & n19287 ;
  assign n19289 = n19286 | n19288 ;
  assign n19290 = n19285 | n19289 ;
  assign n19291 = n3317 | n19290 ;
  assign n19292 = ( n9118 & n19290 ) | ( n9118 & n19291 ) | ( n19290 & n19291 ) ;
  assign n19293 = x32 & n19292 ;
  assign n19294 = x32 & ~n19293 ;
  assign n19295 = ( n19292 & ~n19293 ) | ( n19292 & n19294 ) | ( ~n19293 & n19294 ) ;
  assign n19296 = n19284 | n19295 ;
  assign n19297 = n19284 & n19295 ;
  assign n19298 = n19296 & ~n19297 ;
  assign n19299 = ( n19028 & n19168 ) | ( n19028 & n19169 ) | ( n19168 & n19169 ) ;
  assign n19300 = n19135 | n19150 ;
  assign n19301 = x93 & n9853 ;
  assign n19302 = x92 & n9848 ;
  assign n19303 = x91 & ~n9847 ;
  assign n19304 = n10165 & n19303 ;
  assign n19305 = n19302 | n19304 ;
  assign n19306 = n19301 | n19305 ;
  assign n19307 = n9856 | n19306 ;
  assign n19308 = ( n2931 & n19306 ) | ( n2931 & n19307 ) | ( n19306 & n19307 ) ;
  assign n19309 = x56 & n19308 ;
  assign n19310 = x56 & ~n19309 ;
  assign n19311 = ( n19308 & ~n19309 ) | ( n19308 & n19310 ) | ( ~n19309 & n19310 ) ;
  assign n19312 = n19080 | n19085 ;
  assign n19313 = x84 & n12808 ;
  assign n19314 = x63 & x83 ;
  assign n19315 = ~n12808 & n19314 ;
  assign n19316 = n19313 | n19315 ;
  assign n19317 = n19077 & ~n19316 ;
  assign n19318 = ~n19077 & n19316 ;
  assign n19319 = n19317 | n19318 ;
  assign n19320 = x87 & n11984 ;
  assign n19321 = x86 & n11979 ;
  assign n19322 = x85 & ~n11978 ;
  assign n19323 = n12430 & n19322 ;
  assign n19324 = n19321 | n19323 ;
  assign n19325 = n19320 | n19324 ;
  assign n19326 = n11987 | n19325 ;
  assign n19327 = ( n2067 & n19325 ) | ( n2067 & n19326 ) | ( n19325 & n19326 ) ;
  assign n19328 = x62 & n19327 ;
  assign n19329 = x62 & ~n19328 ;
  assign n19330 = ( n19327 & ~n19328 ) | ( n19327 & n19329 ) | ( ~n19328 & n19329 ) ;
  assign n19331 = ~n19319 & n19330 ;
  assign n19332 = n19319 & ~n19330 ;
  assign n19333 = n19331 | n19332 ;
  assign n19334 = n19312 & ~n19333 ;
  assign n19335 = ~n19312 & n19333 ;
  assign n19336 = n19334 | n19335 ;
  assign n19337 = x90 & n10876 ;
  assign n19338 = x89 & n10871 ;
  assign n19339 = x88 & ~n10870 ;
  assign n19340 = n11305 & n19339 ;
  assign n19341 = n19338 | n19340 ;
  assign n19342 = n19337 | n19341 ;
  assign n19343 = n10879 | n19342 ;
  assign n19344 = ( n2410 & n19342 ) | ( n2410 & n19343 ) | ( n19342 & n19343 ) ;
  assign n19345 = x59 & n19344 ;
  assign n19346 = x59 & ~n19345 ;
  assign n19347 = ( n19344 & ~n19345 ) | ( n19344 & n19346 ) | ( ~n19345 & n19346 ) ;
  assign n19348 = ~n19336 & n19347 ;
  assign n19349 = n19336 & ~n19347 ;
  assign n19350 = n19348 | n19349 ;
  assign n19351 = ( ~n19089 & n19311 ) | ( ~n19089 & n19350 ) | ( n19311 & n19350 ) ;
  assign n19352 = ( n19089 & ~n19350 ) | ( n19089 & n19351 ) | ( ~n19350 & n19351 ) ;
  assign n19353 = ( ~n19311 & n19351 ) | ( ~n19311 & n19352 ) | ( n19351 & n19352 ) ;
  assign n19354 = n19092 & ~n19353 ;
  assign n19355 = n19353 | n19354 ;
  assign n19356 = n19092 & ~n19354 ;
  assign n19357 = n19355 & ~n19356 ;
  assign n19358 = x96 & n8834 ;
  assign n19359 = x95 & n8829 ;
  assign n19360 = x94 & ~n8828 ;
  assign n19361 = n9159 & n19360 ;
  assign n19362 = n19359 | n19361 ;
  assign n19363 = n19358 | n19362 ;
  assign n19364 = n8837 | n19363 ;
  assign n19365 = ( n3509 & n19363 ) | ( n3509 & n19364 ) | ( n19363 & n19364 ) ;
  assign n19366 = x53 & n19365 ;
  assign n19367 = x53 & ~n19366 ;
  assign n19368 = ( n19365 & ~n19366 ) | ( n19365 & n19367 ) | ( ~n19366 & n19367 ) ;
  assign n19369 = n19357 | n19368 ;
  assign n19370 = n19357 & n19368 ;
  assign n19371 = n19369 & ~n19370 ;
  assign n19372 = n19095 & ~n19371 ;
  assign n19373 = ~n19095 & n19371 ;
  assign n19374 = n19372 | n19373 ;
  assign n19375 = x99 & n7812 ;
  assign n19376 = x98 & n7807 ;
  assign n19377 = x97 & ~n7806 ;
  assign n19378 = n8136 & n19377 ;
  assign n19379 = n19376 | n19378 ;
  assign n19380 = n19375 | n19379 ;
  assign n19381 = n7815 | n19380 ;
  assign n19382 = ( n4325 & n19380 ) | ( n4325 & n19381 ) | ( n19380 & n19381 ) ;
  assign n19383 = x50 & n19382 ;
  assign n19384 = x50 & ~n19383 ;
  assign n19385 = ( n19382 & ~n19383 ) | ( n19382 & n19384 ) | ( ~n19383 & n19384 ) ;
  assign n19386 = ~n19374 & n19385 ;
  assign n19387 = n19374 & ~n19385 ;
  assign n19388 = n19386 | n19387 ;
  assign n19389 = n19112 & ~n19388 ;
  assign n19390 = ~n19112 & n19388 ;
  assign n19391 = n19389 | n19390 ;
  assign n19392 = x102 & n6937 ;
  assign n19393 = x101 & n6932 ;
  assign n19394 = x100 & ~n6931 ;
  assign n19395 = n7216 & n19394 ;
  assign n19396 = n19393 | n19395 ;
  assign n19397 = n19392 | n19396 ;
  assign n19398 = n6940 | n19397 ;
  assign n19399 = ( n5025 & n19397 ) | ( n5025 & n19398 ) | ( n19397 & n19398 ) ;
  assign n19400 = x47 & n19399 ;
  assign n19401 = x47 & ~n19400 ;
  assign n19402 = ( n19399 & ~n19400 ) | ( n19399 & n19401 ) | ( ~n19400 & n19401 ) ;
  assign n19403 = ~n19391 & n19402 ;
  assign n19404 = n19391 & ~n19402 ;
  assign n19405 = n19403 | n19404 ;
  assign n19406 = n19117 | n19131 ;
  assign n19407 = ~n19405 & n19406 ;
  assign n19408 = n19405 & ~n19406 ;
  assign n19409 = n19407 | n19408 ;
  assign n19410 = x105 & n6068 ;
  assign n19411 = x104 & n6063 ;
  assign n19412 = x103 & ~n6062 ;
  assign n19413 = n6398 & n19412 ;
  assign n19414 = n19411 | n19413 ;
  assign n19415 = n19410 | n19414 ;
  assign n19416 = n6071 | n19415 ;
  assign n19417 = ( n5788 & n19415 ) | ( n5788 & n19416 ) | ( n19415 & n19416 ) ;
  assign n19418 = x44 & n19417 ;
  assign n19419 = x44 & ~n19418 ;
  assign n19420 = ( n19417 & ~n19418 ) | ( n19417 & n19419 ) | ( ~n19418 & n19419 ) ;
  assign n19421 = ~n19409 & n19420 ;
  assign n19422 = n19409 & ~n19420 ;
  assign n19423 = n19421 | n19422 ;
  assign n19424 = n19300 & ~n19423 ;
  assign n19425 = ~n19300 & n19423 ;
  assign n19426 = n19424 | n19425 ;
  assign n19427 = x108 & n5340 ;
  assign n19428 = x107 & n5335 ;
  assign n19429 = x106 & ~n5334 ;
  assign n19430 = n5580 & n19429 ;
  assign n19431 = n19428 | n19430 ;
  assign n19432 = n19427 | n19431 ;
  assign n19433 = n5343 | n19432 ;
  assign n19434 = ( n6358 & n19432 ) | ( n6358 & n19433 ) | ( n19432 & n19433 ) ;
  assign n19435 = x41 & n19434 ;
  assign n19436 = x41 & ~n19435 ;
  assign n19437 = ( n19434 & ~n19435 ) | ( n19434 & n19436 ) | ( ~n19435 & n19436 ) ;
  assign n19438 = ~n19426 & n19437 ;
  assign n19439 = n19426 & ~n19437 ;
  assign n19440 = n19438 | n19439 ;
  assign n19441 = ( n18862 & n19151 ) | ( n18862 & n19166 ) | ( n19151 & n19166 ) ;
  assign n19442 = n19440 | n19441 ;
  assign n19443 = n19440 & n19441 ;
  assign n19444 = n19442 & ~n19443 ;
  assign n19445 = x111 & n4572 ;
  assign n19446 = x110 & n4567 ;
  assign n19447 = x109 & ~n4566 ;
  assign n19448 = n4828 & n19447 ;
  assign n19449 = n19446 | n19448 ;
  assign n19450 = n19445 | n19449 ;
  assign n19451 = n4575 | n19450 ;
  assign n19452 = ( n7492 & n19450 ) | ( n7492 & n19451 ) | ( n19450 & n19451 ) ;
  assign n19453 = x38 & n19452 ;
  assign n19454 = x38 & ~n19453 ;
  assign n19455 = ( n19452 & ~n19453 ) | ( n19452 & n19454 ) | ( ~n19453 & n19454 ) ;
  assign n19456 = n19444 & ~n19455 ;
  assign n19457 = n19455 | n19456 ;
  assign n19458 = ( ~n19444 & n19456 ) | ( ~n19444 & n19457 ) | ( n19456 & n19457 ) ;
  assign n19459 = n19299 | n19458 ;
  assign n19460 = n19299 & n19458 ;
  assign n19461 = n19459 & ~n19460 ;
  assign n19462 = ( n19283 & n19298 ) | ( n19283 & ~n19461 ) | ( n19298 & ~n19461 ) ;
  assign n19463 = ( ~n19298 & n19461 ) | ( ~n19298 & n19462 ) | ( n19461 & n19462 ) ;
  assign n19464 = ( ~n19283 & n19462 ) | ( ~n19283 & n19463 ) | ( n19462 & n19463 ) ;
  assign n19465 = x120 & n2775 ;
  assign n19466 = x119 & n2770 ;
  assign n19467 = x118 & ~n2769 ;
  assign n19468 = n2978 & n19467 ;
  assign n19469 = n19466 | n19468 ;
  assign n19470 = n19465 | n19469 ;
  assign n19471 = n2778 | n19470 ;
  assign n19472 = ( n10460 & n19470 ) | ( n10460 & n19471 ) | ( n19470 & n19471 ) ;
  assign n19473 = x29 & n19472 ;
  assign n19474 = x29 & ~n19473 ;
  assign n19475 = ( n19472 & ~n19473 ) | ( n19472 & n19474 ) | ( ~n19473 & n19474 ) ;
  assign n19476 = n19175 & n19205 ;
  assign n19477 = n19204 | n19476 ;
  assign n19478 = ( n19464 & n19475 ) | ( n19464 & ~n19477 ) | ( n19475 & ~n19477 ) ;
  assign n19479 = ( ~n19475 & n19477 ) | ( ~n19475 & n19478 ) | ( n19477 & n19478 ) ;
  assign n19480 = ( ~n19464 & n19478 ) | ( ~n19464 & n19479 ) | ( n19478 & n19479 ) ;
  assign n19481 = x123 & n2280 ;
  assign n19482 = x122 & n2275 ;
  assign n19483 = x121 & ~n2274 ;
  assign n19484 = n2481 & n19483 ;
  assign n19485 = n19482 | n19484 ;
  assign n19486 = n19481 | n19485 ;
  assign n19487 = n2283 | n19486 ;
  assign n19488 = ( n11219 & n19486 ) | ( n11219 & n19487 ) | ( n19486 & n19487 ) ;
  assign n19489 = x26 & n19488 ;
  assign n19490 = x26 & ~n19489 ;
  assign n19491 = ( n19488 & ~n19489 ) | ( n19488 & n19490 ) | ( ~n19489 & n19490 ) ;
  assign n19492 = ( n19175 & n19190 ) | ( n19175 & n19205 ) | ( n19190 & n19205 ) ;
  assign n19493 = ( n19189 & ~n19476 ) | ( n19189 & n19492 ) | ( ~n19476 & n19492 ) ;
  assign n19494 = ( n19480 & ~n19491 ) | ( n19480 & n19493 ) | ( ~n19491 & n19493 ) ;
  assign n19495 = ( n19491 & ~n19493 ) | ( n19491 & n19494 ) | ( ~n19493 & n19494 ) ;
  assign n19496 = ( ~n19480 & n19494 ) | ( ~n19480 & n19495 ) | ( n19494 & n19495 ) ;
  assign n19497 = n19272 & ~n19496 ;
  assign n19498 = ~n19272 & n19496 ;
  assign n19499 = n19497 | n19498 ;
  assign n19500 = ~n19248 & n19256 ;
  assign n19501 = n19499 | n19500 ;
  assign n19502 = n19258 | n19501 ;
  assign n19503 = ( n19258 & n19499 ) | ( n19258 & n19500 ) | ( n19499 & n19500 ) ;
  assign n19504 = n19502 & ~n19503 ;
  assign n19505 = n19247 & n19504 ;
  assign n19506 = n19247 | n19504 ;
  assign n19507 = ~n19505 & n19506 ;
  assign n19508 = n19237 | n19240 ;
  assign n19509 = n19237 | n19242 ;
  assign n19510 = ( n17506 & n19508 ) | ( n17506 & n19509 ) | ( n19508 & n19509 ) ;
  assign n19511 = n19507 | n19510 ;
  assign n19512 = n19507 & n19508 ;
  assign n19513 = n19507 & n19509 ;
  assign n19514 = ( n17506 & n19512 ) | ( n17506 & n19513 ) | ( n19512 & n19513 ) ;
  assign n19515 = n19511 & ~n19514 ;
  assign n19516 = n19257 | n19503 ;
  assign n19517 = x124 & n2280 ;
  assign n19518 = x123 & n2275 ;
  assign n19519 = x122 & ~n2274 ;
  assign n19520 = n2481 & n19519 ;
  assign n19521 = n19518 | n19520 ;
  assign n19522 = n19517 | n19521 ;
  assign n19523 = n2283 | n19522 ;
  assign n19524 = ( n11916 & n19522 ) | ( n11916 & n19523 ) | ( n19522 & n19523 ) ;
  assign n19525 = x26 & n19524 ;
  assign n19526 = x26 & ~n19525 ;
  assign n19527 = ( n19524 & ~n19525 ) | ( n19524 & n19526 ) | ( ~n19525 & n19526 ) ;
  assign n19528 = ( n19480 & n19491 ) | ( n19480 & n19493 ) | ( n19491 & n19493 ) ;
  assign n19529 = n19527 | n19528 ;
  assign n19530 = n19527 & n19528 ;
  assign n19531 = n19529 & ~n19530 ;
  assign n19532 = ( n19270 & n19272 ) | ( n19270 & ~n19497 ) | ( n19272 & ~n19497 ) ;
  assign n19533 = x127 & n1817 ;
  assign n19534 = x126 & n1812 ;
  assign n19535 = x125 & ~n1811 ;
  assign n19536 = n1977 & n19535 ;
  assign n19537 = n19534 | n19536 ;
  assign n19538 = n19533 | n19537 ;
  assign n19539 = n1820 | n19538 ;
  assign n19540 = ( n12720 & n19538 ) | ( n12720 & n19539 ) | ( n19538 & n19539 ) ;
  assign n19541 = x23 & n19540 ;
  assign n19542 = x23 & ~n19541 ;
  assign n19543 = ( n19540 & ~n19541 ) | ( n19540 & n19542 ) | ( ~n19541 & n19542 ) ;
  assign n19544 = ~n19532 & n19543 ;
  assign n19545 = n19532 & ~n19543 ;
  assign n19546 = n19544 | n19545 ;
  assign n19547 = n19424 | n19438 ;
  assign n19548 = x109 & n5340 ;
  assign n19549 = x108 & n5335 ;
  assign n19550 = x107 & ~n5334 ;
  assign n19551 = n5580 & n19550 ;
  assign n19552 = n19549 | n19551 ;
  assign n19553 = n19548 | n19552 ;
  assign n19554 = n5343 | n19553 ;
  assign n19555 = ( n6884 & n19553 ) | ( n6884 & n19554 ) | ( n19553 & n19554 ) ;
  assign n19556 = x41 & n19555 ;
  assign n19557 = x41 & ~n19556 ;
  assign n19558 = ( n19555 & ~n19556 ) | ( n19555 & n19557 ) | ( ~n19556 & n19557 ) ;
  assign n19559 = n19407 | n19421 ;
  assign n19560 = x106 & n6068 ;
  assign n19561 = x105 & n6063 ;
  assign n19562 = x104 & ~n6062 ;
  assign n19563 = n6398 & n19562 ;
  assign n19564 = n19561 | n19563 ;
  assign n19565 = n19560 | n19564 ;
  assign n19566 = n6071 | n19565 ;
  assign n19567 = ( n5814 & n19565 ) | ( n5814 & n19566 ) | ( n19565 & n19566 ) ;
  assign n19568 = x44 & n19567 ;
  assign n19569 = x44 & ~n19568 ;
  assign n19570 = ( n19567 & ~n19568 ) | ( n19567 & n19569 ) | ( ~n19568 & n19569 ) ;
  assign n19571 = n19389 | n19403 ;
  assign n19572 = x103 & n6937 ;
  assign n19573 = x102 & n6932 ;
  assign n19574 = x101 & ~n6931 ;
  assign n19575 = n7216 & n19574 ;
  assign n19576 = n19573 | n19575 ;
  assign n19577 = n19572 | n19576 ;
  assign n19578 = n6940 | n19577 ;
  assign n19579 = ( n5264 & n19577 ) | ( n5264 & n19578 ) | ( n19577 & n19578 ) ;
  assign n19580 = x47 & n19579 ;
  assign n19581 = x47 & ~n19580 ;
  assign n19582 = ( n19579 & ~n19580 ) | ( n19579 & n19581 ) | ( ~n19580 & n19581 ) ;
  assign n19583 = x85 & n12808 ;
  assign n19584 = x63 & x84 ;
  assign n19585 = ~n12808 & n19584 ;
  assign n19586 = n19583 | n19585 ;
  assign n19587 = ~x20 & n19586 ;
  assign n19588 = x20 & ~n19586 ;
  assign n19589 = n19587 | n19588 ;
  assign n19590 = n19316 & ~n19589 ;
  assign n19591 = ~n19316 & n19589 ;
  assign n19592 = n19590 | n19591 ;
  assign n19593 = x88 & n11984 ;
  assign n19594 = x87 & n11979 ;
  assign n19595 = x86 & ~n11978 ;
  assign n19596 = n12430 & n19595 ;
  assign n19597 = n19594 | n19596 ;
  assign n19598 = n19593 | n19597 ;
  assign n19599 = n11987 | n19598 ;
  assign n19600 = ( n2095 & n19598 ) | ( n2095 & n19599 ) | ( n19598 & n19599 ) ;
  assign n19601 = ~x62 & n19600 ;
  assign n19602 = x62 & ~n19600 ;
  assign n19603 = n19601 | n19602 ;
  assign n19604 = ~n19592 & n19603 ;
  assign n19605 = n19592 & ~n19603 ;
  assign n19606 = n19604 | n19605 ;
  assign n19607 = n19317 | n19331 ;
  assign n19608 = ~n19606 & n19607 ;
  assign n19609 = n19606 | n19608 ;
  assign n19610 = n19606 & n19607 ;
  assign n19611 = n19609 & ~n19610 ;
  assign n19612 = x91 & n10876 ;
  assign n19613 = x90 & n10871 ;
  assign n19614 = x89 & ~n10870 ;
  assign n19615 = n11305 & n19614 ;
  assign n19616 = n19613 | n19615 ;
  assign n19617 = n19612 | n19616 ;
  assign n19618 = n10879 | n19617 ;
  assign n19619 = ( n2714 & n19617 ) | ( n2714 & n19618 ) | ( n19617 & n19618 ) ;
  assign n19620 = x59 & n19619 ;
  assign n19621 = x59 & ~n19620 ;
  assign n19622 = ( n19619 & ~n19620 ) | ( n19619 & n19621 ) | ( ~n19620 & n19621 ) ;
  assign n19623 = ~n19611 & n19622 ;
  assign n19624 = n19611 & ~n19622 ;
  assign n19625 = n19623 | n19624 ;
  assign n19626 = n19334 | n19348 ;
  assign n19627 = n19625 & ~n19626 ;
  assign n19628 = ~n19625 & n19626 ;
  assign n19629 = n19627 | n19628 ;
  assign n19630 = x94 & n9853 ;
  assign n19631 = x93 & n9848 ;
  assign n19632 = x92 & ~n9847 ;
  assign n19633 = n10165 & n19632 ;
  assign n19634 = n19631 | n19633 ;
  assign n19635 = n19630 | n19634 ;
  assign n19636 = n9856 | n19635 ;
  assign n19637 = ( n3271 & n19635 ) | ( n3271 & n19636 ) | ( n19635 & n19636 ) ;
  assign n19638 = x56 & n19637 ;
  assign n19639 = x56 & ~n19638 ;
  assign n19640 = ( n19637 & ~n19638 ) | ( n19637 & n19639 ) | ( ~n19638 & n19639 ) ;
  assign n19641 = ~n19629 & n19640 ;
  assign n19642 = n19629 | n19641 ;
  assign n19643 = n19629 & n19640 ;
  assign n19644 = n19352 | n19643 ;
  assign n19645 = n19642 & ~n19644 ;
  assign n19646 = ( n19352 & ~n19642 ) | ( n19352 & n19643 ) | ( ~n19642 & n19643 ) ;
  assign n19647 = n19645 | n19646 ;
  assign n19648 = x97 & n8834 ;
  assign n19649 = x96 & n8829 ;
  assign n19650 = x95 & ~n8828 ;
  assign n19651 = n9159 & n19650 ;
  assign n19652 = n19649 | n19651 ;
  assign n19653 = n19648 | n19652 ;
  assign n19654 = n8837 | n19653 ;
  assign n19655 = ( n3707 & n19653 ) | ( n3707 & n19654 ) | ( n19653 & n19654 ) ;
  assign n19656 = x53 & n19655 ;
  assign n19657 = x53 & ~n19656 ;
  assign n19658 = ( n19655 & ~n19656 ) | ( n19655 & n19657 ) | ( ~n19656 & n19657 ) ;
  assign n19659 = ( n19354 & ~n19357 ) | ( n19354 & n19369 ) | ( ~n19357 & n19369 ) ;
  assign n19660 = n19658 & n19659 ;
  assign n19661 = n19658 | n19659 ;
  assign n19662 = ~n19660 & n19661 ;
  assign n19663 = n19647 & n19662 ;
  assign n19664 = n19647 | n19662 ;
  assign n19665 = ~n19663 & n19664 ;
  assign n19666 = x100 & n7812 ;
  assign n19667 = x99 & n7807 ;
  assign n19668 = x98 & ~n7806 ;
  assign n19669 = n8136 & n19668 ;
  assign n19670 = n19667 | n19669 ;
  assign n19671 = n19666 | n19670 ;
  assign n19672 = n7815 | n19671 ;
  assign n19673 = ( n4532 & n19671 ) | ( n4532 & n19672 ) | ( n19671 & n19672 ) ;
  assign n19674 = x50 & n19673 ;
  assign n19675 = x50 & ~n19674 ;
  assign n19676 = ( n19673 & ~n19674 ) | ( n19673 & n19675 ) | ( ~n19674 & n19675 ) ;
  assign n19677 = ~n19665 & n19676 ;
  assign n19678 = n19665 & ~n19676 ;
  assign n19679 = n19677 | n19678 ;
  assign n19680 = n19372 | n19386 ;
  assign n19681 = n19679 & ~n19680 ;
  assign n19682 = ~n19679 & n19680 ;
  assign n19683 = n19681 | n19682 ;
  assign n19684 = n19582 & ~n19683 ;
  assign n19685 = n19683 | n19684 ;
  assign n19686 = ( ~n19582 & n19684 ) | ( ~n19582 & n19685 ) | ( n19684 & n19685 ) ;
  assign n19687 = ~n19571 & n19686 ;
  assign n19688 = n19571 & ~n19686 ;
  assign n19689 = n19687 | n19688 ;
  assign n19690 = n19570 & ~n19689 ;
  assign n19691 = n19689 | n19690 ;
  assign n19692 = ( ~n19570 & n19690 ) | ( ~n19570 & n19691 ) | ( n19690 & n19691 ) ;
  assign n19693 = ~n19559 & n19692 ;
  assign n19694 = n19559 & ~n19692 ;
  assign n19695 = n19693 | n19694 ;
  assign n19696 = n19558 & ~n19695 ;
  assign n19697 = n19695 | n19696 ;
  assign n19698 = ( ~n19558 & n19696 ) | ( ~n19558 & n19697 ) | ( n19696 & n19697 ) ;
  assign n19699 = ~n19547 & n19698 ;
  assign n19700 = n19547 & ~n19698 ;
  assign n19701 = n19699 | n19700 ;
  assign n19702 = x112 & n4572 ;
  assign n19703 = x111 & n4567 ;
  assign n19704 = x110 & ~n4566 ;
  assign n19705 = n4828 & n19704 ;
  assign n19706 = n19703 | n19705 ;
  assign n19707 = n19702 | n19706 ;
  assign n19708 = n4575 | n19707 ;
  assign n19709 = ( n7789 & n19707 ) | ( n7789 & n19708 ) | ( n19707 & n19708 ) ;
  assign n19710 = x38 & n19709 ;
  assign n19711 = x38 & ~n19710 ;
  assign n19712 = ( n19709 & ~n19710 ) | ( n19709 & n19711 ) | ( ~n19710 & n19711 ) ;
  assign n19713 = ~n19701 & n19712 ;
  assign n19714 = n19701 | n19713 ;
  assign n19715 = n19701 & n19712 ;
  assign n19716 = ( n19440 & n19441 ) | ( n19440 & n19456 ) | ( n19441 & n19456 ) ;
  assign n19717 = ~n19715 & n19716 ;
  assign n19718 = n19714 & n19717 ;
  assign n19719 = ( n19714 & ~n19715 ) | ( n19714 & n19716 ) | ( ~n19715 & n19716 ) ;
  assign n19720 = ~n19718 & n19719 ;
  assign n19721 = x115 & n3913 ;
  assign n19722 = x114 & n3908 ;
  assign n19723 = x113 & ~n3907 ;
  assign n19724 = n4152 & n19723 ;
  assign n19725 = n19722 | n19724 ;
  assign n19726 = n19721 | n19725 ;
  assign n19727 = n3916 | n19726 ;
  assign n19728 = ( n8749 & n19726 ) | ( n8749 & n19727 ) | ( n19726 & n19727 ) ;
  assign n19729 = x35 & n19728 ;
  assign n19730 = x35 & ~n19729 ;
  assign n19731 = ( n19728 & ~n19729 ) | ( n19728 & n19730 ) | ( ~n19729 & n19730 ) ;
  assign n19732 = n19720 & n19731 ;
  assign n19733 = n19720 | n19731 ;
  assign n19734 = ~n19732 & n19733 ;
  assign n19735 = ( n19283 & n19299 ) | ( n19283 & n19458 ) | ( n19299 & n19458 ) ;
  assign n19736 = n19734 & n19735 ;
  assign n19737 = n19735 & ~n19736 ;
  assign n19738 = ( n19734 & ~n19736 ) | ( n19734 & n19737 ) | ( ~n19736 & n19737 ) ;
  assign n19739 = x121 & n2775 ;
  assign n19740 = x120 & n2770 ;
  assign n19741 = x119 & ~n2769 ;
  assign n19742 = n2978 & n19741 ;
  assign n19743 = n19740 | n19742 ;
  assign n19744 = n19739 | n19743 ;
  assign n19745 = n2778 | n19744 ;
  assign n19746 = ( n10811 & n19744 ) | ( n10811 & n19745 ) | ( n19744 & n19745 ) ;
  assign n19747 = x29 & n19746 ;
  assign n19748 = x29 & ~n19747 ;
  assign n19749 = ( n19746 & ~n19747 ) | ( n19746 & n19748 ) | ( ~n19747 & n19748 ) ;
  assign n19750 = ( n19464 & n19475 ) | ( n19464 & n19477 ) | ( n19475 & n19477 ) ;
  assign n19751 = ~n19749 & n19750 ;
  assign n19752 = n19749 & ~n19750 ;
  assign n19753 = n19751 | n19752 ;
  assign n19754 = x118 & n3314 ;
  assign n19755 = x117 & n3309 ;
  assign n19756 = x116 & ~n3308 ;
  assign n19757 = n3570 & n19756 ;
  assign n19758 = n19755 | n19757 ;
  assign n19759 = n19754 | n19758 ;
  assign n19760 = n3317 | n19759 ;
  assign n19761 = ( n9760 & n19759 ) | ( n9760 & n19760 ) | ( n19759 & n19760 ) ;
  assign n19762 = x32 & n19761 ;
  assign n19763 = x32 & ~n19762 ;
  assign n19764 = ( n19761 & ~n19762 ) | ( n19761 & n19763 ) | ( ~n19762 & n19763 ) ;
  assign n19765 = ( n19284 & n19295 ) | ( n19284 & ~n19464 ) | ( n19295 & ~n19464 ) ;
  assign n19766 = n19764 | n19765 ;
  assign n19767 = n19764 & n19765 ;
  assign n19768 = n19766 & ~n19767 ;
  assign n19769 = ( n19738 & n19753 ) | ( n19738 & ~n19768 ) | ( n19753 & ~n19768 ) ;
  assign n19770 = ( ~n19753 & n19768 ) | ( ~n19753 & n19769 ) | ( n19768 & n19769 ) ;
  assign n19771 = ( ~n19738 & n19769 ) | ( ~n19738 & n19770 ) | ( n19769 & n19770 ) ;
  assign n19772 = ( n19531 & ~n19546 ) | ( n19531 & n19771 ) | ( ~n19546 & n19771 ) ;
  assign n19773 = ( n19546 & ~n19771 ) | ( n19546 & n19772 ) | ( ~n19771 & n19772 ) ;
  assign n19774 = ( ~n19531 & n19772 ) | ( ~n19531 & n19773 ) | ( n19772 & n19773 ) ;
  assign n19775 = n19516 | n19774 ;
  assign n19776 = n19516 & n19774 ;
  assign n19777 = n19775 & ~n19776 ;
  assign n19778 = n19505 | n19512 ;
  assign n19779 = n19505 | n19513 ;
  assign n19780 = ( n17506 & n19778 ) | ( n17506 & n19779 ) | ( n19778 & n19779 ) ;
  assign n19781 = n19777 | n19780 ;
  assign n19782 = n19777 & n19778 ;
  assign n19783 = n19777 & n19779 ;
  assign n19784 = ( n17506 & n19782 ) | ( n17506 & n19783 ) | ( n19782 & n19783 ) ;
  assign n19785 = n19781 & ~n19784 ;
  assign n19786 = x116 & n3913 ;
  assign n19787 = x115 & n3908 ;
  assign n19788 = x114 & ~n3907 ;
  assign n19789 = n4152 & n19788 ;
  assign n19790 = n19787 | n19789 ;
  assign n19791 = n19786 | n19790 ;
  assign n19792 = n3916 | n19791 ;
  assign n19793 = ( n8778 & n19791 ) | ( n8778 & n19792 ) | ( n19791 & n19792 ) ;
  assign n19794 = x35 & n19793 ;
  assign n19795 = x35 & ~n19794 ;
  assign n19796 = ( n19793 & ~n19794 ) | ( n19793 & n19795 ) | ( ~n19794 & n19795 ) ;
  assign n19797 = n19690 | n19694 ;
  assign n19798 = x107 & n6068 ;
  assign n19799 = x106 & n6063 ;
  assign n19800 = x105 & ~n6062 ;
  assign n19801 = n6398 & n19800 ;
  assign n19802 = n19799 | n19801 ;
  assign n19803 = n19798 | n19802 ;
  assign n19804 = n6071 | n19803 ;
  assign n19805 = ( n6328 & n19803 ) | ( n6328 & n19804 ) | ( n19803 & n19804 ) ;
  assign n19806 = x44 & n19805 ;
  assign n19807 = x44 & ~n19806 ;
  assign n19808 = ( n19805 & ~n19806 ) | ( n19805 & n19807 ) | ( ~n19806 & n19807 ) ;
  assign n19809 = n19641 | n19646 ;
  assign n19810 = x95 & n9853 ;
  assign n19811 = x94 & n9848 ;
  assign n19812 = x93 & ~n9847 ;
  assign n19813 = n10165 & n19812 ;
  assign n19814 = n19811 | n19813 ;
  assign n19815 = n19810 | n19814 ;
  assign n19816 = n9856 | n19815 ;
  assign n19817 = ( n3479 & n19815 ) | ( n3479 & n19816 ) | ( n19815 & n19816 ) ;
  assign n19818 = x56 & n19817 ;
  assign n19819 = x56 & ~n19818 ;
  assign n19820 = ( n19817 & ~n19818 ) | ( n19817 & n19819 ) | ( ~n19818 & n19819 ) ;
  assign n19821 = x86 & n12808 ;
  assign n19822 = x63 & x85 ;
  assign n19823 = ~n12808 & n19822 ;
  assign n19824 = n19821 | n19823 ;
  assign n19825 = n19587 | n19590 ;
  assign n19826 = n19824 & ~n19825 ;
  assign n19827 = ~n19824 & n19825 ;
  assign n19828 = n19826 | n19827 ;
  assign n19829 = x89 & n11984 ;
  assign n19830 = x88 & n11979 ;
  assign n19831 = x87 & ~n11978 ;
  assign n19832 = n12430 & n19831 ;
  assign n19833 = n19830 | n19832 ;
  assign n19834 = n19829 | n19833 ;
  assign n19835 = n11987 | n19834 ;
  assign n19836 = ( n2244 & n19834 ) | ( n2244 & n19835 ) | ( n19834 & n19835 ) ;
  assign n19837 = x62 & n19836 ;
  assign n19838 = x62 & ~n19837 ;
  assign n19839 = ( n19836 & ~n19837 ) | ( n19836 & n19838 ) | ( ~n19837 & n19838 ) ;
  assign n19840 = ~n19828 & n19839 ;
  assign n19841 = n19828 & ~n19839 ;
  assign n19842 = n19840 | n19841 ;
  assign n19843 = n19604 | n19608 ;
  assign n19844 = ~n19842 & n19843 ;
  assign n19845 = n19842 & ~n19843 ;
  assign n19846 = n19844 | n19845 ;
  assign n19847 = x92 & n10876 ;
  assign n19848 = x91 & n10871 ;
  assign n19849 = x90 & ~n10870 ;
  assign n19850 = n11305 & n19849 ;
  assign n19851 = n19848 | n19850 ;
  assign n19852 = n19847 | n19851 ;
  assign n19853 = n10879 | n19852 ;
  assign n19854 = ( n2904 & n19852 ) | ( n2904 & n19853 ) | ( n19852 & n19853 ) ;
  assign n19855 = x59 & n19854 ;
  assign n19856 = x59 & ~n19855 ;
  assign n19857 = ( n19854 & ~n19855 ) | ( n19854 & n19856 ) | ( ~n19855 & n19856 ) ;
  assign n19858 = ~n19846 & n19857 ;
  assign n19859 = n19846 & ~n19857 ;
  assign n19860 = n19858 | n19859 ;
  assign n19861 = n19623 | n19628 ;
  assign n19862 = ( n19820 & n19860 ) | ( n19820 & ~n19861 ) | ( n19860 & ~n19861 ) ;
  assign n19863 = ( ~n19860 & n19861 ) | ( ~n19860 & n19862 ) | ( n19861 & n19862 ) ;
  assign n19864 = ( ~n19820 & n19862 ) | ( ~n19820 & n19863 ) | ( n19862 & n19863 ) ;
  assign n19865 = ~n19809 & n19864 ;
  assign n19866 = x98 & n8834 ;
  assign n19867 = x97 & n8829 ;
  assign n19868 = x96 & ~n8828 ;
  assign n19869 = n9159 & n19868 ;
  assign n19870 = n19867 | n19869 ;
  assign n19871 = n19866 | n19870 ;
  assign n19872 = n8837 | n19871 ;
  assign n19873 = ( n4105 & n19871 ) | ( n4105 & n19872 ) | ( n19871 & n19872 ) ;
  assign n19874 = x53 & n19873 ;
  assign n19875 = x53 & ~n19874 ;
  assign n19876 = ( n19873 & ~n19874 ) | ( n19873 & n19875 ) | ( ~n19874 & n19875 ) ;
  assign n19877 = ( n19809 & ~n19864 ) | ( n19809 & n19876 ) | ( ~n19864 & n19876 ) ;
  assign n19878 = n19865 | n19877 ;
  assign n19879 = ( n19660 & n19662 ) | ( n19660 & ~n19663 ) | ( n19662 & ~n19663 ) ;
  assign n19880 = n19809 & ~n19864 ;
  assign n19881 = n19865 | n19880 ;
  assign n19882 = n19876 & n19881 ;
  assign n19883 = n19879 | n19882 ;
  assign n19884 = n19878 & ~n19883 ;
  assign n19885 = ( ~n19878 & n19879 ) | ( ~n19878 & n19882 ) | ( n19879 & n19882 ) ;
  assign n19886 = n19884 | n19885 ;
  assign n19887 = x101 & n7812 ;
  assign n19888 = x100 & n7807 ;
  assign n19889 = x99 & ~n7806 ;
  assign n19890 = n8136 & n19889 ;
  assign n19891 = n19888 | n19890 ;
  assign n19892 = n19887 | n19891 ;
  assign n19893 = n7815 | n19892 ;
  assign n19894 = ( n4783 & n19892 ) | ( n4783 & n19893 ) | ( n19892 & n19893 ) ;
  assign n19895 = x50 & n19894 ;
  assign n19896 = x50 & ~n19895 ;
  assign n19897 = ( n19894 & ~n19895 ) | ( n19894 & n19896 ) | ( ~n19895 & n19896 ) ;
  assign n19898 = n19886 & ~n19897 ;
  assign n19899 = ~n19886 & n19897 ;
  assign n19900 = n19898 | n19899 ;
  assign n19901 = n19677 | n19682 ;
  assign n19902 = n19900 & n19901 ;
  assign n19903 = ~n19900 & n19901 ;
  assign n19904 = n19900 | n19903 ;
  assign n19905 = x104 & n6937 ;
  assign n19906 = x103 & n6932 ;
  assign n19907 = x102 & ~n6931 ;
  assign n19908 = n7216 & n19907 ;
  assign n19909 = n19906 | n19908 ;
  assign n19910 = n19905 | n19909 ;
  assign n19911 = n6940 | n19910 ;
  assign n19912 = ( n5295 & n19910 ) | ( n5295 & n19911 ) | ( n19910 & n19911 ) ;
  assign n19913 = x47 & n19912 ;
  assign n19914 = x47 & ~n19913 ;
  assign n19915 = ( n19912 & ~n19913 ) | ( n19912 & n19914 ) | ( ~n19913 & n19914 ) ;
  assign n19916 = n19904 & ~n19915 ;
  assign n19917 = ~n19902 & n19916 ;
  assign n19918 = ( n19902 & ~n19904 ) | ( n19902 & n19915 ) | ( ~n19904 & n19915 ) ;
  assign n19919 = n19917 | n19918 ;
  assign n19920 = n19684 | n19688 ;
  assign n19921 = ( n19808 & n19919 ) | ( n19808 & ~n19920 ) | ( n19919 & ~n19920 ) ;
  assign n19922 = ( ~n19919 & n19920 ) | ( ~n19919 & n19921 ) | ( n19920 & n19921 ) ;
  assign n19923 = ( ~n19808 & n19921 ) | ( ~n19808 & n19922 ) | ( n19921 & n19922 ) ;
  assign n19924 = ~n19797 & n19923 ;
  assign n19925 = n19797 & ~n19923 ;
  assign n19926 = n19924 | n19925 ;
  assign n19927 = x110 & n5340 ;
  assign n19928 = x109 & n5335 ;
  assign n19929 = x108 & ~n5334 ;
  assign n19930 = n5580 & n19929 ;
  assign n19931 = n19928 | n19930 ;
  assign n19932 = n19927 | n19931 ;
  assign n19933 = n5343 | n19932 ;
  assign n19934 = ( n7189 & n19932 ) | ( n7189 & n19933 ) | ( n19932 & n19933 ) ;
  assign n19935 = x41 & n19934 ;
  assign n19936 = x41 & ~n19935 ;
  assign n19937 = ( n19934 & ~n19935 ) | ( n19934 & n19936 ) | ( ~n19935 & n19936 ) ;
  assign n19938 = n19926 & n19937 ;
  assign n19939 = ( n19797 & ~n19923 ) | ( n19797 & n19937 ) | ( ~n19923 & n19937 ) ;
  assign n19940 = n19924 | n19939 ;
  assign n19941 = ~n19938 & n19940 ;
  assign n19942 = n19696 | n19700 ;
  assign n19943 = n19941 & ~n19942 ;
  assign n19944 = ~n19941 & n19942 ;
  assign n19945 = n19943 | n19944 ;
  assign n19946 = x113 & n4572 ;
  assign n19947 = x112 & n4567 ;
  assign n19948 = x111 & ~n4566 ;
  assign n19949 = n4828 & n19948 ;
  assign n19950 = n19947 | n19949 ;
  assign n19951 = n19946 | n19950 ;
  assign n19952 = n4575 | n19951 ;
  assign n19953 = ( n8113 & n19951 ) | ( n8113 & n19952 ) | ( n19951 & n19952 ) ;
  assign n19954 = x38 & n19953 ;
  assign n19955 = x38 & ~n19954 ;
  assign n19956 = ( n19953 & ~n19954 ) | ( n19953 & n19955 ) | ( ~n19954 & n19955 ) ;
  assign n19957 = n19945 & n19956 ;
  assign n19958 = ( ~n19941 & n19942 ) | ( ~n19941 & n19956 ) | ( n19942 & n19956 ) ;
  assign n19959 = n19943 | n19958 ;
  assign n19960 = ~n19957 & n19959 ;
  assign n19961 = ~n19713 & n19719 ;
  assign n19962 = ( n19796 & n19960 ) | ( n19796 & ~n19961 ) | ( n19960 & ~n19961 ) ;
  assign n19963 = ( ~n19960 & n19961 ) | ( ~n19960 & n19962 ) | ( n19961 & n19962 ) ;
  assign n19964 = ( ~n19796 & n19962 ) | ( ~n19796 & n19963 ) | ( n19962 & n19963 ) ;
  assign n19965 = x122 & n2775 ;
  assign n19966 = x121 & n2770 ;
  assign n19967 = x120 & ~n2769 ;
  assign n19968 = n2978 & n19967 ;
  assign n19969 = n19966 | n19968 ;
  assign n19970 = n19965 | n19969 ;
  assign n19971 = n2778 | n19970 ;
  assign n19972 = ( n11188 & n19970 ) | ( n11188 & n19971 ) | ( n19970 & n19971 ) ;
  assign n19973 = x29 & n19972 ;
  assign n19974 = x29 & ~n19973 ;
  assign n19975 = ( n19972 & ~n19973 ) | ( n19972 & n19974 ) | ( ~n19973 & n19974 ) ;
  assign n19976 = ( n19738 & n19764 ) | ( n19738 & n19765 ) | ( n19764 & n19765 ) ;
  assign n19977 = n19975 | n19976 ;
  assign n19978 = n19975 & n19976 ;
  assign n19979 = n19977 & ~n19978 ;
  assign n19980 = n19732 | n19736 ;
  assign n19981 = x119 & n3314 ;
  assign n19982 = x118 & n3309 ;
  assign n19983 = x117 & ~n3308 ;
  assign n19984 = n3570 & n19983 ;
  assign n19985 = n19982 | n19984 ;
  assign n19986 = n19981 | n19985 ;
  assign n19987 = n3317 | n19986 ;
  assign n19988 = ( n9789 & n19986 ) | ( n9789 & n19987 ) | ( n19986 & n19987 ) ;
  assign n19989 = x32 & n19988 ;
  assign n19990 = x32 & ~n19989 ;
  assign n19991 = ( n19988 & ~n19989 ) | ( n19988 & n19990 ) | ( ~n19989 & n19990 ) ;
  assign n19992 = n19980 | n19991 ;
  assign n19993 = ~n19991 & n19992 ;
  assign n19994 = ( ~n19980 & n19992 ) | ( ~n19980 & n19993 ) | ( n19992 & n19993 ) ;
  assign n19995 = ( n19964 & n19979 ) | ( n19964 & ~n19994 ) | ( n19979 & ~n19994 ) ;
  assign n19996 = ( ~n19979 & n19994 ) | ( ~n19979 & n19995 ) | ( n19994 & n19995 ) ;
  assign n19997 = ( ~n19964 & n19995 ) | ( ~n19964 & n19996 ) | ( n19995 & n19996 ) ;
  assign n19998 = x127 & n1812 ;
  assign n19999 = x126 & ~n1811 ;
  assign n20000 = n1977 & n19999 ;
  assign n20001 = n19998 | n20000 ;
  assign n20002 = n1820 | n20001 ;
  assign n20003 = ( n13461 & n20001 ) | ( n13461 & n20002 ) | ( n20001 & n20002 ) ;
  assign n20004 = x23 & n20003 ;
  assign n20005 = x23 & ~n20004 ;
  assign n20006 = ( n20003 & ~n20004 ) | ( n20003 & n20005 ) | ( ~n20004 & n20005 ) ;
  assign n20007 = ( n19527 & n19528 ) | ( n19527 & n19771 ) | ( n19528 & n19771 ) ;
  assign n20008 = n20006 | n20007 ;
  assign n20009 = n20006 & n20007 ;
  assign n20010 = n20008 & ~n20009 ;
  assign n20011 = x125 & n2280 ;
  assign n20012 = x124 & n2275 ;
  assign n20013 = x123 & ~n2274 ;
  assign n20014 = n2481 & n20013 ;
  assign n20015 = n20012 | n20014 ;
  assign n20016 = n20011 | n20015 ;
  assign n20017 = n2283 | n20016 ;
  assign n20018 = ( n12310 & n20016 ) | ( n12310 & n20017 ) | ( n20016 & n20017 ) ;
  assign n20019 = x26 & n20018 ;
  assign n20020 = x26 & ~n20019 ;
  assign n20021 = ( n20018 & ~n20019 ) | ( n20018 & n20020 ) | ( ~n20019 & n20020 ) ;
  assign n20022 = ( n19749 & n19750 ) | ( n19749 & ~n19771 ) | ( n19750 & ~n19771 ) ;
  assign n20023 = n20021 | n20022 ;
  assign n20024 = n20021 & n20022 ;
  assign n20025 = n20023 & ~n20024 ;
  assign n20026 = ( n19997 & n20010 ) | ( n19997 & ~n20025 ) | ( n20010 & ~n20025 ) ;
  assign n20027 = ( ~n20010 & n20025 ) | ( ~n20010 & n20026 ) | ( n20025 & n20026 ) ;
  assign n20028 = ( ~n19997 & n20026 ) | ( ~n19997 & n20027 ) | ( n20026 & n20027 ) ;
  assign n20029 = ( n19532 & n19543 ) | ( n19532 & ~n19774 ) | ( n19543 & ~n19774 ) ;
  assign n20030 = n20028 | n20029 ;
  assign n20031 = n20028 & n20029 ;
  assign n20032 = n20030 & ~n20031 ;
  assign n20033 = n19776 | n19782 ;
  assign n20034 = n19776 | n19783 ;
  assign n20035 = ( n17506 & n20033 ) | ( n17506 & n20034 ) | ( n20033 & n20034 ) ;
  assign n20036 = n20032 | n20035 ;
  assign n20037 = n20032 & n20033 ;
  assign n20038 = n20032 & n20034 ;
  assign n20039 = ( n17506 & n20037 ) | ( n17506 & n20038 ) | ( n20037 & n20038 ) ;
  assign n20040 = n20036 & ~n20039 ;
  assign n20041 = ( n20006 & n20007 ) | ( n20006 & ~n20028 ) | ( n20007 & ~n20028 ) ;
  assign n20042 = x123 & n2775 ;
  assign n20043 = x122 & n2770 ;
  assign n20044 = x121 & ~n2769 ;
  assign n20045 = n2978 & n20044 ;
  assign n20046 = n20043 | n20045 ;
  assign n20047 = n20042 | n20046 ;
  assign n20048 = n2778 | n20047 ;
  assign n20049 = ( n11219 & n20047 ) | ( n11219 & n20048 ) | ( n20047 & n20048 ) ;
  assign n20050 = x29 & n20049 ;
  assign n20051 = x29 & ~n20050 ;
  assign n20052 = ( n20049 & ~n20050 ) | ( n20049 & n20051 ) | ( ~n20050 & n20051 ) ;
  assign n20053 = ( n19964 & n19980 ) | ( n19964 & n19991 ) | ( n19980 & n19991 ) ;
  assign n20054 = ~n20052 & n20053 ;
  assign n20055 = n20052 & n20053 ;
  assign n20056 = ( n20052 & n20054 ) | ( n20052 & ~n20055 ) | ( n20054 & ~n20055 ) ;
  assign n20057 = x117 & n3913 ;
  assign n20058 = x116 & n3908 ;
  assign n20059 = x115 & ~n3907 ;
  assign n20060 = n4152 & n20059 ;
  assign n20061 = n20058 | n20060 ;
  assign n20062 = n20057 | n20061 ;
  assign n20063 = n3916 | n20062 ;
  assign n20064 = ( n9118 & n20062 ) | ( n9118 & n20063 ) | ( n20062 & n20063 ) ;
  assign n20065 = x35 & n20064 ;
  assign n20066 = x35 & ~n20065 ;
  assign n20067 = ( n20064 & ~n20065 ) | ( n20064 & n20066 ) | ( ~n20065 & n20066 ) ;
  assign n20068 = x111 & n5340 ;
  assign n20069 = x110 & n5335 ;
  assign n20070 = x109 & ~n5334 ;
  assign n20071 = n5580 & n20070 ;
  assign n20072 = n20069 | n20071 ;
  assign n20073 = n20068 | n20072 ;
  assign n20074 = n5343 | n20073 ;
  assign n20075 = ( n7492 & n20073 ) | ( n7492 & n20074 ) | ( n20073 & n20074 ) ;
  assign n20076 = x41 & n20075 ;
  assign n20077 = x41 & ~n20076 ;
  assign n20078 = ( n20075 & ~n20076 ) | ( n20075 & n20077 ) | ( ~n20076 & n20077 ) ;
  assign n20079 = n19903 | n19918 ;
  assign n20080 = x105 & n6937 ;
  assign n20081 = x104 & n6932 ;
  assign n20082 = x103 & ~n6931 ;
  assign n20083 = n7216 & n20082 ;
  assign n20084 = n20081 | n20083 ;
  assign n20085 = n20080 | n20084 ;
  assign n20086 = n6940 | n20085 ;
  assign n20087 = ( n5788 & n20085 ) | ( n5788 & n20086 ) | ( n20085 & n20086 ) ;
  assign n20088 = x47 & n20087 ;
  assign n20089 = x47 & ~n20088 ;
  assign n20090 = ( n20087 & ~n20088 ) | ( n20087 & n20089 ) | ( ~n20088 & n20089 ) ;
  assign n20091 = n19885 | n19899 ;
  assign n20092 = x102 & n7812 ;
  assign n20093 = x101 & n7807 ;
  assign n20094 = x100 & ~n7806 ;
  assign n20095 = n8136 & n20094 ;
  assign n20096 = n20093 | n20095 ;
  assign n20097 = n20092 | n20096 ;
  assign n20098 = n7815 | n20097 ;
  assign n20099 = ( n5025 & n20097 ) | ( n5025 & n20098 ) | ( n20097 & n20098 ) ;
  assign n20100 = x50 & n20099 ;
  assign n20101 = x50 & ~n20100 ;
  assign n20102 = ( n20099 & ~n20100 ) | ( n20099 & n20101 ) | ( ~n20100 & n20101 ) ;
  assign n20103 = n19844 | n19858 ;
  assign n20104 = x93 & n10876 ;
  assign n20105 = x92 & n10871 ;
  assign n20106 = x91 & ~n10870 ;
  assign n20107 = n11305 & n20106 ;
  assign n20108 = n20105 | n20107 ;
  assign n20109 = n20104 | n20108 ;
  assign n20110 = n10879 | n20109 ;
  assign n20111 = ( n2931 & n20109 ) | ( n2931 & n20110 ) | ( n20109 & n20110 ) ;
  assign n20112 = x59 & n20111 ;
  assign n20113 = x59 & ~n20112 ;
  assign n20114 = ( n20111 & ~n20112 ) | ( n20111 & n20113 ) | ( ~n20112 & n20113 ) ;
  assign n20115 = x87 & n12808 ;
  assign n20116 = x63 & x86 ;
  assign n20117 = ~n12808 & n20116 ;
  assign n20118 = n20115 | n20117 ;
  assign n20119 = n19824 & ~n20118 ;
  assign n20120 = ~n19824 & n20118 ;
  assign n20121 = n20119 | n20120 ;
  assign n20122 = x90 & n11984 ;
  assign n20123 = x89 & n11979 ;
  assign n20124 = x88 & ~n11978 ;
  assign n20125 = n12430 & n20124 ;
  assign n20126 = n20123 | n20125 ;
  assign n20127 = n20122 | n20126 ;
  assign n20128 = n11987 | n20127 ;
  assign n20129 = ( n2410 & n20127 ) | ( n2410 & n20128 ) | ( n20127 & n20128 ) ;
  assign n20130 = x62 & n20129 ;
  assign n20131 = x62 & ~n20130 ;
  assign n20132 = ( n20129 & ~n20130 ) | ( n20129 & n20131 ) | ( ~n20130 & n20131 ) ;
  assign n20133 = ~n20121 & n20132 ;
  assign n20134 = n20121 & ~n20132 ;
  assign n20135 = n20133 | n20134 ;
  assign n20136 = n19827 | n19840 ;
  assign n20137 = ( n20114 & n20135 ) | ( n20114 & ~n20136 ) | ( n20135 & ~n20136 ) ;
  assign n20138 = ( ~n20135 & n20136 ) | ( ~n20135 & n20137 ) | ( n20136 & n20137 ) ;
  assign n20139 = ( ~n20114 & n20137 ) | ( ~n20114 & n20138 ) | ( n20137 & n20138 ) ;
  assign n20140 = ~n20103 & n20139 ;
  assign n20141 = n20103 & ~n20139 ;
  assign n20142 = n20140 | n20141 ;
  assign n20143 = x96 & n9853 ;
  assign n20144 = x95 & n9848 ;
  assign n20145 = x94 & ~n9847 ;
  assign n20146 = n10165 & n20145 ;
  assign n20147 = n20144 | n20146 ;
  assign n20148 = n20143 | n20147 ;
  assign n20149 = n9856 | n20148 ;
  assign n20150 = ( n3509 & n20148 ) | ( n3509 & n20149 ) | ( n20148 & n20149 ) ;
  assign n20151 = x56 & n20150 ;
  assign n20152 = x56 & ~n20151 ;
  assign n20153 = ( n20150 & ~n20151 ) | ( n20150 & n20152 ) | ( ~n20151 & n20152 ) ;
  assign n20154 = n20142 & ~n20153 ;
  assign n20155 = ~n20142 & n20153 ;
  assign n20156 = n20154 | n20155 ;
  assign n20157 = n19863 & ~n20156 ;
  assign n20158 = ~n19863 & n20156 ;
  assign n20159 = n20157 | n20158 ;
  assign n20160 = x99 & n8834 ;
  assign n20161 = x98 & n8829 ;
  assign n20162 = x97 & ~n8828 ;
  assign n20163 = n9159 & n20162 ;
  assign n20164 = n20161 | n20163 ;
  assign n20165 = n20160 | n20164 ;
  assign n20166 = n8837 | n20165 ;
  assign n20167 = ( n4325 & n20165 ) | ( n4325 & n20166 ) | ( n20165 & n20166 ) ;
  assign n20168 = x53 & n20167 ;
  assign n20169 = x53 & ~n20168 ;
  assign n20170 = ( n20167 & ~n20168 ) | ( n20167 & n20169 ) | ( ~n20168 & n20169 ) ;
  assign n20171 = ~n20159 & n20170 ;
  assign n20172 = n20159 & ~n20170 ;
  assign n20173 = n20171 | n20172 ;
  assign n20174 = ( n19877 & n20102 ) | ( n19877 & ~n20173 ) | ( n20102 & ~n20173 ) ;
  assign n20175 = ( ~n19877 & n20173 ) | ( ~n19877 & n20174 ) | ( n20173 & n20174 ) ;
  assign n20176 = ( ~n20102 & n20174 ) | ( ~n20102 & n20175 ) | ( n20174 & n20175 ) ;
  assign n20177 = ( n20090 & ~n20091 ) | ( n20090 & n20176 ) | ( ~n20091 & n20176 ) ;
  assign n20178 = ( n20091 & ~n20176 ) | ( n20091 & n20177 ) | ( ~n20176 & n20177 ) ;
  assign n20179 = ( ~n20090 & n20177 ) | ( ~n20090 & n20178 ) | ( n20177 & n20178 ) ;
  assign n20180 = n20079 & ~n20179 ;
  assign n20181 = ~n20079 & n20179 ;
  assign n20182 = n20180 | n20181 ;
  assign n20183 = x108 & n6068 ;
  assign n20184 = x107 & n6063 ;
  assign n20185 = x106 & ~n6062 ;
  assign n20186 = n6398 & n20185 ;
  assign n20187 = n20184 | n20186 ;
  assign n20188 = n20183 | n20187 ;
  assign n20189 = n6071 | n20188 ;
  assign n20190 = ( n6358 & n20188 ) | ( n6358 & n20189 ) | ( n20188 & n20189 ) ;
  assign n20191 = x44 & n20190 ;
  assign n20192 = x44 & ~n20191 ;
  assign n20193 = ( n20190 & ~n20191 ) | ( n20190 & n20192 ) | ( ~n20191 & n20192 ) ;
  assign n20194 = ~n20182 & n20193 ;
  assign n20195 = n20182 & ~n20193 ;
  assign n20196 = n20194 | n20195 ;
  assign n20197 = ( ~n19922 & n20078 ) | ( ~n19922 & n20196 ) | ( n20078 & n20196 ) ;
  assign n20198 = ( n19922 & ~n20196 ) | ( n19922 & n20197 ) | ( ~n20196 & n20197 ) ;
  assign n20199 = ( ~n20078 & n20197 ) | ( ~n20078 & n20198 ) | ( n20197 & n20198 ) ;
  assign n20200 = ~n19939 & n20199 ;
  assign n20201 = n19939 & ~n20199 ;
  assign n20202 = n20200 | n20201 ;
  assign n20203 = x114 & n4572 ;
  assign n20204 = x113 & n4567 ;
  assign n20205 = x112 & ~n4566 ;
  assign n20206 = n4828 & n20205 ;
  assign n20207 = n20204 | n20206 ;
  assign n20208 = n20203 | n20207 ;
  assign n20209 = n4575 | n20208 ;
  assign n20210 = ( n8437 & n20208 ) | ( n8437 & n20209 ) | ( n20208 & n20209 ) ;
  assign n20211 = x38 & n20210 ;
  assign n20212 = x38 & ~n20211 ;
  assign n20213 = ( n20210 & ~n20211 ) | ( n20210 & n20212 ) | ( ~n20211 & n20212 ) ;
  assign n20214 = n20202 & ~n20213 ;
  assign n20215 = ~n20202 & n20213 ;
  assign n20216 = n20214 | n20215 ;
  assign n20217 = ( n19958 & n20067 ) | ( n19958 & ~n20216 ) | ( n20067 & ~n20216 ) ;
  assign n20218 = ( ~n19958 & n20216 ) | ( ~n19958 & n20217 ) | ( n20216 & n20217 ) ;
  assign n20219 = ( ~n20067 & n20217 ) | ( ~n20067 & n20218 ) | ( n20217 & n20218 ) ;
  assign n20220 = ( ~n19796 & n19960 ) | ( ~n19796 & n19961 ) | ( n19960 & n19961 ) ;
  assign n20221 = x120 & n3314 ;
  assign n20222 = x119 & n3309 ;
  assign n20223 = x118 & ~n3308 ;
  assign n20224 = n3570 & n20223 ;
  assign n20225 = n20222 | n20224 ;
  assign n20226 = n20221 | n20225 ;
  assign n20227 = n3317 | n20226 ;
  assign n20228 = ( n10460 & n20226 ) | ( n10460 & n20227 ) | ( n20226 & n20227 ) ;
  assign n20229 = x32 & n20228 ;
  assign n20230 = x32 & ~n20229 ;
  assign n20231 = ( n20228 & ~n20229 ) | ( n20228 & n20230 ) | ( ~n20229 & n20230 ) ;
  assign n20232 = ( n20219 & n20220 ) | ( n20219 & ~n20231 ) | ( n20220 & ~n20231 ) ;
  assign n20233 = ( ~n20220 & n20231 ) | ( ~n20220 & n20232 ) | ( n20231 & n20232 ) ;
  assign n20234 = ( ~n20219 & n20232 ) | ( ~n20219 & n20233 ) | ( n20232 & n20233 ) ;
  assign n20235 = n20056 & ~n20234 ;
  assign n20236 = ~n20056 & n20234 ;
  assign n20237 = n20235 | n20236 ;
  assign n20238 = x126 & n2280 ;
  assign n20239 = x125 & n2275 ;
  assign n20240 = x124 & ~n2274 ;
  assign n20241 = n2481 & n20240 ;
  assign n20242 = n20239 | n20241 ;
  assign n20243 = n20238 | n20242 ;
  assign n20244 = n2283 | n20243 ;
  assign n20245 = ( n12687 & n20243 ) | ( n12687 & n20244 ) | ( n20243 & n20244 ) ;
  assign n20246 = x26 & n20245 ;
  assign n20247 = x26 & ~n20246 ;
  assign n20248 = ( n20245 & ~n20246 ) | ( n20245 & n20247 ) | ( ~n20246 & n20247 ) ;
  assign n20249 = ( n19975 & n19976 ) | ( n19975 & ~n19997 ) | ( n19976 & ~n19997 ) ;
  assign n20250 = ( n20237 & n20248 ) | ( n20237 & ~n20249 ) | ( n20248 & ~n20249 ) ;
  assign n20251 = ( ~n20248 & n20249 ) | ( ~n20248 & n20250 ) | ( n20249 & n20250 ) ;
  assign n20252 = ( ~n20237 & n20250 ) | ( ~n20237 & n20251 ) | ( n20250 & n20251 ) ;
  assign n20253 = x127 & ~n1811 ;
  assign n20254 = n1977 & n20253 ;
  assign n20255 = ( x127 & n1820 ) | ( x127 & n20254 ) | ( n1820 & n20254 ) ;
  assign n20256 = ( x126 & n20254 ) | ( x126 & n20255 ) | ( n20254 & n20255 ) ;
  assign n20257 = ( n12685 & n20255 ) | ( n12685 & n20256 ) | ( n20255 & n20256 ) ;
  assign n20258 = x23 & n20257 ;
  assign n20259 = x23 & ~n20258 ;
  assign n20260 = ( n20257 & ~n20258 ) | ( n20257 & n20259 ) | ( ~n20258 & n20259 ) ;
  assign n20261 = ( n19997 & n20021 ) | ( n19997 & n20022 ) | ( n20021 & n20022 ) ;
  assign n20262 = ( n20252 & n20260 ) | ( n20252 & ~n20261 ) | ( n20260 & ~n20261 ) ;
  assign n20263 = ( ~n20260 & n20261 ) | ( ~n20260 & n20262 ) | ( n20261 & n20262 ) ;
  assign n20264 = ( ~n20252 & n20262 ) | ( ~n20252 & n20263 ) | ( n20262 & n20263 ) ;
  assign n20265 = n20041 & n20264 ;
  assign n20266 = n20041 & ~n20265 ;
  assign n20267 = n20264 & ~n20265 ;
  assign n20268 = n20266 | n20267 ;
  assign n20269 = n20031 | n20037 ;
  assign n20270 = n20268 & n20269 ;
  assign n20271 = n20031 | n20038 ;
  assign n20272 = n20268 & n20271 ;
  assign n20273 = ( n17506 & n20270 ) | ( n17506 & n20272 ) | ( n20270 & n20272 ) ;
  assign n20274 = ( n17506 & n20269 ) | ( n17506 & n20271 ) | ( n20269 & n20271 ) ;
  assign n20275 = ~n20273 & n20274 ;
  assign n20276 = ( n20268 & ~n20273 ) | ( n20268 & n20275 ) | ( ~n20273 & n20275 ) ;
  assign n20277 = n20201 | n20215 ;
  assign n20278 = x109 & n6068 ;
  assign n20279 = x108 & n6063 ;
  assign n20280 = x107 & ~n6062 ;
  assign n20281 = n6398 & n20280 ;
  assign n20282 = n20279 | n20281 ;
  assign n20283 = n20278 | n20282 ;
  assign n20284 = n6071 | n20283 ;
  assign n20285 = ( n6884 & n20283 ) | ( n6884 & n20284 ) | ( n20283 & n20284 ) ;
  assign n20286 = x44 & n20285 ;
  assign n20287 = x44 & ~n20286 ;
  assign n20288 = ( n20285 & ~n20286 ) | ( n20285 & n20287 ) | ( ~n20286 & n20287 ) ;
  assign n20289 = x106 & n6937 ;
  assign n20290 = x105 & n6932 ;
  assign n20291 = x104 & ~n6931 ;
  assign n20292 = n7216 & n20291 ;
  assign n20293 = n20290 | n20292 ;
  assign n20294 = n20289 | n20293 ;
  assign n20295 = n6940 | n20294 ;
  assign n20296 = ( n5814 & n20294 ) | ( n5814 & n20295 ) | ( n20294 & n20295 ) ;
  assign n20297 = x47 & n20296 ;
  assign n20298 = x47 & ~n20297 ;
  assign n20299 = ( n20296 & ~n20297 ) | ( n20296 & n20298 ) | ( ~n20297 & n20298 ) ;
  assign n20300 = x88 & n12808 ;
  assign n20301 = x63 & x87 ;
  assign n20302 = ~n12808 & n20301 ;
  assign n20303 = n20300 | n20302 ;
  assign n20304 = ~x23 & n20303 ;
  assign n20305 = x23 & ~n20303 ;
  assign n20306 = n20304 | n20305 ;
  assign n20307 = n20118 & ~n20306 ;
  assign n20308 = ~n20118 & n20306 ;
  assign n20309 = n20307 | n20308 ;
  assign n20310 = x91 & n11984 ;
  assign n20311 = x90 & n11979 ;
  assign n20312 = x89 & ~n11978 ;
  assign n20313 = n12430 & n20312 ;
  assign n20314 = n20311 | n20313 ;
  assign n20315 = n20310 | n20314 ;
  assign n20316 = n11987 | n20315 ;
  assign n20317 = ( n2714 & n20315 ) | ( n2714 & n20316 ) | ( n20315 & n20316 ) ;
  assign n20318 = ~x62 & n20317 ;
  assign n20319 = x62 & ~n20317 ;
  assign n20320 = n20318 | n20319 ;
  assign n20321 = ~n20309 & n20320 ;
  assign n20322 = n20309 & ~n20320 ;
  assign n20323 = n20321 | n20322 ;
  assign n20324 = n20119 | n20133 ;
  assign n20325 = n20323 & n20324 ;
  assign n20326 = n20323 | n20324 ;
  assign n20327 = ~n20325 & n20326 ;
  assign n20328 = x94 & n10876 ;
  assign n20329 = x93 & n10871 ;
  assign n20330 = x92 & ~n10870 ;
  assign n20331 = n11305 & n20330 ;
  assign n20332 = n20329 | n20331 ;
  assign n20333 = n20328 | n20332 ;
  assign n20334 = n10879 | n20333 ;
  assign n20335 = ( n3271 & n20333 ) | ( n3271 & n20334 ) | ( n20333 & n20334 ) ;
  assign n20336 = x59 & n20335 ;
  assign n20337 = x59 & ~n20336 ;
  assign n20338 = ( n20335 & ~n20336 ) | ( n20335 & n20337 ) | ( ~n20336 & n20337 ) ;
  assign n20339 = ~n20327 & n20338 ;
  assign n20340 = n20327 & ~n20338 ;
  assign n20341 = n20339 | n20340 ;
  assign n20342 = ~n20138 & n20341 ;
  assign n20343 = n20138 & ~n20341 ;
  assign n20344 = n20342 | n20343 ;
  assign n20345 = x97 & n9853 ;
  assign n20346 = x96 & n9848 ;
  assign n20347 = x95 & ~n9847 ;
  assign n20348 = n10165 & n20347 ;
  assign n20349 = n20346 | n20348 ;
  assign n20350 = n20345 | n20349 ;
  assign n20351 = n9856 | n20350 ;
  assign n20352 = ( n3707 & n20350 ) | ( n3707 & n20351 ) | ( n20350 & n20351 ) ;
  assign n20353 = x56 & n20352 ;
  assign n20354 = x56 & ~n20353 ;
  assign n20355 = ( n20352 & ~n20353 ) | ( n20352 & n20354 ) | ( ~n20353 & n20354 ) ;
  assign n20356 = n20141 | n20155 ;
  assign n20357 = n20355 & n20356 ;
  assign n20358 = n20355 | n20356 ;
  assign n20359 = ~n20357 & n20358 ;
  assign n20360 = ~n20344 & n20359 ;
  assign n20361 = n20344 & ~n20359 ;
  assign n20362 = n20360 | n20361 ;
  assign n20363 = x100 & n8834 ;
  assign n20364 = x99 & n8829 ;
  assign n20365 = x98 & ~n8828 ;
  assign n20366 = n9159 & n20365 ;
  assign n20367 = n20364 | n20366 ;
  assign n20368 = n20363 | n20367 ;
  assign n20369 = n8837 | n20368 ;
  assign n20370 = ( n4532 & n20368 ) | ( n4532 & n20369 ) | ( n20368 & n20369 ) ;
  assign n20371 = x53 & n20370 ;
  assign n20372 = x53 & ~n20371 ;
  assign n20373 = ( n20370 & ~n20371 ) | ( n20370 & n20372 ) | ( ~n20371 & n20372 ) ;
  assign n20374 = ~n20362 & n20373 ;
  assign n20375 = n20362 | n20374 ;
  assign n20376 = n20362 & n20373 ;
  assign n20377 = n20157 | n20171 ;
  assign n20378 = n20376 | n20377 ;
  assign n20379 = n20375 & ~n20378 ;
  assign n20380 = ( ~n20375 & n20376 ) | ( ~n20375 & n20377 ) | ( n20376 & n20377 ) ;
  assign n20381 = n20379 | n20380 ;
  assign n20382 = x103 & n7812 ;
  assign n20383 = x102 & n7807 ;
  assign n20384 = x101 & ~n7806 ;
  assign n20385 = n8136 & n20384 ;
  assign n20386 = n20383 | n20385 ;
  assign n20387 = n20382 | n20386 ;
  assign n20388 = n7815 | n20387 ;
  assign n20389 = ( n5264 & n20387 ) | ( n5264 & n20388 ) | ( n20387 & n20388 ) ;
  assign n20390 = x50 & n20389 ;
  assign n20391 = x50 & ~n20390 ;
  assign n20392 = ( n20389 & ~n20390 ) | ( n20389 & n20391 ) | ( ~n20390 & n20391 ) ;
  assign n20393 = ~n20381 & n20392 ;
  assign n20394 = n20381 | n20393 ;
  assign n20395 = n20381 & n20392 ;
  assign n20396 = n20174 | n20395 ;
  assign n20397 = n20394 & ~n20396 ;
  assign n20398 = ( n20174 & ~n20394 ) | ( n20174 & n20395 ) | ( ~n20394 & n20395 ) ;
  assign n20399 = n20397 | n20398 ;
  assign n20400 = ( n20178 & n20299 ) | ( n20178 & ~n20399 ) | ( n20299 & ~n20399 ) ;
  assign n20401 = ( ~n20178 & n20399 ) | ( ~n20178 & n20400 ) | ( n20399 & n20400 ) ;
  assign n20402 = ( ~n20299 & n20400 ) | ( ~n20299 & n20401 ) | ( n20400 & n20401 ) ;
  assign n20403 = n20288 & ~n20402 ;
  assign n20404 = ~n20288 & n20402 ;
  assign n20405 = n20403 | n20404 ;
  assign n20406 = n20180 | n20194 ;
  assign n20407 = n20405 & ~n20406 ;
  assign n20408 = ~n20405 & n20406 ;
  assign n20409 = n20407 | n20408 ;
  assign n20410 = x112 & n5340 ;
  assign n20411 = x111 & n5335 ;
  assign n20412 = x110 & ~n5334 ;
  assign n20413 = n5580 & n20412 ;
  assign n20414 = n20411 | n20413 ;
  assign n20415 = n20410 | n20414 ;
  assign n20416 = n5343 | n20415 ;
  assign n20417 = ( n7789 & n20415 ) | ( n7789 & n20416 ) | ( n20415 & n20416 ) ;
  assign n20418 = x41 & n20417 ;
  assign n20419 = x41 & ~n20418 ;
  assign n20420 = ( n20417 & ~n20418 ) | ( n20417 & n20419 ) | ( ~n20418 & n20419 ) ;
  assign n20421 = ~n20409 & n20420 ;
  assign n20422 = n20409 | n20421 ;
  assign n20423 = n20409 & n20420 ;
  assign n20424 = n20198 | n20423 ;
  assign n20425 = n20422 & ~n20424 ;
  assign n20426 = ( n20198 & ~n20422 ) | ( n20198 & n20423 ) | ( ~n20422 & n20423 ) ;
  assign n20427 = n20425 | n20426 ;
  assign n20428 = x115 & n4572 ;
  assign n20429 = x114 & n4567 ;
  assign n20430 = x113 & ~n4566 ;
  assign n20431 = n4828 & n20430 ;
  assign n20432 = n20429 | n20431 ;
  assign n20433 = n20428 | n20432 ;
  assign n20434 = n4575 | n20433 ;
  assign n20435 = ( n8749 & n20433 ) | ( n8749 & n20434 ) | ( n20433 & n20434 ) ;
  assign n20436 = x38 & n20435 ;
  assign n20437 = x38 & ~n20436 ;
  assign n20438 = ( n20435 & ~n20436 ) | ( n20435 & n20437 ) | ( ~n20436 & n20437 ) ;
  assign n20439 = ~n20427 & n20438 ;
  assign n20440 = n20427 & ~n20438 ;
  assign n20441 = n20439 | n20440 ;
  assign n20442 = n20277 & ~n20441 ;
  assign n20443 = n20277 & ~n20442 ;
  assign n20444 = n20441 | n20442 ;
  assign n20445 = ~n20443 & n20444 ;
  assign n20446 = x118 & n3913 ;
  assign n20447 = x117 & n3908 ;
  assign n20448 = x116 & ~n3907 ;
  assign n20449 = n4152 & n20448 ;
  assign n20450 = n20447 | n20449 ;
  assign n20451 = n20446 | n20450 ;
  assign n20452 = n3916 | n20451 ;
  assign n20453 = ( n9760 & n20451 ) | ( n9760 & n20452 ) | ( n20451 & n20452 ) ;
  assign n20454 = x35 & n20453 ;
  assign n20455 = x35 & ~n20454 ;
  assign n20456 = ( n20453 & ~n20454 ) | ( n20453 & n20455 ) | ( ~n20454 & n20455 ) ;
  assign n20457 = n20445 & ~n20456 ;
  assign n20458 = ~n20445 & n20456 ;
  assign n20459 = n20457 | n20458 ;
  assign n20460 = n20217 & ~n20459 ;
  assign n20461 = ~n20217 & n20459 ;
  assign n20462 = n20460 | n20461 ;
  assign n20463 = x121 & n3314 ;
  assign n20464 = x120 & n3309 ;
  assign n20465 = x119 & ~n3308 ;
  assign n20466 = n3570 & n20465 ;
  assign n20467 = n20464 | n20466 ;
  assign n20468 = n20463 | n20467 ;
  assign n20469 = n3317 | n20468 ;
  assign n20470 = ( n10811 & n20468 ) | ( n10811 & n20469 ) | ( n20468 & n20469 ) ;
  assign n20471 = x32 & n20470 ;
  assign n20472 = x32 & ~n20471 ;
  assign n20473 = ( n20470 & ~n20471 ) | ( n20470 & n20472 ) | ( ~n20471 & n20472 ) ;
  assign n20474 = n20232 & ~n20473 ;
  assign n20475 = ~n20232 & n20473 ;
  assign n20476 = n20474 | n20475 ;
  assign n20477 = ( n20055 & n20056 ) | ( n20055 & ~n20235 ) | ( n20056 & ~n20235 ) ;
  assign n20478 = x124 & n2775 ;
  assign n20479 = x123 & n2770 ;
  assign n20480 = x122 & ~n2769 ;
  assign n20481 = n2978 & n20480 ;
  assign n20482 = n20479 | n20481 ;
  assign n20483 = n20478 | n20482 ;
  assign n20484 = n2778 | n20483 ;
  assign n20485 = ( n11916 & n20483 ) | ( n11916 & n20484 ) | ( n20483 & n20484 ) ;
  assign n20486 = x29 & n20485 ;
  assign n20487 = x29 & ~n20486 ;
  assign n20488 = ( n20485 & ~n20486 ) | ( n20485 & n20487 ) | ( ~n20486 & n20487 ) ;
  assign n20489 = n20477 & n20488 ;
  assign n20490 = n20488 & ~n20489 ;
  assign n20491 = ( n20477 & ~n20489 ) | ( n20477 & n20490 ) | ( ~n20489 & n20490 ) ;
  assign n20492 = ( n20462 & ~n20476 ) | ( n20462 & n20491 ) | ( ~n20476 & n20491 ) ;
  assign n20493 = ( n20462 & n20476 ) | ( n20462 & ~n20491 ) | ( n20476 & ~n20491 ) ;
  assign n20494 = ( ~n20462 & n20492 ) | ( ~n20462 & n20493 ) | ( n20492 & n20493 ) ;
  assign n20495 = x127 & n2280 ;
  assign n20496 = x126 & n2275 ;
  assign n20497 = x125 & ~n2274 ;
  assign n20498 = n2481 & n20497 ;
  assign n20499 = n20496 | n20498 ;
  assign n20500 = n20495 | n20499 ;
  assign n20501 = n2283 | n20500 ;
  assign n20502 = ( n12720 & n20500 ) | ( n12720 & n20501 ) | ( n20500 & n20501 ) ;
  assign n20503 = x26 & n20502 ;
  assign n20504 = x26 & ~n20503 ;
  assign n20505 = ( n20502 & ~n20503 ) | ( n20502 & n20504 ) | ( ~n20503 & n20504 ) ;
  assign n20506 = ( n20237 & n20248 ) | ( n20237 & n20249 ) | ( n20248 & n20249 ) ;
  assign n20507 = ( n20494 & n20505 ) | ( n20494 & ~n20506 ) | ( n20505 & ~n20506 ) ;
  assign n20508 = ( ~n20505 & n20506 ) | ( ~n20505 & n20507 ) | ( n20506 & n20507 ) ;
  assign n20509 = ( ~n20494 & n20507 ) | ( ~n20494 & n20508 ) | ( n20507 & n20508 ) ;
  assign n20510 = ( n20252 & n20260 ) | ( n20252 & n20261 ) | ( n20260 & n20261 ) ;
  assign n20511 = n20509 & ~n20510 ;
  assign n20512 = n20265 | n20273 ;
  assign n20513 = ( ~n20509 & n20510 ) | ( ~n20509 & n20512 ) | ( n20510 & n20512 ) ;
  assign n20514 = ( n20510 & n20511 ) | ( n20510 & n20512 ) | ( n20511 & n20512 ) ;
  assign n20515 = ( ~n20509 & n20511 ) | ( ~n20509 & n20514 ) | ( n20511 & n20514 ) ;
  assign n20516 = ( n20511 & n20513 ) | ( n20511 & ~n20515 ) | ( n20513 & ~n20515 ) ;
  assign n20517 = n20462 | n20476 ;
  assign n20518 = ( n20489 & ~n20493 ) | ( n20489 & n20517 ) | ( ~n20493 & n20517 ) ;
  assign n20519 = x127 & n2275 ;
  assign n20520 = x126 & ~n2274 ;
  assign n20521 = n2481 & n20520 ;
  assign n20522 = n20519 | n20521 ;
  assign n20523 = n2283 | n20522 ;
  assign n20524 = ( n13461 & n20522 ) | ( n13461 & n20523 ) | ( n20522 & n20523 ) ;
  assign n20525 = x26 & n20524 ;
  assign n20526 = x26 & ~n20525 ;
  assign n20527 = ( n20524 & ~n20525 ) | ( n20524 & n20526 ) | ( ~n20525 & n20526 ) ;
  assign n20528 = n20518 & n20527 ;
  assign n20529 = n20518 & ~n20528 ;
  assign n20530 = ~n20518 & n20527 ;
  assign n20531 = x122 & n3314 ;
  assign n20532 = x121 & n3309 ;
  assign n20533 = x120 & ~n3308 ;
  assign n20534 = n3570 & n20533 ;
  assign n20535 = n20532 | n20534 ;
  assign n20536 = n20531 | n20535 ;
  assign n20537 = n3317 | n20536 ;
  assign n20538 = ( n11188 & n20536 ) | ( n11188 & n20537 ) | ( n20536 & n20537 ) ;
  assign n20539 = x32 & n20538 ;
  assign n20540 = x32 & ~n20539 ;
  assign n20541 = ( n20538 & ~n20539 ) | ( n20538 & n20540 ) | ( ~n20539 & n20540 ) ;
  assign n20542 = n20458 | n20541 ;
  assign n20543 = n20460 | n20542 ;
  assign n20544 = ( n20458 & n20460 ) | ( n20458 & n20541 ) | ( n20460 & n20541 ) ;
  assign n20545 = n20543 & ~n20544 ;
  assign n20546 = n20439 | n20442 ;
  assign n20547 = n20421 | n20426 ;
  assign n20548 = x107 & n6937 ;
  assign n20549 = x106 & n6932 ;
  assign n20550 = x105 & ~n6931 ;
  assign n20551 = n7216 & n20550 ;
  assign n20552 = n20549 | n20551 ;
  assign n20553 = n20548 | n20552 ;
  assign n20554 = n6940 | n20553 ;
  assign n20555 = ( n6328 & n20553 ) | ( n6328 & n20554 ) | ( n20553 & n20554 ) ;
  assign n20556 = x47 & n20555 ;
  assign n20557 = x47 & ~n20556 ;
  assign n20558 = ( n20555 & ~n20556 ) | ( n20555 & n20557 ) | ( ~n20556 & n20557 ) ;
  assign n20559 = n20393 | n20398 ;
  assign n20560 = x104 & n7812 ;
  assign n20561 = x103 & n7807 ;
  assign n20562 = x102 & ~n7806 ;
  assign n20563 = n8136 & n20562 ;
  assign n20564 = n20561 | n20563 ;
  assign n20565 = n20560 | n20564 ;
  assign n20566 = n7815 | n20565 ;
  assign n20567 = ( n5295 & n20565 ) | ( n5295 & n20566 ) | ( n20565 & n20566 ) ;
  assign n20568 = x50 & n20567 ;
  assign n20569 = x50 & ~n20568 ;
  assign n20570 = ( n20567 & ~n20568 ) | ( n20567 & n20569 ) | ( ~n20568 & n20569 ) ;
  assign n20571 = n20374 | n20380 ;
  assign n20572 = n20339 | n20343 ;
  assign n20573 = x95 & n10876 ;
  assign n20574 = x94 & n10871 ;
  assign n20575 = x93 & ~n10870 ;
  assign n20576 = n11305 & n20575 ;
  assign n20577 = n20574 | n20576 ;
  assign n20578 = n20573 | n20577 ;
  assign n20579 = n10879 | n20578 ;
  assign n20580 = ( n3479 & n20578 ) | ( n3479 & n20579 ) | ( n20578 & n20579 ) ;
  assign n20581 = x59 & n20580 ;
  assign n20582 = x59 & ~n20581 ;
  assign n20583 = ( n20580 & ~n20581 ) | ( n20580 & n20582 ) | ( ~n20581 & n20582 ) ;
  assign n20584 = x89 & n12808 ;
  assign n20585 = x63 & x88 ;
  assign n20586 = ~n12808 & n20585 ;
  assign n20587 = n20584 | n20586 ;
  assign n20588 = n20304 | n20307 ;
  assign n20589 = n20587 & ~n20588 ;
  assign n20590 = ~n20587 & n20588 ;
  assign n20591 = n20589 | n20590 ;
  assign n20592 = x92 & n11984 ;
  assign n20593 = x91 & n11979 ;
  assign n20594 = x90 & ~n11978 ;
  assign n20595 = n12430 & n20594 ;
  assign n20596 = n20593 | n20595 ;
  assign n20597 = n20592 | n20596 ;
  assign n20598 = n11987 | n20597 ;
  assign n20599 = ( n2904 & n20597 ) | ( n2904 & n20598 ) | ( n20597 & n20598 ) ;
  assign n20600 = x62 & n20599 ;
  assign n20601 = x62 & ~n20600 ;
  assign n20602 = ( n20599 & ~n20600 ) | ( n20599 & n20601 ) | ( ~n20600 & n20601 ) ;
  assign n20603 = ~n20591 & n20602 ;
  assign n20604 = n20591 & ~n20602 ;
  assign n20605 = n20603 | n20604 ;
  assign n20606 = ( n20321 & ~n20323 ) | ( n20321 & n20326 ) | ( ~n20323 & n20326 ) ;
  assign n20607 = ( n20583 & n20605 ) | ( n20583 & ~n20606 ) | ( n20605 & ~n20606 ) ;
  assign n20608 = ( ~n20605 & n20606 ) | ( ~n20605 & n20607 ) | ( n20606 & n20607 ) ;
  assign n20609 = ( ~n20583 & n20607 ) | ( ~n20583 & n20608 ) | ( n20607 & n20608 ) ;
  assign n20610 = ~n20572 & n20609 ;
  assign n20611 = n20572 & ~n20609 ;
  assign n20612 = n20610 | n20611 ;
  assign n20613 = x98 & n9853 ;
  assign n20614 = x97 & n9848 ;
  assign n20615 = x96 & ~n9847 ;
  assign n20616 = n10165 & n20615 ;
  assign n20617 = n20614 | n20616 ;
  assign n20618 = n20613 | n20617 ;
  assign n20619 = n9856 | n20618 ;
  assign n20620 = ( n4105 & n20618 ) | ( n4105 & n20619 ) | ( n20618 & n20619 ) ;
  assign n20621 = x56 & n20620 ;
  assign n20622 = x56 & ~n20621 ;
  assign n20623 = ( n20620 & ~n20621 ) | ( n20620 & n20622 ) | ( ~n20621 & n20622 ) ;
  assign n20624 = n20612 & n20623 ;
  assign n20625 = ( n20572 & ~n20609 ) | ( n20572 & n20623 ) | ( ~n20609 & n20623 ) ;
  assign n20626 = n20610 | n20625 ;
  assign n20627 = ~n20624 & n20626 ;
  assign n20628 = n20357 | n20360 ;
  assign n20629 = n20627 & ~n20628 ;
  assign n20630 = ~n20627 & n20628 ;
  assign n20631 = n20629 | n20630 ;
  assign n20632 = x101 & n8834 ;
  assign n20633 = x100 & n8829 ;
  assign n20634 = x99 & ~n8828 ;
  assign n20635 = n9159 & n20634 ;
  assign n20636 = n20633 | n20635 ;
  assign n20637 = n20632 | n20636 ;
  assign n20638 = n8837 | n20637 ;
  assign n20639 = ( n4783 & n20637 ) | ( n4783 & n20638 ) | ( n20637 & n20638 ) ;
  assign n20640 = x53 & n20639 ;
  assign n20641 = x53 & ~n20640 ;
  assign n20642 = ( n20639 & ~n20640 ) | ( n20639 & n20641 ) | ( ~n20640 & n20641 ) ;
  assign n20643 = n20631 & ~n20642 ;
  assign n20644 = ~n20631 & n20642 ;
  assign n20645 = n20643 | n20644 ;
  assign n20646 = ( n20570 & n20571 ) | ( n20570 & ~n20645 ) | ( n20571 & ~n20645 ) ;
  assign n20647 = ( ~n20571 & n20645 ) | ( ~n20571 & n20646 ) | ( n20645 & n20646 ) ;
  assign n20648 = ( ~n20570 & n20646 ) | ( ~n20570 & n20647 ) | ( n20646 & n20647 ) ;
  assign n20649 = ( n20558 & n20559 ) | ( n20558 & ~n20648 ) | ( n20559 & ~n20648 ) ;
  assign n20650 = ( ~n20559 & n20648 ) | ( ~n20559 & n20649 ) | ( n20648 & n20649 ) ;
  assign n20651 = ( ~n20558 & n20649 ) | ( ~n20558 & n20650 ) | ( n20649 & n20650 ) ;
  assign n20652 = ~n20400 & n20651 ;
  assign n20653 = n20400 & ~n20651 ;
  assign n20654 = n20652 | n20653 ;
  assign n20655 = x110 & n6068 ;
  assign n20656 = x109 & n6063 ;
  assign n20657 = x108 & ~n6062 ;
  assign n20658 = n6398 & n20657 ;
  assign n20659 = n20656 | n20658 ;
  assign n20660 = n20655 | n20659 ;
  assign n20661 = n6071 | n20660 ;
  assign n20662 = ( n7189 & n20660 ) | ( n7189 & n20661 ) | ( n20660 & n20661 ) ;
  assign n20663 = x44 & n20662 ;
  assign n20664 = x44 & ~n20663 ;
  assign n20665 = ( n20662 & ~n20663 ) | ( n20662 & n20664 ) | ( ~n20663 & n20664 ) ;
  assign n20666 = n20654 & n20665 ;
  assign n20667 = n20403 | n20408 ;
  assign n20668 = n20666 | n20667 ;
  assign n20669 = ( n20400 & ~n20651 ) | ( n20400 & n20665 ) | ( ~n20651 & n20665 ) ;
  assign n20670 = n20652 | n20669 ;
  assign n20671 = ~n20668 & n20670 ;
  assign n20672 = ( n20666 & n20667 ) | ( n20666 & ~n20670 ) | ( n20667 & ~n20670 ) ;
  assign n20673 = n20671 | n20672 ;
  assign n20674 = x113 & n5340 ;
  assign n20675 = x112 & n5335 ;
  assign n20676 = x111 & ~n5334 ;
  assign n20677 = n5580 & n20676 ;
  assign n20678 = n20675 | n20677 ;
  assign n20679 = n20674 | n20678 ;
  assign n20680 = n5343 | n20679 ;
  assign n20681 = ( n8113 & n20679 ) | ( n8113 & n20680 ) | ( n20679 & n20680 ) ;
  assign n20682 = x41 & n20681 ;
  assign n20683 = x41 & ~n20682 ;
  assign n20684 = ( n20681 & ~n20682 ) | ( n20681 & n20683 ) | ( ~n20682 & n20683 ) ;
  assign n20685 = n20673 | n20684 ;
  assign n20686 = ~n20684 & n20685 ;
  assign n20687 = ( ~n20673 & n20685 ) | ( ~n20673 & n20686 ) | ( n20685 & n20686 ) ;
  assign n20688 = ~n20547 & n20687 ;
  assign n20689 = n20547 & ~n20687 ;
  assign n20690 = n20688 | n20689 ;
  assign n20691 = x116 & n4572 ;
  assign n20692 = x115 & n4567 ;
  assign n20693 = x114 & ~n4566 ;
  assign n20694 = n4828 & n20693 ;
  assign n20695 = n20692 | n20694 ;
  assign n20696 = n20691 | n20695 ;
  assign n20697 = n4575 | n20696 ;
  assign n20698 = ( n8778 & n20696 ) | ( n8778 & n20697 ) | ( n20696 & n20697 ) ;
  assign n20699 = x38 & n20698 ;
  assign n20700 = x38 & ~n20699 ;
  assign n20701 = ( n20698 & ~n20699 ) | ( n20698 & n20700 ) | ( ~n20699 & n20700 ) ;
  assign n20702 = ( n20546 & n20690 ) | ( n20546 & ~n20701 ) | ( n20690 & ~n20701 ) ;
  assign n20703 = ( ~n20690 & n20701 ) | ( ~n20690 & n20702 ) | ( n20701 & n20702 ) ;
  assign n20704 = ( ~n20546 & n20702 ) | ( ~n20546 & n20703 ) | ( n20702 & n20703 ) ;
  assign n20705 = x119 & n3913 ;
  assign n20706 = x118 & n3908 ;
  assign n20707 = x117 & ~n3907 ;
  assign n20708 = n4152 & n20707 ;
  assign n20709 = n20706 | n20708 ;
  assign n20710 = n20705 | n20709 ;
  assign n20711 = n3916 | n20710 ;
  assign n20712 = ( n9789 & n20710 ) | ( n9789 & n20711 ) | ( n20710 & n20711 ) ;
  assign n20713 = x35 & n20712 ;
  assign n20714 = x35 & ~n20713 ;
  assign n20715 = ( n20712 & ~n20713 ) | ( n20712 & n20714 ) | ( ~n20713 & n20714 ) ;
  assign n20716 = ~n20704 & n20715 ;
  assign n20717 = n20704 & ~n20715 ;
  assign n20718 = n20716 | n20717 ;
  assign n20719 = n20545 & ~n20718 ;
  assign n20720 = ~n20545 & n20718 ;
  assign n20721 = n20719 | n20720 ;
  assign n20722 = x125 & n2775 ;
  assign n20723 = x124 & n2770 ;
  assign n20724 = x123 & ~n2769 ;
  assign n20725 = n2978 & n20724 ;
  assign n20726 = n20723 | n20725 ;
  assign n20727 = n20722 | n20726 ;
  assign n20728 = n2778 | n20727 ;
  assign n20729 = ( n12310 & n20727 ) | ( n12310 & n20728 ) | ( n20727 & n20728 ) ;
  assign n20730 = x29 & n20729 ;
  assign n20731 = x29 & ~n20730 ;
  assign n20732 = ( n20729 & ~n20730 ) | ( n20729 & n20731 ) | ( ~n20730 & n20731 ) ;
  assign n20733 = ~n20475 & n20517 ;
  assign n20734 = n20732 & ~n20733 ;
  assign n20735 = n20733 | n20734 ;
  assign n20736 = ( ~n20732 & n20734 ) | ( ~n20732 & n20735 ) | ( n20734 & n20735 ) ;
  assign n20737 = n20721 | n20736 ;
  assign n20738 = n20721 & n20736 ;
  assign n20739 = n20737 & ~n20738 ;
  assign n20740 = n20530 | n20739 ;
  assign n20741 = n20529 | n20740 ;
  assign n20742 = ( n20529 & n20530 ) | ( n20529 & n20739 ) | ( n20530 & n20739 ) ;
  assign n20743 = n20741 & ~n20742 ;
  assign n20744 = ( n20494 & n20505 ) | ( n20494 & n20506 ) | ( n20505 & n20506 ) ;
  assign n20745 = n20509 & n20510 ;
  assign n20746 = n20515 | n20745 ;
  assign n20747 = ( n20743 & n20744 ) | ( n20743 & ~n20746 ) | ( n20744 & ~n20746 ) ;
  assign n20748 = ( ~n20744 & n20746 ) | ( ~n20744 & n20747 ) | ( n20746 & n20747 ) ;
  assign n20749 = ( ~n20743 & n20747 ) | ( ~n20743 & n20748 ) | ( n20747 & n20748 ) ;
  assign n20750 = n20528 | n20742 ;
  assign n20751 = x126 & n2775 ;
  assign n20752 = x125 & n2770 ;
  assign n20753 = x124 & ~n2769 ;
  assign n20754 = n2978 & n20753 ;
  assign n20755 = n20752 | n20754 ;
  assign n20756 = n20751 | n20755 ;
  assign n20757 = n2778 | n20756 ;
  assign n20758 = ( n12687 & n20756 ) | ( n12687 & n20757 ) | ( n20756 & n20757 ) ;
  assign n20759 = x29 & n20758 ;
  assign n20760 = x29 & ~n20759 ;
  assign n20761 = ( n20758 & ~n20759 ) | ( n20758 & n20760 ) | ( ~n20759 & n20760 ) ;
  assign n20762 = n20544 | n20719 ;
  assign n20763 = n20761 | n20762 ;
  assign n20764 = n20761 & n20762 ;
  assign n20765 = n20763 & ~n20764 ;
  assign n20766 = x123 & n3314 ;
  assign n20767 = x122 & n3309 ;
  assign n20768 = x121 & ~n3308 ;
  assign n20769 = n3570 & n20768 ;
  assign n20770 = n20767 | n20769 ;
  assign n20771 = n20766 | n20770 ;
  assign n20772 = n3317 | n20771 ;
  assign n20773 = ( n11219 & n20771 ) | ( n11219 & n20772 ) | ( n20771 & n20772 ) ;
  assign n20774 = x32 & n20773 ;
  assign n20775 = x32 & ~n20774 ;
  assign n20776 = ( n20773 & ~n20774 ) | ( n20773 & n20775 ) | ( ~n20774 & n20775 ) ;
  assign n20777 = ( n20546 & n20715 ) | ( n20546 & n20718 ) | ( n20715 & n20718 ) ;
  assign n20778 = n20776 | n20777 ;
  assign n20779 = n20776 & n20777 ;
  assign n20780 = n20778 & ~n20779 ;
  assign n20781 = x120 & n3913 ;
  assign n20782 = x119 & n3908 ;
  assign n20783 = x118 & ~n3907 ;
  assign n20784 = n4152 & n20783 ;
  assign n20785 = n20782 | n20784 ;
  assign n20786 = n20781 | n20785 ;
  assign n20787 = n3916 | n20786 ;
  assign n20788 = ( n10460 & n20786 ) | ( n10460 & n20787 ) | ( n20786 & n20787 ) ;
  assign n20789 = x35 & n20788 ;
  assign n20790 = x35 & ~n20789 ;
  assign n20791 = ( n20788 & ~n20789 ) | ( n20788 & n20790 ) | ( ~n20789 & n20790 ) ;
  assign n20792 = x111 & n6068 ;
  assign n20793 = x110 & n6063 ;
  assign n20794 = x109 & ~n6062 ;
  assign n20795 = n6398 & n20794 ;
  assign n20796 = n20793 | n20795 ;
  assign n20797 = n20792 | n20796 ;
  assign n20798 = n6071 | n20797 ;
  assign n20799 = ( n7492 & n20797 ) | ( n7492 & n20798 ) | ( n20797 & n20798 ) ;
  assign n20800 = x44 & n20799 ;
  assign n20801 = x44 & ~n20800 ;
  assign n20802 = ( n20799 & ~n20800 ) | ( n20799 & n20801 ) | ( ~n20800 & n20801 ) ;
  assign n20803 = x105 & n7812 ;
  assign n20804 = x104 & n7807 ;
  assign n20805 = x103 & ~n7806 ;
  assign n20806 = n8136 & n20805 ;
  assign n20807 = n20804 | n20806 ;
  assign n20808 = n20803 | n20807 ;
  assign n20809 = n7815 | n20808 ;
  assign n20810 = ( n5788 & n20808 ) | ( n5788 & n20809 ) | ( n20808 & n20809 ) ;
  assign n20811 = x50 & n20810 ;
  assign n20812 = x50 & ~n20811 ;
  assign n20813 = ( n20810 & ~n20811 ) | ( n20810 & n20812 ) | ( ~n20811 & n20812 ) ;
  assign n20814 = n20630 | n20644 ;
  assign n20815 = x102 & n8834 ;
  assign n20816 = x101 & n8829 ;
  assign n20817 = x100 & ~n8828 ;
  assign n20818 = n9159 & n20817 ;
  assign n20819 = n20816 | n20818 ;
  assign n20820 = n20815 | n20819 ;
  assign n20821 = n8837 | n20820 ;
  assign n20822 = ( n5025 & n20820 ) | ( n5025 & n20821 ) | ( n20820 & n20821 ) ;
  assign n20823 = x53 & n20822 ;
  assign n20824 = x53 & ~n20823 ;
  assign n20825 = ( n20822 & ~n20823 ) | ( n20822 & n20824 ) | ( ~n20823 & n20824 ) ;
  assign n20826 = x90 & n12808 ;
  assign n20827 = x63 & x89 ;
  assign n20828 = ~n12808 & n20827 ;
  assign n20829 = n20826 | n20828 ;
  assign n20830 = n20587 & ~n20829 ;
  assign n20831 = ~n20587 & n20829 ;
  assign n20832 = n20830 | n20831 ;
  assign n20833 = x93 & n11984 ;
  assign n20834 = x92 & n11979 ;
  assign n20835 = x91 & ~n11978 ;
  assign n20836 = n12430 & n20835 ;
  assign n20837 = n20834 | n20836 ;
  assign n20838 = n20833 | n20837 ;
  assign n20839 = n11987 | n20838 ;
  assign n20840 = ( n2931 & n20838 ) | ( n2931 & n20839 ) | ( n20838 & n20839 ) ;
  assign n20841 = x62 & n20840 ;
  assign n20842 = x62 & ~n20841 ;
  assign n20843 = ( n20840 & ~n20841 ) | ( n20840 & n20842 ) | ( ~n20841 & n20842 ) ;
  assign n20844 = ~n20832 & n20843 ;
  assign n20845 = n20832 & ~n20843 ;
  assign n20846 = n20844 | n20845 ;
  assign n20847 = n20590 | n20603 ;
  assign n20848 = ~n20846 & n20847 ;
  assign n20849 = n20846 & ~n20847 ;
  assign n20850 = n20848 | n20849 ;
  assign n20851 = x96 & n10876 ;
  assign n20852 = x95 & n10871 ;
  assign n20853 = x94 & ~n10870 ;
  assign n20854 = n11305 & n20853 ;
  assign n20855 = n20852 | n20854 ;
  assign n20856 = n20851 | n20855 ;
  assign n20857 = n10879 | n20856 ;
  assign n20858 = ( n3509 & n20856 ) | ( n3509 & n20857 ) | ( n20856 & n20857 ) ;
  assign n20859 = x59 & n20858 ;
  assign n20860 = x59 & ~n20859 ;
  assign n20861 = ( n20858 & ~n20859 ) | ( n20858 & n20860 ) | ( ~n20859 & n20860 ) ;
  assign n20862 = ~n20850 & n20861 ;
  assign n20863 = n20850 & ~n20861 ;
  assign n20864 = n20862 | n20863 ;
  assign n20865 = n20608 & ~n20864 ;
  assign n20866 = ~n20608 & n20864 ;
  assign n20867 = n20865 | n20866 ;
  assign n20868 = x99 & n9853 ;
  assign n20869 = x98 & n9848 ;
  assign n20870 = x97 & ~n9847 ;
  assign n20871 = n10165 & n20870 ;
  assign n20872 = n20869 | n20871 ;
  assign n20873 = n20868 | n20872 ;
  assign n20874 = n9856 | n20873 ;
  assign n20875 = ( n4325 & n20873 ) | ( n4325 & n20874 ) | ( n20873 & n20874 ) ;
  assign n20876 = x56 & n20875 ;
  assign n20877 = x56 & ~n20876 ;
  assign n20878 = ( n20875 & ~n20876 ) | ( n20875 & n20877 ) | ( ~n20876 & n20877 ) ;
  assign n20879 = ~n20867 & n20878 ;
  assign n20880 = n20867 & ~n20878 ;
  assign n20881 = n20879 | n20880 ;
  assign n20882 = ( n20625 & n20825 ) | ( n20625 & ~n20881 ) | ( n20825 & ~n20881 ) ;
  assign n20883 = ( ~n20625 & n20881 ) | ( ~n20625 & n20882 ) | ( n20881 & n20882 ) ;
  assign n20884 = ( ~n20825 & n20882 ) | ( ~n20825 & n20883 ) | ( n20882 & n20883 ) ;
  assign n20885 = ( n20813 & ~n20814 ) | ( n20813 & n20884 ) | ( ~n20814 & n20884 ) ;
  assign n20886 = ( n20813 & n20814 ) | ( n20813 & ~n20884 ) | ( n20814 & ~n20884 ) ;
  assign n20887 = ( ~n20813 & n20885 ) | ( ~n20813 & n20886 ) | ( n20885 & n20886 ) ;
  assign n20888 = n20646 & ~n20887 ;
  assign n20889 = ~n20646 & n20887 ;
  assign n20890 = n20888 | n20889 ;
  assign n20891 = x108 & n6937 ;
  assign n20892 = x107 & n6932 ;
  assign n20893 = x106 & ~n6931 ;
  assign n20894 = n7216 & n20893 ;
  assign n20895 = n20892 | n20894 ;
  assign n20896 = n20891 | n20895 ;
  assign n20897 = n6940 | n20896 ;
  assign n20898 = ( n6358 & n20896 ) | ( n6358 & n20897 ) | ( n20896 & n20897 ) ;
  assign n20899 = x47 & n20898 ;
  assign n20900 = x47 & ~n20899 ;
  assign n20901 = ( n20898 & ~n20899 ) | ( n20898 & n20900 ) | ( ~n20899 & n20900 ) ;
  assign n20902 = ~n20890 & n20901 ;
  assign n20903 = n20890 & ~n20901 ;
  assign n20904 = n20902 | n20903 ;
  assign n20905 = ( ~n20649 & n20802 ) | ( ~n20649 & n20904 ) | ( n20802 & n20904 ) ;
  assign n20906 = ( n20649 & ~n20904 ) | ( n20649 & n20905 ) | ( ~n20904 & n20905 ) ;
  assign n20907 = ( ~n20802 & n20905 ) | ( ~n20802 & n20906 ) | ( n20905 & n20906 ) ;
  assign n20908 = ~n20669 & n20907 ;
  assign n20909 = n20669 & ~n20907 ;
  assign n20910 = n20908 | n20909 ;
  assign n20911 = x114 & n5340 ;
  assign n20912 = x113 & n5335 ;
  assign n20913 = x112 & ~n5334 ;
  assign n20914 = n5580 & n20913 ;
  assign n20915 = n20912 | n20914 ;
  assign n20916 = n20911 | n20915 ;
  assign n20917 = n5343 | n20916 ;
  assign n20918 = ( n8437 & n20916 ) | ( n8437 & n20917 ) | ( n20916 & n20917 ) ;
  assign n20919 = x41 & n20918 ;
  assign n20920 = x41 & ~n20919 ;
  assign n20921 = ( n20918 & ~n20919 ) | ( n20918 & n20920 ) | ( ~n20919 & n20920 ) ;
  assign n20922 = n20910 & ~n20921 ;
  assign n20923 = ~n20910 & n20921 ;
  assign n20924 = n20922 | n20923 ;
  assign n20925 = ( n20668 & n20684 ) | ( n20668 & n20687 ) | ( n20684 & n20687 ) ;
  assign n20926 = n20924 & n20925 ;
  assign n20927 = ~n20924 & n20925 ;
  assign n20928 = n20924 | n20927 ;
  assign n20929 = x117 & n4572 ;
  assign n20930 = x116 & n4567 ;
  assign n20931 = x115 & ~n4566 ;
  assign n20932 = n4828 & n20931 ;
  assign n20933 = n20930 | n20932 ;
  assign n20934 = n20929 | n20933 ;
  assign n20935 = n4575 | n20934 ;
  assign n20936 = ( n9118 & n20934 ) | ( n9118 & n20935 ) | ( n20934 & n20935 ) ;
  assign n20937 = x38 & n20936 ;
  assign n20938 = x38 & ~n20937 ;
  assign n20939 = ( n20936 & ~n20937 ) | ( n20936 & n20938 ) | ( ~n20937 & n20938 ) ;
  assign n20940 = n20928 & ~n20939 ;
  assign n20941 = ~n20926 & n20940 ;
  assign n20942 = ( n20926 & ~n20928 ) | ( n20926 & n20939 ) | ( ~n20928 & n20939 ) ;
  assign n20943 = n20941 | n20942 ;
  assign n20944 = ( n20547 & ~n20687 ) | ( n20547 & n20701 ) | ( ~n20687 & n20701 ) ;
  assign n20945 = ( n20791 & n20943 ) | ( n20791 & ~n20944 ) | ( n20943 & ~n20944 ) ;
  assign n20946 = ( ~n20943 & n20944 ) | ( ~n20943 & n20945 ) | ( n20944 & n20945 ) ;
  assign n20947 = ( ~n20791 & n20945 ) | ( ~n20791 & n20946 ) | ( n20945 & n20946 ) ;
  assign n20948 = n20780 | n20947 ;
  assign n20949 = ( n20776 & n20777 ) | ( n20776 & ~n20947 ) | ( n20777 & ~n20947 ) ;
  assign n20950 = n20778 & ~n20949 ;
  assign n20951 = n20948 & ~n20950 ;
  assign n20952 = ~n20765 & n20951 ;
  assign n20953 = n20765 & ~n20951 ;
  assign n20954 = n20952 | n20953 ;
  assign n20955 = x127 & ~n2274 ;
  assign n20956 = n2481 & n20955 ;
  assign n20957 = ( x127 & n2283 ) | ( x127 & n20956 ) | ( n2283 & n20956 ) ;
  assign n20958 = ( x126 & n20956 ) | ( x126 & n20957 ) | ( n20956 & n20957 ) ;
  assign n20959 = ( n12685 & n20957 ) | ( n12685 & n20958 ) | ( n20957 & n20958 ) ;
  assign n20960 = x26 & n20959 ;
  assign n20961 = x26 & ~n20960 ;
  assign n20962 = ( n20959 & ~n20960 ) | ( n20959 & n20961 ) | ( ~n20960 & n20961 ) ;
  assign n20963 = n20734 & n20962 ;
  assign n20964 = n20962 & ~n20963 ;
  assign n20965 = n20737 & n20964 ;
  assign n20966 = n20954 & ~n20965 ;
  assign n20967 = ( ~n20737 & n20962 ) | ( ~n20737 & n20963 ) | ( n20962 & n20963 ) ;
  assign n20968 = ( ~n20734 & n20737 ) | ( ~n20734 & n20967 ) | ( n20737 & n20967 ) ;
  assign n20969 = n20966 & n20968 ;
  assign n20970 = ( n20954 & ~n20965 ) | ( n20954 & n20968 ) | ( ~n20965 & n20968 ) ;
  assign n20971 = ~n20969 & n20970 ;
  assign n20972 = n20750 & n20971 ;
  assign n20973 = n20750 | n20971 ;
  assign n20974 = ~n20972 & n20973 ;
  assign n20975 = ( n20743 & n20744 ) | ( n20743 & n20745 ) | ( n20744 & n20745 ) ;
  assign n20976 = ( n20741 & ~n20742 ) | ( n20741 & n20744 ) | ( ~n20742 & n20744 ) ;
  assign n20977 = ( n20741 & n20744 ) | ( n20741 & n20976 ) | ( n20744 & n20976 ) ;
  assign n20978 = ( n20515 & n20975 ) | ( n20515 & n20977 ) | ( n20975 & n20977 ) ;
  assign n20979 = n20974 | n20978 ;
  assign n20980 = n20974 & n20975 ;
  assign n20981 = n20974 & n20977 ;
  assign n20982 = ( n20515 & n20980 ) | ( n20515 & n20981 ) | ( n20980 & n20981 ) ;
  assign n20983 = n20979 & ~n20982 ;
  assign n20984 = x127 & n2775 ;
  assign n20985 = x126 & n2770 ;
  assign n20986 = x125 & ~n2769 ;
  assign n20987 = n2978 & n20986 ;
  assign n20988 = n20985 | n20987 ;
  assign n20989 = n20984 | n20988 ;
  assign n20990 = n2778 | n20989 ;
  assign n20991 = ( n12720 & n20989 ) | ( n12720 & n20990 ) | ( n20989 & n20990 ) ;
  assign n20992 = x29 & n20991 ;
  assign n20993 = x29 & ~n20992 ;
  assign n20994 = ( n20991 & ~n20992 ) | ( n20991 & n20993 ) | ( ~n20992 & n20993 ) ;
  assign n20995 = n20764 & n20994 ;
  assign n20996 = n20994 & ~n20995 ;
  assign n20997 = ~n20953 & n20996 ;
  assign n20998 = x124 & n3314 ;
  assign n20999 = x123 & n3309 ;
  assign n21000 = x122 & ~n3308 ;
  assign n21001 = n3570 & n21000 ;
  assign n21002 = n20999 | n21001 ;
  assign n21003 = n20998 | n21002 ;
  assign n21004 = n3317 | n21003 ;
  assign n21005 = ( n11916 & n21003 ) | ( n11916 & n21004 ) | ( n21003 & n21004 ) ;
  assign n21006 = x32 & n21005 ;
  assign n21007 = x32 & ~n21006 ;
  assign n21008 = ( n21005 & ~n21006 ) | ( n21005 & n21007 ) | ( ~n21006 & n21007 ) ;
  assign n21009 = n20927 | n20942 ;
  assign n21010 = n20909 | n20923 ;
  assign n21011 = x112 & n6068 ;
  assign n21012 = x111 & n6063 ;
  assign n21013 = x110 & ~n6062 ;
  assign n21014 = n6398 & n21013 ;
  assign n21015 = n21012 | n21014 ;
  assign n21016 = n21011 | n21015 ;
  assign n21017 = n6071 | n21016 ;
  assign n21018 = ( n7789 & n21016 ) | ( n7789 & n21017 ) | ( n21016 & n21017 ) ;
  assign n21019 = x44 & n21018 ;
  assign n21020 = x44 & ~n21019 ;
  assign n21021 = ( n21018 & ~n21019 ) | ( n21018 & n21020 ) | ( ~n21019 & n21020 ) ;
  assign n21022 = x109 & n6937 ;
  assign n21023 = x108 & n6932 ;
  assign n21024 = x107 & ~n6931 ;
  assign n21025 = n7216 & n21024 ;
  assign n21026 = n21023 | n21025 ;
  assign n21027 = n21022 | n21026 ;
  assign n21028 = n6940 | n21027 ;
  assign n21029 = ( n6884 & n21027 ) | ( n6884 & n21028 ) | ( n21027 & n21028 ) ;
  assign n21030 = x47 & n21029 ;
  assign n21031 = x47 & ~n21030 ;
  assign n21032 = ( n21029 & ~n21030 ) | ( n21029 & n21031 ) | ( ~n21030 & n21031 ) ;
  assign n21033 = x106 & n7812 ;
  assign n21034 = x105 & n7807 ;
  assign n21035 = x104 & ~n7806 ;
  assign n21036 = n8136 & n21035 ;
  assign n21037 = n21034 | n21036 ;
  assign n21038 = n21033 | n21037 ;
  assign n21039 = n7815 | n21038 ;
  assign n21040 = ( n5814 & n21038 ) | ( n5814 & n21039 ) | ( n21038 & n21039 ) ;
  assign n21041 = x50 & n21040 ;
  assign n21042 = x50 & ~n21041 ;
  assign n21043 = ( n21040 & ~n21041 ) | ( n21040 & n21042 ) | ( ~n21041 & n21042 ) ;
  assign n21044 = x97 & n10876 ;
  assign n21045 = x96 & n10871 ;
  assign n21046 = x95 & ~n10870 ;
  assign n21047 = n11305 & n21046 ;
  assign n21048 = n21045 | n21047 ;
  assign n21049 = n21044 | n21048 ;
  assign n21050 = n10879 | n21049 ;
  assign n21051 = ( n3707 & n21049 ) | ( n3707 & n21050 ) | ( n21049 & n21050 ) ;
  assign n21052 = x59 & n21051 ;
  assign n21053 = x59 & ~n21052 ;
  assign n21054 = ( n21051 & ~n21052 ) | ( n21051 & n21053 ) | ( ~n21052 & n21053 ) ;
  assign n21055 = n20848 | n20862 ;
  assign n21056 = n21054 | n21055 ;
  assign n21057 = n21054 & n21055 ;
  assign n21058 = n21056 & ~n21057 ;
  assign n21059 = x94 & n11984 ;
  assign n21060 = x93 & n11979 ;
  assign n21061 = x92 & ~n11978 ;
  assign n21062 = n12430 & n21061 ;
  assign n21063 = n21060 | n21062 ;
  assign n21064 = n21059 | n21063 ;
  assign n21065 = n11987 | n21064 ;
  assign n21066 = ( n3271 & n21064 ) | ( n3271 & n21065 ) | ( n21064 & n21065 ) ;
  assign n21067 = x62 & n21066 ;
  assign n21068 = x62 & ~n21067 ;
  assign n21069 = ( n21066 & ~n21067 ) | ( n21066 & n21068 ) | ( ~n21067 & n21068 ) ;
  assign n21070 = x91 & n12808 ;
  assign n21071 = x63 & x90 ;
  assign n21072 = ~n12808 & n21071 ;
  assign n21073 = n21070 | n21072 ;
  assign n21074 = ~x26 & n21073 ;
  assign n21075 = x26 & ~n21073 ;
  assign n21076 = n21074 | n21075 ;
  assign n21077 = n20829 & ~n21076 ;
  assign n21078 = ~n20829 & n21076 ;
  assign n21079 = n21077 | n21078 ;
  assign n21080 = ( n20830 & n20844 ) | ( n20830 & ~n21079 ) | ( n20844 & ~n21079 ) ;
  assign n21081 = ( n20830 & ~n20831 ) | ( n20830 & n20843 ) | ( ~n20831 & n20843 ) ;
  assign n21082 = n21079 & ~n21081 ;
  assign n21083 = n21080 | n21082 ;
  assign n21084 = n21069 & ~n21083 ;
  assign n21085 = n21083 | n21084 ;
  assign n21086 = ( ~n21069 & n21084 ) | ( ~n21069 & n21085 ) | ( n21084 & n21085 ) ;
  assign n21087 = ~n21058 & n21086 ;
  assign n21088 = n21058 & ~n21086 ;
  assign n21089 = n21087 | n21088 ;
  assign n21090 = x100 & n9853 ;
  assign n21091 = x99 & n9848 ;
  assign n21092 = x98 & ~n9847 ;
  assign n21093 = n10165 & n21092 ;
  assign n21094 = n21091 | n21093 ;
  assign n21095 = n21090 | n21094 ;
  assign n21096 = n9856 | n21095 ;
  assign n21097 = ( n4532 & n21095 ) | ( n4532 & n21096 ) | ( n21095 & n21096 ) ;
  assign n21098 = x56 & n21097 ;
  assign n21099 = x56 & ~n21098 ;
  assign n21100 = ( n21097 & ~n21098 ) | ( n21097 & n21099 ) | ( ~n21098 & n21099 ) ;
  assign n21101 = ~n21089 & n21100 ;
  assign n21102 = n21089 | n21101 ;
  assign n21103 = n21089 & n21100 ;
  assign n21104 = n20865 | n20879 ;
  assign n21105 = n21103 | n21104 ;
  assign n21106 = n21102 & ~n21105 ;
  assign n21107 = ( ~n21102 & n21103 ) | ( ~n21102 & n21104 ) | ( n21103 & n21104 ) ;
  assign n21108 = n21106 | n21107 ;
  assign n21109 = x103 & n8834 ;
  assign n21110 = x102 & n8829 ;
  assign n21111 = x101 & ~n8828 ;
  assign n21112 = n9159 & n21111 ;
  assign n21113 = n21110 | n21112 ;
  assign n21114 = n21109 | n21113 ;
  assign n21115 = n8837 | n21114 ;
  assign n21116 = ( n5264 & n21114 ) | ( n5264 & n21115 ) | ( n21114 & n21115 ) ;
  assign n21117 = x53 & n21116 ;
  assign n21118 = x53 & ~n21117 ;
  assign n21119 = ( n21116 & ~n21117 ) | ( n21116 & n21118 ) | ( ~n21117 & n21118 ) ;
  assign n21120 = ~n21108 & n21119 ;
  assign n21121 = n21108 | n21120 ;
  assign n21122 = n21108 & n21119 ;
  assign n21123 = n20882 | n21122 ;
  assign n21124 = n21121 & ~n21123 ;
  assign n21125 = ( n20882 & ~n21121 ) | ( n20882 & n21122 ) | ( ~n21121 & n21122 ) ;
  assign n21126 = n21124 | n21125 ;
  assign n21127 = ( n20886 & n21043 ) | ( n20886 & ~n21126 ) | ( n21043 & ~n21126 ) ;
  assign n21128 = ( ~n20886 & n21126 ) | ( ~n20886 & n21127 ) | ( n21126 & n21127 ) ;
  assign n21129 = ( ~n21043 & n21127 ) | ( ~n21043 & n21128 ) | ( n21127 & n21128 ) ;
  assign n21130 = n21032 & ~n21129 ;
  assign n21131 = ~n21032 & n21129 ;
  assign n21132 = n21130 | n21131 ;
  assign n21133 = n20888 | n20902 ;
  assign n21134 = n21132 & ~n21133 ;
  assign n21135 = ~n21132 & n21133 ;
  assign n21136 = n21134 | n21135 ;
  assign n21137 = n21021 & ~n21136 ;
  assign n21138 = n21136 | n21137 ;
  assign n21139 = ( ~n21021 & n21137 ) | ( ~n21021 & n21138 ) | ( n21137 & n21138 ) ;
  assign n21140 = ~n20906 & n21139 ;
  assign n21141 = n20906 & ~n21139 ;
  assign n21142 = n21140 | n21141 ;
  assign n21143 = x115 & n5340 ;
  assign n21144 = x114 & n5335 ;
  assign n21145 = x113 & ~n5334 ;
  assign n21146 = n5580 & n21145 ;
  assign n21147 = n21144 | n21146 ;
  assign n21148 = n21143 | n21147 ;
  assign n21149 = n5343 | n21148 ;
  assign n21150 = ( n8749 & n21148 ) | ( n8749 & n21149 ) | ( n21148 & n21149 ) ;
  assign n21151 = x41 & n21150 ;
  assign n21152 = x41 & ~n21151 ;
  assign n21153 = ( n21150 & ~n21151 ) | ( n21150 & n21152 ) | ( ~n21151 & n21152 ) ;
  assign n21154 = ~n21142 & n21153 ;
  assign n21155 = n21142 & ~n21153 ;
  assign n21156 = n21154 | n21155 ;
  assign n21157 = n21010 & ~n21156 ;
  assign n21158 = n21010 & ~n21157 ;
  assign n21159 = n21156 | n21157 ;
  assign n21160 = ~n21158 & n21159 ;
  assign n21161 = x118 & n4572 ;
  assign n21162 = x117 & n4567 ;
  assign n21163 = x116 & ~n4566 ;
  assign n21164 = n4828 & n21163 ;
  assign n21165 = n21162 | n21164 ;
  assign n21166 = n21161 | n21165 ;
  assign n21167 = n4575 | n21166 ;
  assign n21168 = ( n9760 & n21166 ) | ( n9760 & n21167 ) | ( n21166 & n21167 ) ;
  assign n21169 = x38 & n21168 ;
  assign n21170 = x38 & ~n21169 ;
  assign n21171 = ( n21168 & ~n21169 ) | ( n21168 & n21170 ) | ( ~n21169 & n21170 ) ;
  assign n21172 = n21160 & ~n21171 ;
  assign n21173 = ~n21160 & n21171 ;
  assign n21174 = n21172 | n21173 ;
  assign n21175 = n21009 & ~n21174 ;
  assign n21176 = ~n21009 & n21174 ;
  assign n21177 = n21175 | n21176 ;
  assign n21178 = x121 & n3913 ;
  assign n21179 = x120 & n3908 ;
  assign n21180 = x119 & ~n3907 ;
  assign n21181 = n4152 & n21180 ;
  assign n21182 = n21179 | n21181 ;
  assign n21183 = n21178 | n21182 ;
  assign n21184 = n3916 | n21183 ;
  assign n21185 = ( n10811 & n21183 ) | ( n10811 & n21184 ) | ( n21183 & n21184 ) ;
  assign n21186 = x35 & n21185 ;
  assign n21187 = x35 & ~n21186 ;
  assign n21188 = ( n21185 & ~n21186 ) | ( n21185 & n21187 ) | ( ~n21186 & n21187 ) ;
  assign n21189 = ~n21177 & n21188 ;
  assign n21190 = n21177 | n21189 ;
  assign n21191 = n21177 & n21188 ;
  assign n21192 = n20946 | n21191 ;
  assign n21193 = n21190 & ~n21192 ;
  assign n21194 = ( n20946 & ~n21190 ) | ( n20946 & n21191 ) | ( ~n21190 & n21191 ) ;
  assign n21195 = n21193 | n21194 ;
  assign n21196 = ( n20949 & n21008 ) | ( n20949 & ~n21195 ) | ( n21008 & ~n21195 ) ;
  assign n21197 = ( ~n20949 & n21195 ) | ( ~n20949 & n21196 ) | ( n21195 & n21196 ) ;
  assign n21198 = ( ~n21008 & n21196 ) | ( ~n21008 & n21197 ) | ( n21196 & n21197 ) ;
  assign n21199 = ~n20997 & n21198 ;
  assign n21200 = ( n20764 & n20953 ) | ( n20764 & ~n20994 ) | ( n20953 & ~n20994 ) ;
  assign n21201 = n21199 & ~n21200 ;
  assign n21202 = ( n20997 & ~n21198 ) | ( n20997 & n21200 ) | ( ~n21198 & n21200 ) ;
  assign n21203 = n21201 | n21202 ;
  assign n21204 = n20967 & ~n21203 ;
  assign n21205 = ( n20970 & n21203 ) | ( n20970 & ~n21204 ) | ( n21203 & ~n21204 ) ;
  assign n21206 = ~n20967 & n21203 ;
  assign n21207 = n20970 & n21206 ;
  assign n21208 = n21205 & ~n21207 ;
  assign n21209 = n20972 | n20980 ;
  assign n21210 = n20972 | n20981 ;
  assign n21211 = ( n20515 & n21209 ) | ( n20515 & n21210 ) | ( n21209 & n21210 ) ;
  assign n21212 = n21208 | n21211 ;
  assign n21213 = n21208 & n21209 ;
  assign n21214 = n21208 & n21210 ;
  assign n21215 = ( n20515 & n21213 ) | ( n20515 & n21214 ) | ( n21213 & n21214 ) ;
  assign n21216 = n21212 & ~n21215 ;
  assign n21217 = ( n20953 & n20994 ) | ( n20953 & n20995 ) | ( n20994 & n20995 ) ;
  assign n21218 = n21202 | n21217 ;
  assign n21219 = x127 & n2770 ;
  assign n21220 = x126 & ~n2769 ;
  assign n21221 = n2978 & n21220 ;
  assign n21222 = n21219 | n21221 ;
  assign n21223 = n2778 | n21222 ;
  assign n21224 = ( n13461 & n21222 ) | ( n13461 & n21223 ) | ( n21222 & n21223 ) ;
  assign n21225 = x29 & n21224 ;
  assign n21226 = x29 & ~n21225 ;
  assign n21227 = ( n21224 & ~n21225 ) | ( n21224 & n21226 ) | ( ~n21225 & n21226 ) ;
  assign n21228 = x125 & n3314 ;
  assign n21229 = x124 & n3309 ;
  assign n21230 = x123 & ~n3308 ;
  assign n21231 = n3570 & n21230 ;
  assign n21232 = n21229 | n21231 ;
  assign n21233 = n21228 | n21232 ;
  assign n21234 = n3317 | n21233 ;
  assign n21235 = ( n12310 & n21233 ) | ( n12310 & n21234 ) | ( n21233 & n21234 ) ;
  assign n21236 = x32 & n21235 ;
  assign n21237 = x32 & ~n21236 ;
  assign n21238 = ( n21235 & ~n21236 ) | ( n21235 & n21237 ) | ( ~n21236 & n21237 ) ;
  assign n21239 = n21189 | n21238 ;
  assign n21240 = n21194 | n21239 ;
  assign n21241 = ( n21189 & n21194 ) | ( n21189 & n21238 ) | ( n21194 & n21238 ) ;
  assign n21242 = n21240 & ~n21241 ;
  assign n21243 = x122 & n3913 ;
  assign n21244 = x121 & n3908 ;
  assign n21245 = x120 & ~n3907 ;
  assign n21246 = n4152 & n21245 ;
  assign n21247 = n21244 | n21246 ;
  assign n21248 = n21243 | n21247 ;
  assign n21249 = n3916 | n21248 ;
  assign n21250 = ( n11188 & n21248 ) | ( n11188 & n21249 ) | ( n21248 & n21249 ) ;
  assign n21251 = x35 & n21250 ;
  assign n21252 = x35 & ~n21251 ;
  assign n21253 = ( n21250 & ~n21251 ) | ( n21250 & n21252 ) | ( ~n21251 & n21252 ) ;
  assign n21254 = n21173 | n21175 ;
  assign n21255 = x119 & n4572 ;
  assign n21256 = x118 & n4567 ;
  assign n21257 = x117 & ~n4566 ;
  assign n21258 = n4828 & n21257 ;
  assign n21259 = n21256 | n21258 ;
  assign n21260 = n21255 | n21259 ;
  assign n21261 = n4575 | n21260 ;
  assign n21262 = ( n9789 & n21260 ) | ( n9789 & n21261 ) | ( n21260 & n21261 ) ;
  assign n21263 = x38 & n21262 ;
  assign n21264 = x38 & ~n21263 ;
  assign n21265 = ( n21262 & ~n21263 ) | ( n21262 & n21264 ) | ( ~n21263 & n21264 ) ;
  assign n21266 = n21154 | n21157 ;
  assign n21267 = n21137 | n21141 ;
  assign n21268 = x113 & n6068 ;
  assign n21269 = x112 & n6063 ;
  assign n21270 = x111 & ~n6062 ;
  assign n21271 = n6398 & n21270 ;
  assign n21272 = n21269 | n21271 ;
  assign n21273 = n21268 | n21272 ;
  assign n21274 = n6071 | n21273 ;
  assign n21275 = ( n8113 & n21273 ) | ( n8113 & n21274 ) | ( n21273 & n21274 ) ;
  assign n21276 = x44 & n21275 ;
  assign n21277 = x44 & ~n21276 ;
  assign n21278 = ( n21275 & ~n21276 ) | ( n21275 & n21277 ) | ( ~n21276 & n21277 ) ;
  assign n21279 = n21130 | n21135 ;
  assign n21280 = x107 & n7812 ;
  assign n21281 = x106 & n7807 ;
  assign n21282 = x105 & ~n7806 ;
  assign n21283 = n8136 & n21282 ;
  assign n21284 = n21281 | n21283 ;
  assign n21285 = n21280 | n21284 ;
  assign n21286 = n7815 | n21285 ;
  assign n21287 = ( n6328 & n21285 ) | ( n6328 & n21286 ) | ( n21285 & n21286 ) ;
  assign n21288 = x50 & n21287 ;
  assign n21289 = x50 & ~n21288 ;
  assign n21290 = ( n21287 & ~n21288 ) | ( n21287 & n21289 ) | ( ~n21288 & n21289 ) ;
  assign n21291 = n21120 | n21125 ;
  assign n21292 = x101 & n9853 ;
  assign n21293 = x100 & n9848 ;
  assign n21294 = x99 & ~n9847 ;
  assign n21295 = n10165 & n21294 ;
  assign n21296 = n21293 | n21295 ;
  assign n21297 = n21292 | n21296 ;
  assign n21298 = n9856 | n21297 ;
  assign n21299 = ( n4783 & n21297 ) | ( n4783 & n21298 ) | ( n21297 & n21298 ) ;
  assign n21300 = x56 & n21299 ;
  assign n21301 = x56 & ~n21300 ;
  assign n21302 = ( n21299 & ~n21300 ) | ( n21299 & n21301 ) | ( ~n21300 & n21301 ) ;
  assign n21303 = n21057 | n21088 ;
  assign n21304 = x98 & n10876 ;
  assign n21305 = x97 & n10871 ;
  assign n21306 = x96 & ~n10870 ;
  assign n21307 = n11305 & n21306 ;
  assign n21308 = n21305 | n21307 ;
  assign n21309 = n21304 | n21308 ;
  assign n21310 = n10879 | n21309 ;
  assign n21311 = ( n4105 & n21309 ) | ( n4105 & n21310 ) | ( n21309 & n21310 ) ;
  assign n21312 = x59 & n21311 ;
  assign n21313 = x59 & ~n21312 ;
  assign n21314 = ( n21311 & ~n21312 ) | ( n21311 & n21313 ) | ( ~n21312 & n21313 ) ;
  assign n21315 = x95 & n11984 ;
  assign n21316 = x94 & n11979 ;
  assign n21317 = x93 & ~n11978 ;
  assign n21318 = n12430 & n21317 ;
  assign n21319 = n21316 | n21318 ;
  assign n21320 = n21315 | n21319 ;
  assign n21321 = n11987 | n21320 ;
  assign n21322 = ( n3479 & n21320 ) | ( n3479 & n21321 ) | ( n21320 & n21321 ) ;
  assign n21323 = ~x62 & n21322 ;
  assign n21324 = x92 & n12808 ;
  assign n21325 = x63 & x91 ;
  assign n21326 = ~n12808 & n21325 ;
  assign n21327 = n21324 | n21326 ;
  assign n21328 = n21074 | n21077 ;
  assign n21329 = n21327 & ~n21328 ;
  assign n21330 = ~n21327 & n21328 ;
  assign n21331 = n21329 | n21330 ;
  assign n21332 = x62 & ~n21322 ;
  assign n21333 = n21331 & ~n21332 ;
  assign n21334 = ~n21323 & n21333 ;
  assign n21335 = ( n21323 & ~n21331 ) | ( n21323 & n21332 ) | ( ~n21331 & n21332 ) ;
  assign n21336 = n21334 | n21335 ;
  assign n21337 = n21080 | n21084 ;
  assign n21338 = ( n21314 & n21336 ) | ( n21314 & ~n21337 ) | ( n21336 & ~n21337 ) ;
  assign n21339 = ( ~n21336 & n21337 ) | ( ~n21336 & n21338 ) | ( n21337 & n21338 ) ;
  assign n21340 = ( ~n21314 & n21338 ) | ( ~n21314 & n21339 ) | ( n21338 & n21339 ) ;
  assign n21341 = ( n21302 & ~n21303 ) | ( n21302 & n21340 ) | ( ~n21303 & n21340 ) ;
  assign n21342 = ( n21303 & ~n21340 ) | ( n21303 & n21341 ) | ( ~n21340 & n21341 ) ;
  assign n21343 = ( ~n21302 & n21341 ) | ( ~n21302 & n21342 ) | ( n21341 & n21342 ) ;
  assign n21344 = n21101 | n21107 ;
  assign n21345 = x104 & n8834 ;
  assign n21346 = x103 & n8829 ;
  assign n21347 = x102 & ~n8828 ;
  assign n21348 = n9159 & n21347 ;
  assign n21349 = n21346 | n21348 ;
  assign n21350 = n21345 | n21349 ;
  assign n21351 = n8837 | n21350 ;
  assign n21352 = ( n5295 & n21350 ) | ( n5295 & n21351 ) | ( n21350 & n21351 ) ;
  assign n21353 = x53 & n21352 ;
  assign n21354 = x53 & ~n21353 ;
  assign n21355 = ( n21352 & ~n21353 ) | ( n21352 & n21354 ) | ( ~n21353 & n21354 ) ;
  assign n21356 = ( n21343 & ~n21344 ) | ( n21343 & n21355 ) | ( ~n21344 & n21355 ) ;
  assign n21357 = ( n21344 & ~n21355 ) | ( n21344 & n21356 ) | ( ~n21355 & n21356 ) ;
  assign n21358 = ( ~n21343 & n21356 ) | ( ~n21343 & n21357 ) | ( n21356 & n21357 ) ;
  assign n21359 = ( n21290 & n21291 ) | ( n21290 & ~n21358 ) | ( n21291 & ~n21358 ) ;
  assign n21360 = ( ~n21291 & n21358 ) | ( ~n21291 & n21359 ) | ( n21358 & n21359 ) ;
  assign n21361 = ( ~n21290 & n21359 ) | ( ~n21290 & n21360 ) | ( n21359 & n21360 ) ;
  assign n21362 = ~n21127 & n21361 ;
  assign n21363 = n21127 & ~n21361 ;
  assign n21364 = n21362 | n21363 ;
  assign n21365 = x110 & n6937 ;
  assign n21366 = x109 & n6932 ;
  assign n21367 = x108 & ~n6931 ;
  assign n21368 = n7216 & n21367 ;
  assign n21369 = n21366 | n21368 ;
  assign n21370 = n21365 | n21369 ;
  assign n21371 = n6940 | n21370 ;
  assign n21372 = ( n7189 & n21370 ) | ( n7189 & n21371 ) | ( n21370 & n21371 ) ;
  assign n21373 = x47 & n21372 ;
  assign n21374 = x47 & ~n21373 ;
  assign n21375 = ( n21372 & ~n21373 ) | ( n21372 & n21374 ) | ( ~n21373 & n21374 ) ;
  assign n21376 = n21364 & n21375 ;
  assign n21377 = ( n21127 & ~n21361 ) | ( n21127 & n21375 ) | ( ~n21361 & n21375 ) ;
  assign n21378 = n21362 | n21377 ;
  assign n21379 = ~n21376 & n21378 ;
  assign n21380 = ( n21278 & ~n21279 ) | ( n21278 & n21379 ) | ( ~n21279 & n21379 ) ;
  assign n21381 = ( n21279 & ~n21379 ) | ( n21279 & n21380 ) | ( ~n21379 & n21380 ) ;
  assign n21382 = ( ~n21278 & n21380 ) | ( ~n21278 & n21381 ) | ( n21380 & n21381 ) ;
  assign n21383 = ~n21267 & n21382 ;
  assign n21384 = n21267 & ~n21382 ;
  assign n21385 = n21383 | n21384 ;
  assign n21386 = x116 & n5340 ;
  assign n21387 = x115 & n5335 ;
  assign n21388 = x114 & ~n5334 ;
  assign n21389 = n5580 & n21388 ;
  assign n21390 = n21387 | n21389 ;
  assign n21391 = n21386 | n21390 ;
  assign n21392 = n5343 | n21391 ;
  assign n21393 = ( n8778 & n21391 ) | ( n8778 & n21392 ) | ( n21391 & n21392 ) ;
  assign n21394 = x41 & n21393 ;
  assign n21395 = x41 & ~n21394 ;
  assign n21396 = ( n21393 & ~n21394 ) | ( n21393 & n21395 ) | ( ~n21394 & n21395 ) ;
  assign n21397 = n21385 & n21396 ;
  assign n21398 = ( n21267 & ~n21382 ) | ( n21267 & n21396 ) | ( ~n21382 & n21396 ) ;
  assign n21399 = n21383 | n21398 ;
  assign n21400 = ~n21397 & n21399 ;
  assign n21401 = ( n21265 & n21266 ) | ( n21265 & ~n21400 ) | ( n21266 & ~n21400 ) ;
  assign n21402 = ( ~n21266 & n21400 ) | ( ~n21266 & n21401 ) | ( n21400 & n21401 ) ;
  assign n21403 = ( ~n21265 & n21401 ) | ( ~n21265 & n21402 ) | ( n21401 & n21402 ) ;
  assign n21404 = ( n21253 & n21254 ) | ( n21253 & ~n21403 ) | ( n21254 & ~n21403 ) ;
  assign n21405 = ( ~n21254 & n21403 ) | ( ~n21254 & n21404 ) | ( n21403 & n21404 ) ;
  assign n21406 = ( ~n21253 & n21404 ) | ( ~n21253 & n21405 ) | ( n21404 & n21405 ) ;
  assign n21407 = n21242 & ~n21406 ;
  assign n21408 = ~n21242 & n21406 ;
  assign n21409 = n21407 | n21408 ;
  assign n21410 = ( ~n21196 & n21227 ) | ( ~n21196 & n21409 ) | ( n21227 & n21409 ) ;
  assign n21411 = ( n21196 & ~n21409 ) | ( n21196 & n21410 ) | ( ~n21409 & n21410 ) ;
  assign n21412 = ( ~n21227 & n21410 ) | ( ~n21227 & n21411 ) | ( n21410 & n21411 ) ;
  assign n21413 = ~n21218 & n21412 ;
  assign n21414 = n21218 & ~n21412 ;
  assign n21415 = n21413 | n21414 ;
  assign n21416 = n21205 & ~n21213 ;
  assign n21417 = n21205 & ~n21214 ;
  assign n21418 = ( ~n20515 & n21416 ) | ( ~n20515 & n21417 ) | ( n21416 & n21417 ) ;
  assign n21419 = n21415 & n21418 ;
  assign n21420 = n21415 | n21416 ;
  assign n21421 = n21415 | n21417 ;
  assign n21422 = ( ~n20515 & n21420 ) | ( ~n20515 & n21421 ) | ( n21420 & n21421 ) ;
  assign n21423 = ~n21419 & n21422 ;
  assign n21424 = x127 & ~n2769 ;
  assign n21425 = n2978 & n21424 ;
  assign n21426 = ( x127 & n2778 ) | ( x127 & n21425 ) | ( n2778 & n21425 ) ;
  assign n21427 = ( x126 & n21425 ) | ( x126 & n21426 ) | ( n21425 & n21426 ) ;
  assign n21428 = ( n12685 & n21426 ) | ( n12685 & n21427 ) | ( n21426 & n21427 ) ;
  assign n21429 = x29 & n21428 ;
  assign n21430 = x29 & ~n21429 ;
  assign n21431 = ( n21428 & ~n21429 ) | ( n21428 & n21430 ) | ( ~n21429 & n21430 ) ;
  assign n21432 = n21241 & n21431 ;
  assign n21433 = ( n21407 & n21431 ) | ( n21407 & n21432 ) | ( n21431 & n21432 ) ;
  assign n21434 = ( n21241 & n21407 ) | ( n21241 & ~n21433 ) | ( n21407 & ~n21433 ) ;
  assign n21435 = x126 & n3314 ;
  assign n21436 = x125 & n3309 ;
  assign n21437 = x124 & ~n3308 ;
  assign n21438 = n3570 & n21437 ;
  assign n21439 = n21436 | n21438 ;
  assign n21440 = n21435 | n21439 ;
  assign n21441 = n3317 | n21440 ;
  assign n21442 = ( n12687 & n21440 ) | ( n12687 & n21441 ) | ( n21440 & n21441 ) ;
  assign n21443 = x32 & n21442 ;
  assign n21444 = x32 & ~n21443 ;
  assign n21445 = ( n21442 & ~n21443 ) | ( n21442 & n21444 ) | ( ~n21443 & n21444 ) ;
  assign n21446 = n21404 | n21445 ;
  assign n21447 = n21404 & n21445 ;
  assign n21448 = n21446 & ~n21447 ;
  assign n21449 = x123 & n3913 ;
  assign n21450 = x122 & n3908 ;
  assign n21451 = x121 & ~n3907 ;
  assign n21452 = n4152 & n21451 ;
  assign n21453 = n21450 | n21452 ;
  assign n21454 = n21449 | n21453 ;
  assign n21455 = n3916 | n21454 ;
  assign n21456 = ( n11219 & n21454 ) | ( n11219 & n21455 ) | ( n21454 & n21455 ) ;
  assign n21457 = x35 & n21456 ;
  assign n21458 = x35 & ~n21457 ;
  assign n21459 = ( n21456 & ~n21457 ) | ( n21456 & n21458 ) | ( ~n21457 & n21458 ) ;
  assign n21460 = x111 & n6937 ;
  assign n21461 = x110 & n6932 ;
  assign n21462 = x109 & ~n6931 ;
  assign n21463 = n7216 & n21462 ;
  assign n21464 = n21461 | n21463 ;
  assign n21465 = n21460 | n21464 ;
  assign n21466 = n6940 | n21465 ;
  assign n21467 = ( n7492 & n21465 ) | ( n7492 & n21466 ) | ( n21465 & n21466 ) ;
  assign n21468 = x47 & n21467 ;
  assign n21469 = x47 & ~n21468 ;
  assign n21470 = ( n21467 & ~n21468 ) | ( n21467 & n21469 ) | ( ~n21468 & n21469 ) ;
  assign n21471 = ( n21344 & n21355 ) | ( n21344 & n21358 ) | ( n21355 & n21358 ) ;
  assign n21472 = x105 & n8834 ;
  assign n21473 = x104 & n8829 ;
  assign n21474 = x103 & ~n8828 ;
  assign n21475 = n9159 & n21474 ;
  assign n21476 = n21473 | n21475 ;
  assign n21477 = n21472 | n21476 ;
  assign n21478 = n8837 | n21477 ;
  assign n21479 = ( n5788 & n21477 ) | ( n5788 & n21478 ) | ( n21477 & n21478 ) ;
  assign n21480 = x53 & n21479 ;
  assign n21481 = x53 & ~n21480 ;
  assign n21482 = ( n21479 & ~n21480 ) | ( n21479 & n21481 ) | ( ~n21480 & n21481 ) ;
  assign n21483 = x102 & n9853 ;
  assign n21484 = x101 & n9848 ;
  assign n21485 = x100 & ~n9847 ;
  assign n21486 = n10165 & n21485 ;
  assign n21487 = n21484 | n21486 ;
  assign n21488 = n21483 | n21487 ;
  assign n21489 = n9856 | n21488 ;
  assign n21490 = ( n5025 & n21488 ) | ( n5025 & n21489 ) | ( n21488 & n21489 ) ;
  assign n21491 = x56 & n21490 ;
  assign n21492 = x56 & ~n21491 ;
  assign n21493 = ( n21490 & ~n21491 ) | ( n21490 & n21492 ) | ( ~n21491 & n21492 ) ;
  assign n21494 = x99 & n10876 ;
  assign n21495 = x98 & n10871 ;
  assign n21496 = x97 & ~n10870 ;
  assign n21497 = n11305 & n21496 ;
  assign n21498 = n21495 | n21497 ;
  assign n21499 = n21494 | n21498 ;
  assign n21500 = n10879 | n21499 ;
  assign n21501 = ( n4325 & n21499 ) | ( n4325 & n21500 ) | ( n21499 & n21500 ) ;
  assign n21502 = x59 & n21501 ;
  assign n21503 = x59 & ~n21502 ;
  assign n21504 = ( n21501 & ~n21502 ) | ( n21501 & n21503 ) | ( ~n21502 & n21503 ) ;
  assign n21505 = x96 & n11984 ;
  assign n21506 = x95 & n11979 ;
  assign n21507 = x94 & ~n11978 ;
  assign n21508 = n12430 & n21507 ;
  assign n21509 = n21506 | n21508 ;
  assign n21510 = n21505 | n21509 ;
  assign n21511 = n11987 | n21510 ;
  assign n21512 = ( n3509 & n21510 ) | ( n3509 & n21511 ) | ( n21510 & n21511 ) ;
  assign n21513 = x62 & n21512 ;
  assign n21514 = x62 & ~n21513 ;
  assign n21515 = ( n21512 & ~n21513 ) | ( n21512 & n21514 ) | ( ~n21513 & n21514 ) ;
  assign n21516 = x93 & n12808 ;
  assign n21517 = x63 & x92 ;
  assign n21518 = ~n12808 & n21517 ;
  assign n21519 = n21516 | n21518 ;
  assign n21520 = ~n21327 & n21519 ;
  assign n21521 = n21327 & ~n21519 ;
  assign n21522 = ( n21328 & ~n21519 ) | ( n21328 & n21521 ) | ( ~n21519 & n21521 ) ;
  assign n21523 = n21520 | n21522 ;
  assign n21524 = n21335 | n21523 ;
  assign n21525 = n21520 | n21521 ;
  assign n21526 = ( n21330 & n21335 ) | ( n21330 & n21525 ) | ( n21335 & n21525 ) ;
  assign n21527 = n21524 & ~n21526 ;
  assign n21528 = ( n21504 & ~n21515 ) | ( n21504 & n21527 ) | ( ~n21515 & n21527 ) ;
  assign n21529 = ( n21515 & ~n21527 ) | ( n21515 & n21528 ) | ( ~n21527 & n21528 ) ;
  assign n21530 = ( ~n21504 & n21528 ) | ( ~n21504 & n21529 ) | ( n21528 & n21529 ) ;
  assign n21531 = ( ~n21339 & n21493 ) | ( ~n21339 & n21530 ) | ( n21493 & n21530 ) ;
  assign n21532 = ( n21339 & ~n21530 ) | ( n21339 & n21531 ) | ( ~n21530 & n21531 ) ;
  assign n21533 = ( ~n21493 & n21531 ) | ( ~n21493 & n21532 ) | ( n21531 & n21532 ) ;
  assign n21534 = ( n21342 & n21482 ) | ( n21342 & ~n21533 ) | ( n21482 & ~n21533 ) ;
  assign n21535 = ( ~n21342 & n21533 ) | ( ~n21342 & n21534 ) | ( n21533 & n21534 ) ;
  assign n21536 = ( ~n21482 & n21534 ) | ( ~n21482 & n21535 ) | ( n21534 & n21535 ) ;
  assign n21537 = n21471 & ~n21536 ;
  assign n21538 = ~n21471 & n21536 ;
  assign n21539 = n21537 | n21538 ;
  assign n21540 = x108 & n7812 ;
  assign n21541 = x107 & n7807 ;
  assign n21542 = x106 & ~n7806 ;
  assign n21543 = n8136 & n21542 ;
  assign n21544 = n21541 | n21543 ;
  assign n21545 = n21540 | n21544 ;
  assign n21546 = n7815 | n21545 ;
  assign n21547 = ( n6358 & n21545 ) | ( n6358 & n21546 ) | ( n21545 & n21546 ) ;
  assign n21548 = x50 & n21547 ;
  assign n21549 = x50 & ~n21548 ;
  assign n21550 = ( n21547 & ~n21548 ) | ( n21547 & n21549 ) | ( ~n21548 & n21549 ) ;
  assign n21551 = ~n21539 & n21550 ;
  assign n21552 = n21539 & ~n21550 ;
  assign n21553 = n21551 | n21552 ;
  assign n21554 = ( ~n21359 & n21470 ) | ( ~n21359 & n21553 ) | ( n21470 & n21553 ) ;
  assign n21555 = ( n21359 & ~n21553 ) | ( n21359 & n21554 ) | ( ~n21553 & n21554 ) ;
  assign n21556 = ( ~n21470 & n21554 ) | ( ~n21470 & n21555 ) | ( n21554 & n21555 ) ;
  assign n21557 = ~n21377 & n21556 ;
  assign n21558 = n21377 & ~n21556 ;
  assign n21559 = n21557 | n21558 ;
  assign n21560 = x114 & n6068 ;
  assign n21561 = x113 & n6063 ;
  assign n21562 = x112 & ~n6062 ;
  assign n21563 = n6398 & n21562 ;
  assign n21564 = n21561 | n21563 ;
  assign n21565 = n21560 | n21564 ;
  assign n21566 = n6071 | n21565 ;
  assign n21567 = ( n8437 & n21565 ) | ( n8437 & n21566 ) | ( n21565 & n21566 ) ;
  assign n21568 = x44 & n21567 ;
  assign n21569 = x44 & ~n21568 ;
  assign n21570 = ( n21567 & ~n21568 ) | ( n21567 & n21569 ) | ( ~n21568 & n21569 ) ;
  assign n21571 = n21559 & ~n21570 ;
  assign n21572 = ~n21559 & n21570 ;
  assign n21573 = n21571 | n21572 ;
  assign n21574 = n21381 & n21573 ;
  assign n21575 = n21381 & ~n21573 ;
  assign n21576 = n21573 | n21575 ;
  assign n21577 = x117 & n5340 ;
  assign n21578 = x116 & n5335 ;
  assign n21579 = x115 & ~n5334 ;
  assign n21580 = n5580 & n21579 ;
  assign n21581 = n21578 | n21580 ;
  assign n21582 = n21577 | n21581 ;
  assign n21583 = n5343 | n21582 ;
  assign n21584 = ( n9118 & n21582 ) | ( n9118 & n21583 ) | ( n21582 & n21583 ) ;
  assign n21585 = x41 & n21584 ;
  assign n21586 = x41 & ~n21585 ;
  assign n21587 = ( n21584 & ~n21585 ) | ( n21584 & n21586 ) | ( ~n21585 & n21586 ) ;
  assign n21588 = n21576 & ~n21587 ;
  assign n21589 = ~n21574 & n21588 ;
  assign n21590 = ( n21574 & ~n21576 ) | ( n21574 & n21587 ) | ( ~n21576 & n21587 ) ;
  assign n21591 = n21589 | n21590 ;
  assign n21592 = n21398 & ~n21591 ;
  assign n21593 = ~n21398 & n21591 ;
  assign n21594 = n21592 | n21593 ;
  assign n21595 = x120 & n4572 ;
  assign n21596 = x119 & n4567 ;
  assign n21597 = x118 & ~n4566 ;
  assign n21598 = n4828 & n21597 ;
  assign n21599 = n21596 | n21598 ;
  assign n21600 = n21595 | n21599 ;
  assign n21601 = n4575 | n21600 ;
  assign n21602 = ( n10460 & n21600 ) | ( n10460 & n21601 ) | ( n21600 & n21601 ) ;
  assign n21603 = x38 & n21602 ;
  assign n21604 = x38 & ~n21603 ;
  assign n21605 = ( n21602 & ~n21603 ) | ( n21602 & n21604 ) | ( ~n21603 & n21604 ) ;
  assign n21606 = ~n21594 & n21605 ;
  assign n21607 = n21594 & ~n21605 ;
  assign n21608 = n21606 | n21607 ;
  assign n21609 = ( ~n21401 & n21459 ) | ( ~n21401 & n21608 ) | ( n21459 & n21608 ) ;
  assign n21610 = ( n21401 & ~n21608 ) | ( n21401 & n21609 ) | ( ~n21608 & n21609 ) ;
  assign n21611 = ( ~n21459 & n21609 ) | ( ~n21459 & n21610 ) | ( n21609 & n21610 ) ;
  assign n21612 = ~n21448 & n21611 ;
  assign n21613 = n21448 & ~n21611 ;
  assign n21614 = n21612 | n21613 ;
  assign n21615 = n21431 & ~n21432 ;
  assign n21616 = ~n21407 & n21615 ;
  assign n21617 = n21614 & ~n21616 ;
  assign n21618 = ~n21434 & n21617 ;
  assign n21619 = ( n21434 & ~n21614 ) | ( n21434 & n21616 ) | ( ~n21614 & n21616 ) ;
  assign n21620 = n21618 | n21619 ;
  assign n21621 = n21411 & ~n21620 ;
  assign n21622 = n21411 & ~n21621 ;
  assign n21623 = ~n21414 & n21420 ;
  assign n21624 = ~n21414 & n21421 ;
  assign n21625 = ( ~n20515 & n21623 ) | ( ~n20515 & n21624 ) | ( n21623 & n21624 ) ;
  assign n21626 = n21411 | n21620 ;
  assign n21627 = n21625 & n21626 ;
  assign n21628 = ~n21622 & n21627 ;
  assign n21629 = ~n21622 & n21626 ;
  assign n21630 = n21623 | n21629 ;
  assign n21631 = n21624 | n21629 ;
  assign n21632 = ( ~n20515 & n21630 ) | ( ~n20515 & n21631 ) | ( n21630 & n21631 ) ;
  assign n21633 = ~n21628 & n21632 ;
  assign n21634 = n21433 | n21619 ;
  assign n21635 = n21447 | n21613 ;
  assign n21636 = x127 & n3314 ;
  assign n21637 = x126 & n3309 ;
  assign n21638 = x125 & ~n3308 ;
  assign n21639 = n3570 & n21638 ;
  assign n21640 = n21637 | n21639 ;
  assign n21641 = n21636 | n21640 ;
  assign n21642 = n3317 | n21641 ;
  assign n21643 = ( n12720 & n21641 ) | ( n12720 & n21642 ) | ( n21641 & n21642 ) ;
  assign n21644 = x32 & n21643 ;
  assign n21645 = x32 & ~n21644 ;
  assign n21646 = ( n21643 & ~n21644 ) | ( n21643 & n21645 ) | ( ~n21644 & n21645 ) ;
  assign n21647 = n21635 & n21646 ;
  assign n21648 = n21635 & ~n21647 ;
  assign n21649 = x124 & n3913 ;
  assign n21650 = x123 & n3908 ;
  assign n21651 = x122 & ~n3907 ;
  assign n21652 = n4152 & n21651 ;
  assign n21653 = n21650 | n21652 ;
  assign n21654 = n21649 | n21653 ;
  assign n21655 = n3916 | n21654 ;
  assign n21656 = ( n11916 & n21654 ) | ( n11916 & n21655 ) | ( n21654 & n21655 ) ;
  assign n21657 = x35 & n21656 ;
  assign n21658 = x35 & ~n21657 ;
  assign n21659 = ( n21656 & ~n21657 ) | ( n21656 & n21658 ) | ( ~n21657 & n21658 ) ;
  assign n21660 = n21575 | n21590 ;
  assign n21661 = n21558 | n21572 ;
  assign n21662 = x112 & n6937 ;
  assign n21663 = x111 & n6932 ;
  assign n21664 = x110 & ~n6931 ;
  assign n21665 = n7216 & n21664 ;
  assign n21666 = n21663 | n21665 ;
  assign n21667 = n21662 | n21666 ;
  assign n21668 = n6940 | n21667 ;
  assign n21669 = ( n7789 & n21667 ) | ( n7789 & n21668 ) | ( n21667 & n21668 ) ;
  assign n21670 = x47 & n21669 ;
  assign n21671 = x47 & ~n21670 ;
  assign n21672 = ( n21669 & ~n21670 ) | ( n21669 & n21671 ) | ( ~n21670 & n21671 ) ;
  assign n21673 = x109 & n7812 ;
  assign n21674 = x108 & n7807 ;
  assign n21675 = x107 & ~n7806 ;
  assign n21676 = n8136 & n21675 ;
  assign n21677 = n21674 | n21676 ;
  assign n21678 = n21673 | n21677 ;
  assign n21679 = n7815 | n21678 ;
  assign n21680 = ( n6884 & n21678 ) | ( n6884 & n21679 ) | ( n21678 & n21679 ) ;
  assign n21681 = x50 & n21680 ;
  assign n21682 = x50 & ~n21681 ;
  assign n21683 = ( n21680 & ~n21681 ) | ( n21680 & n21682 ) | ( ~n21681 & n21682 ) ;
  assign n21684 = x106 & n8834 ;
  assign n21685 = x105 & n8829 ;
  assign n21686 = x104 & ~n8828 ;
  assign n21687 = n9159 & n21686 ;
  assign n21688 = n21685 | n21687 ;
  assign n21689 = n21684 | n21688 ;
  assign n21690 = n8837 | n21689 ;
  assign n21691 = ( n5814 & n21689 ) | ( n5814 & n21690 ) | ( n21689 & n21690 ) ;
  assign n21692 = x53 & n21691 ;
  assign n21693 = x53 & ~n21692 ;
  assign n21694 = ( n21691 & ~n21692 ) | ( n21691 & n21693 ) | ( ~n21692 & n21693 ) ;
  assign n21695 = ( n21335 & ~n21520 ) | ( n21335 & n21522 ) | ( ~n21520 & n21522 ) ;
  assign n21696 = x94 & n12808 ;
  assign n21697 = x63 & x93 ;
  assign n21698 = ~n12808 & n21697 ;
  assign n21699 = n21696 | n21698 ;
  assign n21700 = ~x29 & n21699 ;
  assign n21701 = x29 & ~n21699 ;
  assign n21702 = n21700 | n21701 ;
  assign n21703 = n21519 | n21702 ;
  assign n21704 = n21519 & ~n21702 ;
  assign n21705 = ( ~n21519 & n21703 ) | ( ~n21519 & n21704 ) | ( n21703 & n21704 ) ;
  assign n21706 = n21695 & ~n21705 ;
  assign n21707 = n21695 & ~n21706 ;
  assign n21708 = n21695 | n21705 ;
  assign n21709 = ~n21707 & n21708 ;
  assign n21710 = x97 & n11984 ;
  assign n21711 = x96 & n11979 ;
  assign n21712 = x95 & ~n11978 ;
  assign n21713 = n12430 & n21712 ;
  assign n21714 = n21711 | n21713 ;
  assign n21715 = n21710 | n21714 ;
  assign n21716 = n11987 | n21715 ;
  assign n21717 = ( n3707 & n21715 ) | ( n3707 & n21716 ) | ( n21715 & n21716 ) ;
  assign n21718 = x62 & n21717 ;
  assign n21719 = x62 & ~n21718 ;
  assign n21720 = ( n21717 & ~n21718 ) | ( n21717 & n21719 ) | ( ~n21718 & n21719 ) ;
  assign n21721 = n21709 & n21720 ;
  assign n21722 = ( n21707 & ~n21708 ) | ( n21707 & n21720 ) | ( ~n21708 & n21720 ) ;
  assign n21723 = ( n21709 & ~n21721 ) | ( n21709 & n21722 ) | ( ~n21721 & n21722 ) ;
  assign n21724 = x100 & n10876 ;
  assign n21725 = x99 & n10871 ;
  assign n21726 = x98 & ~n10870 ;
  assign n21727 = n11305 & n21726 ;
  assign n21728 = n21725 | n21727 ;
  assign n21729 = n21724 | n21728 ;
  assign n21730 = n10879 | n21729 ;
  assign n21731 = ( n4532 & n21729 ) | ( n4532 & n21730 ) | ( n21729 & n21730 ) ;
  assign n21732 = x59 & n21731 ;
  assign n21733 = x59 & ~n21732 ;
  assign n21734 = ( n21731 & ~n21732 ) | ( n21731 & n21733 ) | ( ~n21732 & n21733 ) ;
  assign n21735 = ~n21723 & n21734 ;
  assign n21736 = n21723 & ~n21734 ;
  assign n21737 = n21735 | n21736 ;
  assign n21738 = n21529 & ~n21737 ;
  assign n21739 = ~n21529 & n21737 ;
  assign n21740 = n21738 | n21739 ;
  assign n21741 = x103 & n9853 ;
  assign n21742 = x102 & n9848 ;
  assign n21743 = x101 & ~n9847 ;
  assign n21744 = n10165 & n21743 ;
  assign n21745 = n21742 | n21744 ;
  assign n21746 = n21741 | n21745 ;
  assign n21747 = n9856 | n21746 ;
  assign n21748 = ( n5264 & n21746 ) | ( n5264 & n21747 ) | ( n21746 & n21747 ) ;
  assign n21749 = x56 & n21748 ;
  assign n21750 = x56 & ~n21749 ;
  assign n21751 = ( n21748 & ~n21749 ) | ( n21748 & n21750 ) | ( ~n21749 & n21750 ) ;
  assign n21752 = ~n21740 & n21751 ;
  assign n21753 = n21740 | n21752 ;
  assign n21754 = n21740 & n21751 ;
  assign n21755 = n21532 | n21754 ;
  assign n21756 = n21753 & ~n21755 ;
  assign n21757 = ( n21532 & ~n21753 ) | ( n21532 & n21754 ) | ( ~n21753 & n21754 ) ;
  assign n21758 = n21756 | n21757 ;
  assign n21759 = ( n21534 & n21694 ) | ( n21534 & ~n21758 ) | ( n21694 & ~n21758 ) ;
  assign n21760 = ( ~n21534 & n21758 ) | ( ~n21534 & n21759 ) | ( n21758 & n21759 ) ;
  assign n21761 = ( ~n21694 & n21759 ) | ( ~n21694 & n21760 ) | ( n21759 & n21760 ) ;
  assign n21762 = n21683 & ~n21761 ;
  assign n21763 = ~n21683 & n21761 ;
  assign n21764 = n21762 | n21763 ;
  assign n21765 = n21537 | n21551 ;
  assign n21766 = n21764 & ~n21765 ;
  assign n21767 = ~n21764 & n21765 ;
  assign n21768 = n21766 | n21767 ;
  assign n21769 = n21672 & ~n21768 ;
  assign n21770 = n21768 | n21769 ;
  assign n21771 = ( ~n21672 & n21769 ) | ( ~n21672 & n21770 ) | ( n21769 & n21770 ) ;
  assign n21772 = ~n21555 & n21771 ;
  assign n21773 = n21555 & ~n21771 ;
  assign n21774 = n21772 | n21773 ;
  assign n21775 = x115 & n6068 ;
  assign n21776 = x114 & n6063 ;
  assign n21777 = x113 & ~n6062 ;
  assign n21778 = n6398 & n21777 ;
  assign n21779 = n21776 | n21778 ;
  assign n21780 = n21775 | n21779 ;
  assign n21781 = n6071 | n21780 ;
  assign n21782 = ( n8749 & n21780 ) | ( n8749 & n21781 ) | ( n21780 & n21781 ) ;
  assign n21783 = x44 & n21782 ;
  assign n21784 = x44 & ~n21783 ;
  assign n21785 = ( n21782 & ~n21783 ) | ( n21782 & n21784 ) | ( ~n21783 & n21784 ) ;
  assign n21786 = ~n21774 & n21785 ;
  assign n21787 = n21774 & ~n21785 ;
  assign n21788 = n21786 | n21787 ;
  assign n21789 = n21661 & ~n21788 ;
  assign n21790 = n21661 & ~n21789 ;
  assign n21791 = n21788 | n21789 ;
  assign n21792 = ~n21790 & n21791 ;
  assign n21793 = x118 & n5340 ;
  assign n21794 = x117 & n5335 ;
  assign n21795 = x116 & ~n5334 ;
  assign n21796 = n5580 & n21795 ;
  assign n21797 = n21794 | n21796 ;
  assign n21798 = n21793 | n21797 ;
  assign n21799 = n5343 | n21798 ;
  assign n21800 = ( n9760 & n21798 ) | ( n9760 & n21799 ) | ( n21798 & n21799 ) ;
  assign n21801 = x41 & n21800 ;
  assign n21802 = x41 & ~n21801 ;
  assign n21803 = ( n21800 & ~n21801 ) | ( n21800 & n21802 ) | ( ~n21801 & n21802 ) ;
  assign n21804 = n21792 & ~n21803 ;
  assign n21805 = ~n21792 & n21803 ;
  assign n21806 = n21804 | n21805 ;
  assign n21807 = n21660 & ~n21806 ;
  assign n21808 = ~n21660 & n21806 ;
  assign n21809 = n21807 | n21808 ;
  assign n21810 = x121 & n4572 ;
  assign n21811 = x120 & n4567 ;
  assign n21812 = x119 & ~n4566 ;
  assign n21813 = n4828 & n21812 ;
  assign n21814 = n21811 | n21813 ;
  assign n21815 = n21810 | n21814 ;
  assign n21816 = n4575 | n21815 ;
  assign n21817 = ( n10811 & n21815 ) | ( n10811 & n21816 ) | ( n21815 & n21816 ) ;
  assign n21818 = x38 & n21817 ;
  assign n21819 = x38 & ~n21818 ;
  assign n21820 = ( n21817 & ~n21818 ) | ( n21817 & n21819 ) | ( ~n21818 & n21819 ) ;
  assign n21821 = ~n21809 & n21820 ;
  assign n21822 = n21809 | n21821 ;
  assign n21823 = n21809 & n21820 ;
  assign n21824 = n21592 | n21606 ;
  assign n21825 = n21823 | n21824 ;
  assign n21826 = n21822 & ~n21825 ;
  assign n21827 = ( ~n21822 & n21823 ) | ( ~n21822 & n21824 ) | ( n21823 & n21824 ) ;
  assign n21828 = n21826 | n21827 ;
  assign n21829 = n21659 & ~n21828 ;
  assign n21830 = n21828 | n21829 ;
  assign n21831 = ( ~n21659 & n21829 ) | ( ~n21659 & n21830 ) | ( n21829 & n21830 ) ;
  assign n21832 = ~n21610 & n21831 ;
  assign n21833 = n21610 & ~n21831 ;
  assign n21834 = n21832 | n21833 ;
  assign n21835 = ~n21635 & n21646 ;
  assign n21836 = n21834 & ~n21835 ;
  assign n21837 = ~n21648 & n21836 ;
  assign n21838 = ( n21648 & ~n21834 ) | ( n21648 & n21835 ) | ( ~n21834 & n21835 ) ;
  assign n21839 = n21837 | n21838 ;
  assign n21840 = n21634 & ~n21839 ;
  assign n21841 = ~n21634 & n21839 ;
  assign n21842 = n21840 | n21841 ;
  assign n21843 = ~n21621 & n21630 ;
  assign n21844 = ~n21621 & n21631 ;
  assign n21845 = ( ~n20515 & n21843 ) | ( ~n20515 & n21844 ) | ( n21843 & n21844 ) ;
  assign n21846 = n21842 & n21845 ;
  assign n21847 = n21842 | n21843 ;
  assign n21848 = n21842 | n21844 ;
  assign n21849 = ( ~n20515 & n21847 ) | ( ~n20515 & n21848 ) | ( n21847 & n21848 ) ;
  assign n21850 = ~n21846 & n21849 ;
  assign n21851 = n21647 | n21838 ;
  assign n21852 = x125 & n3913 ;
  assign n21853 = x124 & n3908 ;
  assign n21854 = x123 & ~n3907 ;
  assign n21855 = n4152 & n21854 ;
  assign n21856 = n21853 | n21855 ;
  assign n21857 = n21852 | n21856 ;
  assign n21858 = n3916 | n21857 ;
  assign n21859 = ( n12310 & n21857 ) | ( n12310 & n21858 ) | ( n21857 & n21858 ) ;
  assign n21860 = x35 & n21859 ;
  assign n21861 = x35 & ~n21860 ;
  assign n21862 = ( n21859 & ~n21860 ) | ( n21859 & n21861 ) | ( ~n21860 & n21861 ) ;
  assign n21863 = x127 & n3309 ;
  assign n21864 = x126 & ~n3308 ;
  assign n21865 = n3570 & n21864 ;
  assign n21866 = n21863 | n21865 ;
  assign n21867 = n3317 | n21866 ;
  assign n21868 = ( n13461 & n21866 ) | ( n13461 & n21867 ) | ( n21866 & n21867 ) ;
  assign n21869 = x32 & n21868 ;
  assign n21870 = x32 & ~n21869 ;
  assign n21871 = ( n21868 & ~n21869 ) | ( n21868 & n21870 ) | ( ~n21869 & n21870 ) ;
  assign n21872 = n21829 | n21833 ;
  assign n21873 = n21871 & n21872 ;
  assign n21874 = n21871 | n21872 ;
  assign n21875 = ~n21873 & n21874 ;
  assign n21876 = n21821 | n21827 ;
  assign n21877 = x122 & n4572 ;
  assign n21878 = x121 & n4567 ;
  assign n21879 = x120 & ~n4566 ;
  assign n21880 = n4828 & n21879 ;
  assign n21881 = n21878 | n21880 ;
  assign n21882 = n21877 | n21881 ;
  assign n21883 = n4575 | n21882 ;
  assign n21884 = ( n11188 & n21882 ) | ( n11188 & n21883 ) | ( n21882 & n21883 ) ;
  assign n21885 = x38 & n21884 ;
  assign n21886 = x38 & ~n21885 ;
  assign n21887 = ( n21884 & ~n21885 ) | ( n21884 & n21886 ) | ( ~n21885 & n21886 ) ;
  assign n21888 = n21805 | n21807 ;
  assign n21889 = x119 & n5340 ;
  assign n21890 = x118 & n5335 ;
  assign n21891 = x117 & ~n5334 ;
  assign n21892 = n5580 & n21891 ;
  assign n21893 = n21890 | n21892 ;
  assign n21894 = n21889 | n21893 ;
  assign n21895 = n5343 | n21894 ;
  assign n21896 = ( n9789 & n21894 ) | ( n9789 & n21895 ) | ( n21894 & n21895 ) ;
  assign n21897 = x41 & n21896 ;
  assign n21898 = x41 & ~n21897 ;
  assign n21899 = ( n21896 & ~n21897 ) | ( n21896 & n21898 ) | ( ~n21897 & n21898 ) ;
  assign n21900 = n21786 | n21789 ;
  assign n21901 = x116 & n6068 ;
  assign n21902 = x115 & n6063 ;
  assign n21903 = x114 & ~n6062 ;
  assign n21904 = n6398 & n21903 ;
  assign n21905 = n21902 | n21904 ;
  assign n21906 = n21901 | n21905 ;
  assign n21907 = n6071 | n21906 ;
  assign n21908 = ( n8778 & n21906 ) | ( n8778 & n21907 ) | ( n21906 & n21907 ) ;
  assign n21909 = x44 & n21908 ;
  assign n21910 = x44 & ~n21909 ;
  assign n21911 = ( n21908 & ~n21909 ) | ( n21908 & n21910 ) | ( ~n21909 & n21910 ) ;
  assign n21912 = n21769 | n21773 ;
  assign n21913 = x107 & n8834 ;
  assign n21914 = x106 & n8829 ;
  assign n21915 = x105 & ~n8828 ;
  assign n21916 = n9159 & n21915 ;
  assign n21917 = n21914 | n21916 ;
  assign n21918 = n21913 | n21917 ;
  assign n21919 = n8837 | n21918 ;
  assign n21920 = ( n6328 & n21918 ) | ( n6328 & n21919 ) | ( n21918 & n21919 ) ;
  assign n21921 = x53 & n21920 ;
  assign n21922 = x53 & ~n21921 ;
  assign n21923 = ( n21920 & ~n21921 ) | ( n21920 & n21922 ) | ( ~n21921 & n21922 ) ;
  assign n21924 = n21752 | n21757 ;
  assign n21925 = n21735 | n21738 ;
  assign n21926 = x98 & n11984 ;
  assign n21927 = x97 & n11979 ;
  assign n21928 = x96 & ~n11978 ;
  assign n21929 = n12430 & n21928 ;
  assign n21930 = n21927 | n21929 ;
  assign n21931 = n21926 | n21930 ;
  assign n21932 = n11987 | n21931 ;
  assign n21933 = ( n4105 & n21931 ) | ( n4105 & n21932 ) | ( n21931 & n21932 ) ;
  assign n21934 = ~x62 & n21933 ;
  assign n21935 = x95 & n12808 ;
  assign n21936 = x63 & x94 ;
  assign n21937 = ~n12808 & n21936 ;
  assign n21938 = n21935 | n21937 ;
  assign n21939 = n21700 | n21704 ;
  assign n21940 = n21938 & ~n21939 ;
  assign n21941 = ~n21938 & n21939 ;
  assign n21942 = n21940 | n21941 ;
  assign n21943 = x62 & ~n21933 ;
  assign n21944 = n21942 & ~n21943 ;
  assign n21945 = ~n21934 & n21944 ;
  assign n21946 = ( n21934 & ~n21942 ) | ( n21934 & n21943 ) | ( ~n21942 & n21943 ) ;
  assign n21947 = n21945 | n21946 ;
  assign n21948 = n21706 & ~n21947 ;
  assign n21949 = n21947 | n21948 ;
  assign n21950 = n21722 | n21949 ;
  assign n21951 = x101 & n10876 ;
  assign n21952 = x100 & n10871 ;
  assign n21953 = x99 & ~n10870 ;
  assign n21954 = n11305 & n21953 ;
  assign n21955 = n21952 | n21954 ;
  assign n21956 = n21951 | n21955 ;
  assign n21957 = n10879 | n21956 ;
  assign n21958 = ( n4783 & n21956 ) | ( n4783 & n21957 ) | ( n21956 & n21957 ) ;
  assign n21959 = x59 & n21958 ;
  assign n21960 = x59 & ~n21959 ;
  assign n21961 = ( n21958 & ~n21959 ) | ( n21958 & n21960 ) | ( ~n21959 & n21960 ) ;
  assign n21962 = n21950 & ~n21961 ;
  assign n21963 = ( n21706 & n21722 ) | ( n21706 & n21947 ) | ( n21722 & n21947 ) ;
  assign n21964 = n21962 & ~n21963 ;
  assign n21965 = ( ~n21950 & n21961 ) | ( ~n21950 & n21963 ) | ( n21961 & n21963 ) ;
  assign n21966 = n21964 | n21965 ;
  assign n21967 = x104 & n9853 ;
  assign n21968 = x103 & n9848 ;
  assign n21969 = x102 & ~n9847 ;
  assign n21970 = n10165 & n21969 ;
  assign n21971 = n21968 | n21970 ;
  assign n21972 = n21967 | n21971 ;
  assign n21973 = n9856 | n21972 ;
  assign n21974 = ( n5295 & n21972 ) | ( n5295 & n21973 ) | ( n21972 & n21973 ) ;
  assign n21975 = x56 & n21974 ;
  assign n21976 = x56 & ~n21975 ;
  assign n21977 = ( n21974 & ~n21975 ) | ( n21974 & n21976 ) | ( ~n21975 & n21976 ) ;
  assign n21978 = ( n21925 & ~n21966 ) | ( n21925 & n21977 ) | ( ~n21966 & n21977 ) ;
  assign n21979 = ( n21966 & ~n21977 ) | ( n21966 & n21978 ) | ( ~n21977 & n21978 ) ;
  assign n21980 = ( ~n21925 & n21978 ) | ( ~n21925 & n21979 ) | ( n21978 & n21979 ) ;
  assign n21981 = ( n21923 & n21924 ) | ( n21923 & ~n21980 ) | ( n21924 & ~n21980 ) ;
  assign n21982 = ( ~n21924 & n21980 ) | ( ~n21924 & n21981 ) | ( n21980 & n21981 ) ;
  assign n21983 = ( ~n21923 & n21981 ) | ( ~n21923 & n21982 ) | ( n21981 & n21982 ) ;
  assign n21984 = ~n21759 & n21983 ;
  assign n21985 = n21759 & ~n21983 ;
  assign n21986 = n21984 | n21985 ;
  assign n21987 = x110 & n7812 ;
  assign n21988 = x109 & n7807 ;
  assign n21989 = x108 & ~n7806 ;
  assign n21990 = n8136 & n21989 ;
  assign n21991 = n21988 | n21990 ;
  assign n21992 = n21987 | n21991 ;
  assign n21993 = n7815 | n21992 ;
  assign n21994 = ( n7189 & n21992 ) | ( n7189 & n21993 ) | ( n21992 & n21993 ) ;
  assign n21995 = x50 & n21994 ;
  assign n21996 = x50 & ~n21995 ;
  assign n21997 = ( n21994 & ~n21995 ) | ( n21994 & n21996 ) | ( ~n21995 & n21996 ) ;
  assign n21998 = n21986 & n21997 ;
  assign n21999 = ( n21759 & ~n21983 ) | ( n21759 & n21997 ) | ( ~n21983 & n21997 ) ;
  assign n22000 = n21984 | n21999 ;
  assign n22001 = ~n21998 & n22000 ;
  assign n22002 = n21762 | n21767 ;
  assign n22003 = n22001 & ~n22002 ;
  assign n22004 = ~n22001 & n22002 ;
  assign n22005 = n22003 | n22004 ;
  assign n22006 = x113 & n6937 ;
  assign n22007 = x112 & n6932 ;
  assign n22008 = x111 & ~n6931 ;
  assign n22009 = n7216 & n22008 ;
  assign n22010 = n22007 | n22009 ;
  assign n22011 = n22006 | n22010 ;
  assign n22012 = n6940 | n22011 ;
  assign n22013 = ( n8113 & n22011 ) | ( n8113 & n22012 ) | ( n22011 & n22012 ) ;
  assign n22014 = x47 & n22013 ;
  assign n22015 = x47 & ~n22014 ;
  assign n22016 = ( n22013 & ~n22014 ) | ( n22013 & n22015 ) | ( ~n22014 & n22015 ) ;
  assign n22017 = n22005 & n22016 ;
  assign n22018 = ( ~n22001 & n22002 ) | ( ~n22001 & n22016 ) | ( n22002 & n22016 ) ;
  assign n22019 = n22003 | n22018 ;
  assign n22020 = ~n22017 & n22019 ;
  assign n22021 = ( n21911 & ~n21912 ) | ( n21911 & n22020 ) | ( ~n21912 & n22020 ) ;
  assign n22022 = ( n21912 & ~n22020 ) | ( n21912 & n22021 ) | ( ~n22020 & n22021 ) ;
  assign n22023 = ( ~n21911 & n22021 ) | ( ~n21911 & n22022 ) | ( n22021 & n22022 ) ;
  assign n22024 = ( n21899 & n21900 ) | ( n21899 & ~n22023 ) | ( n21900 & ~n22023 ) ;
  assign n22025 = ( ~n21900 & n22023 ) | ( ~n21900 & n22024 ) | ( n22023 & n22024 ) ;
  assign n22026 = ( ~n21899 & n22024 ) | ( ~n21899 & n22025 ) | ( n22024 & n22025 ) ;
  assign n22027 = ( n21887 & n21888 ) | ( n21887 & ~n22026 ) | ( n21888 & ~n22026 ) ;
  assign n22028 = ( ~n21888 & n22026 ) | ( ~n21888 & n22027 ) | ( n22026 & n22027 ) ;
  assign n22029 = ( ~n21887 & n22027 ) | ( ~n21887 & n22028 ) | ( n22027 & n22028 ) ;
  assign n22030 = ~n21876 & n22029 ;
  assign n22031 = n21876 & ~n22029 ;
  assign n22032 = n22030 | n22031 ;
  assign n22033 = ( n21862 & n21875 ) | ( n21862 & ~n22032 ) | ( n21875 & ~n22032 ) ;
  assign n22034 = ( ~n21875 & n22032 ) | ( ~n21875 & n22033 ) | ( n22032 & n22033 ) ;
  assign n22035 = ( ~n21862 & n22033 ) | ( ~n21862 & n22034 ) | ( n22033 & n22034 ) ;
  assign n22036 = n21851 & ~n22035 ;
  assign n22037 = n21851 & ~n22036 ;
  assign n22038 = n21851 | n22035 ;
  assign n22039 = ~n22037 & n22038 ;
  assign n22040 = ~n21840 & n21847 ;
  assign n22041 = ~n21840 & n21848 ;
  assign n22042 = ( ~n20515 & n22040 ) | ( ~n20515 & n22041 ) | ( n22040 & n22041 ) ;
  assign n22043 = n22039 & n22042 ;
  assign n22044 = n22039 | n22040 ;
  assign n22045 = n22039 | n22041 ;
  assign n22046 = ( ~n20515 & n22044 ) | ( ~n20515 & n22045 ) | ( n22044 & n22045 ) ;
  assign n22047 = ~n22043 & n22046 ;
  assign n22048 = x123 & n4572 ;
  assign n22049 = x122 & n4567 ;
  assign n22050 = x121 & ~n4566 ;
  assign n22051 = n4828 & n22050 ;
  assign n22052 = n22049 | n22051 ;
  assign n22053 = n22048 | n22052 ;
  assign n22054 = n4575 | n22053 ;
  assign n22055 = ( n11219 & n22053 ) | ( n11219 & n22054 ) | ( n22053 & n22054 ) ;
  assign n22056 = x38 & n22055 ;
  assign n22057 = x38 & ~n22056 ;
  assign n22058 = ( n22055 & ~n22056 ) | ( n22055 & n22057 ) | ( ~n22056 & n22057 ) ;
  assign n22059 = x111 & n7812 ;
  assign n22060 = x110 & n7807 ;
  assign n22061 = x109 & ~n7806 ;
  assign n22062 = n8136 & n22061 ;
  assign n22063 = n22060 | n22062 ;
  assign n22064 = n22059 | n22063 ;
  assign n22065 = n7815 | n22064 ;
  assign n22066 = ( n7492 & n22064 ) | ( n7492 & n22065 ) | ( n22064 & n22065 ) ;
  assign n22067 = x50 & n22066 ;
  assign n22068 = x50 & ~n22067 ;
  assign n22069 = ( n22066 & ~n22067 ) | ( n22066 & n22068 ) | ( ~n22067 & n22068 ) ;
  assign n22070 = x99 & n11984 ;
  assign n22071 = x98 & n11979 ;
  assign n22072 = x97 & ~n11978 ;
  assign n22073 = n12430 & n22072 ;
  assign n22074 = n22071 | n22073 ;
  assign n22075 = n22070 | n22074 ;
  assign n22076 = n11987 | n22075 ;
  assign n22077 = ( n4325 & n22075 ) | ( n4325 & n22076 ) | ( n22075 & n22076 ) ;
  assign n22078 = x62 & n22077 ;
  assign n22079 = x62 & ~n22078 ;
  assign n22080 = ( n22077 & ~n22078 ) | ( n22077 & n22079 ) | ( ~n22078 & n22079 ) ;
  assign n22081 = x96 & n12808 ;
  assign n22082 = x63 & x95 ;
  assign n22083 = ~n12808 & n22082 ;
  assign n22084 = n22081 | n22083 ;
  assign n22085 = ( n21938 & n21946 ) | ( n21938 & n22084 ) | ( n21946 & n22084 ) ;
  assign n22086 = n21938 | n21939 ;
  assign n22087 = ( n21946 & n22084 ) | ( n21946 & ~n22086 ) | ( n22084 & ~n22086 ) ;
  assign n22088 = ~n21938 & n22084 ;
  assign n22089 = ( n21939 & n21940 ) | ( n21939 & ~n22084 ) | ( n21940 & ~n22084 ) ;
  assign n22090 = ( n21946 & ~n22088 ) | ( n21946 & n22089 ) | ( ~n22088 & n22089 ) ;
  assign n22091 = ( ~n22085 & n22087 ) | ( ~n22085 & n22090 ) | ( n22087 & n22090 ) ;
  assign n22092 = n22080 & ~n22091 ;
  assign n22093 = ~n22080 & n22091 ;
  assign n22094 = n22092 | n22093 ;
  assign n22095 = x102 & n10876 ;
  assign n22096 = x101 & n10871 ;
  assign n22097 = x100 & ~n10870 ;
  assign n22098 = n11305 & n22097 ;
  assign n22099 = n22096 | n22098 ;
  assign n22100 = n22095 | n22099 ;
  assign n22101 = n10879 | n22100 ;
  assign n22102 = ( n5025 & n22100 ) | ( n5025 & n22101 ) | ( n22100 & n22101 ) ;
  assign n22103 = x59 & n22102 ;
  assign n22104 = x59 & ~n22103 ;
  assign n22105 = ( n22102 & ~n22103 ) | ( n22102 & n22104 ) | ( ~n22103 & n22104 ) ;
  assign n22106 = n22094 | n22105 ;
  assign n22107 = n22094 & n22105 ;
  assign n22108 = n22106 & ~n22107 ;
  assign n22109 = ( ~n21947 & n21950 ) | ( ~n21947 & n21965 ) | ( n21950 & n21965 ) ;
  assign n22110 = ~n22108 & n22109 ;
  assign n22111 = n22108 & ~n22109 ;
  assign n22112 = n22110 | n22111 ;
  assign n22113 = x105 & n9853 ;
  assign n22114 = x104 & n9848 ;
  assign n22115 = x103 & ~n9847 ;
  assign n22116 = n10165 & n22115 ;
  assign n22117 = n22114 | n22116 ;
  assign n22118 = n22113 | n22117 ;
  assign n22119 = n9856 | n22118 ;
  assign n22120 = ( n5788 & n22118 ) | ( n5788 & n22119 ) | ( n22118 & n22119 ) ;
  assign n22121 = x56 & n22120 ;
  assign n22122 = x56 & ~n22121 ;
  assign n22123 = ( n22120 & ~n22121 ) | ( n22120 & n22122 ) | ( ~n22121 & n22122 ) ;
  assign n22124 = ~n22112 & n22123 ;
  assign n22125 = n22112 & ~n22123 ;
  assign n22126 = n22124 | n22125 ;
  assign n22127 = n21978 & ~n22126 ;
  assign n22128 = ~n21978 & n22126 ;
  assign n22129 = n22127 | n22128 ;
  assign n22130 = x108 & n8834 ;
  assign n22131 = x107 & n8829 ;
  assign n22132 = x106 & ~n8828 ;
  assign n22133 = n9159 & n22132 ;
  assign n22134 = n22131 | n22133 ;
  assign n22135 = n22130 | n22134 ;
  assign n22136 = n8837 | n22135 ;
  assign n22137 = ( n6358 & n22135 ) | ( n6358 & n22136 ) | ( n22135 & n22136 ) ;
  assign n22138 = x53 & n22137 ;
  assign n22139 = x53 & ~n22138 ;
  assign n22140 = ( n22137 & ~n22138 ) | ( n22137 & n22139 ) | ( ~n22138 & n22139 ) ;
  assign n22141 = ~n22129 & n22140 ;
  assign n22142 = n22129 & ~n22140 ;
  assign n22143 = n22141 | n22142 ;
  assign n22144 = ( ~n21981 & n22069 ) | ( ~n21981 & n22143 ) | ( n22069 & n22143 ) ;
  assign n22145 = ( n21981 & ~n22143 ) | ( n21981 & n22144 ) | ( ~n22143 & n22144 ) ;
  assign n22146 = ( ~n22069 & n22144 ) | ( ~n22069 & n22145 ) | ( n22144 & n22145 ) ;
  assign n22147 = ~n21999 & n22146 ;
  assign n22148 = n21999 & ~n22146 ;
  assign n22149 = n22147 | n22148 ;
  assign n22150 = x114 & n6937 ;
  assign n22151 = x113 & n6932 ;
  assign n22152 = x112 & ~n6931 ;
  assign n22153 = n7216 & n22152 ;
  assign n22154 = n22151 | n22153 ;
  assign n22155 = n22150 | n22154 ;
  assign n22156 = n6940 | n22155 ;
  assign n22157 = ( n8437 & n22155 ) | ( n8437 & n22156 ) | ( n22155 & n22156 ) ;
  assign n22158 = x47 & n22157 ;
  assign n22159 = x47 & ~n22158 ;
  assign n22160 = ( n22157 & ~n22158 ) | ( n22157 & n22159 ) | ( ~n22158 & n22159 ) ;
  assign n22161 = n22149 & ~n22160 ;
  assign n22162 = ~n22149 & n22160 ;
  assign n22163 = n22161 | n22162 ;
  assign n22164 = n22018 & ~n22163 ;
  assign n22165 = n22018 & ~n22164 ;
  assign n22166 = n22018 | n22163 ;
  assign n22167 = x117 & n6068 ;
  assign n22168 = x116 & n6063 ;
  assign n22169 = x115 & ~n6062 ;
  assign n22170 = n6398 & n22169 ;
  assign n22171 = n22168 | n22170 ;
  assign n22172 = n22167 | n22171 ;
  assign n22173 = n6071 | n22172 ;
  assign n22174 = ( n9118 & n22172 ) | ( n9118 & n22173 ) | ( n22172 & n22173 ) ;
  assign n22175 = x44 & n22174 ;
  assign n22176 = x44 & ~n22175 ;
  assign n22177 = ( n22174 & ~n22175 ) | ( n22174 & n22176 ) | ( ~n22175 & n22176 ) ;
  assign n22178 = n22166 & ~n22177 ;
  assign n22179 = ~n22165 & n22178 ;
  assign n22180 = ( n22165 & ~n22166 ) | ( n22165 & n22177 ) | ( ~n22166 & n22177 ) ;
  assign n22181 = n22179 | n22180 ;
  assign n22182 = n22022 & ~n22181 ;
  assign n22183 = ~n22022 & n22181 ;
  assign n22184 = n22182 | n22183 ;
  assign n22185 = x120 & n5340 ;
  assign n22186 = x119 & n5335 ;
  assign n22187 = x118 & ~n5334 ;
  assign n22188 = n5580 & n22187 ;
  assign n22189 = n22186 | n22188 ;
  assign n22190 = n22185 | n22189 ;
  assign n22191 = n5343 | n22190 ;
  assign n22192 = ( n10460 & n22190 ) | ( n10460 & n22191 ) | ( n22190 & n22191 ) ;
  assign n22193 = x41 & n22192 ;
  assign n22194 = x41 & ~n22193 ;
  assign n22195 = ( n22192 & ~n22193 ) | ( n22192 & n22194 ) | ( ~n22193 & n22194 ) ;
  assign n22196 = ~n22184 & n22195 ;
  assign n22197 = n22184 & ~n22195 ;
  assign n22198 = n22196 | n22197 ;
  assign n22199 = ( ~n22024 & n22058 ) | ( ~n22024 & n22198 ) | ( n22058 & n22198 ) ;
  assign n22200 = ( n22024 & ~n22198 ) | ( n22024 & n22199 ) | ( ~n22198 & n22199 ) ;
  assign n22201 = ( ~n22058 & n22199 ) | ( ~n22058 & n22200 ) | ( n22199 & n22200 ) ;
  assign n22202 = ~n22027 & n22201 ;
  assign n22203 = n22027 & ~n22201 ;
  assign n22204 = n22202 | n22203 ;
  assign n22205 = x126 & n3913 ;
  assign n22206 = x125 & n3908 ;
  assign n22207 = x124 & ~n3907 ;
  assign n22208 = n4152 & n22207 ;
  assign n22209 = n22206 | n22208 ;
  assign n22210 = n22205 | n22209 ;
  assign n22211 = n3916 | n22210 ;
  assign n22212 = ( n12687 & n22210 ) | ( n12687 & n22211 ) | ( n22210 & n22211 ) ;
  assign n22213 = x35 & n22212 ;
  assign n22214 = x35 & ~n22213 ;
  assign n22215 = ( n22212 & ~n22213 ) | ( n22212 & n22214 ) | ( ~n22213 & n22214 ) ;
  assign n22216 = n22204 & n22215 ;
  assign n22217 = ( n22027 & ~n22201 ) | ( n22027 & n22215 ) | ( ~n22201 & n22215 ) ;
  assign n22218 = n22202 | n22217 ;
  assign n22219 = ~n22216 & n22218 ;
  assign n22220 = x127 & ~n3308 ;
  assign n22221 = n3570 & n22220 ;
  assign n22222 = ( x127 & n3317 ) | ( x127 & n22221 ) | ( n3317 & n22221 ) ;
  assign n22223 = ( x126 & n22221 ) | ( x126 & n22222 ) | ( n22221 & n22222 ) ;
  assign n22224 = ( n12685 & n22222 ) | ( n12685 & n22223 ) | ( n22222 & n22223 ) ;
  assign n22225 = x32 & n22224 ;
  assign n22226 = x32 & ~n22225 ;
  assign n22227 = ( n22224 & ~n22225 ) | ( n22224 & n22226 ) | ( ~n22225 & n22226 ) ;
  assign n22228 = ( n21862 & n21876 ) | ( n21862 & ~n22029 ) | ( n21876 & ~n22029 ) ;
  assign n22229 = ( n22219 & n22227 ) | ( n22219 & ~n22228 ) | ( n22227 & ~n22228 ) ;
  assign n22230 = ( ~n22227 & n22228 ) | ( ~n22227 & n22229 ) | ( n22228 & n22229 ) ;
  assign n22231 = ( ~n22219 & n22229 ) | ( ~n22219 & n22230 ) | ( n22229 & n22230 ) ;
  assign n22232 = ( n21871 & n21872 ) | ( n21871 & n22035 ) | ( n21872 & n22035 ) ;
  assign n22233 = n22231 & n22232 ;
  assign n22234 = ~n22036 & n22044 ;
  assign n22235 = ~n22231 & n22232 ;
  assign n22236 = n22231 | n22235 ;
  assign n22237 = ~n22233 & n22236 ;
  assign n22238 = n22234 | n22237 ;
  assign n22239 = ~n22036 & n22045 ;
  assign n22240 = n22237 | n22239 ;
  assign n22241 = ( ~n20515 & n22238 ) | ( ~n20515 & n22240 ) | ( n22238 & n22240 ) ;
  assign n22242 = ( ~n20515 & n22234 ) | ( ~n20515 & n22239 ) | ( n22234 & n22239 ) ;
  assign n22243 = ( n22231 & n22232 ) | ( n22231 & n22242 ) | ( n22232 & n22242 ) ;
  assign n22244 = ( n22233 & n22241 ) | ( n22233 & ~n22243 ) | ( n22241 & ~n22243 ) ;
  assign n22245 = x127 & n3913 ;
  assign n22246 = x126 & n3908 ;
  assign n22247 = x125 & ~n3907 ;
  assign n22248 = n4152 & n22247 ;
  assign n22249 = n22246 | n22248 ;
  assign n22250 = n22245 | n22249 ;
  assign n22251 = n3916 | n22250 ;
  assign n22252 = ( n12720 & n22250 ) | ( n12720 & n22251 ) | ( n22250 & n22251 ) ;
  assign n22253 = x35 & n22252 ;
  assign n22254 = x35 & ~n22253 ;
  assign n22255 = ( n22252 & ~n22253 ) | ( n22252 & n22254 ) | ( ~n22253 & n22254 ) ;
  assign n22256 = n22217 & n22255 ;
  assign n22257 = n22217 & ~n22256 ;
  assign n22258 = x124 & n4572 ;
  assign n22259 = x123 & n4567 ;
  assign n22260 = x122 & ~n4566 ;
  assign n22261 = n4828 & n22260 ;
  assign n22262 = n22259 | n22261 ;
  assign n22263 = n22258 | n22262 ;
  assign n22264 = n4575 | n22263 ;
  assign n22265 = ( n11916 & n22263 ) | ( n11916 & n22264 ) | ( n22263 & n22264 ) ;
  assign n22266 = x38 & n22265 ;
  assign n22267 = x38 & ~n22266 ;
  assign n22268 = ( n22265 & ~n22266 ) | ( n22265 & n22267 ) | ( ~n22266 & n22267 ) ;
  assign n22269 = n22164 | n22180 ;
  assign n22270 = n22148 | n22162 ;
  assign n22271 = n22110 | n22124 ;
  assign n22272 = x106 & n9853 ;
  assign n22273 = x105 & n9848 ;
  assign n22274 = x104 & ~n9847 ;
  assign n22275 = n10165 & n22274 ;
  assign n22276 = n22273 | n22275 ;
  assign n22277 = n22272 | n22276 ;
  assign n22278 = n9856 | n22277 ;
  assign n22279 = ( n5814 & n22277 ) | ( n5814 & n22278 ) | ( n22277 & n22278 ) ;
  assign n22280 = x56 & n22279 ;
  assign n22281 = x56 & ~n22280 ;
  assign n22282 = ( n22279 & ~n22280 ) | ( n22279 & n22281 ) | ( ~n22280 & n22281 ) ;
  assign n22283 = x97 & n12808 ;
  assign n22284 = x63 & x96 ;
  assign n22285 = ~n12808 & n22284 ;
  assign n22286 = n22283 | n22285 ;
  assign n22287 = ~x32 & n22286 ;
  assign n22288 = x32 & ~n22286 ;
  assign n22289 = n22287 | n22288 ;
  assign n22290 = n22084 | n22289 ;
  assign n22291 = n22084 & ~n22289 ;
  assign n22292 = ( ~n22084 & n22290 ) | ( ~n22084 & n22291 ) | ( n22290 & n22291 ) ;
  assign n22293 = n22090 & ~n22292 ;
  assign n22294 = n22090 & ~n22293 ;
  assign n22295 = n22090 | n22292 ;
  assign n22296 = ~n22294 & n22295 ;
  assign n22297 = x100 & n11984 ;
  assign n22298 = x99 & n11979 ;
  assign n22299 = x98 & ~n11978 ;
  assign n22300 = n12430 & n22299 ;
  assign n22301 = n22298 | n22300 ;
  assign n22302 = n22297 | n22301 ;
  assign n22303 = n11987 | n22302 ;
  assign n22304 = ( n4532 & n22302 ) | ( n4532 & n22303 ) | ( n22302 & n22303 ) ;
  assign n22305 = x62 & n22304 ;
  assign n22306 = x62 & ~n22305 ;
  assign n22307 = ( n22304 & ~n22305 ) | ( n22304 & n22306 ) | ( ~n22305 & n22306 ) ;
  assign n22308 = n22296 & n22307 ;
  assign n22309 = ( n22294 & ~n22295 ) | ( n22294 & n22307 ) | ( ~n22295 & n22307 ) ;
  assign n22310 = ( n22296 & ~n22308 ) | ( n22296 & n22309 ) | ( ~n22308 & n22309 ) ;
  assign n22311 = x103 & n10876 ;
  assign n22312 = x102 & n10871 ;
  assign n22313 = x101 & ~n10870 ;
  assign n22314 = n11305 & n22313 ;
  assign n22315 = n22312 | n22314 ;
  assign n22316 = n22311 | n22315 ;
  assign n22317 = n10879 | n22316 ;
  assign n22318 = ( n5264 & n22316 ) | ( n5264 & n22317 ) | ( n22316 & n22317 ) ;
  assign n22319 = x59 & n22318 ;
  assign n22320 = x59 & ~n22319 ;
  assign n22321 = ( n22318 & ~n22319 ) | ( n22318 & n22320 ) | ( ~n22319 & n22320 ) ;
  assign n22322 = ~n22310 & n22321 ;
  assign n22323 = n22310 & ~n22321 ;
  assign n22324 = n22322 | n22323 ;
  assign n22325 = ( n22092 & ~n22094 ) | ( n22092 & n22106 ) | ( ~n22094 & n22106 ) ;
  assign n22326 = ~n22324 & n22325 ;
  assign n22327 = n22324 & ~n22325 ;
  assign n22328 = n22326 | n22327 ;
  assign n22329 = n22282 & ~n22328 ;
  assign n22330 = n22328 | n22329 ;
  assign n22331 = ( ~n22282 & n22329 ) | ( ~n22282 & n22330 ) | ( n22329 & n22330 ) ;
  assign n22332 = ~n22271 & n22331 ;
  assign n22333 = n22271 & ~n22331 ;
  assign n22334 = n22332 | n22333 ;
  assign n22335 = x109 & n8834 ;
  assign n22336 = x108 & n8829 ;
  assign n22337 = x107 & ~n8828 ;
  assign n22338 = n9159 & n22337 ;
  assign n22339 = n22336 | n22338 ;
  assign n22340 = n22335 | n22339 ;
  assign n22341 = n8837 | n22340 ;
  assign n22342 = ( n6884 & n22340 ) | ( n6884 & n22341 ) | ( n22340 & n22341 ) ;
  assign n22343 = x53 & n22342 ;
  assign n22344 = x53 & ~n22343 ;
  assign n22345 = ( n22342 & ~n22343 ) | ( n22342 & n22344 ) | ( ~n22343 & n22344 ) ;
  assign n22346 = ~n22334 & n22345 ;
  assign n22347 = n22334 | n22346 ;
  assign n22348 = n22334 & n22345 ;
  assign n22349 = n22127 | n22141 ;
  assign n22350 = n22348 | n22349 ;
  assign n22351 = n22347 & ~n22350 ;
  assign n22352 = ( ~n22347 & n22348 ) | ( ~n22347 & n22349 ) | ( n22348 & n22349 ) ;
  assign n22353 = n22351 | n22352 ;
  assign n22354 = x112 & n7812 ;
  assign n22355 = x111 & n7807 ;
  assign n22356 = x110 & ~n7806 ;
  assign n22357 = n8136 & n22356 ;
  assign n22358 = n22355 | n22357 ;
  assign n22359 = n22354 | n22358 ;
  assign n22360 = n7815 | n22359 ;
  assign n22361 = ( n7789 & n22359 ) | ( n7789 & n22360 ) | ( n22359 & n22360 ) ;
  assign n22362 = x50 & n22361 ;
  assign n22363 = x50 & ~n22362 ;
  assign n22364 = ( n22361 & ~n22362 ) | ( n22361 & n22363 ) | ( ~n22362 & n22363 ) ;
  assign n22365 = ~n22353 & n22364 ;
  assign n22366 = n22353 | n22365 ;
  assign n22367 = n22353 & n22364 ;
  assign n22368 = n22145 | n22367 ;
  assign n22369 = n22366 & ~n22368 ;
  assign n22370 = ( n22145 & ~n22366 ) | ( n22145 & n22367 ) | ( ~n22366 & n22367 ) ;
  assign n22371 = n22369 | n22370 ;
  assign n22372 = x115 & n6937 ;
  assign n22373 = x114 & n6932 ;
  assign n22374 = x113 & ~n6931 ;
  assign n22375 = n7216 & n22374 ;
  assign n22376 = n22373 | n22375 ;
  assign n22377 = n22372 | n22376 ;
  assign n22378 = n6940 | n22377 ;
  assign n22379 = ( n8749 & n22377 ) | ( n8749 & n22378 ) | ( n22377 & n22378 ) ;
  assign n22380 = x47 & n22379 ;
  assign n22381 = x47 & ~n22380 ;
  assign n22382 = ( n22379 & ~n22380 ) | ( n22379 & n22381 ) | ( ~n22380 & n22381 ) ;
  assign n22383 = ~n22371 & n22382 ;
  assign n22384 = n22371 & ~n22382 ;
  assign n22385 = n22383 | n22384 ;
  assign n22386 = n22270 & ~n22385 ;
  assign n22387 = n22270 & ~n22386 ;
  assign n22388 = n22385 | n22386 ;
  assign n22389 = ~n22387 & n22388 ;
  assign n22390 = x118 & n6068 ;
  assign n22391 = x117 & n6063 ;
  assign n22392 = x116 & ~n6062 ;
  assign n22393 = n6398 & n22392 ;
  assign n22394 = n22391 | n22393 ;
  assign n22395 = n22390 | n22394 ;
  assign n22396 = n6071 | n22395 ;
  assign n22397 = ( n9760 & n22395 ) | ( n9760 & n22396 ) | ( n22395 & n22396 ) ;
  assign n22398 = x44 & n22397 ;
  assign n22399 = x44 & ~n22398 ;
  assign n22400 = ( n22397 & ~n22398 ) | ( n22397 & n22399 ) | ( ~n22398 & n22399 ) ;
  assign n22401 = n22389 & ~n22400 ;
  assign n22402 = ~n22389 & n22400 ;
  assign n22403 = n22401 | n22402 ;
  assign n22404 = n22269 & ~n22403 ;
  assign n22405 = ~n22269 & n22403 ;
  assign n22406 = n22404 | n22405 ;
  assign n22407 = x121 & n5340 ;
  assign n22408 = x120 & n5335 ;
  assign n22409 = x119 & ~n5334 ;
  assign n22410 = n5580 & n22409 ;
  assign n22411 = n22408 | n22410 ;
  assign n22412 = n22407 | n22411 ;
  assign n22413 = n5343 | n22412 ;
  assign n22414 = ( n10811 & n22412 ) | ( n10811 & n22413 ) | ( n22412 & n22413 ) ;
  assign n22415 = x41 & n22414 ;
  assign n22416 = x41 & ~n22415 ;
  assign n22417 = ( n22414 & ~n22415 ) | ( n22414 & n22416 ) | ( ~n22415 & n22416 ) ;
  assign n22418 = ~n22406 & n22417 ;
  assign n22419 = n22406 | n22418 ;
  assign n22420 = n22406 & n22417 ;
  assign n22421 = n22182 | n22196 ;
  assign n22422 = n22420 | n22421 ;
  assign n22423 = n22419 & ~n22422 ;
  assign n22424 = ( ~n22419 & n22420 ) | ( ~n22419 & n22421 ) | ( n22420 & n22421 ) ;
  assign n22425 = n22423 | n22424 ;
  assign n22426 = n22268 & ~n22425 ;
  assign n22427 = n22425 | n22426 ;
  assign n22428 = ( ~n22268 & n22426 ) | ( ~n22268 & n22427 ) | ( n22426 & n22427 ) ;
  assign n22429 = ~n22200 & n22428 ;
  assign n22430 = n22200 & ~n22428 ;
  assign n22431 = n22429 | n22430 ;
  assign n22432 = ~n22217 & n22255 ;
  assign n22433 = n22431 & ~n22432 ;
  assign n22434 = ~n22257 & n22433 ;
  assign n22435 = ( n22257 & ~n22431 ) | ( n22257 & n22432 ) | ( ~n22431 & n22432 ) ;
  assign n22436 = n22434 | n22435 ;
  assign n22437 = ( ~n22219 & n22227 ) | ( ~n22219 & n22228 ) | ( n22227 & n22228 ) ;
  assign n22438 = ~n22436 & n22437 ;
  assign n22439 = n22436 & ~n22437 ;
  assign n22440 = n22438 | n22439 ;
  assign n22441 = ~n22235 & n22238 ;
  assign n22442 = ~n22235 & n22240 ;
  assign n22443 = ( ~n20515 & n22441 ) | ( ~n20515 & n22442 ) | ( n22441 & n22442 ) ;
  assign n22444 = n22440 & n22443 ;
  assign n22445 = n22440 | n22441 ;
  assign n22446 = n22440 | n22442 ;
  assign n22447 = ( ~n20515 & n22445 ) | ( ~n20515 & n22446 ) | ( n22445 & n22446 ) ;
  assign n22448 = ~n22444 & n22447 ;
  assign n22449 = ~n22438 & n22445 ;
  assign n22450 = ~n22438 & n22446 ;
  assign n22451 = ( ~n20515 & n22449 ) | ( ~n20515 & n22450 ) | ( n22449 & n22450 ) ;
  assign n22452 = n22256 | n22435 ;
  assign n22453 = x125 & n4572 ;
  assign n22454 = x124 & n4567 ;
  assign n22455 = x123 & ~n4566 ;
  assign n22456 = n4828 & n22455 ;
  assign n22457 = n22454 | n22456 ;
  assign n22458 = n22453 | n22457 ;
  assign n22459 = n4575 | n22458 ;
  assign n22460 = ( n12310 & n22458 ) | ( n12310 & n22459 ) | ( n22458 & n22459 ) ;
  assign n22461 = x38 & n22460 ;
  assign n22462 = x38 & ~n22461 ;
  assign n22463 = ( n22460 & ~n22461 ) | ( n22460 & n22462 ) | ( ~n22461 & n22462 ) ;
  assign n22464 = x127 & n3908 ;
  assign n22465 = x126 & ~n3907 ;
  assign n22466 = n4152 & n22465 ;
  assign n22467 = n22464 | n22466 ;
  assign n22468 = n3916 | n22467 ;
  assign n22469 = ( n13461 & n22467 ) | ( n13461 & n22468 ) | ( n22467 & n22468 ) ;
  assign n22470 = x35 & n22469 ;
  assign n22471 = x35 & ~n22470 ;
  assign n22472 = ( n22469 & ~n22470 ) | ( n22469 & n22471 ) | ( ~n22470 & n22471 ) ;
  assign n22473 = n22426 | n22430 ;
  assign n22474 = n22472 & n22473 ;
  assign n22475 = n22472 | n22473 ;
  assign n22476 = ~n22474 & n22475 ;
  assign n22477 = n22418 | n22424 ;
  assign n22478 = x122 & n5340 ;
  assign n22479 = x121 & n5335 ;
  assign n22480 = x120 & ~n5334 ;
  assign n22481 = n5580 & n22480 ;
  assign n22482 = n22479 | n22481 ;
  assign n22483 = n22478 | n22482 ;
  assign n22484 = n5343 | n22483 ;
  assign n22485 = ( n11188 & n22483 ) | ( n11188 & n22484 ) | ( n22483 & n22484 ) ;
  assign n22486 = x41 & n22485 ;
  assign n22487 = x41 & ~n22486 ;
  assign n22488 = ( n22485 & ~n22486 ) | ( n22485 & n22487 ) | ( ~n22486 & n22487 ) ;
  assign n22489 = n22383 | n22386 ;
  assign n22490 = n22329 | n22333 ;
  assign n22491 = x107 & n9853 ;
  assign n22492 = x106 & n9848 ;
  assign n22493 = x105 & ~n9847 ;
  assign n22494 = n10165 & n22493 ;
  assign n22495 = n22492 | n22494 ;
  assign n22496 = n22491 | n22495 ;
  assign n22497 = n9856 | n22496 ;
  assign n22498 = ( n6328 & n22496 ) | ( n6328 & n22497 ) | ( n22496 & n22497 ) ;
  assign n22499 = x56 & n22498 ;
  assign n22500 = x56 & ~n22499 ;
  assign n22501 = ( n22498 & ~n22499 ) | ( n22498 & n22500 ) | ( ~n22499 & n22500 ) ;
  assign n22502 = n22322 | n22326 ;
  assign n22503 = x101 & n11984 ;
  assign n22504 = x100 & n11979 ;
  assign n22505 = x99 & ~n11978 ;
  assign n22506 = n12430 & n22505 ;
  assign n22507 = n22504 | n22506 ;
  assign n22508 = n22503 | n22507 ;
  assign n22509 = n11987 | n22508 ;
  assign n22510 = ( n4783 & n22508 ) | ( n4783 & n22509 ) | ( n22508 & n22509 ) ;
  assign n22511 = ~x62 & n22510 ;
  assign n22512 = x98 & n12808 ;
  assign n22513 = x63 & x97 ;
  assign n22514 = ~n12808 & n22513 ;
  assign n22515 = n22512 | n22514 ;
  assign n22516 = n22287 | n22291 ;
  assign n22517 = n22515 & ~n22516 ;
  assign n22518 = ~n22515 & n22516 ;
  assign n22519 = n22517 | n22518 ;
  assign n22520 = x62 & ~n22510 ;
  assign n22521 = n22519 & ~n22520 ;
  assign n22522 = ~n22511 & n22521 ;
  assign n22523 = ( n22511 & ~n22519 ) | ( n22511 & n22520 ) | ( ~n22519 & n22520 ) ;
  assign n22524 = n22522 | n22523 ;
  assign n22525 = n22293 | n22309 ;
  assign n22526 = x104 & n10876 ;
  assign n22527 = x103 & n10871 ;
  assign n22528 = x102 & ~n10870 ;
  assign n22529 = n11305 & n22528 ;
  assign n22530 = n22527 | n22529 ;
  assign n22531 = n22526 | n22530 ;
  assign n22532 = n10879 | n22531 ;
  assign n22533 = ( n5295 & n22531 ) | ( n5295 & n22532 ) | ( n22531 & n22532 ) ;
  assign n22534 = x59 & n22533 ;
  assign n22535 = x59 & ~n22534 ;
  assign n22536 = ( n22533 & ~n22534 ) | ( n22533 & n22535 ) | ( ~n22534 & n22535 ) ;
  assign n22537 = ( n22524 & ~n22525 ) | ( n22524 & n22536 ) | ( ~n22525 & n22536 ) ;
  assign n22538 = ( n22525 & ~n22536 ) | ( n22525 & n22537 ) | ( ~n22536 & n22537 ) ;
  assign n22539 = ( ~n22524 & n22537 ) | ( ~n22524 & n22538 ) | ( n22537 & n22538 ) ;
  assign n22540 = ( n22501 & n22502 ) | ( n22501 & ~n22539 ) | ( n22502 & ~n22539 ) ;
  assign n22541 = ( ~n22502 & n22539 ) | ( ~n22502 & n22540 ) | ( n22539 & n22540 ) ;
  assign n22542 = ( ~n22501 & n22540 ) | ( ~n22501 & n22541 ) | ( n22540 & n22541 ) ;
  assign n22543 = ~n22490 & n22542 ;
  assign n22544 = n22490 & ~n22542 ;
  assign n22545 = n22543 | n22544 ;
  assign n22546 = x110 & n8834 ;
  assign n22547 = x109 & n8829 ;
  assign n22548 = x108 & ~n8828 ;
  assign n22549 = n9159 & n22548 ;
  assign n22550 = n22547 | n22549 ;
  assign n22551 = n22546 | n22550 ;
  assign n22552 = n8837 | n22551 ;
  assign n22553 = ( n7189 & n22551 ) | ( n7189 & n22552 ) | ( n22551 & n22552 ) ;
  assign n22554 = x53 & n22553 ;
  assign n22555 = x53 & ~n22554 ;
  assign n22556 = ( n22553 & ~n22554 ) | ( n22553 & n22555 ) | ( ~n22554 & n22555 ) ;
  assign n22557 = n22545 & n22556 ;
  assign n22558 = ( n22490 & ~n22542 ) | ( n22490 & n22556 ) | ( ~n22542 & n22556 ) ;
  assign n22559 = n22543 | n22558 ;
  assign n22560 = ~n22557 & n22559 ;
  assign n22561 = n22346 | n22352 ;
  assign n22562 = n22560 & ~n22561 ;
  assign n22563 = x113 & n7812 ;
  assign n22564 = x112 & n7807 ;
  assign n22565 = x111 & ~n7806 ;
  assign n22566 = n8136 & n22565 ;
  assign n22567 = n22564 | n22566 ;
  assign n22568 = n22563 | n22567 ;
  assign n22569 = n7815 | n22568 ;
  assign n22570 = ( n8113 & n22568 ) | ( n8113 & n22569 ) | ( n22568 & n22569 ) ;
  assign n22571 = x50 & n22570 ;
  assign n22572 = x50 & ~n22571 ;
  assign n22573 = ( n22570 & ~n22571 ) | ( n22570 & n22572 ) | ( ~n22571 & n22572 ) ;
  assign n22574 = ( ~n22560 & n22561 ) | ( ~n22560 & n22573 ) | ( n22561 & n22573 ) ;
  assign n22575 = n22562 | n22574 ;
  assign n22576 = n22365 | n22370 ;
  assign n22577 = ~n22560 & n22561 ;
  assign n22578 = n22562 | n22577 ;
  assign n22579 = n22573 & n22578 ;
  assign n22580 = n22576 | n22579 ;
  assign n22581 = n22575 & ~n22580 ;
  assign n22582 = ( ~n22575 & n22576 ) | ( ~n22575 & n22579 ) | ( n22576 & n22579 ) ;
  assign n22583 = n22581 | n22582 ;
  assign n22584 = x116 & n6937 ;
  assign n22585 = x115 & n6932 ;
  assign n22586 = x114 & ~n6931 ;
  assign n22587 = n7216 & n22586 ;
  assign n22588 = n22585 | n22587 ;
  assign n22589 = n22584 | n22588 ;
  assign n22590 = n6940 | n22589 ;
  assign n22591 = ( n8778 & n22589 ) | ( n8778 & n22590 ) | ( n22589 & n22590 ) ;
  assign n22592 = x47 & n22591 ;
  assign n22593 = x47 & ~n22592 ;
  assign n22594 = ( n22591 & ~n22592 ) | ( n22591 & n22593 ) | ( ~n22592 & n22593 ) ;
  assign n22595 = ( n22489 & n22583 ) | ( n22489 & ~n22594 ) | ( n22583 & ~n22594 ) ;
  assign n22596 = ( ~n22583 & n22594 ) | ( ~n22583 & n22595 ) | ( n22594 & n22595 ) ;
  assign n22597 = ( ~n22489 & n22595 ) | ( ~n22489 & n22596 ) | ( n22595 & n22596 ) ;
  assign n22598 = x119 & n6068 ;
  assign n22599 = x118 & n6063 ;
  assign n22600 = x117 & ~n6062 ;
  assign n22601 = n6398 & n22600 ;
  assign n22602 = n22599 | n22601 ;
  assign n22603 = n22598 | n22602 ;
  assign n22604 = n6071 | n22603 ;
  assign n22605 = ( n9789 & n22603 ) | ( n9789 & n22604 ) | ( n22603 & n22604 ) ;
  assign n22606 = x44 & n22605 ;
  assign n22607 = x44 & ~n22606 ;
  assign n22608 = ( n22605 & ~n22606 ) | ( n22605 & n22607 ) | ( ~n22606 & n22607 ) ;
  assign n22609 = ~n22597 & n22608 ;
  assign n22610 = n22597 & ~n22608 ;
  assign n22611 = n22609 | n22610 ;
  assign n22612 = n22402 | n22404 ;
  assign n22613 = ( n22488 & n22611 ) | ( n22488 & ~n22612 ) | ( n22611 & ~n22612 ) ;
  assign n22614 = ( ~n22611 & n22612 ) | ( ~n22611 & n22613 ) | ( n22612 & n22613 ) ;
  assign n22615 = ( ~n22488 & n22613 ) | ( ~n22488 & n22614 ) | ( n22613 & n22614 ) ;
  assign n22616 = ~n22477 & n22615 ;
  assign n22617 = n22477 & ~n22615 ;
  assign n22618 = n22616 | n22617 ;
  assign n22619 = ( n22463 & n22476 ) | ( n22463 & ~n22618 ) | ( n22476 & ~n22618 ) ;
  assign n22620 = ( ~n22476 & n22618 ) | ( ~n22476 & n22619 ) | ( n22618 & n22619 ) ;
  assign n22621 = ( ~n22463 & n22619 ) | ( ~n22463 & n22620 ) | ( n22619 & n22620 ) ;
  assign n22622 = n22452 & ~n22621 ;
  assign n22623 = ~n22452 & n22621 ;
  assign n22624 = n22622 | n22623 ;
  assign n22625 = n22451 & n22624 ;
  assign n22626 = n22449 | n22624 ;
  assign n22627 = n22450 | n22624 ;
  assign n22628 = ( ~n20515 & n22626 ) | ( ~n20515 & n22627 ) | ( n22626 & n22627 ) ;
  assign n22629 = ~n22625 & n22628 ;
  assign n22630 = ~n22583 & n22594 ;
  assign n22631 = n22582 | n22630 ;
  assign n22632 = x111 & n8834 ;
  assign n22633 = x110 & n8829 ;
  assign n22634 = x109 & ~n8828 ;
  assign n22635 = n9159 & n22634 ;
  assign n22636 = n22633 | n22635 ;
  assign n22637 = n22632 | n22636 ;
  assign n22638 = n8837 | n22637 ;
  assign n22639 = ( n7492 & n22637 ) | ( n7492 & n22638 ) | ( n22637 & n22638 ) ;
  assign n22640 = x53 & n22639 ;
  assign n22641 = x53 & ~n22640 ;
  assign n22642 = ( n22639 & ~n22640 ) | ( n22639 & n22641 ) | ( ~n22640 & n22641 ) ;
  assign n22643 = x102 & n11984 ;
  assign n22644 = x101 & n11979 ;
  assign n22645 = x100 & ~n11978 ;
  assign n22646 = n12430 & n22645 ;
  assign n22647 = n22644 | n22646 ;
  assign n22648 = n22643 | n22647 ;
  assign n22649 = n11987 | n22648 ;
  assign n22650 = ( n5025 & n22648 ) | ( n5025 & n22649 ) | ( n22648 & n22649 ) ;
  assign n22651 = x62 & n22650 ;
  assign n22652 = x62 & ~n22651 ;
  assign n22653 = ( n22650 & ~n22651 ) | ( n22650 & n22652 ) | ( ~n22651 & n22652 ) ;
  assign n22654 = x99 & n12808 ;
  assign n22655 = x63 & x98 ;
  assign n22656 = ~n12808 & n22655 ;
  assign n22657 = n22654 | n22656 ;
  assign n22658 = ( n22515 & n22523 ) | ( n22515 & n22657 ) | ( n22523 & n22657 ) ;
  assign n22659 = n22515 | n22516 ;
  assign n22660 = ( n22523 & n22657 ) | ( n22523 & ~n22659 ) | ( n22657 & ~n22659 ) ;
  assign n22661 = ~n22515 & n22657 ;
  assign n22662 = ( n22516 & n22517 ) | ( n22516 & ~n22657 ) | ( n22517 & ~n22657 ) ;
  assign n22663 = ( n22523 & ~n22661 ) | ( n22523 & n22662 ) | ( ~n22661 & n22662 ) ;
  assign n22664 = ( ~n22658 & n22660 ) | ( ~n22658 & n22663 ) | ( n22660 & n22663 ) ;
  assign n22665 = n22653 & ~n22664 ;
  assign n22666 = ~n22653 & n22664 ;
  assign n22667 = n22665 | n22666 ;
  assign n22668 = x105 & n10876 ;
  assign n22669 = x104 & n10871 ;
  assign n22670 = x103 & ~n10870 ;
  assign n22671 = n11305 & n22670 ;
  assign n22672 = n22669 | n22671 ;
  assign n22673 = n22668 | n22672 ;
  assign n22674 = n10879 | n22673 ;
  assign n22675 = ( n5788 & n22673 ) | ( n5788 & n22674 ) | ( n22673 & n22674 ) ;
  assign n22676 = x59 & n22675 ;
  assign n22677 = x59 & ~n22676 ;
  assign n22678 = ( n22675 & ~n22676 ) | ( n22675 & n22677 ) | ( ~n22676 & n22677 ) ;
  assign n22679 = n22667 | n22678 ;
  assign n22680 = n22667 & n22678 ;
  assign n22681 = n22679 & ~n22680 ;
  assign n22682 = ( n22525 & n22536 ) | ( n22525 & n22539 ) | ( n22536 & n22539 ) ;
  assign n22683 = ~n22681 & n22682 ;
  assign n22684 = n22681 & ~n22682 ;
  assign n22685 = n22683 | n22684 ;
  assign n22686 = x108 & n9853 ;
  assign n22687 = x107 & n9848 ;
  assign n22688 = x106 & ~n9847 ;
  assign n22689 = n10165 & n22688 ;
  assign n22690 = n22687 | n22689 ;
  assign n22691 = n22686 | n22690 ;
  assign n22692 = n9856 | n22691 ;
  assign n22693 = ( n6358 & n22691 ) | ( n6358 & n22692 ) | ( n22691 & n22692 ) ;
  assign n22694 = x56 & n22693 ;
  assign n22695 = x56 & ~n22694 ;
  assign n22696 = ( n22693 & ~n22694 ) | ( n22693 & n22695 ) | ( ~n22694 & n22695 ) ;
  assign n22697 = ~n22685 & n22696 ;
  assign n22698 = n22685 & ~n22696 ;
  assign n22699 = n22697 | n22698 ;
  assign n22700 = ( ~n22540 & n22642 ) | ( ~n22540 & n22699 ) | ( n22642 & n22699 ) ;
  assign n22701 = ( n22540 & ~n22699 ) | ( n22540 & n22700 ) | ( ~n22699 & n22700 ) ;
  assign n22702 = ( ~n22642 & n22700 ) | ( ~n22642 & n22701 ) | ( n22700 & n22701 ) ;
  assign n22703 = ~n22558 & n22702 ;
  assign n22704 = n22558 & ~n22702 ;
  assign n22705 = n22703 | n22704 ;
  assign n22706 = x114 & n7812 ;
  assign n22707 = x113 & n7807 ;
  assign n22708 = x112 & ~n7806 ;
  assign n22709 = n8136 & n22708 ;
  assign n22710 = n22707 | n22709 ;
  assign n22711 = n22706 | n22710 ;
  assign n22712 = n7815 | n22711 ;
  assign n22713 = ( n8437 & n22711 ) | ( n8437 & n22712 ) | ( n22711 & n22712 ) ;
  assign n22714 = x50 & n22713 ;
  assign n22715 = x50 & ~n22714 ;
  assign n22716 = ( n22713 & ~n22714 ) | ( n22713 & n22715 ) | ( ~n22714 & n22715 ) ;
  assign n22717 = n22705 & ~n22716 ;
  assign n22718 = ~n22705 & n22716 ;
  assign n22719 = n22717 | n22718 ;
  assign n22720 = x117 & n6937 ;
  assign n22721 = x116 & n6932 ;
  assign n22722 = x115 & ~n6931 ;
  assign n22723 = n7216 & n22722 ;
  assign n22724 = n22721 | n22723 ;
  assign n22725 = n22720 | n22724 ;
  assign n22726 = n6940 | n22725 ;
  assign n22727 = ( n9118 & n22725 ) | ( n9118 & n22726 ) | ( n22725 & n22726 ) ;
  assign n22728 = x47 & n22727 ;
  assign n22729 = x47 & ~n22728 ;
  assign n22730 = ( n22727 & ~n22728 ) | ( n22727 & n22729 ) | ( ~n22728 & n22729 ) ;
  assign n22731 = ( n22574 & ~n22719 ) | ( n22574 & n22730 ) | ( ~n22719 & n22730 ) ;
  assign n22732 = ( n22719 & ~n22730 ) | ( n22719 & n22731 ) | ( ~n22730 & n22731 ) ;
  assign n22733 = ( ~n22574 & n22731 ) | ( ~n22574 & n22732 ) | ( n22731 & n22732 ) ;
  assign n22734 = n22631 & ~n22733 ;
  assign n22735 = ~n22631 & n22733 ;
  assign n22736 = n22734 | n22735 ;
  assign n22737 = x120 & n6068 ;
  assign n22738 = x119 & n6063 ;
  assign n22739 = x118 & ~n6062 ;
  assign n22740 = n6398 & n22739 ;
  assign n22741 = n22738 | n22740 ;
  assign n22742 = n22737 | n22741 ;
  assign n22743 = n6071 | n22742 ;
  assign n22744 = ( n10460 & n22742 ) | ( n10460 & n22743 ) | ( n22742 & n22743 ) ;
  assign n22745 = x44 & n22744 ;
  assign n22746 = x44 & ~n22745 ;
  assign n22747 = ( n22744 & ~n22745 ) | ( n22744 & n22746 ) | ( ~n22745 & n22746 ) ;
  assign n22748 = ~n22736 & n22747 ;
  assign n22749 = n22736 & ~n22747 ;
  assign n22750 = n22748 | n22749 ;
  assign n22751 = ( n22489 & n22608 ) | ( n22489 & n22611 ) | ( n22608 & n22611 ) ;
  assign n22752 = ~n22750 & n22751 ;
  assign n22753 = n22750 & ~n22751 ;
  assign n22754 = n22752 | n22753 ;
  assign n22755 = x123 & n5340 ;
  assign n22756 = x122 & n5335 ;
  assign n22757 = x121 & ~n5334 ;
  assign n22758 = n5580 & n22757 ;
  assign n22759 = n22756 | n22758 ;
  assign n22760 = n22755 | n22759 ;
  assign n22761 = n5343 | n22760 ;
  assign n22762 = ( n11219 & n22760 ) | ( n11219 & n22761 ) | ( n22760 & n22761 ) ;
  assign n22763 = x41 & n22762 ;
  assign n22764 = x41 & ~n22763 ;
  assign n22765 = ( n22762 & ~n22763 ) | ( n22762 & n22764 ) | ( ~n22763 & n22764 ) ;
  assign n22766 = ( n22614 & n22754 ) | ( n22614 & ~n22765 ) | ( n22754 & ~n22765 ) ;
  assign n22767 = ( ~n22754 & n22765 ) | ( ~n22754 & n22766 ) | ( n22765 & n22766 ) ;
  assign n22768 = ( ~n22614 & n22766 ) | ( ~n22614 & n22767 ) | ( n22766 & n22767 ) ;
  assign n22769 = x126 & n4572 ;
  assign n22770 = x125 & n4567 ;
  assign n22771 = x124 & ~n4566 ;
  assign n22772 = n4828 & n22771 ;
  assign n22773 = n22770 | n22772 ;
  assign n22774 = n22769 | n22773 ;
  assign n22775 = n4575 | n22774 ;
  assign n22776 = ( n12687 & n22774 ) | ( n12687 & n22775 ) | ( n22774 & n22775 ) ;
  assign n22777 = x38 & n22776 ;
  assign n22778 = x38 & ~n22777 ;
  assign n22779 = ( n22776 & ~n22777 ) | ( n22776 & n22778 ) | ( ~n22777 & n22778 ) ;
  assign n22780 = n22768 | n22779 ;
  assign n22781 = ~n22779 & n22780 ;
  assign n22782 = ( ~n22768 & n22780 ) | ( ~n22768 & n22781 ) | ( n22780 & n22781 ) ;
  assign n22783 = x127 & ~n3907 ;
  assign n22784 = n4152 & n22783 ;
  assign n22785 = ( x127 & n3916 ) | ( x127 & n22784 ) | ( n3916 & n22784 ) ;
  assign n22786 = ( x126 & n22784 ) | ( x126 & n22785 ) | ( n22784 & n22785 ) ;
  assign n22787 = ( n12685 & n22785 ) | ( n12685 & n22786 ) | ( n22785 & n22786 ) ;
  assign n22788 = x35 & n22787 ;
  assign n22789 = x35 & ~n22788 ;
  assign n22790 = ( n22787 & ~n22788 ) | ( n22787 & n22789 ) | ( ~n22788 & n22789 ) ;
  assign n22791 = ( n22463 & n22477 ) | ( n22463 & ~n22615 ) | ( n22477 & ~n22615 ) ;
  assign n22792 = ( n22782 & n22790 ) | ( n22782 & ~n22791 ) | ( n22790 & ~n22791 ) ;
  assign n22793 = ( ~n22790 & n22791 ) | ( ~n22790 & n22792 ) | ( n22791 & n22792 ) ;
  assign n22794 = ( ~n22782 & n22792 ) | ( ~n22782 & n22793 ) | ( n22792 & n22793 ) ;
  assign n22795 = ( n22472 & n22473 ) | ( n22472 & n22621 ) | ( n22473 & n22621 ) ;
  assign n22796 = ~n22794 & n22795 ;
  assign n22797 = n22794 & ~n22795 ;
  assign n22798 = n22796 | n22797 ;
  assign n22799 = ~n22622 & n22626 ;
  assign n22800 = ~n22622 & n22627 ;
  assign n22801 = ( ~n20515 & n22799 ) | ( ~n20515 & n22800 ) | ( n22799 & n22800 ) ;
  assign n22802 = n22798 & n22801 ;
  assign n22803 = n22798 | n22799 ;
  assign n22804 = n22798 | n22800 ;
  assign n22805 = ( ~n20515 & n22803 ) | ( ~n20515 & n22804 ) | ( n22803 & n22804 ) ;
  assign n22806 = ~n22802 & n22805 ;
  assign n22807 = n22734 | n22748 ;
  assign n22808 = x121 & n6068 ;
  assign n22809 = x120 & n6063 ;
  assign n22810 = x119 & ~n6062 ;
  assign n22811 = n6398 & n22810 ;
  assign n22812 = n22809 | n22811 ;
  assign n22813 = n22808 | n22812 ;
  assign n22814 = n6071 | n22813 ;
  assign n22815 = ( n10811 & n22813 ) | ( n10811 & n22814 ) | ( n22813 & n22814 ) ;
  assign n22816 = x44 & n22815 ;
  assign n22817 = x44 & ~n22816 ;
  assign n22818 = ( n22815 & ~n22816 ) | ( n22815 & n22817 ) | ( ~n22816 & n22817 ) ;
  assign n22819 = x109 & n9853 ;
  assign n22820 = x108 & n9848 ;
  assign n22821 = x107 & ~n9847 ;
  assign n22822 = n10165 & n22821 ;
  assign n22823 = n22820 | n22822 ;
  assign n22824 = n22819 | n22823 ;
  assign n22825 = n9856 | n22824 ;
  assign n22826 = ( n6884 & n22824 ) | ( n6884 & n22825 ) | ( n22824 & n22825 ) ;
  assign n22827 = x56 & n22826 ;
  assign n22828 = x56 & ~n22827 ;
  assign n22829 = ( n22826 & ~n22827 ) | ( n22826 & n22828 ) | ( ~n22827 & n22828 ) ;
  assign n22830 = ( n22665 & ~n22667 ) | ( n22665 & n22679 ) | ( ~n22667 & n22679 ) ;
  assign n22831 = x100 & n12808 ;
  assign n22832 = x63 & x99 ;
  assign n22833 = ~n12808 & n22832 ;
  assign n22834 = n22831 | n22833 ;
  assign n22835 = ( x35 & ~n22657 ) | ( x35 & n22834 ) | ( ~n22657 & n22834 ) ;
  assign n22836 = ( ~x35 & n22657 ) | ( ~x35 & n22834 ) | ( n22657 & n22834 ) ;
  assign n22837 = ( ~n22834 & n22835 ) | ( ~n22834 & n22836 ) | ( n22835 & n22836 ) ;
  assign n22838 = n22663 & ~n22837 ;
  assign n22839 = ~n22663 & n22837 ;
  assign n22840 = n22838 | n22839 ;
  assign n22841 = x103 & n11984 ;
  assign n22842 = x102 & n11979 ;
  assign n22843 = x101 & ~n11978 ;
  assign n22844 = n12430 & n22843 ;
  assign n22845 = n22842 | n22844 ;
  assign n22846 = n22841 | n22845 ;
  assign n22847 = n11987 | n22846 ;
  assign n22848 = ( n5264 & n22846 ) | ( n5264 & n22847 ) | ( n22846 & n22847 ) ;
  assign n22849 = x62 & n22848 ;
  assign n22850 = x62 & ~n22849 ;
  assign n22851 = ( n22848 & ~n22849 ) | ( n22848 & n22850 ) | ( ~n22849 & n22850 ) ;
  assign n22852 = n22840 & ~n22851 ;
  assign n22853 = ~n22840 & n22851 ;
  assign n22854 = n22852 | n22853 ;
  assign n22855 = x106 & n10876 ;
  assign n22856 = x105 & n10871 ;
  assign n22857 = x104 & ~n10870 ;
  assign n22858 = n11305 & n22857 ;
  assign n22859 = n22856 | n22858 ;
  assign n22860 = n22855 | n22859 ;
  assign n22861 = n10879 | n22860 ;
  assign n22862 = ( n5814 & n22860 ) | ( n5814 & n22861 ) | ( n22860 & n22861 ) ;
  assign n22863 = x59 & n22862 ;
  assign n22864 = x59 & ~n22863 ;
  assign n22865 = ( n22862 & ~n22863 ) | ( n22862 & n22864 ) | ( ~n22863 & n22864 ) ;
  assign n22866 = ( n22830 & n22854 ) | ( n22830 & ~n22865 ) | ( n22854 & ~n22865 ) ;
  assign n22867 = ( ~n22854 & n22865 ) | ( ~n22854 & n22866 ) | ( n22865 & n22866 ) ;
  assign n22868 = ( ~n22830 & n22866 ) | ( ~n22830 & n22867 ) | ( n22866 & n22867 ) ;
  assign n22869 = n22829 & ~n22868 ;
  assign n22870 = ~n22829 & n22868 ;
  assign n22871 = n22869 | n22870 ;
  assign n22872 = n22683 | n22697 ;
  assign n22873 = n22871 & ~n22872 ;
  assign n22874 = ~n22871 & n22872 ;
  assign n22875 = n22873 | n22874 ;
  assign n22876 = x112 & n8834 ;
  assign n22877 = x111 & n8829 ;
  assign n22878 = x110 & ~n8828 ;
  assign n22879 = n9159 & n22878 ;
  assign n22880 = n22877 | n22879 ;
  assign n22881 = n22876 | n22880 ;
  assign n22882 = n8837 | n22881 ;
  assign n22883 = ( n7789 & n22881 ) | ( n7789 & n22882 ) | ( n22881 & n22882 ) ;
  assign n22884 = x53 & n22883 ;
  assign n22885 = x53 & ~n22884 ;
  assign n22886 = ( n22883 & ~n22884 ) | ( n22883 & n22885 ) | ( ~n22884 & n22885 ) ;
  assign n22887 = ~n22875 & n22886 ;
  assign n22888 = n22875 | n22887 ;
  assign n22889 = n22875 & n22886 ;
  assign n22890 = n22701 | n22889 ;
  assign n22891 = n22888 & ~n22890 ;
  assign n22892 = ( n22701 & ~n22888 ) | ( n22701 & n22889 ) | ( ~n22888 & n22889 ) ;
  assign n22893 = n22891 | n22892 ;
  assign n22894 = x115 & n7812 ;
  assign n22895 = x114 & n7807 ;
  assign n22896 = x113 & ~n7806 ;
  assign n22897 = n8136 & n22896 ;
  assign n22898 = n22895 | n22897 ;
  assign n22899 = n22894 | n22898 ;
  assign n22900 = n7815 | n22899 ;
  assign n22901 = ( n8749 & n22899 ) | ( n8749 & n22900 ) | ( n22899 & n22900 ) ;
  assign n22902 = x50 & n22901 ;
  assign n22903 = x50 & ~n22902 ;
  assign n22904 = ( n22901 & ~n22902 ) | ( n22901 & n22903 ) | ( ~n22902 & n22903 ) ;
  assign n22905 = n22893 & ~n22904 ;
  assign n22906 = ~n22893 & n22904 ;
  assign n22907 = n22905 | n22906 ;
  assign n22908 = n22704 | n22718 ;
  assign n22909 = ~n22907 & n22908 ;
  assign n22910 = n22907 & ~n22908 ;
  assign n22911 = n22909 | n22910 ;
  assign n22912 = x118 & n6937 ;
  assign n22913 = x117 & n6932 ;
  assign n22914 = x116 & ~n6931 ;
  assign n22915 = n7216 & n22914 ;
  assign n22916 = n22913 | n22915 ;
  assign n22917 = n22912 | n22916 ;
  assign n22918 = n6940 | n22917 ;
  assign n22919 = ( n9760 & n22917 ) | ( n9760 & n22918 ) | ( n22917 & n22918 ) ;
  assign n22920 = x47 & n22919 ;
  assign n22921 = x47 & ~n22920 ;
  assign n22922 = ( n22919 & ~n22920 ) | ( n22919 & n22921 ) | ( ~n22920 & n22921 ) ;
  assign n22923 = ~n22911 & n22922 ;
  assign n22924 = n22911 & ~n22922 ;
  assign n22925 = n22923 | n22924 ;
  assign n22926 = n22731 & ~n22925 ;
  assign n22927 = ~n22731 & n22925 ;
  assign n22928 = n22926 | n22927 ;
  assign n22929 = n22818 & ~n22928 ;
  assign n22930 = n22928 | n22929 ;
  assign n22931 = ( ~n22818 & n22929 ) | ( ~n22818 & n22930 ) | ( n22929 & n22930 ) ;
  assign n22932 = ~n22807 & n22931 ;
  assign n22933 = n22807 & ~n22931 ;
  assign n22934 = n22932 | n22933 ;
  assign n22935 = x124 & n5340 ;
  assign n22936 = x123 & n5335 ;
  assign n22937 = x122 & ~n5334 ;
  assign n22938 = n5580 & n22937 ;
  assign n22939 = n22936 | n22938 ;
  assign n22940 = n22935 | n22939 ;
  assign n22941 = n5343 | n22940 ;
  assign n22942 = ( n11916 & n22940 ) | ( n11916 & n22941 ) | ( n22940 & n22941 ) ;
  assign n22943 = x41 & n22942 ;
  assign n22944 = x41 & ~n22943 ;
  assign n22945 = ( n22942 & ~n22943 ) | ( n22942 & n22944 ) | ( ~n22943 & n22944 ) ;
  assign n22946 = ~n22934 & n22945 ;
  assign n22947 = n22934 | n22946 ;
  assign n22948 = n22934 & n22945 ;
  assign n22949 = ~n22754 & n22765 ;
  assign n22950 = n22752 | n22949 ;
  assign n22951 = n22948 | n22950 ;
  assign n22952 = n22947 & ~n22951 ;
  assign n22953 = ( ~n22947 & n22948 ) | ( ~n22947 & n22950 ) | ( n22948 & n22950 ) ;
  assign n22954 = n22952 | n22953 ;
  assign n22955 = x127 & n4572 ;
  assign n22956 = x126 & n4567 ;
  assign n22957 = x125 & ~n4566 ;
  assign n22958 = n4828 & n22957 ;
  assign n22959 = n22956 | n22958 ;
  assign n22960 = n22955 | n22959 ;
  assign n22961 = n4575 | n22960 ;
  assign n22962 = ( n12720 & n22960 ) | ( n12720 & n22961 ) | ( n22960 & n22961 ) ;
  assign n22963 = x38 & n22962 ;
  assign n22964 = x38 & ~n22963 ;
  assign n22965 = ( n22962 & ~n22963 ) | ( n22962 & n22964 ) | ( ~n22963 & n22964 ) ;
  assign n22966 = ~n22954 & n22965 ;
  assign n22967 = n22954 | n22966 ;
  assign n22968 = n22954 & n22965 ;
  assign n22969 = ( n22614 & n22779 ) | ( n22614 & n22782 ) | ( n22779 & n22782 ) ;
  assign n22970 = n22968 | n22969 ;
  assign n22971 = n22967 & ~n22970 ;
  assign n22972 = ( ~n22967 & n22968 ) | ( ~n22967 & n22969 ) | ( n22968 & n22969 ) ;
  assign n22973 = n22971 | n22972 ;
  assign n22974 = n22790 & n22791 ;
  assign n22975 = ~n22973 & n22974 ;
  assign n22976 = n22791 & ~n22974 ;
  assign n22977 = ( ~n22782 & n22792 ) | ( ~n22782 & n22976 ) | ( n22792 & n22976 ) ;
  assign n22978 = ( ~n22973 & n22975 ) | ( ~n22973 & n22977 ) | ( n22975 & n22977 ) ;
  assign n22979 = n22973 & ~n22974 ;
  assign n22980 = ~n22977 & n22979 ;
  assign n22981 = n22978 | n22980 ;
  assign n22982 = ~n22796 & n22803 ;
  assign n22983 = ~n22796 & n22804 ;
  assign n22984 = ( ~n20515 & n22982 ) | ( ~n20515 & n22983 ) | ( n22982 & n22983 ) ;
  assign n22985 = n22981 & n22984 ;
  assign n22986 = n22981 | n22982 ;
  assign n22987 = n22981 | n22983 ;
  assign n22988 = ( ~n20515 & n22986 ) | ( ~n20515 & n22987 ) | ( n22986 & n22987 ) ;
  assign n22989 = ~n22985 & n22988 ;
  assign n22990 = n22966 | n22972 ;
  assign n22991 = x125 & n5340 ;
  assign n22992 = x124 & n5335 ;
  assign n22993 = x123 & ~n5334 ;
  assign n22994 = n5580 & n22993 ;
  assign n22995 = n22992 | n22994 ;
  assign n22996 = n22991 | n22995 ;
  assign n22997 = n5343 | n22996 ;
  assign n22998 = ( n12310 & n22996 ) | ( n12310 & n22997 ) | ( n22996 & n22997 ) ;
  assign n22999 = x41 & n22998 ;
  assign n23000 = x41 & ~n22999 ;
  assign n23001 = ( n22998 & ~n22999 ) | ( n22998 & n23000 ) | ( ~n22999 & n23000 ) ;
  assign n23002 = x127 & n4567 ;
  assign n23003 = x126 & ~n4566 ;
  assign n23004 = n4828 & n23003 ;
  assign n23005 = n23002 | n23004 ;
  assign n23006 = n4575 | n23005 ;
  assign n23007 = ( n13461 & n23005 ) | ( n13461 & n23006 ) | ( n23005 & n23006 ) ;
  assign n23008 = x38 & n23007 ;
  assign n23009 = x38 & ~n23008 ;
  assign n23010 = ( n23007 & ~n23008 ) | ( n23007 & n23009 ) | ( ~n23008 & n23009 ) ;
  assign n23011 = n22946 | n23010 ;
  assign n23012 = n22953 | n23011 ;
  assign n23013 = ( n22946 & n22953 ) | ( n22946 & n23010 ) | ( n22953 & n23010 ) ;
  assign n23014 = n23012 & ~n23013 ;
  assign n23015 = n22838 | n22853 ;
  assign n23016 = x104 & n11984 ;
  assign n23017 = x103 & n11979 ;
  assign n23018 = x102 & ~n11978 ;
  assign n23019 = n12430 & n23018 ;
  assign n23020 = n23017 | n23019 ;
  assign n23021 = n23016 | n23020 ;
  assign n23022 = n11987 | n23021 ;
  assign n23023 = ( n5295 & n23021 ) | ( n5295 & n23022 ) | ( n23021 & n23022 ) ;
  assign n23024 = ~x62 & n23023 ;
  assign n23025 = x62 & ~n23023 ;
  assign n23026 = n23024 | n23025 ;
  assign n23027 = x101 & n12808 ;
  assign n23028 = x63 & x100 ;
  assign n23029 = ~n12808 & n23028 ;
  assign n23030 = n23027 | n23029 ;
  assign n23031 = n22836 & ~n23030 ;
  assign n23032 = n22836 & ~n23031 ;
  assign n23033 = n22836 | n23030 ;
  assign n23034 = ~n23032 & n23033 ;
  assign n23035 = n23026 & ~n23034 ;
  assign n23036 = ~n23026 & n23034 ;
  assign n23037 = n23035 | n23036 ;
  assign n23038 = x107 & n10876 ;
  assign n23039 = x106 & n10871 ;
  assign n23040 = x105 & ~n10870 ;
  assign n23041 = n11305 & n23040 ;
  assign n23042 = n23039 | n23041 ;
  assign n23043 = n23038 | n23042 ;
  assign n23044 = n10879 | n23043 ;
  assign n23045 = ( n6328 & n23043 ) | ( n6328 & n23044 ) | ( n23043 & n23044 ) ;
  assign n23046 = x59 & n23045 ;
  assign n23047 = x59 & ~n23046 ;
  assign n23048 = ( n23045 & ~n23046 ) | ( n23045 & n23047 ) | ( ~n23046 & n23047 ) ;
  assign n23049 = ( n23015 & ~n23037 ) | ( n23015 & n23048 ) | ( ~n23037 & n23048 ) ;
  assign n23050 = ( n23037 & ~n23048 ) | ( n23037 & n23049 ) | ( ~n23048 & n23049 ) ;
  assign n23051 = ( ~n23015 & n23049 ) | ( ~n23015 & n23050 ) | ( n23049 & n23050 ) ;
  assign n23052 = ~n22867 & n23051 ;
  assign n23053 = n22867 & ~n23051 ;
  assign n23054 = n23052 | n23053 ;
  assign n23055 = x110 & n9853 ;
  assign n23056 = x109 & n9848 ;
  assign n23057 = x108 & ~n9847 ;
  assign n23058 = n10165 & n23057 ;
  assign n23059 = n23056 | n23058 ;
  assign n23060 = n23055 | n23059 ;
  assign n23061 = n9856 | n23060 ;
  assign n23062 = ( n7189 & n23060 ) | ( n7189 & n23061 ) | ( n23060 & n23061 ) ;
  assign n23063 = x56 & n23062 ;
  assign n23064 = x56 & ~n23063 ;
  assign n23065 = ( n23062 & ~n23063 ) | ( n23062 & n23064 ) | ( ~n23063 & n23064 ) ;
  assign n23066 = n23054 & n23065 ;
  assign n23067 = ( n22867 & ~n23051 ) | ( n22867 & n23065 ) | ( ~n23051 & n23065 ) ;
  assign n23068 = n23052 | n23067 ;
  assign n23069 = ~n23066 & n23068 ;
  assign n23070 = n22869 | n22874 ;
  assign n23071 = n23069 & ~n23070 ;
  assign n23072 = ~n23069 & n23070 ;
  assign n23073 = n23071 | n23072 ;
  assign n23074 = x113 & n8834 ;
  assign n23075 = x112 & n8829 ;
  assign n23076 = x111 & ~n8828 ;
  assign n23077 = n9159 & n23076 ;
  assign n23078 = n23075 | n23077 ;
  assign n23079 = n23074 | n23078 ;
  assign n23080 = n8837 | n23079 ;
  assign n23081 = ( n8113 & n23079 ) | ( n8113 & n23080 ) | ( n23079 & n23080 ) ;
  assign n23082 = x53 & n23081 ;
  assign n23083 = x53 & ~n23082 ;
  assign n23084 = ( n23081 & ~n23082 ) | ( n23081 & n23083 ) | ( ~n23082 & n23083 ) ;
  assign n23085 = n23073 & n23084 ;
  assign n23086 = ( ~n23069 & n23070 ) | ( ~n23069 & n23084 ) | ( n23070 & n23084 ) ;
  assign n23087 = n23071 | n23086 ;
  assign n23088 = ~n23085 & n23087 ;
  assign n23089 = n22887 | n22892 ;
  assign n23090 = n23088 & ~n23089 ;
  assign n23091 = ~n23088 & n23089 ;
  assign n23092 = n23090 | n23091 ;
  assign n23093 = x116 & n7812 ;
  assign n23094 = x115 & n7807 ;
  assign n23095 = x114 & ~n7806 ;
  assign n23096 = n8136 & n23095 ;
  assign n23097 = n23094 | n23096 ;
  assign n23098 = n23093 | n23097 ;
  assign n23099 = n7815 | n23098 ;
  assign n23100 = ( n8778 & n23098 ) | ( n8778 & n23099 ) | ( n23098 & n23099 ) ;
  assign n23101 = x50 & n23100 ;
  assign n23102 = x50 & ~n23101 ;
  assign n23103 = ( n23100 & ~n23101 ) | ( n23100 & n23102 ) | ( ~n23101 & n23102 ) ;
  assign n23104 = n23092 & n23103 ;
  assign n23105 = ( ~n23088 & n23089 ) | ( ~n23088 & n23103 ) | ( n23089 & n23103 ) ;
  assign n23106 = n23090 | n23105 ;
  assign n23107 = ~n23104 & n23106 ;
  assign n23108 = n22906 | n22909 ;
  assign n23109 = ~n23107 & n23108 ;
  assign n23110 = n23107 & ~n23108 ;
  assign n23111 = n23109 | n23110 ;
  assign n23112 = x119 & n6937 ;
  assign n23113 = x118 & n6932 ;
  assign n23114 = x117 & ~n6931 ;
  assign n23115 = n7216 & n23114 ;
  assign n23116 = n23113 | n23115 ;
  assign n23117 = n23112 | n23116 ;
  assign n23118 = n6940 | n23117 ;
  assign n23119 = ( n9789 & n23117 ) | ( n9789 & n23118 ) | ( n23117 & n23118 ) ;
  assign n23120 = x47 & n23119 ;
  assign n23121 = x47 & ~n23120 ;
  assign n23122 = ( n23119 & ~n23120 ) | ( n23119 & n23121 ) | ( ~n23120 & n23121 ) ;
  assign n23123 = ~n23111 & n23122 ;
  assign n23124 = n23111 | n23123 ;
  assign n23125 = n22923 | n22926 ;
  assign n23126 = n23111 & n23122 ;
  assign n23127 = n23125 | n23126 ;
  assign n23128 = n23124 & ~n23127 ;
  assign n23129 = ( ~n23124 & n23125 ) | ( ~n23124 & n23126 ) | ( n23125 & n23126 ) ;
  assign n23130 = n23128 | n23129 ;
  assign n23131 = x122 & n6068 ;
  assign n23132 = x121 & n6063 ;
  assign n23133 = x120 & ~n6062 ;
  assign n23134 = n6398 & n23133 ;
  assign n23135 = n23132 | n23134 ;
  assign n23136 = n23131 | n23135 ;
  assign n23137 = n6071 | n23136 ;
  assign n23138 = ( n11188 & n23136 ) | ( n11188 & n23137 ) | ( n23136 & n23137 ) ;
  assign n23139 = x44 & n23138 ;
  assign n23140 = x44 & ~n23139 ;
  assign n23141 = ( n23138 & ~n23139 ) | ( n23138 & n23140 ) | ( ~n23139 & n23140 ) ;
  assign n23142 = ~n23130 & n23141 ;
  assign n23143 = n23130 | n23142 ;
  assign n23144 = n23130 & n23141 ;
  assign n23145 = n22929 | n22933 ;
  assign n23146 = n23144 | n23145 ;
  assign n23147 = n23143 & ~n23146 ;
  assign n23148 = ( ~n23143 & n23144 ) | ( ~n23143 & n23145 ) | ( n23144 & n23145 ) ;
  assign n23149 = n23147 | n23148 ;
  assign n23150 = ( n23001 & n23014 ) | ( n23001 & ~n23149 ) | ( n23014 & ~n23149 ) ;
  assign n23151 = ( ~n23014 & n23149 ) | ( ~n23014 & n23150 ) | ( n23149 & n23150 ) ;
  assign n23152 = ( ~n23001 & n23150 ) | ( ~n23001 & n23151 ) | ( n23150 & n23151 ) ;
  assign n23153 = ~n22990 & n23152 ;
  assign n23154 = n22990 & ~n23152 ;
  assign n23155 = n23153 | n23154 ;
  assign n23156 = ~n22978 & n22986 ;
  assign n23157 = ~n22978 & n22987 ;
  assign n23158 = ( ~n20515 & n23156 ) | ( ~n20515 & n23157 ) | ( n23156 & n23157 ) ;
  assign n23159 = n23155 & n23158 ;
  assign n23160 = n23155 | n23156 ;
  assign n23161 = n23155 | n23157 ;
  assign n23162 = ( ~n20515 & n23160 ) | ( ~n20515 & n23161 ) | ( n23160 & n23161 ) ;
  assign n23163 = ~n23159 & n23162 ;
  assign n23164 = ( n23012 & n23013 ) | ( n23012 & n23152 ) | ( n23013 & n23152 ) ;
  assign n23165 = n23129 | n23142 ;
  assign n23166 = x123 & n6068 ;
  assign n23167 = x122 & n6063 ;
  assign n23168 = x121 & ~n6062 ;
  assign n23169 = n6398 & n23168 ;
  assign n23170 = n23167 | n23169 ;
  assign n23171 = n23166 | n23170 ;
  assign n23172 = n6071 | n23171 ;
  assign n23173 = ( n11219 & n23171 ) | ( n11219 & n23172 ) | ( n23171 & n23172 ) ;
  assign n23174 = x44 & n23173 ;
  assign n23175 = x44 & ~n23174 ;
  assign n23176 = ( n23173 & ~n23174 ) | ( n23173 & n23175 ) | ( ~n23174 & n23175 ) ;
  assign n23177 = x102 & n12808 ;
  assign n23178 = x63 & x101 ;
  assign n23179 = ~n12808 & n23178 ;
  assign n23180 = n23177 | n23179 ;
  assign n23181 = ~n23030 & n23180 ;
  assign n23182 = n23030 | n23181 ;
  assign n23183 = n23180 & ~n23181 ;
  assign n23184 = n23182 & ~n23183 ;
  assign n23185 = n23031 | n23184 ;
  assign n23186 = n23035 | n23185 ;
  assign n23187 = n23031 | n23035 ;
  assign n23188 = n23184 & n23187 ;
  assign n23189 = n23186 & ~n23188 ;
  assign n23190 = x105 & n11984 ;
  assign n23191 = x104 & n11979 ;
  assign n23192 = x103 & ~n11978 ;
  assign n23193 = n12430 & n23192 ;
  assign n23194 = n23191 | n23193 ;
  assign n23195 = n23190 | n23194 ;
  assign n23196 = n11987 | n23195 ;
  assign n23197 = ( n5788 & n23195 ) | ( n5788 & n23196 ) | ( n23195 & n23196 ) ;
  assign n23198 = x62 & n23197 ;
  assign n23199 = x62 & ~n23198 ;
  assign n23200 = ( n23197 & ~n23198 ) | ( n23197 & n23199 ) | ( ~n23198 & n23199 ) ;
  assign n23201 = ~n23189 & n23200 ;
  assign n23202 = n23189 & ~n23200 ;
  assign n23203 = n23201 | n23202 ;
  assign n23204 = x108 & n10876 ;
  assign n23205 = x107 & n10871 ;
  assign n23206 = x106 & ~n10870 ;
  assign n23207 = n11305 & n23206 ;
  assign n23208 = n23205 | n23207 ;
  assign n23209 = n23204 | n23208 ;
  assign n23210 = n10879 | n23209 ;
  assign n23211 = ( n6358 & n23209 ) | ( n6358 & n23210 ) | ( n23209 & n23210 ) ;
  assign n23212 = x59 & n23211 ;
  assign n23213 = x59 & ~n23212 ;
  assign n23214 = ( n23211 & ~n23212 ) | ( n23211 & n23213 ) | ( ~n23212 & n23213 ) ;
  assign n23215 = n23203 | n23214 ;
  assign n23216 = n23203 & n23214 ;
  assign n23217 = n23215 & ~n23216 ;
  assign n23218 = ~n23049 & n23217 ;
  assign n23219 = n23049 & ~n23217 ;
  assign n23220 = n23218 | n23219 ;
  assign n23221 = x111 & n9853 ;
  assign n23222 = x110 & n9848 ;
  assign n23223 = x109 & ~n9847 ;
  assign n23224 = n10165 & n23223 ;
  assign n23225 = n23222 | n23224 ;
  assign n23226 = n23221 | n23225 ;
  assign n23227 = n9856 | n23226 ;
  assign n23228 = ( n7492 & n23226 ) | ( n7492 & n23227 ) | ( n23226 & n23227 ) ;
  assign n23229 = x56 & n23228 ;
  assign n23230 = x56 & ~n23229 ;
  assign n23231 = ( n23228 & ~n23229 ) | ( n23228 & n23230 ) | ( ~n23229 & n23230 ) ;
  assign n23232 = n23220 & n23231 ;
  assign n23233 = ( n23049 & ~n23217 ) | ( n23049 & n23231 ) | ( ~n23217 & n23231 ) ;
  assign n23234 = n23218 | n23233 ;
  assign n23235 = ~n23232 & n23234 ;
  assign n23236 = ~n23067 & n23235 ;
  assign n23237 = n23067 & ~n23235 ;
  assign n23238 = n23236 | n23237 ;
  assign n23239 = x114 & n8834 ;
  assign n23240 = x113 & n8829 ;
  assign n23241 = x112 & ~n8828 ;
  assign n23242 = n9159 & n23241 ;
  assign n23243 = n23240 | n23242 ;
  assign n23244 = n23239 | n23243 ;
  assign n23245 = n8837 | n23244 ;
  assign n23246 = ( n8437 & n23244 ) | ( n8437 & n23245 ) | ( n23244 & n23245 ) ;
  assign n23247 = x53 & n23246 ;
  assign n23248 = x53 & ~n23247 ;
  assign n23249 = ( n23246 & ~n23247 ) | ( n23246 & n23248 ) | ( ~n23247 & n23248 ) ;
  assign n23250 = n23238 & ~n23249 ;
  assign n23251 = ~n23238 & n23249 ;
  assign n23252 = n23250 | n23251 ;
  assign n23253 = x117 & n7812 ;
  assign n23254 = x116 & n7807 ;
  assign n23255 = x115 & ~n7806 ;
  assign n23256 = n8136 & n23255 ;
  assign n23257 = n23254 | n23256 ;
  assign n23258 = n23253 | n23257 ;
  assign n23259 = n7815 | n23258 ;
  assign n23260 = ( n9118 & n23258 ) | ( n9118 & n23259 ) | ( n23258 & n23259 ) ;
  assign n23261 = x50 & n23260 ;
  assign n23262 = x50 & ~n23261 ;
  assign n23263 = ( n23260 & ~n23261 ) | ( n23260 & n23262 ) | ( ~n23261 & n23262 ) ;
  assign n23264 = ( n23086 & ~n23252 ) | ( n23086 & n23263 ) | ( ~n23252 & n23263 ) ;
  assign n23265 = ( n23252 & ~n23263 ) | ( n23252 & n23264 ) | ( ~n23263 & n23264 ) ;
  assign n23266 = ( ~n23086 & n23264 ) | ( ~n23086 & n23265 ) | ( n23264 & n23265 ) ;
  assign n23267 = n23105 & ~n23266 ;
  assign n23268 = ~n23105 & n23266 ;
  assign n23269 = n23267 | n23268 ;
  assign n23270 = x120 & n6937 ;
  assign n23271 = x119 & n6932 ;
  assign n23272 = x118 & ~n6931 ;
  assign n23273 = n7216 & n23272 ;
  assign n23274 = n23271 | n23273 ;
  assign n23275 = n23270 | n23274 ;
  assign n23276 = n6940 | n23275 ;
  assign n23277 = ( n10460 & n23275 ) | ( n10460 & n23276 ) | ( n23275 & n23276 ) ;
  assign n23278 = x47 & n23277 ;
  assign n23279 = x47 & ~n23278 ;
  assign n23280 = ( n23277 & ~n23278 ) | ( n23277 & n23279 ) | ( ~n23278 & n23279 ) ;
  assign n23281 = ~n23269 & n23280 ;
  assign n23282 = n23269 & ~n23280 ;
  assign n23283 = n23281 | n23282 ;
  assign n23284 = n23109 | n23123 ;
  assign n23285 = ( n23176 & n23283 ) | ( n23176 & ~n23284 ) | ( n23283 & ~n23284 ) ;
  assign n23286 = ( ~n23283 & n23284 ) | ( ~n23283 & n23285 ) | ( n23284 & n23285 ) ;
  assign n23287 = ( ~n23176 & n23285 ) | ( ~n23176 & n23286 ) | ( n23285 & n23286 ) ;
  assign n23288 = ~n23165 & n23287 ;
  assign n23289 = n23165 & ~n23287 ;
  assign n23290 = n23288 | n23289 ;
  assign n23291 = x126 & n5340 ;
  assign n23292 = x125 & n5335 ;
  assign n23293 = x124 & ~n5334 ;
  assign n23294 = n5580 & n23293 ;
  assign n23295 = n23292 | n23294 ;
  assign n23296 = n23291 | n23295 ;
  assign n23297 = n5343 | n23296 ;
  assign n23298 = ( n12687 & n23296 ) | ( n12687 & n23297 ) | ( n23296 & n23297 ) ;
  assign n23299 = x41 & n23298 ;
  assign n23300 = x41 & ~n23299 ;
  assign n23301 = ( n23298 & ~n23299 ) | ( n23298 & n23300 ) | ( ~n23299 & n23300 ) ;
  assign n23302 = n23290 & n23301 ;
  assign n23303 = ( n23165 & ~n23287 ) | ( n23165 & n23301 ) | ( ~n23287 & n23301 ) ;
  assign n23304 = n23288 | n23303 ;
  assign n23305 = ~n23302 & n23304 ;
  assign n23306 = x127 & ~n4566 ;
  assign n23307 = n4828 & n23306 ;
  assign n23308 = ( x127 & n4575 ) | ( x127 & n23307 ) | ( n4575 & n23307 ) ;
  assign n23309 = ( x126 & n23307 ) | ( x126 & n23308 ) | ( n23307 & n23308 ) ;
  assign n23310 = ( n12685 & n23308 ) | ( n12685 & n23309 ) | ( n23308 & n23309 ) ;
  assign n23311 = x38 & n23310 ;
  assign n23312 = x38 & ~n23311 ;
  assign n23313 = ( n23310 & ~n23311 ) | ( n23310 & n23312 ) | ( ~n23311 & n23312 ) ;
  assign n23314 = n23001 & ~n23149 ;
  assign n23315 = n23148 | n23314 ;
  assign n23316 = ( n23305 & n23313 ) | ( n23305 & ~n23315 ) | ( n23313 & ~n23315 ) ;
  assign n23317 = ( ~n23313 & n23315 ) | ( ~n23313 & n23316 ) | ( n23315 & n23316 ) ;
  assign n23318 = ( ~n23305 & n23316 ) | ( ~n23305 & n23317 ) | ( n23316 & n23317 ) ;
  assign n23319 = n23164 & ~n23318 ;
  assign n23320 = ~n23164 & n23318 ;
  assign n23321 = n23319 | n23320 ;
  assign n23322 = ~n23154 & n23160 ;
  assign n23323 = ~n23154 & n23161 ;
  assign n23324 = ( ~n20515 & n23322 ) | ( ~n20515 & n23323 ) | ( n23322 & n23323 ) ;
  assign n23325 = n23321 & n23324 ;
  assign n23326 = n23321 | n23322 ;
  assign n23327 = n23321 | n23323 ;
  assign n23328 = ( ~n20515 & n23326 ) | ( ~n20515 & n23327 ) | ( n23326 & n23327 ) ;
  assign n23329 = ~n23325 & n23328 ;
  assign n23330 = x127 & n5340 ;
  assign n23331 = x126 & n5335 ;
  assign n23332 = x125 & ~n5334 ;
  assign n23333 = n5580 & n23332 ;
  assign n23334 = n23331 | n23333 ;
  assign n23335 = n23330 | n23334 ;
  assign n23336 = n5343 | n23335 ;
  assign n23337 = ( n12720 & n23335 ) | ( n12720 & n23336 ) | ( n23335 & n23336 ) ;
  assign n23338 = x41 & n23337 ;
  assign n23339 = x41 & ~n23338 ;
  assign n23340 = ( n23337 & ~n23338 ) | ( n23337 & n23339 ) | ( ~n23338 & n23339 ) ;
  assign n23341 = x124 & n6068 ;
  assign n23342 = x123 & n6063 ;
  assign n23343 = x122 & ~n6062 ;
  assign n23344 = n6398 & n23343 ;
  assign n23345 = n23342 | n23344 ;
  assign n23346 = n23341 | n23345 ;
  assign n23347 = n6071 | n23346 ;
  assign n23348 = ( n11916 & n23346 ) | ( n11916 & n23347 ) | ( n23346 & n23347 ) ;
  assign n23349 = x44 & n23348 ;
  assign n23350 = x44 & ~n23349 ;
  assign n23351 = ( n23348 & ~n23349 ) | ( n23348 & n23350 ) | ( ~n23349 & n23350 ) ;
  assign n23352 = n23267 | n23281 ;
  assign n23353 = x121 & n6937 ;
  assign n23354 = x120 & n6932 ;
  assign n23355 = x119 & ~n6931 ;
  assign n23356 = n7216 & n23355 ;
  assign n23357 = n23354 | n23356 ;
  assign n23358 = n23353 | n23357 ;
  assign n23359 = n6940 | n23358 ;
  assign n23360 = ( n10811 & n23358 ) | ( n10811 & n23359 ) | ( n23358 & n23359 ) ;
  assign n23361 = x47 & n23360 ;
  assign n23362 = x47 & ~n23361 ;
  assign n23363 = ( n23360 & ~n23361 ) | ( n23360 & n23362 ) | ( ~n23361 & n23362 ) ;
  assign n23364 = x112 & n9853 ;
  assign n23365 = x111 & n9848 ;
  assign n23366 = x110 & ~n9847 ;
  assign n23367 = n10165 & n23366 ;
  assign n23368 = n23365 | n23367 ;
  assign n23369 = n23364 | n23368 ;
  assign n23370 = n9856 | n23369 ;
  assign n23371 = ( n7789 & n23369 ) | ( n7789 & n23370 ) | ( n23369 & n23370 ) ;
  assign n23372 = x56 & n23371 ;
  assign n23373 = x56 & ~n23372 ;
  assign n23374 = ( n23371 & ~n23372 ) | ( n23371 & n23373 ) | ( ~n23372 & n23373 ) ;
  assign n23375 = ( n23201 & ~n23203 ) | ( n23201 & n23215 ) | ( ~n23203 & n23215 ) ;
  assign n23376 = x109 & n10876 ;
  assign n23377 = x108 & n10871 ;
  assign n23378 = x107 & ~n10870 ;
  assign n23379 = n11305 & n23378 ;
  assign n23380 = n23377 | n23379 ;
  assign n23381 = n23376 | n23380 ;
  assign n23382 = n10879 | n23381 ;
  assign n23383 = ( n6884 & n23381 ) | ( n6884 & n23382 ) | ( n23381 & n23382 ) ;
  assign n23384 = x59 & n23383 ;
  assign n23385 = x59 & ~n23384 ;
  assign n23386 = ( n23383 & ~n23384 ) | ( n23383 & n23385 ) | ( ~n23384 & n23385 ) ;
  assign n23387 = x106 & n11984 ;
  assign n23388 = x105 & n11979 ;
  assign n23389 = x104 & ~n11978 ;
  assign n23390 = n12430 & n23389 ;
  assign n23391 = n23388 | n23390 ;
  assign n23392 = n23387 | n23391 ;
  assign n23393 = n11987 | n23392 ;
  assign n23394 = ( n5814 & n23392 ) | ( n5814 & n23393 ) | ( n23392 & n23393 ) ;
  assign n23395 = x62 & n23394 ;
  assign n23396 = x62 & ~n23395 ;
  assign n23397 = ( n23394 & ~n23395 ) | ( n23394 & n23396 ) | ( ~n23395 & n23396 ) ;
  assign n23398 = x103 & n12808 ;
  assign n23399 = x63 & x102 ;
  assign n23400 = ~n12808 & n23399 ;
  assign n23401 = n23398 | n23400 ;
  assign n23402 = ( x38 & ~n23030 ) | ( x38 & n23401 ) | ( ~n23030 & n23401 ) ;
  assign n23403 = ( ~x38 & n23030 ) | ( ~x38 & n23401 ) | ( n23030 & n23401 ) ;
  assign n23404 = ( ~n23401 & n23402 ) | ( ~n23401 & n23403 ) | ( n23402 & n23403 ) ;
  assign n23405 = ( ~n23030 & n23180 ) | ( ~n23030 & n23187 ) | ( n23180 & n23187 ) ;
  assign n23406 = ~n23404 & n23405 ;
  assign n23407 = n23404 & ~n23405 ;
  assign n23408 = n23406 | n23407 ;
  assign n23409 = n23397 & ~n23408 ;
  assign n23410 = n23408 | n23409 ;
  assign n23411 = ( ~n23397 & n23409 ) | ( ~n23397 & n23410 ) | ( n23409 & n23410 ) ;
  assign n23412 = ( n23375 & ~n23386 ) | ( n23375 & n23411 ) | ( ~n23386 & n23411 ) ;
  assign n23413 = ( n23386 & ~n23411 ) | ( n23386 & n23412 ) | ( ~n23411 & n23412 ) ;
  assign n23414 = ( ~n23375 & n23412 ) | ( ~n23375 & n23413 ) | ( n23412 & n23413 ) ;
  assign n23415 = n23374 & ~n23414 ;
  assign n23416 = ~n23374 & n23414 ;
  assign n23417 = n23415 | n23416 ;
  assign n23418 = ~n23233 & n23417 ;
  assign n23419 = n23233 & ~n23417 ;
  assign n23420 = n23418 | n23419 ;
  assign n23421 = x115 & n8834 ;
  assign n23422 = x114 & n8829 ;
  assign n23423 = x113 & ~n8828 ;
  assign n23424 = n9159 & n23423 ;
  assign n23425 = n23422 | n23424 ;
  assign n23426 = n23421 | n23425 ;
  assign n23427 = n8837 | n23426 ;
  assign n23428 = ( n8749 & n23426 ) | ( n8749 & n23427 ) | ( n23426 & n23427 ) ;
  assign n23429 = x53 & n23428 ;
  assign n23430 = x53 & ~n23429 ;
  assign n23431 = ( n23428 & ~n23429 ) | ( n23428 & n23430 ) | ( ~n23429 & n23430 ) ;
  assign n23432 = n23420 & ~n23431 ;
  assign n23433 = ~n23420 & n23431 ;
  assign n23434 = n23432 | n23433 ;
  assign n23435 = n23237 | n23251 ;
  assign n23436 = ~n23434 & n23435 ;
  assign n23437 = n23434 & ~n23435 ;
  assign n23438 = n23436 | n23437 ;
  assign n23439 = x118 & n7812 ;
  assign n23440 = x117 & n7807 ;
  assign n23441 = x116 & ~n7806 ;
  assign n23442 = n8136 & n23441 ;
  assign n23443 = n23440 | n23442 ;
  assign n23444 = n23439 | n23443 ;
  assign n23445 = n7815 | n23444 ;
  assign n23446 = ( n9760 & n23444 ) | ( n9760 & n23445 ) | ( n23444 & n23445 ) ;
  assign n23447 = x50 & n23446 ;
  assign n23448 = x50 & ~n23447 ;
  assign n23449 = ( n23446 & ~n23447 ) | ( n23446 & n23448 ) | ( ~n23447 & n23448 ) ;
  assign n23450 = ~n23438 & n23449 ;
  assign n23451 = n23438 & ~n23449 ;
  assign n23452 = n23450 | n23451 ;
  assign n23453 = n23264 & ~n23452 ;
  assign n23454 = ~n23264 & n23452 ;
  assign n23455 = n23453 | n23454 ;
  assign n23456 = n23363 & ~n23455 ;
  assign n23457 = n23455 | n23456 ;
  assign n23458 = ( ~n23363 & n23456 ) | ( ~n23363 & n23457 ) | ( n23456 & n23457 ) ;
  assign n23459 = ~n23352 & n23458 ;
  assign n23460 = n23352 & ~n23458 ;
  assign n23461 = n23459 | n23460 ;
  assign n23462 = n23351 & ~n23461 ;
  assign n23463 = n23461 | n23462 ;
  assign n23464 = ( ~n23351 & n23462 ) | ( ~n23351 & n23463 ) | ( n23462 & n23463 ) ;
  assign n23465 = ~n23286 & n23464 ;
  assign n23466 = n23286 & ~n23464 ;
  assign n23467 = n23465 | n23466 ;
  assign n23468 = n23340 & ~n23467 ;
  assign n23469 = n23467 | n23468 ;
  assign n23470 = ( ~n23340 & n23468 ) | ( ~n23340 & n23469 ) | ( n23468 & n23469 ) ;
  assign n23471 = ~n23303 & n23470 ;
  assign n23472 = n23303 & ~n23470 ;
  assign n23473 = n23471 | n23472 ;
  assign n23474 = ( ~n23305 & n23313 ) | ( ~n23305 & n23315 ) | ( n23313 & n23315 ) ;
  assign n23475 = ~n23473 & n23474 ;
  assign n23476 = n23473 & ~n23474 ;
  assign n23477 = n23475 | n23476 ;
  assign n23478 = ~n23319 & n23326 ;
  assign n23479 = ~n23319 & n23327 ;
  assign n23480 = ( ~n20515 & n23478 ) | ( ~n20515 & n23479 ) | ( n23478 & n23479 ) ;
  assign n23481 = n23477 & n23480 ;
  assign n23482 = n23477 | n23478 ;
  assign n23483 = n23477 | n23479 ;
  assign n23484 = ( ~n20515 & n23482 ) | ( ~n20515 & n23483 ) | ( n23482 & n23483 ) ;
  assign n23485 = ~n23481 & n23484 ;
  assign n23486 = x125 & n6068 ;
  assign n23487 = x124 & n6063 ;
  assign n23488 = x123 & ~n6062 ;
  assign n23489 = n6398 & n23488 ;
  assign n23490 = n23487 | n23489 ;
  assign n23491 = n23486 | n23490 ;
  assign n23492 = n6071 | n23491 ;
  assign n23493 = ( n12310 & n23491 ) | ( n12310 & n23492 ) | ( n23491 & n23492 ) ;
  assign n23494 = x44 & n23493 ;
  assign n23495 = x44 & ~n23494 ;
  assign n23496 = ( n23493 & ~n23494 ) | ( n23493 & n23495 ) | ( ~n23494 & n23495 ) ;
  assign n23497 = x127 & n5335 ;
  assign n23498 = x126 & ~n5334 ;
  assign n23499 = n5580 & n23498 ;
  assign n23500 = n23497 | n23499 ;
  assign n23501 = n5343 | n23500 ;
  assign n23502 = ( n13461 & n23500 ) | ( n13461 & n23501 ) | ( n23500 & n23501 ) ;
  assign n23503 = x41 & n23502 ;
  assign n23504 = x41 & ~n23503 ;
  assign n23505 = ( n23502 & ~n23503 ) | ( n23502 & n23504 ) | ( ~n23503 & n23504 ) ;
  assign n23506 = n23462 | n23466 ;
  assign n23507 = n23505 & n23506 ;
  assign n23508 = n23505 | n23506 ;
  assign n23509 = ~n23507 & n23508 ;
  assign n23510 = n23450 | n23453 ;
  assign n23511 = x110 & n10876 ;
  assign n23512 = x109 & n10871 ;
  assign n23513 = x108 & ~n10870 ;
  assign n23514 = n11305 & n23513 ;
  assign n23515 = n23512 | n23514 ;
  assign n23516 = n23511 | n23515 ;
  assign n23517 = n10879 | n23516 ;
  assign n23518 = ( n7189 & n23516 ) | ( n7189 & n23517 ) | ( n23516 & n23517 ) ;
  assign n23519 = x59 & n23518 ;
  assign n23520 = x59 & ~n23519 ;
  assign n23521 = ( n23518 & ~n23519 ) | ( n23518 & n23520 ) | ( ~n23519 & n23520 ) ;
  assign n23522 = x104 & n12808 ;
  assign n23523 = x63 & x103 ;
  assign n23524 = ~n12808 & n23523 ;
  assign n23525 = n23522 | n23524 ;
  assign n23526 = n23403 & ~n23525 ;
  assign n23527 = ~n23403 & n23525 ;
  assign n23528 = n23526 | n23527 ;
  assign n23529 = x107 & n11984 ;
  assign n23530 = x106 & n11979 ;
  assign n23531 = x105 & ~n11978 ;
  assign n23532 = n12430 & n23531 ;
  assign n23533 = n23530 | n23532 ;
  assign n23534 = n23529 | n23533 ;
  assign n23535 = n11987 | n23534 ;
  assign n23536 = ( n6328 & n23534 ) | ( n6328 & n23535 ) | ( n23534 & n23535 ) ;
  assign n23537 = x62 & n23536 ;
  assign n23538 = x62 & ~n23537 ;
  assign n23539 = ( n23536 & ~n23537 ) | ( n23536 & n23538 ) | ( ~n23537 & n23538 ) ;
  assign n23540 = ~n23528 & n23539 ;
  assign n23541 = n23528 & ~n23539 ;
  assign n23542 = n23540 | n23541 ;
  assign n23543 = n23406 | n23409 ;
  assign n23544 = ( n23521 & n23542 ) | ( n23521 & ~n23543 ) | ( n23542 & ~n23543 ) ;
  assign n23545 = ( ~n23542 & n23543 ) | ( ~n23542 & n23544 ) | ( n23543 & n23544 ) ;
  assign n23546 = ( ~n23521 & n23544 ) | ( ~n23521 & n23545 ) | ( n23544 & n23545 ) ;
  assign n23547 = ~n23413 & n23546 ;
  assign n23548 = n23413 & ~n23546 ;
  assign n23549 = n23547 | n23548 ;
  assign n23550 = x113 & n9853 ;
  assign n23551 = x112 & n9848 ;
  assign n23552 = x111 & ~n9847 ;
  assign n23553 = n10165 & n23552 ;
  assign n23554 = n23551 | n23553 ;
  assign n23555 = n23550 | n23554 ;
  assign n23556 = n9856 | n23555 ;
  assign n23557 = ( n8113 & n23555 ) | ( n8113 & n23556 ) | ( n23555 & n23556 ) ;
  assign n23558 = x56 & n23557 ;
  assign n23559 = x56 & ~n23558 ;
  assign n23560 = ( n23557 & ~n23558 ) | ( n23557 & n23559 ) | ( ~n23558 & n23559 ) ;
  assign n23561 = n23549 & n23560 ;
  assign n23562 = ( n23413 & ~n23546 ) | ( n23413 & n23560 ) | ( ~n23546 & n23560 ) ;
  assign n23563 = n23547 | n23562 ;
  assign n23564 = ~n23561 & n23563 ;
  assign n23565 = n23415 | n23419 ;
  assign n23566 = n23564 & ~n23565 ;
  assign n23567 = ~n23564 & n23565 ;
  assign n23568 = n23566 | n23567 ;
  assign n23569 = x116 & n8834 ;
  assign n23570 = x115 & n8829 ;
  assign n23571 = x114 & ~n8828 ;
  assign n23572 = n9159 & n23571 ;
  assign n23573 = n23570 | n23572 ;
  assign n23574 = n23569 | n23573 ;
  assign n23575 = n8837 | n23574 ;
  assign n23576 = ( n8778 & n23574 ) | ( n8778 & n23575 ) | ( n23574 & n23575 ) ;
  assign n23577 = x53 & n23576 ;
  assign n23578 = x53 & ~n23577 ;
  assign n23579 = ( n23576 & ~n23577 ) | ( n23576 & n23578 ) | ( ~n23577 & n23578 ) ;
  assign n23580 = n23568 & n23579 ;
  assign n23581 = ( ~n23564 & n23565 ) | ( ~n23564 & n23579 ) | ( n23565 & n23579 ) ;
  assign n23582 = n23566 | n23581 ;
  assign n23583 = ~n23580 & n23582 ;
  assign n23584 = n23433 | n23436 ;
  assign n23585 = ~n23583 & n23584 ;
  assign n23586 = n23583 | n23585 ;
  assign n23587 = n23583 & n23584 ;
  assign n23588 = n23586 & ~n23587 ;
  assign n23589 = x119 & n7812 ;
  assign n23590 = x118 & n7807 ;
  assign n23591 = x117 & ~n7806 ;
  assign n23592 = n8136 & n23591 ;
  assign n23593 = n23590 | n23592 ;
  assign n23594 = n23589 | n23593 ;
  assign n23595 = n7815 | n23594 ;
  assign n23596 = ( n9789 & n23594 ) | ( n9789 & n23595 ) | ( n23594 & n23595 ) ;
  assign n23597 = x50 & n23596 ;
  assign n23598 = x50 & ~n23597 ;
  assign n23599 = ( n23596 & ~n23597 ) | ( n23596 & n23598 ) | ( ~n23597 & n23598 ) ;
  assign n23600 = ~n23588 & n23599 ;
  assign n23601 = n23588 & ~n23599 ;
  assign n23602 = n23600 | n23601 ;
  assign n23603 = ~n23510 & n23602 ;
  assign n23604 = x122 & n6937 ;
  assign n23605 = x121 & n6932 ;
  assign n23606 = x120 & ~n6931 ;
  assign n23607 = n7216 & n23606 ;
  assign n23608 = n23605 | n23607 ;
  assign n23609 = n23604 | n23608 ;
  assign n23610 = n6940 | n23609 ;
  assign n23611 = ( n11188 & n23609 ) | ( n11188 & n23610 ) | ( n23609 & n23610 ) ;
  assign n23612 = x47 & n23611 ;
  assign n23613 = x47 & ~n23612 ;
  assign n23614 = ( n23611 & ~n23612 ) | ( n23611 & n23613 ) | ( ~n23612 & n23613 ) ;
  assign n23615 = ( n23510 & ~n23602 ) | ( n23510 & n23614 ) | ( ~n23602 & n23614 ) ;
  assign n23616 = n23603 | n23615 ;
  assign n23617 = n23456 | n23460 ;
  assign n23618 = n23510 & ~n23602 ;
  assign n23619 = n23603 | n23618 ;
  assign n23620 = n23614 & n23619 ;
  assign n23621 = n23617 | n23620 ;
  assign n23622 = n23616 & ~n23621 ;
  assign n23623 = ( ~n23616 & n23617 ) | ( ~n23616 & n23620 ) | ( n23617 & n23620 ) ;
  assign n23624 = n23622 | n23623 ;
  assign n23625 = ( n23496 & n23509 ) | ( n23496 & ~n23624 ) | ( n23509 & ~n23624 ) ;
  assign n23626 = ( ~n23509 & n23624 ) | ( ~n23509 & n23625 ) | ( n23624 & n23625 ) ;
  assign n23627 = ( ~n23496 & n23625 ) | ( ~n23496 & n23626 ) | ( n23625 & n23626 ) ;
  assign n23628 = n23468 | n23472 ;
  assign n23629 = n23627 & ~n23628 ;
  assign n23630 = ~n23627 & n23628 ;
  assign n23631 = n23629 | n23630 ;
  assign n23632 = ~n23475 & n23482 ;
  assign n23633 = ~n23475 & n23483 ;
  assign n23634 = ( ~n20515 & n23632 ) | ( ~n20515 & n23633 ) | ( n23632 & n23633 ) ;
  assign n23635 = n23631 & n23634 ;
  assign n23636 = n23631 | n23632 ;
  assign n23637 = n23631 | n23633 ;
  assign n23638 = ( ~n20515 & n23636 ) | ( ~n20515 & n23637 ) | ( n23636 & n23637 ) ;
  assign n23639 = ~n23635 & n23638 ;
  assign n23640 = x111 & n10876 ;
  assign n23641 = x110 & n10871 ;
  assign n23642 = x109 & ~n10870 ;
  assign n23643 = n11305 & n23642 ;
  assign n23644 = n23641 | n23643 ;
  assign n23645 = n23640 | n23644 ;
  assign n23646 = n10879 | n23645 ;
  assign n23647 = ( n7492 & n23645 ) | ( n7492 & n23646 ) | ( n23645 & n23646 ) ;
  assign n23648 = x59 & n23647 ;
  assign n23649 = x59 & ~n23648 ;
  assign n23650 = ( n23647 & ~n23648 ) | ( n23647 & n23649 ) | ( ~n23648 & n23649 ) ;
  assign n23651 = x108 & n11984 ;
  assign n23652 = x107 & n11979 ;
  assign n23653 = x106 & ~n11978 ;
  assign n23654 = n12430 & n23653 ;
  assign n23655 = n23652 | n23654 ;
  assign n23656 = n23651 | n23655 ;
  assign n23657 = n11987 | n23656 ;
  assign n23658 = ( n6358 & n23656 ) | ( n6358 & n23657 ) | ( n23656 & n23657 ) ;
  assign n23659 = x62 & n23658 ;
  assign n23660 = x62 & ~n23659 ;
  assign n23661 = ( n23658 & ~n23659 ) | ( n23658 & n23660 ) | ( ~n23659 & n23660 ) ;
  assign n23662 = x105 & n12808 ;
  assign n23663 = x63 & x104 ;
  assign n23664 = ~n12808 & n23663 ;
  assign n23665 = n23662 | n23664 ;
  assign n23666 = ~n23525 & n23665 ;
  assign n23667 = n23525 | n23666 ;
  assign n23668 = n23665 & ~n23666 ;
  assign n23669 = n23667 & ~n23668 ;
  assign n23670 = ( n23526 & n23540 ) | ( n23526 & ~n23669 ) | ( n23540 & ~n23669 ) ;
  assign n23671 = n23669 | n23670 ;
  assign n23672 = ( n23526 & n23540 ) | ( n23526 & ~n23670 ) | ( n23540 & ~n23670 ) ;
  assign n23673 = n23671 & ~n23672 ;
  assign n23674 = ( n23650 & ~n23661 ) | ( n23650 & n23673 ) | ( ~n23661 & n23673 ) ;
  assign n23675 = ( n23661 & ~n23673 ) | ( n23661 & n23674 ) | ( ~n23673 & n23674 ) ;
  assign n23676 = ( ~n23650 & n23674 ) | ( ~n23650 & n23675 ) | ( n23674 & n23675 ) ;
  assign n23677 = ~n23545 & n23676 ;
  assign n23678 = n23545 & ~n23676 ;
  assign n23679 = n23677 | n23678 ;
  assign n23680 = x114 & n9853 ;
  assign n23681 = x113 & n9848 ;
  assign n23682 = x112 & ~n9847 ;
  assign n23683 = n10165 & n23682 ;
  assign n23684 = n23681 | n23683 ;
  assign n23685 = n23680 | n23684 ;
  assign n23686 = n9856 | n23685 ;
  assign n23687 = ( n8437 & n23685 ) | ( n8437 & n23686 ) | ( n23685 & n23686 ) ;
  assign n23688 = x56 & n23687 ;
  assign n23689 = x56 & ~n23688 ;
  assign n23690 = ( n23687 & ~n23688 ) | ( n23687 & n23689 ) | ( ~n23688 & n23689 ) ;
  assign n23691 = n23679 & ~n23690 ;
  assign n23692 = ~n23679 & n23690 ;
  assign n23693 = n23691 | n23692 ;
  assign n23694 = n23562 & ~n23693 ;
  assign n23695 = n23562 & ~n23694 ;
  assign n23696 = n23562 | n23693 ;
  assign n23697 = x117 & n8834 ;
  assign n23698 = x116 & n8829 ;
  assign n23699 = x115 & ~n8828 ;
  assign n23700 = n9159 & n23699 ;
  assign n23701 = n23698 | n23700 ;
  assign n23702 = n23697 | n23701 ;
  assign n23703 = n8837 | n23702 ;
  assign n23704 = ( n9118 & n23702 ) | ( n9118 & n23703 ) | ( n23702 & n23703 ) ;
  assign n23705 = x53 & n23704 ;
  assign n23706 = x53 & ~n23705 ;
  assign n23707 = ( n23704 & ~n23705 ) | ( n23704 & n23706 ) | ( ~n23705 & n23706 ) ;
  assign n23708 = n23696 & ~n23707 ;
  assign n23709 = ~n23695 & n23708 ;
  assign n23710 = ( n23695 & ~n23696 ) | ( n23695 & n23707 ) | ( ~n23696 & n23707 ) ;
  assign n23711 = n23709 | n23710 ;
  assign n23712 = n23581 & ~n23711 ;
  assign n23713 = n23581 & ~n23712 ;
  assign n23714 = n23581 | n23711 ;
  assign n23715 = x120 & n7812 ;
  assign n23716 = x119 & n7807 ;
  assign n23717 = x118 & ~n7806 ;
  assign n23718 = n8136 & n23717 ;
  assign n23719 = n23716 | n23718 ;
  assign n23720 = n23715 | n23719 ;
  assign n23721 = n7815 | n23720 ;
  assign n23722 = ( n10460 & n23720 ) | ( n10460 & n23721 ) | ( n23720 & n23721 ) ;
  assign n23723 = x50 & n23722 ;
  assign n23724 = x50 & ~n23723 ;
  assign n23725 = ( n23722 & ~n23723 ) | ( n23722 & n23724 ) | ( ~n23723 & n23724 ) ;
  assign n23726 = n23714 & ~n23725 ;
  assign n23727 = ~n23713 & n23726 ;
  assign n23728 = ( n23713 & ~n23714 ) | ( n23713 & n23725 ) | ( ~n23714 & n23725 ) ;
  assign n23729 = n23727 | n23728 ;
  assign n23730 = ~n23585 & n23729 ;
  assign n23731 = ~n23600 & n23730 ;
  assign n23732 = ( n23585 & n23600 ) | ( n23585 & ~n23729 ) | ( n23600 & ~n23729 ) ;
  assign n23733 = n23731 | n23732 ;
  assign n23734 = x123 & n6937 ;
  assign n23735 = x122 & n6932 ;
  assign n23736 = x121 & ~n6931 ;
  assign n23737 = n7216 & n23736 ;
  assign n23738 = n23735 | n23737 ;
  assign n23739 = n23734 | n23738 ;
  assign n23740 = n6940 | n23739 ;
  assign n23741 = ( n11219 & n23739 ) | ( n11219 & n23740 ) | ( n23739 & n23740 ) ;
  assign n23742 = x47 & n23741 ;
  assign n23743 = x47 & ~n23742 ;
  assign n23744 = ( n23741 & ~n23742 ) | ( n23741 & n23743 ) | ( ~n23742 & n23743 ) ;
  assign n23745 = n23733 | n23744 ;
  assign n23746 = ~n23744 & n23745 ;
  assign n23747 = ( ~n23733 & n23745 ) | ( ~n23733 & n23746 ) | ( n23745 & n23746 ) ;
  assign n23748 = ~n23615 & n23747 ;
  assign n23749 = n23615 & ~n23747 ;
  assign n23750 = n23748 | n23749 ;
  assign n23751 = x126 & n6068 ;
  assign n23752 = x125 & n6063 ;
  assign n23753 = x124 & ~n6062 ;
  assign n23754 = n6398 & n23753 ;
  assign n23755 = n23752 | n23754 ;
  assign n23756 = n23751 | n23755 ;
  assign n23757 = n6071 | n23756 ;
  assign n23758 = ( n12687 & n23756 ) | ( n12687 & n23757 ) | ( n23756 & n23757 ) ;
  assign n23759 = x44 & n23758 ;
  assign n23760 = x44 & ~n23759 ;
  assign n23761 = ( n23758 & ~n23759 ) | ( n23758 & n23760 ) | ( ~n23759 & n23760 ) ;
  assign n23762 = n23750 & n23761 ;
  assign n23763 = ( n23615 & ~n23747 ) | ( n23615 & n23761 ) | ( ~n23747 & n23761 ) ;
  assign n23764 = n23748 | n23763 ;
  assign n23765 = ~n23762 & n23764 ;
  assign n23766 = x127 & ~n5334 ;
  assign n23767 = n5580 & n23766 ;
  assign n23768 = ( x127 & n5343 ) | ( x127 & n23767 ) | ( n5343 & n23767 ) ;
  assign n23769 = ( x126 & n23767 ) | ( x126 & n23768 ) | ( n23767 & n23768 ) ;
  assign n23770 = ( n12685 & n23768 ) | ( n12685 & n23769 ) | ( n23768 & n23769 ) ;
  assign n23771 = x41 & n23770 ;
  assign n23772 = x41 & ~n23771 ;
  assign n23773 = ( n23770 & ~n23771 ) | ( n23770 & n23772 ) | ( ~n23771 & n23772 ) ;
  assign n23774 = n23496 & ~n23624 ;
  assign n23775 = n23623 | n23774 ;
  assign n23776 = ( n23765 & n23773 ) | ( n23765 & ~n23775 ) | ( n23773 & ~n23775 ) ;
  assign n23777 = ( ~n23773 & n23775 ) | ( ~n23773 & n23776 ) | ( n23775 & n23776 ) ;
  assign n23778 = ( ~n23765 & n23776 ) | ( ~n23765 & n23777 ) | ( n23776 & n23777 ) ;
  assign n23779 = ( n23505 & n23506 ) | ( n23505 & n23627 ) | ( n23506 & n23627 ) ;
  assign n23780 = ~n23778 & n23779 ;
  assign n23781 = n23778 & ~n23779 ;
  assign n23782 = n23780 | n23781 ;
  assign n23783 = ~n23630 & n23636 ;
  assign n23784 = ~n23630 & n23637 ;
  assign n23785 = ( ~n20515 & n23783 ) | ( ~n20515 & n23784 ) | ( n23783 & n23784 ) ;
  assign n23786 = n23782 & n23785 ;
  assign n23787 = n23782 | n23783 ;
  assign n23788 = n23782 | n23784 ;
  assign n23789 = ( ~n20515 & n23787 ) | ( ~n20515 & n23788 ) | ( n23787 & n23788 ) ;
  assign n23790 = ~n23786 & n23789 ;
  assign n23791 = x127 & n6068 ;
  assign n23792 = x126 & n6063 ;
  assign n23793 = x125 & ~n6062 ;
  assign n23794 = n6398 & n23793 ;
  assign n23795 = n23792 | n23794 ;
  assign n23796 = n23791 | n23795 ;
  assign n23797 = n6071 | n23796 ;
  assign n23798 = ( n12720 & n23796 ) | ( n12720 & n23797 ) | ( n23796 & n23797 ) ;
  assign n23799 = x44 & n23798 ;
  assign n23800 = x44 & ~n23799 ;
  assign n23801 = ( n23798 & ~n23799 ) | ( n23798 & n23800 ) | ( ~n23799 & n23800 ) ;
  assign n23802 = ( n23732 & n23744 ) | ( n23732 & n23747 ) | ( n23744 & n23747 ) ;
  assign n23803 = x124 & n6937 ;
  assign n23804 = x123 & n6932 ;
  assign n23805 = x122 & ~n6931 ;
  assign n23806 = n7216 & n23805 ;
  assign n23807 = n23804 | n23806 ;
  assign n23808 = n23803 | n23807 ;
  assign n23809 = n6940 | n23808 ;
  assign n23810 = ( n11916 & n23808 ) | ( n11916 & n23809 ) | ( n23808 & n23809 ) ;
  assign n23811 = x47 & n23810 ;
  assign n23812 = x47 & ~n23811 ;
  assign n23813 = ( n23810 & ~n23811 ) | ( n23810 & n23812 ) | ( ~n23811 & n23812 ) ;
  assign n23814 = n23712 | n23728 ;
  assign n23815 = n23694 | n23710 ;
  assign n23816 = n23678 | n23692 ;
  assign n23817 = x115 & n9853 ;
  assign n23818 = x114 & n9848 ;
  assign n23819 = x113 & ~n9847 ;
  assign n23820 = n10165 & n23819 ;
  assign n23821 = n23818 | n23820 ;
  assign n23822 = n23817 | n23821 ;
  assign n23823 = n9856 | n23822 ;
  assign n23824 = ( n8749 & n23822 ) | ( n8749 & n23823 ) | ( n23822 & n23823 ) ;
  assign n23825 = x56 & n23824 ;
  assign n23826 = x56 & ~n23825 ;
  assign n23827 = ( n23824 & ~n23825 ) | ( n23824 & n23826 ) | ( ~n23825 & n23826 ) ;
  assign n23828 = n23666 | n23670 ;
  assign n23829 = x109 & n11984 ;
  assign n23830 = x108 & n11979 ;
  assign n23831 = x107 & ~n11978 ;
  assign n23832 = n12430 & n23831 ;
  assign n23833 = n23830 | n23832 ;
  assign n23834 = n23829 | n23833 ;
  assign n23835 = n11987 | n23834 ;
  assign n23836 = ( n6884 & n23834 ) | ( n6884 & n23835 ) | ( n23834 & n23835 ) ;
  assign n23837 = ~x62 & n23836 ;
  assign n23838 = x62 & ~n23836 ;
  assign n23839 = n23837 | n23838 ;
  assign n23840 = x106 & n12808 ;
  assign n23841 = x63 & x105 ;
  assign n23842 = ~n12808 & n23841 ;
  assign n23843 = n23840 | n23842 ;
  assign n23844 = ( x41 & ~n23525 ) | ( x41 & n23843 ) | ( ~n23525 & n23843 ) ;
  assign n23845 = ( ~x41 & n23525 ) | ( ~x41 & n23843 ) | ( n23525 & n23843 ) ;
  assign n23846 = ( ~n23843 & n23844 ) | ( ~n23843 & n23845 ) | ( n23844 & n23845 ) ;
  assign n23847 = ( n23828 & ~n23839 ) | ( n23828 & n23846 ) | ( ~n23839 & n23846 ) ;
  assign n23848 = ( n23839 & ~n23846 ) | ( n23839 & n23847 ) | ( ~n23846 & n23847 ) ;
  assign n23849 = ( ~n23828 & n23847 ) | ( ~n23828 & n23848 ) | ( n23847 & n23848 ) ;
  assign n23850 = x112 & n10876 ;
  assign n23851 = x111 & n10871 ;
  assign n23852 = x110 & ~n10870 ;
  assign n23853 = n11305 & n23852 ;
  assign n23854 = n23851 | n23853 ;
  assign n23855 = n23850 | n23854 ;
  assign n23856 = n10879 | n23855 ;
  assign n23857 = ( n7789 & n23855 ) | ( n7789 & n23856 ) | ( n23855 & n23856 ) ;
  assign n23858 = x59 & n23857 ;
  assign n23859 = x59 & ~n23858 ;
  assign n23860 = ( n23857 & ~n23858 ) | ( n23857 & n23859 ) | ( ~n23858 & n23859 ) ;
  assign n23861 = ~n23849 & n23860 ;
  assign n23862 = n23849 | n23861 ;
  assign n23863 = n23849 & n23860 ;
  assign n23864 = n23675 | n23863 ;
  assign n23865 = n23862 & ~n23864 ;
  assign n23866 = ( n23675 & ~n23862 ) | ( n23675 & n23863 ) | ( ~n23862 & n23863 ) ;
  assign n23867 = n23865 | n23866 ;
  assign n23868 = n23827 & ~n23867 ;
  assign n23869 = n23867 | n23868 ;
  assign n23870 = ( ~n23827 & n23868 ) | ( ~n23827 & n23869 ) | ( n23868 & n23869 ) ;
  assign n23871 = n23816 & ~n23870 ;
  assign n23872 = ~n23816 & n23870 ;
  assign n23873 = n23871 | n23872 ;
  assign n23874 = x118 & n8834 ;
  assign n23875 = x117 & n8829 ;
  assign n23876 = x116 & ~n8828 ;
  assign n23877 = n9159 & n23876 ;
  assign n23878 = n23875 | n23877 ;
  assign n23879 = n23874 | n23878 ;
  assign n23880 = n8837 | n23879 ;
  assign n23881 = ( n9760 & n23879 ) | ( n9760 & n23880 ) | ( n23879 & n23880 ) ;
  assign n23882 = x53 & n23881 ;
  assign n23883 = x53 & ~n23882 ;
  assign n23884 = ( n23881 & ~n23882 ) | ( n23881 & n23883 ) | ( ~n23882 & n23883 ) ;
  assign n23885 = n23873 & ~n23884 ;
  assign n23886 = ~n23873 & n23884 ;
  assign n23887 = n23885 | n23886 ;
  assign n23888 = n23815 & ~n23887 ;
  assign n23889 = ~n23815 & n23887 ;
  assign n23890 = n23888 | n23889 ;
  assign n23891 = x121 & n7812 ;
  assign n23892 = x120 & n7807 ;
  assign n23893 = x119 & ~n7806 ;
  assign n23894 = n8136 & n23893 ;
  assign n23895 = n23892 | n23894 ;
  assign n23896 = n23891 | n23895 ;
  assign n23897 = n7815 | n23896 ;
  assign n23898 = ( n10811 & n23896 ) | ( n10811 & n23897 ) | ( n23896 & n23897 ) ;
  assign n23899 = x50 & n23898 ;
  assign n23900 = x50 & ~n23899 ;
  assign n23901 = ( n23898 & ~n23899 ) | ( n23898 & n23900 ) | ( ~n23899 & n23900 ) ;
  assign n23902 = n23890 & ~n23901 ;
  assign n23903 = ~n23890 & n23901 ;
  assign n23904 = n23902 | n23903 ;
  assign n23905 = n23814 & ~n23904 ;
  assign n23906 = ~n23814 & n23904 ;
  assign n23907 = n23905 | n23906 ;
  assign n23908 = n23813 & ~n23907 ;
  assign n23909 = n23907 | n23908 ;
  assign n23910 = ( ~n23813 & n23908 ) | ( ~n23813 & n23909 ) | ( n23908 & n23909 ) ;
  assign n23911 = ~n23802 & n23910 ;
  assign n23912 = n23802 & ~n23910 ;
  assign n23913 = n23911 | n23912 ;
  assign n23914 = n23801 & ~n23913 ;
  assign n23915 = n23913 | n23914 ;
  assign n23916 = ( ~n23801 & n23914 ) | ( ~n23801 & n23915 ) | ( n23914 & n23915 ) ;
  assign n23917 = ~n23763 & n23916 ;
  assign n23918 = n23763 & ~n23916 ;
  assign n23919 = n23917 | n23918 ;
  assign n23920 = n23773 & n23775 ;
  assign n23921 = n23919 & ~n23920 ;
  assign n23922 = n23775 & ~n23920 ;
  assign n23923 = ( ~n23765 & n23776 ) | ( ~n23765 & n23922 ) | ( n23776 & n23922 ) ;
  assign n23924 = n23921 & ~n23923 ;
  assign n23925 = ( ~n23919 & n23920 ) | ( ~n23919 & n23923 ) | ( n23920 & n23923 ) ;
  assign n23926 = n23924 | n23925 ;
  assign n23927 = ~n23780 & n23787 ;
  assign n23928 = ~n23780 & n23788 ;
  assign n23929 = ( ~n20515 & n23927 ) | ( ~n20515 & n23928 ) | ( n23927 & n23928 ) ;
  assign n23930 = n23926 & n23929 ;
  assign n23931 = n23926 | n23927 ;
  assign n23932 = n23926 | n23928 ;
  assign n23933 = ( ~n20515 & n23931 ) | ( ~n20515 & n23932 ) | ( n23931 & n23932 ) ;
  assign n23934 = ~n23930 & n23933 ;
  assign n23935 = x127 & n6063 ;
  assign n23936 = x126 & ~n6062 ;
  assign n23937 = n6398 & n23936 ;
  assign n23938 = n23935 | n23937 ;
  assign n23939 = n6071 | n23938 ;
  assign n23940 = ( n13461 & n23938 ) | ( n13461 & n23939 ) | ( n23938 & n23939 ) ;
  assign n23941 = x44 & n23940 ;
  assign n23942 = x44 & ~n23941 ;
  assign n23943 = ( n23940 & ~n23941 ) | ( n23940 & n23942 ) | ( ~n23941 & n23942 ) ;
  assign n23944 = n23908 | n23912 ;
  assign n23945 = n23943 & n23944 ;
  assign n23946 = n23943 | n23944 ;
  assign n23947 = ~n23945 & n23946 ;
  assign n23948 = n23903 | n23905 ;
  assign n23949 = n23861 | n23866 ;
  assign n23950 = x113 & n10876 ;
  assign n23951 = x112 & n10871 ;
  assign n23952 = x111 & ~n10870 ;
  assign n23953 = n11305 & n23952 ;
  assign n23954 = n23951 | n23953 ;
  assign n23955 = n23950 | n23954 ;
  assign n23956 = n10879 | n23955 ;
  assign n23957 = ( n8113 & n23955 ) | ( n8113 & n23956 ) | ( n23955 & n23956 ) ;
  assign n23958 = x59 & n23957 ;
  assign n23959 = x59 & ~n23958 ;
  assign n23960 = ( n23957 & ~n23958 ) | ( n23957 & n23959 ) | ( ~n23958 & n23959 ) ;
  assign n23961 = x107 & n12808 ;
  assign n23962 = x63 & x106 ;
  assign n23963 = ~n12808 & n23962 ;
  assign n23964 = n23961 | n23963 ;
  assign n23965 = n23845 & ~n23964 ;
  assign n23966 = n23845 & ~n23965 ;
  assign n23967 = n23845 | n23964 ;
  assign n23968 = ~n23966 & n23967 ;
  assign n23969 = x110 & n11984 ;
  assign n23970 = x109 & n11979 ;
  assign n23971 = x108 & ~n11978 ;
  assign n23972 = n12430 & n23971 ;
  assign n23973 = n23970 | n23972 ;
  assign n23974 = n23969 | n23973 ;
  assign n23975 = n11987 | n23974 ;
  assign n23976 = ( n7189 & n23974 ) | ( n7189 & n23975 ) | ( n23974 & n23975 ) ;
  assign n23977 = x62 & n23976 ;
  assign n23978 = x62 & ~n23977 ;
  assign n23979 = ( n23976 & ~n23977 ) | ( n23976 & n23978 ) | ( ~n23977 & n23978 ) ;
  assign n23980 = ~n23968 & n23979 ;
  assign n23981 = n23968 & ~n23979 ;
  assign n23982 = n23980 | n23981 ;
  assign n23983 = ( ~n23848 & n23960 ) | ( ~n23848 & n23982 ) | ( n23960 & n23982 ) ;
  assign n23984 = ( n23848 & ~n23982 ) | ( n23848 & n23983 ) | ( ~n23982 & n23983 ) ;
  assign n23985 = ( ~n23960 & n23983 ) | ( ~n23960 & n23984 ) | ( n23983 & n23984 ) ;
  assign n23986 = ~n23949 & n23985 ;
  assign n23987 = n23949 & ~n23985 ;
  assign n23988 = n23986 | n23987 ;
  assign n23989 = x116 & n9853 ;
  assign n23990 = x115 & n9848 ;
  assign n23991 = x114 & ~n9847 ;
  assign n23992 = n10165 & n23991 ;
  assign n23993 = n23990 | n23992 ;
  assign n23994 = n23989 | n23993 ;
  assign n23995 = n9856 | n23994 ;
  assign n23996 = ( n8778 & n23994 ) | ( n8778 & n23995 ) | ( n23994 & n23995 ) ;
  assign n23997 = x56 & n23996 ;
  assign n23998 = x56 & ~n23997 ;
  assign n23999 = ( n23996 & ~n23997 ) | ( n23996 & n23998 ) | ( ~n23997 & n23998 ) ;
  assign n24000 = n23988 & n23999 ;
  assign n24001 = ( n23949 & ~n23985 ) | ( n23949 & n23999 ) | ( ~n23985 & n23999 ) ;
  assign n24002 = n23986 | n24001 ;
  assign n24003 = ~n24000 & n24002 ;
  assign n24004 = n23868 | n23871 ;
  assign n24005 = n24003 & ~n24004 ;
  assign n24006 = ~n24003 & n24004 ;
  assign n24007 = n24005 | n24006 ;
  assign n24008 = x119 & n8834 ;
  assign n24009 = x118 & n8829 ;
  assign n24010 = x117 & ~n8828 ;
  assign n24011 = n9159 & n24010 ;
  assign n24012 = n24009 | n24011 ;
  assign n24013 = n24008 | n24012 ;
  assign n24014 = n8837 | n24013 ;
  assign n24015 = ( n9789 & n24013 ) | ( n9789 & n24014 ) | ( n24013 & n24014 ) ;
  assign n24016 = x53 & n24015 ;
  assign n24017 = x53 & ~n24016 ;
  assign n24018 = ( n24015 & ~n24016 ) | ( n24015 & n24017 ) | ( ~n24016 & n24017 ) ;
  assign n24019 = n24007 & n24018 ;
  assign n24020 = ( ~n24003 & n24004 ) | ( ~n24003 & n24018 ) | ( n24004 & n24018 ) ;
  assign n24021 = n24005 | n24020 ;
  assign n24022 = ~n24019 & n24021 ;
  assign n24023 = ( n23886 & n23888 ) | ( n23886 & n24022 ) | ( n23888 & n24022 ) ;
  assign n24024 = n23886 | n23888 ;
  assign n24025 = n24022 | n24024 ;
  assign n24026 = ~n24023 & n24025 ;
  assign n24027 = x122 & n7812 ;
  assign n24028 = x121 & n7807 ;
  assign n24029 = x120 & ~n7806 ;
  assign n24030 = n8136 & n24029 ;
  assign n24031 = n24028 | n24030 ;
  assign n24032 = n24027 | n24031 ;
  assign n24033 = n7815 | n24032 ;
  assign n24034 = ( n11188 & n24032 ) | ( n11188 & n24033 ) | ( n24032 & n24033 ) ;
  assign n24035 = x50 & n24034 ;
  assign n24036 = x50 & ~n24035 ;
  assign n24037 = ( n24034 & ~n24035 ) | ( n24034 & n24036 ) | ( ~n24035 & n24036 ) ;
  assign n24038 = n24026 & ~n24037 ;
  assign n24039 = ~n24026 & n24037 ;
  assign n24040 = n24038 | n24039 ;
  assign n24041 = n23948 & ~n24040 ;
  assign n24042 = n23948 & ~n24041 ;
  assign n24043 = n24040 | n24041 ;
  assign n24044 = ~n24042 & n24043 ;
  assign n24045 = x125 & n6937 ;
  assign n24046 = x124 & n6932 ;
  assign n24047 = x123 & ~n6931 ;
  assign n24048 = n7216 & n24047 ;
  assign n24049 = n24046 | n24048 ;
  assign n24050 = n24045 | n24049 ;
  assign n24051 = n6940 | n24050 ;
  assign n24052 = ( n12310 & n24050 ) | ( n12310 & n24051 ) | ( n24050 & n24051 ) ;
  assign n24053 = x47 & n24052 ;
  assign n24054 = x47 & ~n24053 ;
  assign n24055 = ( n24052 & ~n24053 ) | ( n24052 & n24054 ) | ( ~n24053 & n24054 ) ;
  assign n24056 = n24044 & n24055 ;
  assign n24057 = n24044 | n24055 ;
  assign n24058 = ~n24056 & n24057 ;
  assign n24059 = n23947 & ~n24058 ;
  assign n24060 = n24058 | n24059 ;
  assign n24061 = ( ~n23947 & n24059 ) | ( ~n23947 & n24060 ) | ( n24059 & n24060 ) ;
  assign n24062 = n23914 | n23918 ;
  assign n24063 = n24061 & ~n24062 ;
  assign n24064 = ~n24061 & n24062 ;
  assign n24065 = n24063 | n24064 ;
  assign n24066 = ~n23925 & n23931 ;
  assign n24067 = ~n23925 & n23932 ;
  assign n24068 = ( ~n20515 & n24066 ) | ( ~n20515 & n24067 ) | ( n24066 & n24067 ) ;
  assign n24069 = n24065 & n24068 ;
  assign n24070 = n24065 | n24066 ;
  assign n24071 = n24065 | n24067 ;
  assign n24072 = ( ~n20515 & n24070 ) | ( ~n20515 & n24071 ) | ( n24070 & n24071 ) ;
  assign n24073 = ~n24069 & n24072 ;
  assign n24074 = n23945 | n24059 ;
  assign n24075 = x127 & ~n6062 ;
  assign n24076 = n6398 & n24075 ;
  assign n24077 = ( x127 & n6071 ) | ( x127 & n24076 ) | ( n6071 & n24076 ) ;
  assign n24078 = ( x126 & n24076 ) | ( x126 & n24077 ) | ( n24076 & n24077 ) ;
  assign n24079 = ( n12685 & n24077 ) | ( n12685 & n24078 ) | ( n24077 & n24078 ) ;
  assign n24080 = x44 & n24079 ;
  assign n24081 = x44 & ~n24080 ;
  assign n24082 = ( n24079 & ~n24080 ) | ( n24079 & n24081 ) | ( ~n24080 & n24081 ) ;
  assign n24083 = ( n24041 & ~n24044 ) | ( n24041 & n24057 ) | ( ~n24044 & n24057 ) ;
  assign n24084 = n24082 & n24083 ;
  assign n24085 = n24082 | n24083 ;
  assign n24086 = ~n24084 & n24085 ;
  assign n24087 = x123 & n7812 ;
  assign n24088 = x122 & n7807 ;
  assign n24089 = x121 & ~n7806 ;
  assign n24090 = n8136 & n24089 ;
  assign n24091 = n24088 | n24090 ;
  assign n24092 = n24087 | n24091 ;
  assign n24093 = n7815 | n24092 ;
  assign n24094 = ( n11219 & n24092 ) | ( n11219 & n24093 ) | ( n24092 & n24093 ) ;
  assign n24095 = x50 & n24094 ;
  assign n24096 = x50 & ~n24095 ;
  assign n24097 = ( n24094 & ~n24095 ) | ( n24094 & n24096 ) | ( ~n24095 & n24096 ) ;
  assign n24098 = x108 & n12808 ;
  assign n24099 = x63 & x107 ;
  assign n24100 = ~n12808 & n24099 ;
  assign n24101 = n24098 | n24100 ;
  assign n24102 = ~n23964 & n24101 ;
  assign n24103 = n23964 & ~n24101 ;
  assign n24104 = n24102 | n24103 ;
  assign n24105 = x111 & n11984 ;
  assign n24106 = x110 & n11979 ;
  assign n24107 = x109 & ~n11978 ;
  assign n24108 = n12430 & n24107 ;
  assign n24109 = n24106 | n24108 ;
  assign n24110 = n24105 | n24109 ;
  assign n24111 = n11987 | n24110 ;
  assign n24112 = ( n7492 & n24110 ) | ( n7492 & n24111 ) | ( n24110 & n24111 ) ;
  assign n24113 = x62 & n24112 ;
  assign n24114 = x62 & ~n24113 ;
  assign n24115 = ( n24112 & ~n24113 ) | ( n24112 & n24114 ) | ( ~n24113 & n24114 ) ;
  assign n24116 = ~n24104 & n24115 ;
  assign n24117 = n24104 & ~n24115 ;
  assign n24118 = n24116 | n24117 ;
  assign n24119 = n23965 | n23980 ;
  assign n24120 = n24118 & n24119 ;
  assign n24121 = ~n24118 & n24119 ;
  assign n24122 = n24118 | n24121 ;
  assign n24123 = x114 & n10876 ;
  assign n24124 = x113 & n10871 ;
  assign n24125 = x112 & ~n10870 ;
  assign n24126 = n11305 & n24125 ;
  assign n24127 = n24124 | n24126 ;
  assign n24128 = n24123 | n24127 ;
  assign n24129 = n10879 | n24128 ;
  assign n24130 = ( n8437 & n24128 ) | ( n8437 & n24129 ) | ( n24128 & n24129 ) ;
  assign n24131 = x59 & n24130 ;
  assign n24132 = x59 & ~n24131 ;
  assign n24133 = ( n24130 & ~n24131 ) | ( n24130 & n24132 ) | ( ~n24131 & n24132 ) ;
  assign n24134 = n24122 & ~n24133 ;
  assign n24135 = ~n24120 & n24134 ;
  assign n24136 = ( n24120 & ~n24122 ) | ( n24120 & n24133 ) | ( ~n24122 & n24133 ) ;
  assign n24137 = n24135 | n24136 ;
  assign n24138 = x117 & n9853 ;
  assign n24139 = x116 & n9848 ;
  assign n24140 = x115 & ~n9847 ;
  assign n24141 = n10165 & n24140 ;
  assign n24142 = n24139 | n24141 ;
  assign n24143 = n24138 | n24142 ;
  assign n24144 = n9856 | n24143 ;
  assign n24145 = ( n9118 & n24143 ) | ( n9118 & n24144 ) | ( n24143 & n24144 ) ;
  assign n24146 = x56 & n24145 ;
  assign n24147 = x56 & ~n24146 ;
  assign n24148 = ( n24145 & ~n24146 ) | ( n24145 & n24147 ) | ( ~n24146 & n24147 ) ;
  assign n24149 = ( n23984 & ~n24137 ) | ( n23984 & n24148 ) | ( ~n24137 & n24148 ) ;
  assign n24150 = ( n24137 & ~n24148 ) | ( n24137 & n24149 ) | ( ~n24148 & n24149 ) ;
  assign n24151 = ( ~n23984 & n24149 ) | ( ~n23984 & n24150 ) | ( n24149 & n24150 ) ;
  assign n24152 = n24001 & ~n24151 ;
  assign n24153 = n24001 & ~n24152 ;
  assign n24154 = n24001 | n24151 ;
  assign n24155 = x120 & n8834 ;
  assign n24156 = x119 & n8829 ;
  assign n24157 = x118 & ~n8828 ;
  assign n24158 = n9159 & n24157 ;
  assign n24159 = n24156 | n24158 ;
  assign n24160 = n24155 | n24159 ;
  assign n24161 = n8837 | n24160 ;
  assign n24162 = ( n10460 & n24160 ) | ( n10460 & n24161 ) | ( n24160 & n24161 ) ;
  assign n24163 = x53 & n24162 ;
  assign n24164 = x53 & ~n24163 ;
  assign n24165 = ( n24162 & ~n24163 ) | ( n24162 & n24164 ) | ( ~n24163 & n24164 ) ;
  assign n24166 = n24154 & ~n24165 ;
  assign n24167 = ~n24153 & n24166 ;
  assign n24168 = ( n24153 & ~n24154 ) | ( n24153 & n24165 ) | ( ~n24154 & n24165 ) ;
  assign n24169 = n24167 | n24168 ;
  assign n24170 = ( n24020 & n24097 ) | ( n24020 & ~n24169 ) | ( n24097 & ~n24169 ) ;
  assign n24171 = ( ~n24020 & n24169 ) | ( ~n24020 & n24170 ) | ( n24169 & n24170 ) ;
  assign n24172 = ( ~n24097 & n24170 ) | ( ~n24097 & n24171 ) | ( n24170 & n24171 ) ;
  assign n24173 = ( ~n24022 & n24024 ) | ( ~n24022 & n24037 ) | ( n24024 & n24037 ) ;
  assign n24174 = ~n24172 & n24173 ;
  assign n24175 = n24172 | n24174 ;
  assign n24176 = n24172 & n24173 ;
  assign n24177 = n24175 & ~n24176 ;
  assign n24178 = x126 & n6937 ;
  assign n24179 = x125 & n6932 ;
  assign n24180 = x124 & ~n6931 ;
  assign n24181 = n7216 & n24180 ;
  assign n24182 = n24179 | n24181 ;
  assign n24183 = n24178 | n24182 ;
  assign n24184 = n6940 | n24183 ;
  assign n24185 = ( n12687 & n24183 ) | ( n12687 & n24184 ) | ( n24183 & n24184 ) ;
  assign n24186 = x47 & n24185 ;
  assign n24187 = x47 & ~n24186 ;
  assign n24188 = ( n24185 & ~n24186 ) | ( n24185 & n24187 ) | ( ~n24186 & n24187 ) ;
  assign n24189 = ~n24177 & n24188 ;
  assign n24190 = n24177 & ~n24188 ;
  assign n24191 = n24189 | n24190 ;
  assign n24192 = n24086 & n24191 ;
  assign n24193 = n24086 | n24191 ;
  assign n24194 = ~n24192 & n24193 ;
  assign n24195 = n24074 & ~n24194 ;
  assign n24196 = ~n24074 & n24194 ;
  assign n24197 = n24195 | n24196 ;
  assign n24198 = ~n24064 & n24070 ;
  assign n24199 = ~n24064 & n24071 ;
  assign n24200 = ( ~n20515 & n24198 ) | ( ~n20515 & n24199 ) | ( n24198 & n24199 ) ;
  assign n24201 = n24197 & n24200 ;
  assign n24202 = n24197 | n24198 ;
  assign n24203 = n24197 | n24199 ;
  assign n24204 = ( ~n20515 & n24202 ) | ( ~n20515 & n24203 ) | ( n24202 & n24203 ) ;
  assign n24205 = ~n24201 & n24204 ;
  assign n24206 = n24174 | n24189 ;
  assign n24207 = x127 & n6937 ;
  assign n24208 = x126 & n6932 ;
  assign n24209 = x125 & ~n6931 ;
  assign n24210 = n7216 & n24209 ;
  assign n24211 = n24208 | n24210 ;
  assign n24212 = n24207 | n24211 ;
  assign n24213 = n6940 | n24212 ;
  assign n24214 = ( n12720 & n24212 ) | ( n12720 & n24213 ) | ( n24212 & n24213 ) ;
  assign n24215 = x47 & n24214 ;
  assign n24216 = x47 & ~n24215 ;
  assign n24217 = ( n24214 & ~n24215 ) | ( n24214 & n24216 ) | ( ~n24215 & n24216 ) ;
  assign n24218 = n24152 | n24168 ;
  assign n24219 = n24121 | n24136 ;
  assign n24220 = x109 & n12808 ;
  assign n24221 = x63 & x108 ;
  assign n24222 = ~n12808 & n24221 ;
  assign n24223 = n24220 | n24222 ;
  assign n24224 = ~x44 & n24223 ;
  assign n24225 = x44 & ~n24223 ;
  assign n24226 = n24224 | n24225 ;
  assign n24227 = n23964 | n24226 ;
  assign n24228 = n23964 & ~n24226 ;
  assign n24229 = ( ~n23964 & n24227 ) | ( ~n23964 & n24228 ) | ( n24227 & n24228 ) ;
  assign n24230 = ( n24102 & n24116 ) | ( n24102 & ~n24229 ) | ( n24116 & ~n24229 ) ;
  assign n24231 = ( n24102 & n24116 ) | ( n24102 & ~n24230 ) | ( n24116 & ~n24230 ) ;
  assign n24232 = n24229 | n24230 ;
  assign n24233 = ~n24231 & n24232 ;
  assign n24234 = x112 & n11984 ;
  assign n24235 = x111 & n11979 ;
  assign n24236 = x110 & ~n11978 ;
  assign n24237 = n12430 & n24236 ;
  assign n24238 = n24235 | n24237 ;
  assign n24239 = n24234 | n24238 ;
  assign n24240 = n11987 | n24239 ;
  assign n24241 = ( n7789 & n24239 ) | ( n7789 & n24240 ) | ( n24239 & n24240 ) ;
  assign n24242 = x62 & n24241 ;
  assign n24243 = x62 & ~n24242 ;
  assign n24244 = ( n24241 & ~n24242 ) | ( n24241 & n24243 ) | ( ~n24242 & n24243 ) ;
  assign n24245 = n24233 | n24244 ;
  assign n24246 = n24233 & n24244 ;
  assign n24247 = x115 & n10876 ;
  assign n24248 = x114 & n10871 ;
  assign n24249 = x113 & ~n10870 ;
  assign n24250 = n11305 & n24249 ;
  assign n24251 = n24248 | n24250 ;
  assign n24252 = n24247 | n24251 ;
  assign n24253 = n10879 | n24252 ;
  assign n24254 = ( n8749 & n24252 ) | ( n8749 & n24253 ) | ( n24252 & n24253 ) ;
  assign n24255 = x59 & n24254 ;
  assign n24256 = x59 & ~n24255 ;
  assign n24257 = ( n24254 & ~n24255 ) | ( n24254 & n24256 ) | ( ~n24255 & n24256 ) ;
  assign n24258 = n24246 | n24257 ;
  assign n24259 = n24245 & ~n24258 ;
  assign n24260 = ( ~n24245 & n24246 ) | ( ~n24245 & n24257 ) | ( n24246 & n24257 ) ;
  assign n24261 = n24259 | n24260 ;
  assign n24262 = n24219 & ~n24261 ;
  assign n24263 = ~n24219 & n24261 ;
  assign n24264 = n24262 | n24263 ;
  assign n24265 = x118 & n9853 ;
  assign n24266 = x117 & n9848 ;
  assign n24267 = x116 & ~n9847 ;
  assign n24268 = n10165 & n24267 ;
  assign n24269 = n24266 | n24268 ;
  assign n24270 = n24265 | n24269 ;
  assign n24271 = n9856 | n24270 ;
  assign n24272 = ( n9760 & n24270 ) | ( n9760 & n24271 ) | ( n24270 & n24271 ) ;
  assign n24273 = x56 & n24272 ;
  assign n24274 = x56 & ~n24273 ;
  assign n24275 = ( n24272 & ~n24273 ) | ( n24272 & n24274 ) | ( ~n24273 & n24274 ) ;
  assign n24276 = n24264 & ~n24275 ;
  assign n24277 = ~n24264 & n24275 ;
  assign n24278 = n24276 | n24277 ;
  assign n24279 = n24149 & ~n24278 ;
  assign n24280 = ~n24149 & n24278 ;
  assign n24281 = n24279 | n24280 ;
  assign n24282 = x121 & n8834 ;
  assign n24283 = x120 & n8829 ;
  assign n24284 = x119 & ~n8828 ;
  assign n24285 = n9159 & n24284 ;
  assign n24286 = n24283 | n24285 ;
  assign n24287 = n24282 | n24286 ;
  assign n24288 = n8837 | n24287 ;
  assign n24289 = ( n10811 & n24287 ) | ( n10811 & n24288 ) | ( n24287 & n24288 ) ;
  assign n24290 = x53 & n24289 ;
  assign n24291 = x53 & ~n24290 ;
  assign n24292 = ( n24289 & ~n24290 ) | ( n24289 & n24291 ) | ( ~n24290 & n24291 ) ;
  assign n24293 = n24281 & ~n24292 ;
  assign n24294 = ~n24281 & n24292 ;
  assign n24295 = n24293 | n24294 ;
  assign n24296 = n24218 & ~n24295 ;
  assign n24297 = ~n24218 & n24295 ;
  assign n24298 = n24296 | n24297 ;
  assign n24299 = x124 & n7812 ;
  assign n24300 = x123 & n7807 ;
  assign n24301 = x122 & ~n7806 ;
  assign n24302 = n8136 & n24301 ;
  assign n24303 = n24300 | n24302 ;
  assign n24304 = n24299 | n24303 ;
  assign n24305 = n7815 | n24304 ;
  assign n24306 = ( n11916 & n24304 ) | ( n11916 & n24305 ) | ( n24304 & n24305 ) ;
  assign n24307 = x50 & n24306 ;
  assign n24308 = x50 & ~n24307 ;
  assign n24309 = ( n24306 & ~n24307 ) | ( n24306 & n24308 ) | ( ~n24307 & n24308 ) ;
  assign n24310 = n24298 & ~n24309 ;
  assign n24311 = ~n24298 & n24309 ;
  assign n24312 = n24310 | n24311 ;
  assign n24313 = n24170 & ~n24312 ;
  assign n24314 = ~n24170 & n24312 ;
  assign n24315 = n24313 | n24314 ;
  assign n24316 = n24217 & ~n24315 ;
  assign n24317 = n24315 | n24316 ;
  assign n24318 = ( ~n24217 & n24316 ) | ( ~n24217 & n24317 ) | ( n24316 & n24317 ) ;
  assign n24319 = ~n24206 & n24318 ;
  assign n24320 = n24206 & ~n24318 ;
  assign n24321 = n24319 | n24320 ;
  assign n24322 = ( n24084 & n24086 ) | ( n24084 & ~n24192 ) | ( n24086 & ~n24192 ) ;
  assign n24323 = ~n24321 & n24322 ;
  assign n24324 = n24321 & ~n24322 ;
  assign n24325 = n24323 | n24324 ;
  assign n24326 = ~n24195 & n24204 ;
  assign n24327 = n24325 & n24326 ;
  assign n24328 = n24325 | n24326 ;
  assign n24329 = ~n24327 & n24328 ;
  assign n24330 = x127 & n6932 ;
  assign n24331 = x126 & ~n6931 ;
  assign n24332 = n7216 & n24331 ;
  assign n24333 = n24330 | n24332 ;
  assign n24334 = n6940 | n24333 ;
  assign n24335 = ( n13461 & n24333 ) | ( n13461 & n24334 ) | ( n24333 & n24334 ) ;
  assign n24336 = x47 & n24335 ;
  assign n24337 = x47 & ~n24336 ;
  assign n24338 = ( n24335 & ~n24336 ) | ( n24335 & n24337 ) | ( ~n24336 & n24337 ) ;
  assign n24339 = n24311 | n24338 ;
  assign n24340 = n24313 | n24339 ;
  assign n24341 = ( n24311 & n24313 ) | ( n24311 & n24338 ) | ( n24313 & n24338 ) ;
  assign n24342 = n24340 & ~n24341 ;
  assign n24343 = n24294 | n24296 ;
  assign n24344 = x122 & n8834 ;
  assign n24345 = x121 & n8829 ;
  assign n24346 = x120 & ~n8828 ;
  assign n24347 = n9159 & n24346 ;
  assign n24348 = n24345 | n24347 ;
  assign n24349 = n24344 | n24348 ;
  assign n24350 = n8837 | n24349 ;
  assign n24351 = ( n11188 & n24349 ) | ( n11188 & n24350 ) | ( n24349 & n24350 ) ;
  assign n24352 = x53 & n24351 ;
  assign n24353 = x53 & ~n24352 ;
  assign n24354 = ( n24351 & ~n24352 ) | ( n24351 & n24353 ) | ( ~n24352 & n24353 ) ;
  assign n24355 = n24277 | n24279 ;
  assign n24356 = x119 & n9853 ;
  assign n24357 = x118 & n9848 ;
  assign n24358 = x117 & ~n9847 ;
  assign n24359 = n10165 & n24358 ;
  assign n24360 = n24357 | n24359 ;
  assign n24361 = n24356 | n24360 ;
  assign n24362 = n9856 | n24361 ;
  assign n24363 = ( n9789 & n24361 ) | ( n9789 & n24362 ) | ( n24361 & n24362 ) ;
  assign n24364 = x56 & n24363 ;
  assign n24365 = x56 & ~n24364 ;
  assign n24366 = ( n24363 & ~n24364 ) | ( n24363 & n24365 ) | ( ~n24364 & n24365 ) ;
  assign n24389 = ( ~n24229 & n24231 ) | ( ~n24229 & n24245 ) | ( n24231 & n24245 ) ;
  assign n24367 = x113 & n11984 ;
  assign n24368 = x112 & n11979 ;
  assign n24369 = x111 & ~n11978 ;
  assign n24370 = n12430 & n24369 ;
  assign n24371 = n24368 | n24370 ;
  assign n24372 = n24367 | n24371 ;
  assign n24373 = n11987 | n24372 ;
  assign n24374 = ( n8113 & n24372 ) | ( n8113 & n24373 ) | ( n24372 & n24373 ) ;
  assign n24375 = ~x62 & n24374 ;
  assign n24376 = x110 & n12808 ;
  assign n24377 = x63 & x109 ;
  assign n24378 = ~n12808 & n24377 ;
  assign n24379 = n24376 | n24378 ;
  assign n24380 = n24224 | n24228 ;
  assign n24381 = n24379 & ~n24380 ;
  assign n24382 = ~n24379 & n24380 ;
  assign n24383 = n24381 | n24382 ;
  assign n24384 = x62 & ~n24374 ;
  assign n24385 = n24383 & ~n24384 ;
  assign n24386 = ~n24375 & n24385 ;
  assign n24387 = ( n24375 & ~n24383 ) | ( n24375 & n24384 ) | ( ~n24383 & n24384 ) ;
  assign n24388 = n24386 | n24387 ;
  assign n24390 = ~n24388 & n24389 ;
  assign n24391 = n24389 & ~n24390 ;
  assign n24392 = n24388 | n24389 ;
  assign n24393 = x116 & n10876 ;
  assign n24394 = x115 & n10871 ;
  assign n24395 = x114 & ~n10870 ;
  assign n24396 = n11305 & n24395 ;
  assign n24397 = n24394 | n24396 ;
  assign n24398 = n24393 | n24397 ;
  assign n24399 = n10879 | n24398 ;
  assign n24400 = ( n8778 & n24398 ) | ( n8778 & n24399 ) | ( n24398 & n24399 ) ;
  assign n24401 = x59 & n24400 ;
  assign n24402 = x59 & ~n24401 ;
  assign n24403 = ( n24400 & ~n24401 ) | ( n24400 & n24402 ) | ( ~n24401 & n24402 ) ;
  assign n24404 = n24392 & ~n24403 ;
  assign n24405 = ~n24391 & n24404 ;
  assign n24406 = ( n24391 & ~n24392 ) | ( n24391 & n24403 ) | ( ~n24392 & n24403 ) ;
  assign n24407 = n24405 | n24406 ;
  assign n24408 = n24260 | n24262 ;
  assign n24409 = ( n24366 & n24407 ) | ( n24366 & ~n24408 ) | ( n24407 & ~n24408 ) ;
  assign n24410 = ( ~n24407 & n24408 ) | ( ~n24407 & n24409 ) | ( n24408 & n24409 ) ;
  assign n24411 = ( ~n24366 & n24409 ) | ( ~n24366 & n24410 ) | ( n24409 & n24410 ) ;
  assign n24412 = ( n24354 & ~n24355 ) | ( n24354 & n24411 ) | ( ~n24355 & n24411 ) ;
  assign n24413 = ( n24354 & n24355 ) | ( n24354 & ~n24411 ) | ( n24355 & ~n24411 ) ;
  assign n24414 = ( ~n24354 & n24412 ) | ( ~n24354 & n24413 ) | ( n24412 & n24413 ) ;
  assign n24415 = n24343 & ~n24414 ;
  assign n24416 = n24343 & ~n24415 ;
  assign n24417 = n24414 | n24415 ;
  assign n24418 = ~n24416 & n24417 ;
  assign n24419 = x125 & n7812 ;
  assign n24420 = x124 & n7807 ;
  assign n24421 = x123 & ~n7806 ;
  assign n24422 = n8136 & n24421 ;
  assign n24423 = n24420 | n24422 ;
  assign n24424 = n24419 | n24423 ;
  assign n24425 = n7815 | n24424 ;
  assign n24426 = ( n12310 & n24424 ) | ( n12310 & n24425 ) | ( n24424 & n24425 ) ;
  assign n24427 = x50 & n24426 ;
  assign n24428 = x50 & ~n24427 ;
  assign n24429 = ( n24426 & ~n24427 ) | ( n24426 & n24428 ) | ( ~n24427 & n24428 ) ;
  assign n24430 = n24418 & n24429 ;
  assign n24431 = n24418 | n24429 ;
  assign n24432 = ~n24430 & n24431 ;
  assign n24433 = n24342 & ~n24432 ;
  assign n24434 = n24432 | n24433 ;
  assign n24435 = ( ~n24342 & n24433 ) | ( ~n24342 & n24434 ) | ( n24433 & n24434 ) ;
  assign n24436 = n24316 | n24320 ;
  assign n24437 = n24435 & ~n24436 ;
  assign n24438 = ~n24435 & n24436 ;
  assign n24439 = n24437 | n24438 ;
  assign n24440 = ~n24323 & n24328 ;
  assign n24441 = n24439 & n24440 ;
  assign n24442 = n24323 & ~n24439 ;
  assign n24443 = ( n24328 & n24439 ) | ( n24328 & ~n24442 ) | ( n24439 & ~n24442 ) ;
  assign n24444 = ~n24441 & n24443 ;
  assign n24445 = n24390 | n24406 ;
  assign n24446 = x117 & n10876 ;
  assign n24447 = x116 & n10871 ;
  assign n24448 = x115 & ~n10870 ;
  assign n24449 = n11305 & n24448 ;
  assign n24450 = n24447 | n24449 ;
  assign n24451 = n24446 | n24450 ;
  assign n24452 = n10879 | n24451 ;
  assign n24453 = ( n9118 & n24451 ) | ( n9118 & n24452 ) | ( n24451 & n24452 ) ;
  assign n24454 = x59 & n24453 ;
  assign n24455 = x59 & ~n24454 ;
  assign n24456 = ( n24453 & ~n24454 ) | ( n24453 & n24455 ) | ( ~n24454 & n24455 ) ;
  assign n24457 = x114 & n11984 ;
  assign n24458 = x113 & n11979 ;
  assign n24459 = x112 & ~n11978 ;
  assign n24460 = n12430 & n24459 ;
  assign n24461 = n24458 | n24460 ;
  assign n24462 = n24457 | n24461 ;
  assign n24463 = n11987 | n24462 ;
  assign n24464 = ( n8437 & n24462 ) | ( n8437 & n24463 ) | ( n24462 & n24463 ) ;
  assign n24465 = x62 & n24464 ;
  assign n24466 = x62 & ~n24465 ;
  assign n24467 = ( n24464 & ~n24465 ) | ( n24464 & n24466 ) | ( ~n24465 & n24466 ) ;
  assign n24468 = x111 & n12808 ;
  assign n24469 = x63 & x110 ;
  assign n24470 = ~n12808 & n24469 ;
  assign n24471 = n24468 | n24470 ;
  assign n24472 = ~n24379 & n24471 ;
  assign n24473 = n24379 & ~n24471 ;
  assign n24474 = ( n24380 & ~n24471 ) | ( n24380 & n24473 ) | ( ~n24471 & n24473 ) ;
  assign n24475 = n24472 | n24474 ;
  assign n24476 = n24387 | n24475 ;
  assign n24477 = n24472 | n24473 ;
  assign n24478 = ( n24382 & n24387 ) | ( n24382 & n24477 ) | ( n24387 & n24477 ) ;
  assign n24479 = n24476 & ~n24478 ;
  assign n24480 = ( n24456 & ~n24467 ) | ( n24456 & n24479 ) | ( ~n24467 & n24479 ) ;
  assign n24481 = ( n24467 & ~n24479 ) | ( n24467 & n24480 ) | ( ~n24479 & n24480 ) ;
  assign n24482 = ( ~n24456 & n24480 ) | ( ~n24456 & n24481 ) | ( n24480 & n24481 ) ;
  assign n24483 = n24445 & ~n24482 ;
  assign n24484 = n24445 & ~n24483 ;
  assign n24485 = n24482 | n24483 ;
  assign n24486 = ~n24484 & n24485 ;
  assign n24487 = x120 & n9853 ;
  assign n24488 = x119 & n9848 ;
  assign n24489 = x118 & ~n9847 ;
  assign n24490 = n10165 & n24489 ;
  assign n24491 = n24488 | n24490 ;
  assign n24492 = n24487 | n24491 ;
  assign n24493 = n9856 | n24492 ;
  assign n24494 = ( n10460 & n24492 ) | ( n10460 & n24493 ) | ( n24492 & n24493 ) ;
  assign n24495 = x56 & n24494 ;
  assign n24496 = x56 & ~n24495 ;
  assign n24497 = ( n24494 & ~n24495 ) | ( n24494 & n24496 ) | ( ~n24495 & n24496 ) ;
  assign n24498 = ( n24410 & n24486 ) | ( n24410 & ~n24497 ) | ( n24486 & ~n24497 ) ;
  assign n24499 = ( ~n24486 & n24497 ) | ( ~n24486 & n24498 ) | ( n24497 & n24498 ) ;
  assign n24500 = ( ~n24410 & n24498 ) | ( ~n24410 & n24499 ) | ( n24498 & n24499 ) ;
  assign n24501 = x123 & n8834 ;
  assign n24502 = x122 & n8829 ;
  assign n24503 = x121 & ~n8828 ;
  assign n24504 = n9159 & n24503 ;
  assign n24505 = n24502 | n24504 ;
  assign n24506 = n24501 | n24505 ;
  assign n24507 = n8837 | n24506 ;
  assign n24508 = ( n11219 & n24506 ) | ( n11219 & n24507 ) | ( n24506 & n24507 ) ;
  assign n24509 = x53 & n24508 ;
  assign n24510 = x53 & ~n24509 ;
  assign n24511 = ( n24508 & ~n24509 ) | ( n24508 & n24510 ) | ( ~n24509 & n24510 ) ;
  assign n24512 = n24500 | n24511 ;
  assign n24513 = ~n24511 & n24512 ;
  assign n24514 = ( ~n24500 & n24512 ) | ( ~n24500 & n24513 ) | ( n24512 & n24513 ) ;
  assign n24515 = n24413 & ~n24514 ;
  assign n24516 = n24514 | n24515 ;
  assign n24517 = n24413 & n24514 ;
  assign n24518 = n24516 & ~n24517 ;
  assign n24519 = x126 & n7812 ;
  assign n24520 = x125 & n7807 ;
  assign n24521 = x124 & ~n7806 ;
  assign n24522 = n8136 & n24521 ;
  assign n24523 = n24520 | n24522 ;
  assign n24524 = n24519 | n24523 ;
  assign n24525 = n7815 | n24524 ;
  assign n24526 = ( n12687 & n24524 ) | ( n12687 & n24525 ) | ( n24524 & n24525 ) ;
  assign n24527 = x50 & n24526 ;
  assign n24528 = x50 & ~n24527 ;
  assign n24529 = ( n24526 & ~n24527 ) | ( n24526 & n24528 ) | ( ~n24527 & n24528 ) ;
  assign n24530 = ~n24518 & n24529 ;
  assign n24531 = n24518 & ~n24529 ;
  assign n24532 = n24530 | n24531 ;
  assign n24533 = x127 & ~n6931 ;
  assign n24534 = n7216 & n24533 ;
  assign n24535 = ( x127 & n6940 ) | ( x127 & n24534 ) | ( n6940 & n24534 ) ;
  assign n24536 = ( x126 & n24534 ) | ( x126 & n24535 ) | ( n24534 & n24535 ) ;
  assign n24537 = ( n12685 & n24535 ) | ( n12685 & n24536 ) | ( n24535 & n24536 ) ;
  assign n24538 = x47 & n24537 ;
  assign n24539 = x47 & ~n24538 ;
  assign n24540 = ( n24537 & ~n24538 ) | ( n24537 & n24539 ) | ( ~n24538 & n24539 ) ;
  assign n24541 = ( n24415 & ~n24418 ) | ( n24415 & n24431 ) | ( ~n24418 & n24431 ) ;
  assign n24542 = n24540 & n24541 ;
  assign n24543 = n24540 | n24541 ;
  assign n24544 = ~n24542 & n24543 ;
  assign n24545 = ~n24532 & n24544 ;
  assign n24546 = n24532 | n24545 ;
  assign n24547 = n24544 & ~n24545 ;
  assign n24548 = n24546 & ~n24547 ;
  assign n24549 = n24341 | n24433 ;
  assign n24550 = n24548 & ~n24549 ;
  assign n24551 = ~n24548 & n24549 ;
  assign n24552 = n24550 | n24551 ;
  assign n24553 = n24438 | n24442 ;
  assign n24554 = ( n24328 & n24437 ) | ( n24328 & ~n24553 ) | ( n24437 & ~n24553 ) ;
  assign n24555 = n24552 & n24554 ;
  assign n24556 = ~n24552 & n24553 ;
  assign n24557 = n24437 | n24552 ;
  assign n24558 = ( n24328 & ~n24556 ) | ( n24328 & n24557 ) | ( ~n24556 & n24557 ) ;
  assign n24559 = ~n24555 & n24558 ;
  assign n24560 = n24515 | n24530 ;
  assign n24561 = x127 & n7812 ;
  assign n24562 = x126 & n7807 ;
  assign n24563 = x125 & ~n7806 ;
  assign n24564 = n8136 & n24563 ;
  assign n24565 = n24562 | n24564 ;
  assign n24566 = n24561 | n24565 ;
  assign n24567 = n7815 | n24566 ;
  assign n24568 = ( n12720 & n24566 ) | ( n12720 & n24567 ) | ( n24566 & n24567 ) ;
  assign n24569 = x50 & n24568 ;
  assign n24570 = x50 & ~n24569 ;
  assign n24571 = ( n24568 & ~n24569 ) | ( n24568 & n24570 ) | ( ~n24569 & n24570 ) ;
  assign n24572 = ( n24387 & ~n24472 ) | ( n24387 & n24474 ) | ( ~n24472 & n24474 ) ;
  assign n24573 = x115 & n11984 ;
  assign n24574 = x114 & n11979 ;
  assign n24575 = x113 & ~n11978 ;
  assign n24576 = n12430 & n24575 ;
  assign n24577 = n24574 | n24576 ;
  assign n24578 = n24573 | n24577 ;
  assign n24579 = n11987 | n24578 ;
  assign n24580 = ( n8749 & n24578 ) | ( n8749 & n24579 ) | ( n24578 & n24579 ) ;
  assign n24581 = ~x62 & n24580 ;
  assign n24582 = x62 & ~n24580 ;
  assign n24583 = n24581 | n24582 ;
  assign n24584 = x112 & n12808 ;
  assign n24585 = x63 & x111 ;
  assign n24586 = ~n12808 & n24585 ;
  assign n24587 = n24584 | n24586 ;
  assign n24588 = ( x47 & ~n24471 ) | ( x47 & n24587 ) | ( ~n24471 & n24587 ) ;
  assign n24589 = ( ~x47 & n24471 ) | ( ~x47 & n24587 ) | ( n24471 & n24587 ) ;
  assign n24590 = ( ~n24587 & n24588 ) | ( ~n24587 & n24589 ) | ( n24588 & n24589 ) ;
  assign n24591 = n24583 & ~n24590 ;
  assign n24592 = ~n24583 & n24590 ;
  assign n24593 = n24591 | n24592 ;
  assign n24594 = n24572 | n24593 ;
  assign n24595 = n24572 & n24593 ;
  assign n24596 = x118 & n10876 ;
  assign n24597 = x117 & n10871 ;
  assign n24598 = x116 & ~n10870 ;
  assign n24599 = n11305 & n24598 ;
  assign n24600 = n24597 | n24599 ;
  assign n24601 = n24596 | n24600 ;
  assign n24602 = n10879 | n24601 ;
  assign n24603 = ( n9760 & n24601 ) | ( n9760 & n24602 ) | ( n24601 & n24602 ) ;
  assign n24604 = x59 & n24603 ;
  assign n24605 = x59 & ~n24604 ;
  assign n24606 = ( n24603 & ~n24604 ) | ( n24603 & n24605 ) | ( ~n24604 & n24605 ) ;
  assign n24607 = n24595 | n24606 ;
  assign n24608 = n24594 & ~n24607 ;
  assign n24609 = ( ~n24594 & n24595 ) | ( ~n24594 & n24606 ) | ( n24595 & n24606 ) ;
  assign n24610 = n24608 | n24609 ;
  assign n24611 = n24481 & ~n24610 ;
  assign n24612 = ~n24481 & n24610 ;
  assign n24613 = n24611 | n24612 ;
  assign n24614 = x121 & n9853 ;
  assign n24615 = x120 & n9848 ;
  assign n24616 = x119 & ~n9847 ;
  assign n24617 = n10165 & n24616 ;
  assign n24618 = n24615 | n24617 ;
  assign n24619 = n24614 | n24618 ;
  assign n24620 = n9856 | n24619 ;
  assign n24621 = ( n10811 & n24619 ) | ( n10811 & n24620 ) | ( n24619 & n24620 ) ;
  assign n24622 = x56 & n24621 ;
  assign n24623 = x56 & ~n24622 ;
  assign n24624 = ( n24621 & ~n24622 ) | ( n24621 & n24623 ) | ( ~n24622 & n24623 ) ;
  assign n24625 = n24613 & ~n24624 ;
  assign n24626 = ~n24613 & n24624 ;
  assign n24627 = n24625 | n24626 ;
  assign n24628 = ~n24486 & n24497 ;
  assign n24629 = n24483 | n24628 ;
  assign n24630 = ~n24627 & n24629 ;
  assign n24631 = n24627 & ~n24629 ;
  assign n24632 = n24630 | n24631 ;
  assign n24633 = x124 & n8834 ;
  assign n24634 = x123 & n8829 ;
  assign n24635 = x122 & ~n8828 ;
  assign n24636 = n9159 & n24635 ;
  assign n24637 = n24634 | n24636 ;
  assign n24638 = n24633 | n24637 ;
  assign n24639 = n8837 | n24638 ;
  assign n24640 = ( n11916 & n24638 ) | ( n11916 & n24639 ) | ( n24638 & n24639 ) ;
  assign n24641 = x53 & n24640 ;
  assign n24642 = x53 & ~n24641 ;
  assign n24643 = ( n24640 & ~n24641 ) | ( n24640 & n24642 ) | ( ~n24641 & n24642 ) ;
  assign n24644 = n24632 & ~n24643 ;
  assign n24645 = ~n24632 & n24643 ;
  assign n24646 = n24644 | n24645 ;
  assign n24647 = ( n24410 & n24511 ) | ( n24410 & n24514 ) | ( n24511 & n24514 ) ;
  assign n24648 = ~n24646 & n24647 ;
  assign n24649 = n24646 & ~n24647 ;
  assign n24650 = n24648 | n24649 ;
  assign n24651 = n24571 & ~n24650 ;
  assign n24652 = n24650 | n24651 ;
  assign n24653 = ( ~n24571 & n24651 ) | ( ~n24571 & n24652 ) | ( n24651 & n24652 ) ;
  assign n24654 = ~n24560 & n24653 ;
  assign n24655 = n24560 & ~n24653 ;
  assign n24656 = n24654 | n24655 ;
  assign n24657 = n24542 | n24545 ;
  assign n24658 = n24656 & ~n24657 ;
  assign n24659 = ~n24656 & n24657 ;
  assign n24660 = n24658 | n24659 ;
  assign n24661 = n24551 | n24556 ;
  assign n24662 = ~n24551 & n24557 ;
  assign n24663 = ( n24328 & ~n24661 ) | ( n24328 & n24662 ) | ( ~n24661 & n24662 ) ;
  assign n24664 = n24660 & n24663 ;
  assign n24665 = ~n24660 & n24661 ;
  assign n24666 = n24660 | n24662 ;
  assign n24667 = ( n24328 & ~n24665 ) | ( n24328 & n24666 ) | ( ~n24665 & n24666 ) ;
  assign n24668 = ~n24664 & n24667 ;
  assign n24669 = n24651 | n24655 ;
  assign n24670 = x127 & n7807 ;
  assign n24671 = x126 & ~n7806 ;
  assign n24672 = n8136 & n24671 ;
  assign n24673 = n24670 | n24672 ;
  assign n24674 = n7815 | n24673 ;
  assign n24675 = ( n13461 & n24673 ) | ( n13461 & n24674 ) | ( n24673 & n24674 ) ;
  assign n24676 = x50 & n24675 ;
  assign n24677 = x50 & ~n24676 ;
  assign n24678 = ( n24675 & ~n24676 ) | ( n24675 & n24677 ) | ( ~n24676 & n24677 ) ;
  assign n24679 = n24645 | n24648 ;
  assign n24680 = x125 & n8834 ;
  assign n24681 = x124 & n8829 ;
  assign n24682 = x123 & ~n8828 ;
  assign n24683 = n9159 & n24682 ;
  assign n24684 = n24681 | n24683 ;
  assign n24685 = n24680 | n24684 ;
  assign n24686 = n8837 | n24685 ;
  assign n24687 = ( n12310 & n24685 ) | ( n12310 & n24686 ) | ( n24685 & n24686 ) ;
  assign n24688 = x53 & n24687 ;
  assign n24689 = x53 & ~n24688 ;
  assign n24690 = ( n24687 & ~n24688 ) | ( n24687 & n24689 ) | ( ~n24688 & n24689 ) ;
  assign n24691 = n24626 | n24630 ;
  assign n24692 = ( n24572 & n24583 ) | ( n24572 & ~n24590 ) | ( n24583 & ~n24590 ) ;
  assign n24693 = x113 & n12808 ;
  assign n24694 = x63 & x112 ;
  assign n24695 = ~n12808 & n24694 ;
  assign n24696 = n24693 | n24695 ;
  assign n24697 = n24589 & ~n24696 ;
  assign n24698 = ~n24589 & n24696 ;
  assign n24699 = n24697 | n24698 ;
  assign n24700 = x116 & n11984 ;
  assign n24701 = x115 & n11979 ;
  assign n24702 = x114 & ~n11978 ;
  assign n24703 = n12430 & n24702 ;
  assign n24704 = n24701 | n24703 ;
  assign n24705 = n24700 | n24704 ;
  assign n24706 = n11987 | n24705 ;
  assign n24707 = ( n8778 & n24705 ) | ( n8778 & n24706 ) | ( n24705 & n24706 ) ;
  assign n24708 = x62 & n24707 ;
  assign n24709 = x62 & ~n24708 ;
  assign n24710 = ( n24707 & ~n24708 ) | ( n24707 & n24709 ) | ( ~n24708 & n24709 ) ;
  assign n24711 = ~n24699 & n24710 ;
  assign n24712 = n24699 & ~n24710 ;
  assign n24713 = n24711 | n24712 ;
  assign n24714 = n24692 & ~n24713 ;
  assign n24715 = n24692 & ~n24714 ;
  assign n24716 = n24692 | n24713 ;
  assign n24717 = x119 & n10876 ;
  assign n24718 = x118 & n10871 ;
  assign n24719 = x117 & ~n10870 ;
  assign n24720 = n11305 & n24719 ;
  assign n24721 = n24718 | n24720 ;
  assign n24722 = n24717 | n24721 ;
  assign n24723 = n10879 | n24722 ;
  assign n24724 = ( n9789 & n24722 ) | ( n9789 & n24723 ) | ( n24722 & n24723 ) ;
  assign n24725 = x59 & n24724 ;
  assign n24726 = x59 & ~n24725 ;
  assign n24727 = ( n24724 & ~n24725 ) | ( n24724 & n24726 ) | ( ~n24725 & n24726 ) ;
  assign n24728 = n24716 & ~n24727 ;
  assign n24729 = ~n24715 & n24728 ;
  assign n24730 = ( n24715 & ~n24716 ) | ( n24715 & n24727 ) | ( ~n24716 & n24727 ) ;
  assign n24731 = n24729 | n24730 ;
  assign n24732 = n24609 | n24611 ;
  assign n24733 = ~n24731 & n24732 ;
  assign n24734 = n24731 & ~n24732 ;
  assign n24735 = n24733 | n24734 ;
  assign n24736 = x122 & n9853 ;
  assign n24737 = x121 & n9848 ;
  assign n24738 = x120 & ~n9847 ;
  assign n24739 = n10165 & n24738 ;
  assign n24740 = n24737 | n24739 ;
  assign n24741 = n24736 | n24740 ;
  assign n24742 = n9856 | n24741 ;
  assign n24743 = ( n11188 & n24741 ) | ( n11188 & n24742 ) | ( n24741 & n24742 ) ;
  assign n24744 = x56 & n24743 ;
  assign n24745 = x56 & ~n24744 ;
  assign n24746 = ( n24743 & ~n24744 ) | ( n24743 & n24745 ) | ( ~n24744 & n24745 ) ;
  assign n24747 = ~n24735 & n24746 ;
  assign n24748 = n24735 & ~n24746 ;
  assign n24749 = n24747 | n24748 ;
  assign n24750 = ( n24690 & n24691 ) | ( n24690 & ~n24749 ) | ( n24691 & ~n24749 ) ;
  assign n24751 = ( ~n24691 & n24749 ) | ( ~n24691 & n24750 ) | ( n24749 & n24750 ) ;
  assign n24752 = ( ~n24690 & n24750 ) | ( ~n24690 & n24751 ) | ( n24750 & n24751 ) ;
  assign n24753 = ( n24678 & ~n24679 ) | ( n24678 & n24752 ) | ( ~n24679 & n24752 ) ;
  assign n24754 = ( n24679 & ~n24752 ) | ( n24679 & n24753 ) | ( ~n24752 & n24753 ) ;
  assign n24755 = ( ~n24678 & n24753 ) | ( ~n24678 & n24754 ) | ( n24753 & n24754 ) ;
  assign n24756 = ~n24669 & n24755 ;
  assign n24757 = n24669 & ~n24755 ;
  assign n24758 = n24756 | n24757 ;
  assign n24759 = n24659 | n24665 ;
  assign n24760 = ~n24659 & n24666 ;
  assign n24761 = ( n24328 & ~n24759 ) | ( n24328 & n24760 ) | ( ~n24759 & n24760 ) ;
  assign n24762 = n24758 & n24761 ;
  assign n24763 = ~n24758 & n24759 ;
  assign n24764 = n24758 | n24760 ;
  assign n24765 = ( n24328 & ~n24763 ) | ( n24328 & n24764 ) | ( ~n24763 & n24764 ) ;
  assign n24766 = ~n24762 & n24765 ;
  assign n24767 = n24691 & ~n24749 ;
  assign n24768 = n24750 & ~n24767 ;
  assign n24769 = x127 & ~n7806 ;
  assign n24770 = n8136 & n24769 ;
  assign n24771 = ( x127 & n7815 ) | ( x127 & n24770 ) | ( n7815 & n24770 ) ;
  assign n24772 = ( x126 & n24770 ) | ( x126 & n24771 ) | ( n24770 & n24771 ) ;
  assign n24773 = ( n12685 & n24771 ) | ( n12685 & n24772 ) | ( n24771 & n24772 ) ;
  assign n24774 = x50 & n24773 ;
  assign n24775 = x50 & ~n24774 ;
  assign n24776 = ( n24773 & ~n24774 ) | ( n24773 & n24775 ) | ( ~n24774 & n24775 ) ;
  assign n24777 = n24767 | n24776 ;
  assign n24778 = n24768 | n24777 ;
  assign n24779 = ( n24767 & n24768 ) | ( n24767 & n24776 ) | ( n24768 & n24776 ) ;
  assign n24780 = n24778 & ~n24779 ;
  assign n24781 = n24733 | n24747 ;
  assign n24782 = n24714 | n24730 ;
  assign n24783 = x117 & n11984 ;
  assign n24784 = x116 & n11979 ;
  assign n24785 = x115 & ~n11978 ;
  assign n24786 = n12430 & n24785 ;
  assign n24787 = n24784 | n24786 ;
  assign n24788 = n24783 | n24787 ;
  assign n24789 = n11987 | n24788 ;
  assign n24790 = ( n9118 & n24788 ) | ( n9118 & n24789 ) | ( n24788 & n24789 ) ;
  assign n24791 = ~x62 & n24790 ;
  assign n24792 = x62 & ~n24790 ;
  assign n24793 = n24791 | n24792 ;
  assign n24794 = x114 & n12808 ;
  assign n24795 = x63 & x113 ;
  assign n24796 = ~n12808 & n24795 ;
  assign n24797 = n24794 | n24796 ;
  assign n24798 = ~n24696 & n24797 ;
  assign n24799 = n24696 | n24798 ;
  assign n24800 = n24797 & ~n24798 ;
  assign n24801 = n24799 & ~n24800 ;
  assign n24802 = n24793 & ~n24801 ;
  assign n24803 = ~n24793 & n24801 ;
  assign n24804 = n24802 | n24803 ;
  assign n24805 = n24697 | n24711 ;
  assign n24806 = n24804 & ~n24805 ;
  assign n24807 = ~n24804 & n24805 ;
  assign n24808 = n24806 | n24807 ;
  assign n24809 = x120 & n10876 ;
  assign n24810 = x119 & n10871 ;
  assign n24811 = x118 & ~n10870 ;
  assign n24812 = n11305 & n24811 ;
  assign n24813 = n24810 | n24812 ;
  assign n24814 = n24809 | n24813 ;
  assign n24815 = n10879 | n24814 ;
  assign n24816 = ( n10460 & n24814 ) | ( n10460 & n24815 ) | ( n24814 & n24815 ) ;
  assign n24817 = x59 & n24816 ;
  assign n24818 = x59 & ~n24817 ;
  assign n24819 = ( n24816 & ~n24817 ) | ( n24816 & n24818 ) | ( ~n24817 & n24818 ) ;
  assign n24820 = n24808 & ~n24819 ;
  assign n24821 = ~n24808 & n24819 ;
  assign n24822 = n24820 | n24821 ;
  assign n24823 = n24782 & ~n24822 ;
  assign n24824 = ~n24782 & n24822 ;
  assign n24825 = n24823 | n24824 ;
  assign n24826 = x123 & n9853 ;
  assign n24827 = x122 & n9848 ;
  assign n24828 = x121 & ~n9847 ;
  assign n24829 = n10165 & n24828 ;
  assign n24830 = n24827 | n24829 ;
  assign n24831 = n24826 | n24830 ;
  assign n24832 = n9856 | n24831 ;
  assign n24833 = ( n11219 & n24831 ) | ( n11219 & n24832 ) | ( n24831 & n24832 ) ;
  assign n24834 = x56 & n24833 ;
  assign n24835 = x56 & ~n24834 ;
  assign n24836 = ( n24833 & ~n24834 ) | ( n24833 & n24835 ) | ( ~n24834 & n24835 ) ;
  assign n24837 = ( n24781 & n24825 ) | ( n24781 & ~n24836 ) | ( n24825 & ~n24836 ) ;
  assign n24838 = ( ~n24825 & n24836 ) | ( ~n24825 & n24837 ) | ( n24836 & n24837 ) ;
  assign n24839 = ( ~n24781 & n24837 ) | ( ~n24781 & n24838 ) | ( n24837 & n24838 ) ;
  assign n24840 = x126 & n8834 ;
  assign n24841 = x125 & n8829 ;
  assign n24842 = x124 & ~n8828 ;
  assign n24843 = n9159 & n24842 ;
  assign n24844 = n24841 | n24843 ;
  assign n24845 = n24840 | n24844 ;
  assign n24846 = n8837 | n24845 ;
  assign n24847 = ( n12687 & n24845 ) | ( n12687 & n24846 ) | ( n24845 & n24846 ) ;
  assign n24848 = x53 & n24847 ;
  assign n24849 = x53 & ~n24848 ;
  assign n24850 = ( n24847 & ~n24848 ) | ( n24847 & n24849 ) | ( ~n24848 & n24849 ) ;
  assign n24851 = n24839 | n24850 ;
  assign n24852 = ~n24850 & n24851 ;
  assign n24853 = ( ~n24839 & n24851 ) | ( ~n24839 & n24852 ) | ( n24851 & n24852 ) ;
  assign n24854 = n24780 & ~n24853 ;
  assign n24855 = n24853 | n24854 ;
  assign n24856 = ( ~n24780 & n24854 ) | ( ~n24780 & n24855 ) | ( n24854 & n24855 ) ;
  assign n24857 = ~n24754 & n24856 ;
  assign n24858 = n24754 & ~n24856 ;
  assign n24859 = n24857 | n24858 ;
  assign n24860 = n24757 | n24763 ;
  assign n24861 = ~n24757 & n24764 ;
  assign n24862 = ( n24328 & ~n24860 ) | ( n24328 & n24861 ) | ( ~n24860 & n24861 ) ;
  assign n24863 = n24859 & n24862 ;
  assign n24864 = ~n24859 & n24860 ;
  assign n24865 = n24859 | n24861 ;
  assign n24866 = ( n24328 & ~n24864 ) | ( n24328 & n24865 ) | ( ~n24864 & n24865 ) ;
  assign n24867 = ~n24863 & n24866 ;
  assign n24868 = ( n24781 & n24850 ) | ( n24781 & n24853 ) | ( n24850 & n24853 ) ;
  assign n24869 = x127 & n8834 ;
  assign n24870 = x126 & n8829 ;
  assign n24871 = x125 & ~n8828 ;
  assign n24872 = n9159 & n24871 ;
  assign n24873 = n24870 | n24872 ;
  assign n24874 = n24869 | n24873 ;
  assign n24875 = n8837 | n24874 ;
  assign n24876 = ( n12720 & n24874 ) | ( n12720 & n24875 ) | ( n24874 & n24875 ) ;
  assign n24877 = x53 & n24876 ;
  assign n24878 = x53 & ~n24877 ;
  assign n24879 = ( n24876 & ~n24877 ) | ( n24876 & n24878 ) | ( ~n24877 & n24878 ) ;
  assign n24880 = n24798 | n24802 ;
  assign n24881 = x115 & n12808 ;
  assign n24882 = x63 & x114 ;
  assign n24883 = ~n12808 & n24882 ;
  assign n24884 = n24881 | n24883 ;
  assign n24885 = ~x50 & n24884 ;
  assign n24886 = x50 & ~n24884 ;
  assign n24887 = n24885 | n24886 ;
  assign n24888 = n24696 & ~n24887 ;
  assign n24889 = ~n24696 & n24887 ;
  assign n24890 = n24888 | n24889 ;
  assign n24891 = n24798 & ~n24890 ;
  assign n24892 = ( n24802 & ~n24890 ) | ( n24802 & n24891 ) | ( ~n24890 & n24891 ) ;
  assign n24893 = n24880 & ~n24892 ;
  assign n24894 = n24890 | n24891 ;
  assign n24895 = n24802 | n24894 ;
  assign n24896 = x118 & n11984 ;
  assign n24897 = x117 & n11979 ;
  assign n24898 = x116 & ~n11978 ;
  assign n24899 = n12430 & n24898 ;
  assign n24900 = n24897 | n24899 ;
  assign n24901 = n24896 | n24900 ;
  assign n24902 = n11987 | n24901 ;
  assign n24903 = ( n9760 & n24901 ) | ( n9760 & n24902 ) | ( n24901 & n24902 ) ;
  assign n24904 = x62 & n24903 ;
  assign n24905 = x62 & ~n24904 ;
  assign n24906 = ( n24903 & ~n24904 ) | ( n24903 & n24905 ) | ( ~n24904 & n24905 ) ;
  assign n24907 = n24895 & ~n24906 ;
  assign n24908 = ~n24893 & n24907 ;
  assign n24909 = ( n24893 & ~n24895 ) | ( n24893 & n24906 ) | ( ~n24895 & n24906 ) ;
  assign n24910 = n24908 | n24909 ;
  assign n24911 = x121 & n10876 ;
  assign n24912 = x120 & n10871 ;
  assign n24913 = x119 & ~n10870 ;
  assign n24914 = n11305 & n24913 ;
  assign n24915 = n24912 | n24914 ;
  assign n24916 = n24911 | n24915 ;
  assign n24917 = n10879 | n24916 ;
  assign n24918 = ( n10811 & n24916 ) | ( n10811 & n24917 ) | ( n24916 & n24917 ) ;
  assign n24919 = x59 & n24918 ;
  assign n24920 = x59 & ~n24919 ;
  assign n24921 = ( n24918 & ~n24919 ) | ( n24918 & n24920 ) | ( ~n24919 & n24920 ) ;
  assign n24922 = ~n24910 & n24921 ;
  assign n24923 = n24910 | n24922 ;
  assign n24924 = n24910 & n24921 ;
  assign n24925 = n24807 | n24821 ;
  assign n24926 = n24924 | n24925 ;
  assign n24927 = n24923 & ~n24926 ;
  assign n24928 = ( ~n24923 & n24924 ) | ( ~n24923 & n24925 ) | ( n24924 & n24925 ) ;
  assign n24929 = n24927 | n24928 ;
  assign n24930 = x124 & n9853 ;
  assign n24931 = x123 & n9848 ;
  assign n24932 = x122 & ~n9847 ;
  assign n24933 = n10165 & n24932 ;
  assign n24934 = n24931 | n24933 ;
  assign n24935 = n24930 | n24934 ;
  assign n24936 = n9856 | n24935 ;
  assign n24937 = ( n11916 & n24935 ) | ( n11916 & n24936 ) | ( n24935 & n24936 ) ;
  assign n24938 = x56 & n24937 ;
  assign n24939 = x56 & ~n24938 ;
  assign n24940 = ( n24937 & ~n24938 ) | ( n24937 & n24939 ) | ( ~n24938 & n24939 ) ;
  assign n24941 = ~n24929 & n24940 ;
  assign n24942 = n24929 & ~n24940 ;
  assign n24943 = n24941 | n24942 ;
  assign n24944 = ~n24825 & n24836 ;
  assign n24945 = n24823 | n24944 ;
  assign n24946 = ~n24943 & n24945 ;
  assign n24947 = n24943 & ~n24945 ;
  assign n24948 = n24946 | n24947 ;
  assign n24949 = n24879 & ~n24948 ;
  assign n24950 = n24948 | n24949 ;
  assign n24951 = ( ~n24879 & n24949 ) | ( ~n24879 & n24950 ) | ( n24949 & n24950 ) ;
  assign n24952 = ~n24868 & n24951 ;
  assign n24953 = n24868 & ~n24951 ;
  assign n24954 = n24952 | n24953 ;
  assign n24955 = n24779 | n24854 ;
  assign n24956 = n24954 & ~n24955 ;
  assign n24957 = ~n24954 & n24955 ;
  assign n24958 = n24956 | n24957 ;
  assign n24959 = n24858 | n24864 ;
  assign n24960 = ~n24858 & n24865 ;
  assign n24961 = ( n24328 & ~n24959 ) | ( n24328 & n24960 ) | ( ~n24959 & n24960 ) ;
  assign n24962 = n24958 & n24961 ;
  assign n24963 = ~n24958 & n24959 ;
  assign n24964 = n24958 | n24960 ;
  assign n24965 = ( n24328 & ~n24963 ) | ( n24328 & n24964 ) | ( ~n24963 & n24964 ) ;
  assign n24966 = ~n24962 & n24965 ;
  assign n24967 = n24949 | n24953 ;
  assign n24968 = x127 & n8829 ;
  assign n24969 = x126 & ~n8828 ;
  assign n24970 = n9159 & n24969 ;
  assign n24971 = n24968 | n24970 ;
  assign n24972 = n8837 | n24971 ;
  assign n24973 = ( n13461 & n24971 ) | ( n13461 & n24972 ) | ( n24971 & n24972 ) ;
  assign n24974 = x53 & n24973 ;
  assign n24975 = x53 & ~n24974 ;
  assign n24976 = ( n24973 & ~n24974 ) | ( n24973 & n24975 ) | ( ~n24974 & n24975 ) ;
  assign n24977 = n24941 | n24946 ;
  assign n24978 = x125 & n9853 ;
  assign n24979 = x124 & n9848 ;
  assign n24980 = x123 & ~n9847 ;
  assign n24981 = n10165 & n24980 ;
  assign n24982 = n24979 | n24981 ;
  assign n24983 = n24978 | n24982 ;
  assign n24984 = n9856 | n24983 ;
  assign n24985 = ( n12310 & n24983 ) | ( n12310 & n24984 ) | ( n24983 & n24984 ) ;
  assign n24986 = x56 & n24985 ;
  assign n24987 = x56 & ~n24986 ;
  assign n24988 = ( n24985 & ~n24986 ) | ( n24985 & n24987 ) | ( ~n24986 & n24987 ) ;
  assign n24989 = n24922 | n24928 ;
  assign n24990 = x119 & n11984 ;
  assign n24991 = x118 & n11979 ;
  assign n24992 = x117 & ~n11978 ;
  assign n24993 = n12430 & n24992 ;
  assign n24994 = n24991 | n24993 ;
  assign n24995 = n24990 | n24994 ;
  assign n24996 = n11987 | n24995 ;
  assign n24997 = ( n9789 & n24995 ) | ( n9789 & n24996 ) | ( n24995 & n24996 ) ;
  assign n24998 = ~x62 & n24997 ;
  assign n24999 = x116 & n12808 ;
  assign n25000 = x63 & x115 ;
  assign n25001 = ~n12808 & n25000 ;
  assign n25002 = n24999 | n25001 ;
  assign n25003 = n24885 | n24888 ;
  assign n25004 = n25002 & ~n25003 ;
  assign n25005 = ~n25002 & n25003 ;
  assign n25006 = n25004 | n25005 ;
  assign n25007 = x62 & ~n24997 ;
  assign n25008 = n25006 & ~n25007 ;
  assign n25009 = ~n24998 & n25008 ;
  assign n25010 = ( n24998 & ~n25006 ) | ( n24998 & n25007 ) | ( ~n25006 & n25007 ) ;
  assign n25011 = n25009 | n25010 ;
  assign n25012 = n24892 & ~n25011 ;
  assign n25013 = ( n24909 & ~n25011 ) | ( n24909 & n25012 ) | ( ~n25011 & n25012 ) ;
  assign n25014 = ~n24892 & n25011 ;
  assign n25015 = ~n24909 & n25014 ;
  assign n25016 = n25013 | n25015 ;
  assign n25017 = x122 & n10876 ;
  assign n25018 = x121 & n10871 ;
  assign n25019 = x120 & ~n10870 ;
  assign n25020 = n11305 & n25019 ;
  assign n25021 = n25018 | n25020 ;
  assign n25022 = n25017 | n25021 ;
  assign n25023 = n10879 | n25022 ;
  assign n25024 = ( n11188 & n25022 ) | ( n11188 & n25023 ) | ( n25022 & n25023 ) ;
  assign n25025 = x59 & n25024 ;
  assign n25026 = x59 & ~n25025 ;
  assign n25027 = ( n25024 & ~n25025 ) | ( n25024 & n25026 ) | ( ~n25025 & n25026 ) ;
  assign n25028 = ~n25016 & n25027 ;
  assign n25029 = n25016 & ~n25027 ;
  assign n25030 = n25028 | n25029 ;
  assign n25031 = ( n24988 & n24989 ) | ( n24988 & ~n25030 ) | ( n24989 & ~n25030 ) ;
  assign n25032 = ( ~n24989 & n25030 ) | ( ~n24989 & n25031 ) | ( n25030 & n25031 ) ;
  assign n25033 = ( ~n24988 & n25031 ) | ( ~n24988 & n25032 ) | ( n25031 & n25032 ) ;
  assign n25034 = ( n24976 & n24977 ) | ( n24976 & ~n25033 ) | ( n24977 & ~n25033 ) ;
  assign n25035 = ( ~n24977 & n25033 ) | ( ~n24977 & n25034 ) | ( n25033 & n25034 ) ;
  assign n25036 = ( ~n24976 & n25034 ) | ( ~n24976 & n25035 ) | ( n25034 & n25035 ) ;
  assign n25037 = ~n24967 & n25036 ;
  assign n25038 = n24967 & ~n25036 ;
  assign n25039 = n25037 | n25038 ;
  assign n25040 = n24957 | n24963 ;
  assign n25041 = ~n24957 & n24964 ;
  assign n25042 = ( n24328 & ~n25040 ) | ( n24328 & n25041 ) | ( ~n25040 & n25041 ) ;
  assign n25043 = n25039 & n25042 ;
  assign n25044 = ~n25039 & n25040 ;
  assign n25045 = n25039 | n25041 ;
  assign n25046 = ( n24328 & ~n25044 ) | ( n24328 & n25045 ) | ( ~n25044 & n25045 ) ;
  assign n25047 = ~n25043 & n25046 ;
  assign n25048 = n24989 & ~n25030 ;
  assign n25049 = n25031 & ~n25048 ;
  assign n25050 = x127 & ~n8828 ;
  assign n25051 = n9159 & n25050 ;
  assign n25052 = ( x127 & n8837 ) | ( x127 & n25051 ) | ( n8837 & n25051 ) ;
  assign n25053 = ( x126 & n25051 ) | ( x126 & n25052 ) | ( n25051 & n25052 ) ;
  assign n25054 = ( n12685 & n25052 ) | ( n12685 & n25053 ) | ( n25052 & n25053 ) ;
  assign n25055 = x53 & n25054 ;
  assign n25056 = x53 & ~n25055 ;
  assign n25057 = ( n25054 & ~n25055 ) | ( n25054 & n25056 ) | ( ~n25055 & n25056 ) ;
  assign n25058 = n25048 | n25057 ;
  assign n25059 = n25049 | n25058 ;
  assign n25060 = ( n25048 & n25049 ) | ( n25048 & n25057 ) | ( n25049 & n25057 ) ;
  assign n25061 = n25059 & ~n25060 ;
  assign n25062 = n25013 | n25028 ;
  assign n25063 = x123 & n10876 ;
  assign n25064 = x122 & n10871 ;
  assign n25065 = x121 & ~n10870 ;
  assign n25066 = n11305 & n25065 ;
  assign n25067 = n25064 | n25066 ;
  assign n25068 = n25063 | n25067 ;
  assign n25069 = n10879 | n25068 ;
  assign n25070 = ( n11219 & n25068 ) | ( n11219 & n25069 ) | ( n25068 & n25069 ) ;
  assign n25071 = x59 & n25070 ;
  assign n25072 = x59 & ~n25071 ;
  assign n25073 = ( n25070 & ~n25071 ) | ( n25070 & n25072 ) | ( ~n25071 & n25072 ) ;
  assign n25074 = x120 & n11984 ;
  assign n25075 = x119 & n11979 ;
  assign n25076 = x118 & ~n11978 ;
  assign n25077 = n12430 & n25076 ;
  assign n25078 = n25075 | n25077 ;
  assign n25079 = n25074 | n25078 ;
  assign n25080 = n11987 | n25079 ;
  assign n25081 = ( n10460 & n25079 ) | ( n10460 & n25080 ) | ( n25079 & n25080 ) ;
  assign n25082 = x62 & n25081 ;
  assign n25083 = x62 & ~n25082 ;
  assign n25084 = ( n25081 & ~n25082 ) | ( n25081 & n25083 ) | ( ~n25082 & n25083 ) ;
  assign n25085 = x117 & n12808 ;
  assign n25086 = x63 & x116 ;
  assign n25087 = ~n12808 & n25086 ;
  assign n25088 = n25085 | n25087 ;
  assign n25089 = ~n25002 & n25088 ;
  assign n25090 = n25002 & ~n25088 ;
  assign n25091 = ( n25003 & ~n25088 ) | ( n25003 & n25090 ) | ( ~n25088 & n25090 ) ;
  assign n25092 = n25089 | n25091 ;
  assign n25093 = n25010 | n25092 ;
  assign n25094 = n25089 | n25090 ;
  assign n25095 = ( n25005 & n25010 ) | ( n25005 & n25094 ) | ( n25010 & n25094 ) ;
  assign n25096 = n25093 & ~n25095 ;
  assign n25097 = ( n25073 & ~n25084 ) | ( n25073 & n25096 ) | ( ~n25084 & n25096 ) ;
  assign n25098 = ( n25084 & ~n25096 ) | ( n25084 & n25097 ) | ( ~n25096 & n25097 ) ;
  assign n25099 = ( ~n25073 & n25097 ) | ( ~n25073 & n25098 ) | ( n25097 & n25098 ) ;
  assign n25100 = ~n25062 & n25099 ;
  assign n25101 = n25062 & ~n25099 ;
  assign n25102 = n25100 | n25101 ;
  assign n25103 = x126 & n9853 ;
  assign n25104 = x125 & n9848 ;
  assign n25105 = x124 & ~n9847 ;
  assign n25106 = n10165 & n25105 ;
  assign n25107 = n25104 | n25106 ;
  assign n25108 = n25103 | n25107 ;
  assign n25109 = n9856 | n25108 ;
  assign n25110 = ( n12687 & n25108 ) | ( n12687 & n25109 ) | ( n25108 & n25109 ) ;
  assign n25111 = x56 & n25110 ;
  assign n25112 = x56 & ~n25111 ;
  assign n25113 = ( n25110 & ~n25111 ) | ( n25110 & n25112 ) | ( ~n25111 & n25112 ) ;
  assign n25114 = n25102 & n25113 ;
  assign n25115 = ( n25062 & ~n25099 ) | ( n25062 & n25113 ) | ( ~n25099 & n25113 ) ;
  assign n25116 = n25100 | n25115 ;
  assign n25117 = ~n25114 & n25116 ;
  assign n25118 = n25061 & ~n25117 ;
  assign n25119 = n25117 | n25118 ;
  assign n25120 = ( ~n25061 & n25118 ) | ( ~n25061 & n25119 ) | ( n25118 & n25119 ) ;
  assign n25121 = ~n25034 & n25120 ;
  assign n25122 = n25034 & ~n25120 ;
  assign n25123 = n25121 | n25122 ;
  assign n25124 = n25038 | n25044 ;
  assign n25125 = ~n25038 & n25045 ;
  assign n25126 = ( n24328 & ~n25124 ) | ( n24328 & n25125 ) | ( ~n25124 & n25125 ) ;
  assign n25127 = n25123 & n25126 ;
  assign n25128 = ~n25123 & n25124 ;
  assign n25129 = n25123 | n25125 ;
  assign n25130 = ( n24328 & ~n25128 ) | ( n24328 & n25129 ) | ( ~n25128 & n25129 ) ;
  assign n25131 = ~n25127 & n25130 ;
  assign n25132 = x124 & n10876 ;
  assign n25133 = x123 & n10871 ;
  assign n25134 = x122 & ~n10870 ;
  assign n25135 = n11305 & n25134 ;
  assign n25136 = n25133 | n25135 ;
  assign n25137 = n25132 | n25136 ;
  assign n25138 = n10879 | n25137 ;
  assign n25139 = ( n11916 & n25137 ) | ( n11916 & n25138 ) | ( n25137 & n25138 ) ;
  assign n25140 = x59 & n25139 ;
  assign n25141 = x59 & ~n25140 ;
  assign n25142 = ( n25139 & ~n25140 ) | ( n25139 & n25141 ) | ( ~n25140 & n25141 ) ;
  assign n25143 = ( n25010 & ~n25089 ) | ( n25010 & n25091 ) | ( ~n25089 & n25091 ) ;
  assign n25144 = x121 & n11984 ;
  assign n25145 = x120 & n11979 ;
  assign n25146 = x119 & ~n11978 ;
  assign n25147 = n12430 & n25146 ;
  assign n25148 = n25145 | n25147 ;
  assign n25149 = n25144 | n25148 ;
  assign n25150 = n11987 | n25149 ;
  assign n25151 = ( n10811 & n25149 ) | ( n10811 & n25150 ) | ( n25149 & n25150 ) ;
  assign n25152 = ~x62 & n25151 ;
  assign n25153 = x62 & ~n25151 ;
  assign n25154 = n25152 | n25153 ;
  assign n25155 = x118 & n12808 ;
  assign n25156 = x63 & x117 ;
  assign n25157 = ~n12808 & n25156 ;
  assign n25158 = n25155 | n25157 ;
  assign n25159 = ( x53 & ~n25088 ) | ( x53 & n25158 ) | ( ~n25088 & n25158 ) ;
  assign n25160 = ( ~x53 & n25088 ) | ( ~x53 & n25158 ) | ( n25088 & n25158 ) ;
  assign n25161 = ( ~n25158 & n25159 ) | ( ~n25158 & n25160 ) | ( n25159 & n25160 ) ;
  assign n25162 = n25154 & ~n25161 ;
  assign n25163 = ~n25154 & n25161 ;
  assign n25164 = n25162 | n25163 ;
  assign n25165 = n25143 & ~n25164 ;
  assign n25166 = ~n25143 & n25164 ;
  assign n25167 = n25165 | n25166 ;
  assign n25168 = n25142 & ~n25167 ;
  assign n25169 = n25167 | n25168 ;
  assign n25170 = ( ~n25142 & n25168 ) | ( ~n25142 & n25169 ) | ( n25168 & n25169 ) ;
  assign n25171 = n25098 & ~n25170 ;
  assign n25172 = ~n25098 & n25170 ;
  assign n25173 = n25171 | n25172 ;
  assign n25174 = x127 & n9853 ;
  assign n25175 = x126 & n9848 ;
  assign n25176 = x125 & ~n9847 ;
  assign n25177 = n10165 & n25176 ;
  assign n25178 = n25175 | n25177 ;
  assign n25179 = n25174 | n25178 ;
  assign n25180 = n9856 | n25179 ;
  assign n25181 = ( n12720 & n25179 ) | ( n12720 & n25180 ) | ( n25179 & n25180 ) ;
  assign n25182 = x56 & n25181 ;
  assign n25183 = x56 & ~n25182 ;
  assign n25184 = ( n25181 & ~n25182 ) | ( n25181 & n25183 ) | ( ~n25182 & n25183 ) ;
  assign n25185 = ( ~n25115 & n25173 ) | ( ~n25115 & n25184 ) | ( n25173 & n25184 ) ;
  assign n25186 = ( n25115 & ~n25184 ) | ( n25115 & n25185 ) | ( ~n25184 & n25185 ) ;
  assign n25187 = ( ~n25173 & n25185 ) | ( ~n25173 & n25186 ) | ( n25185 & n25186 ) ;
  assign n25188 = n25060 | n25118 ;
  assign n25189 = ~n25187 & n25188 ;
  assign n25190 = n25187 & ~n25188 ;
  assign n25191 = n25189 | n25190 ;
  assign n25192 = n25122 | n25128 ;
  assign n25193 = ~n25122 & n25129 ;
  assign n25194 = ( n24328 & ~n25192 ) | ( n24328 & n25193 ) | ( ~n25192 & n25193 ) ;
  assign n25195 = n25191 & n25194 ;
  assign n25196 = ~n25191 & n25192 ;
  assign n25197 = n25191 | n25193 ;
  assign n25198 = ( n24328 & ~n25196 ) | ( n24328 & n25197 ) | ( ~n25196 & n25197 ) ;
  assign n25199 = ~n25195 & n25198 ;
  assign n25200 = x127 & n9848 ;
  assign n25201 = x126 & ~n9847 ;
  assign n25202 = n10165 & n25201 ;
  assign n25203 = n25200 | n25202 ;
  assign n25204 = n9856 | n25203 ;
  assign n25205 = ( n13461 & n25203 ) | ( n13461 & n25204 ) | ( n25203 & n25204 ) ;
  assign n25206 = x56 & n25205 ;
  assign n25207 = x56 & ~n25206 ;
  assign n25208 = ( n25205 & ~n25206 ) | ( n25205 & n25207 ) | ( ~n25206 & n25207 ) ;
  assign n25209 = n25168 | n25171 ;
  assign n25210 = n25162 | n25165 ;
  assign n25211 = x119 & n12808 ;
  assign n25212 = x63 & x118 ;
  assign n25213 = ~n12808 & n25212 ;
  assign n25214 = n25211 | n25213 ;
  assign n25215 = n25160 & ~n25214 ;
  assign n25216 = ~n25160 & n25214 ;
  assign n25217 = n25215 | n25216 ;
  assign n25218 = x122 & n11984 ;
  assign n25219 = x121 & n11979 ;
  assign n25220 = x120 & ~n11978 ;
  assign n25221 = n12430 & n25220 ;
  assign n25222 = n25219 | n25221 ;
  assign n25223 = n25218 | n25222 ;
  assign n25224 = n11987 | n25223 ;
  assign n25225 = ( n11188 & n25223 ) | ( n11188 & n25224 ) | ( n25223 & n25224 ) ;
  assign n25226 = x62 & n25225 ;
  assign n25227 = x62 & ~n25226 ;
  assign n25228 = ( n25225 & ~n25226 ) | ( n25225 & n25227 ) | ( ~n25226 & n25227 ) ;
  assign n25229 = ~n25217 & n25228 ;
  assign n25230 = n25217 & ~n25228 ;
  assign n25231 = n25229 | n25230 ;
  assign n25232 = n25210 & ~n25231 ;
  assign n25233 = n25210 & ~n25232 ;
  assign n25234 = n25210 | n25231 ;
  assign n25235 = x125 & n10876 ;
  assign n25236 = x124 & n10871 ;
  assign n25237 = x123 & ~n10870 ;
  assign n25238 = n11305 & n25237 ;
  assign n25239 = n25236 | n25238 ;
  assign n25240 = n25235 | n25239 ;
  assign n25241 = n10879 | n25240 ;
  assign n25242 = ( n12310 & n25240 ) | ( n12310 & n25241 ) | ( n25240 & n25241 ) ;
  assign n25243 = x59 & n25242 ;
  assign n25244 = x59 & ~n25243 ;
  assign n25245 = ( n25242 & ~n25243 ) | ( n25242 & n25244 ) | ( ~n25243 & n25244 ) ;
  assign n25246 = n25234 & ~n25245 ;
  assign n25247 = ~n25233 & n25246 ;
  assign n25248 = ( n25233 & ~n25234 ) | ( n25233 & n25245 ) | ( ~n25234 & n25245 ) ;
  assign n25249 = n25247 | n25248 ;
  assign n25250 = ( n25208 & n25209 ) | ( n25208 & ~n25249 ) | ( n25209 & ~n25249 ) ;
  assign n25251 = ( ~n25209 & n25249 ) | ( ~n25209 & n25250 ) | ( n25249 & n25250 ) ;
  assign n25252 = ( ~n25208 & n25250 ) | ( ~n25208 & n25251 ) | ( n25250 & n25251 ) ;
  assign n25253 = ( n25115 & ~n25173 ) | ( n25115 & n25184 ) | ( ~n25173 & n25184 ) ;
  assign n25254 = ~n25252 & n25253 ;
  assign n25255 = n25252 | n25254 ;
  assign n25256 = n25253 & ~n25254 ;
  assign n25257 = n25255 & ~n25256 ;
  assign n25258 = n25189 | n25196 ;
  assign n25259 = ~n25189 & n25197 ;
  assign n25260 = ( n24328 & ~n25258 ) | ( n24328 & n25259 ) | ( ~n25258 & n25259 ) ;
  assign n25261 = n25257 & n25260 ;
  assign n25262 = ~n25257 & n25258 ;
  assign n25263 = n25257 | n25259 ;
  assign n25264 = ( n24328 & ~n25262 ) | ( n24328 & n25263 ) | ( ~n25262 & n25263 ) ;
  assign n25265 = ~n25261 & n25264 ;
  assign n25266 = x127 & ~n9847 ;
  assign n25267 = n10165 & n25266 ;
  assign n25268 = ( x127 & n9856 ) | ( x127 & n25267 ) | ( n9856 & n25267 ) ;
  assign n25269 = ( x126 & n25267 ) | ( x126 & n25268 ) | ( n25267 & n25268 ) ;
  assign n25270 = ( n12685 & n25268 ) | ( n12685 & n25269 ) | ( n25268 & n25269 ) ;
  assign n25271 = x56 & n25270 ;
  assign n25272 = x56 & ~n25271 ;
  assign n25273 = ( n25270 & ~n25271 ) | ( n25270 & n25272 ) | ( ~n25271 & n25272 ) ;
  assign n25274 = n25232 | n25273 ;
  assign n25275 = n25248 | n25274 ;
  assign n25276 = ( n25232 & n25248 ) | ( n25232 & n25273 ) | ( n25248 & n25273 ) ;
  assign n25277 = n25275 & ~n25276 ;
  assign n25278 = n25215 | n25229 ;
  assign n25279 = x123 & n11984 ;
  assign n25280 = x122 & n11979 ;
  assign n25281 = x121 & ~n11978 ;
  assign n25282 = n12430 & n25281 ;
  assign n25283 = n25280 | n25282 ;
  assign n25284 = n25279 | n25283 ;
  assign n25285 = n11987 | n25284 ;
  assign n25286 = ( n11219 & n25284 ) | ( n11219 & n25285 ) | ( n25284 & n25285 ) ;
  assign n25287 = ~x62 & n25286 ;
  assign n25288 = x62 & ~n25286 ;
  assign n25289 = n25287 | n25288 ;
  assign n25290 = x120 & n12808 ;
  assign n25291 = x63 & x119 ;
  assign n25292 = ~n12808 & n25291 ;
  assign n25293 = n25290 | n25292 ;
  assign n25294 = ~n25214 & n25293 ;
  assign n25295 = n25214 | n25294 ;
  assign n25296 = n25293 & ~n25294 ;
  assign n25297 = n25295 & ~n25296 ;
  assign n25298 = n25289 & ~n25297 ;
  assign n25299 = ~n25289 & n25297 ;
  assign n25300 = n25298 | n25299 ;
  assign n25301 = x126 & n10876 ;
  assign n25302 = x125 & n10871 ;
  assign n25303 = x124 & ~n10870 ;
  assign n25304 = n11305 & n25303 ;
  assign n25305 = n25302 | n25304 ;
  assign n25306 = n25301 | n25305 ;
  assign n25307 = n10879 | n25306 ;
  assign n25308 = ( n12687 & n25306 ) | ( n12687 & n25307 ) | ( n25306 & n25307 ) ;
  assign n25309 = x59 & n25308 ;
  assign n25310 = x59 & ~n25309 ;
  assign n25311 = ( n25308 & ~n25309 ) | ( n25308 & n25310 ) | ( ~n25309 & n25310 ) ;
  assign n25312 = ( n25278 & ~n25300 ) | ( n25278 & n25311 ) | ( ~n25300 & n25311 ) ;
  assign n25313 = ( n25300 & ~n25311 ) | ( n25300 & n25312 ) | ( ~n25311 & n25312 ) ;
  assign n25314 = ( ~n25278 & n25312 ) | ( ~n25278 & n25313 ) | ( n25312 & n25313 ) ;
  assign n25315 = n25277 & ~n25314 ;
  assign n25316 = n25314 | n25315 ;
  assign n25317 = ( ~n25277 & n25315 ) | ( ~n25277 & n25316 ) | ( n25315 & n25316 ) ;
  assign n25318 = ~n25250 & n25317 ;
  assign n25319 = n25250 & ~n25317 ;
  assign n25320 = n25318 | n25319 ;
  assign n25321 = n25254 | n25262 ;
  assign n25322 = ~n25254 & n25263 ;
  assign n25323 = ( n24328 & ~n25321 ) | ( n24328 & n25322 ) | ( ~n25321 & n25322 ) ;
  assign n25324 = n25320 & n25323 ;
  assign n25325 = ~n25320 & n25321 ;
  assign n25326 = n25320 | n25322 ;
  assign n25327 = ( n24328 & ~n25325 ) | ( n24328 & n25326 ) | ( ~n25325 & n25326 ) ;
  assign n25328 = ~n25324 & n25327 ;
  assign n25329 = x127 & n10876 ;
  assign n25330 = x126 & n10871 ;
  assign n25331 = x125 & ~n10870 ;
  assign n25332 = n11305 & n25331 ;
  assign n25333 = n25330 | n25332 ;
  assign n25334 = n25329 | n25333 ;
  assign n25335 = n10879 | n25334 ;
  assign n25336 = ( n12720 & n25334 ) | ( n12720 & n25335 ) | ( n25334 & n25335 ) ;
  assign n25337 = x59 & n25336 ;
  assign n25338 = x59 & ~n25337 ;
  assign n25339 = ( n25336 & ~n25337 ) | ( n25336 & n25338 ) | ( ~n25337 & n25338 ) ;
  assign n25340 = n25312 & n25339 ;
  assign n25341 = n25312 & ~n25340 ;
  assign n25342 = ~n25312 & n25339 ;
  assign n25343 = n25341 | n25342 ;
  assign n25344 = x121 & n12808 ;
  assign n25345 = x63 & x120 ;
  assign n25346 = ~n12808 & n25345 ;
  assign n25347 = n25344 | n25346 ;
  assign n25348 = ~x56 & n25347 ;
  assign n25349 = n25347 & ~n25348 ;
  assign n25350 = x56 | n25347 ;
  assign n25351 = ~n25349 & n25350 ;
  assign n25352 = n25214 & ~n25351 ;
  assign n25353 = ~n25214 & n25351 ;
  assign n25354 = n25352 | n25353 ;
  assign n25355 = n25294 & ~n25354 ;
  assign n25356 = ( n25298 & ~n25354 ) | ( n25298 & n25355 ) | ( ~n25354 & n25355 ) ;
  assign n25357 = ~n25294 & n25354 ;
  assign n25358 = ~n25298 & n25357 ;
  assign n25359 = n25356 | n25358 ;
  assign n25360 = x124 & n11984 ;
  assign n25361 = x123 & n11979 ;
  assign n25362 = x122 & ~n11978 ;
  assign n25363 = n12430 & n25362 ;
  assign n25364 = n25361 | n25363 ;
  assign n25365 = n25360 | n25364 ;
  assign n25366 = n11987 | n25365 ;
  assign n25367 = ( n11916 & n25365 ) | ( n11916 & n25366 ) | ( n25365 & n25366 ) ;
  assign n25368 = x62 & n25367 ;
  assign n25369 = x62 & ~n25368 ;
  assign n25370 = ( n25367 & ~n25368 ) | ( n25367 & n25369 ) | ( ~n25368 & n25369 ) ;
  assign n25371 = ~n25359 & n25370 ;
  assign n25372 = n25359 & ~n25370 ;
  assign n25373 = n25343 & ~n25372 ;
  assign n25374 = ~n25371 & n25373 ;
  assign n25375 = n25343 & ~n25374 ;
  assign n25376 = n25276 | n25315 ;
  assign n25377 = n25372 | n25373 ;
  assign n25378 = n25371 | n25377 ;
  assign n25379 = ~n25376 & n25378 ;
  assign n25380 = ~n25375 & n25379 ;
  assign n25381 = ( n25375 & n25376 ) | ( n25375 & ~n25378 ) | ( n25376 & ~n25378 ) ;
  assign n25382 = n25380 | n25381 ;
  assign n25383 = n25319 | n25325 ;
  assign n25384 = ~n25319 & n25326 ;
  assign n25385 = ( n24328 & ~n25383 ) | ( n24328 & n25384 ) | ( ~n25383 & n25384 ) ;
  assign n25386 = n25382 & n25385 ;
  assign n25387 = ~n25382 & n25383 ;
  assign n25388 = n25382 | n25384 ;
  assign n25389 = ( n24328 & ~n25387 ) | ( n24328 & n25388 ) | ( ~n25387 & n25388 ) ;
  assign n25390 = ~n25386 & n25389 ;
  assign n25391 = n25340 | n25374 ;
  assign n25392 = x127 & n10871 ;
  assign n25393 = x126 & ~n10870 ;
  assign n25394 = n11305 & n25393 ;
  assign n25395 = n25392 | n25394 ;
  assign n25396 = n10879 | n25395 ;
  assign n25397 = ( n13461 & n25395 ) | ( n13461 & n25396 ) | ( n25395 & n25396 ) ;
  assign n25398 = x59 & n25397 ;
  assign n25399 = x59 & ~n25398 ;
  assign n25400 = ( n25397 & ~n25398 ) | ( n25397 & n25399 ) | ( ~n25398 & n25399 ) ;
  assign n25401 = x122 & n12808 ;
  assign n25402 = x63 & x121 ;
  assign n25403 = ~n12808 & n25402 ;
  assign n25404 = n25401 | n25403 ;
  assign n25405 = ~n25348 & n25404 ;
  assign n25406 = ~n25352 & n25405 ;
  assign n25407 = ( n25348 & n25352 ) | ( n25348 & ~n25404 ) | ( n25352 & ~n25404 ) ;
  assign n25408 = n25406 | n25407 ;
  assign n25409 = x125 & n11984 ;
  assign n25410 = x124 & n11979 ;
  assign n25411 = x123 & ~n11978 ;
  assign n25412 = n12430 & n25411 ;
  assign n25413 = n25410 | n25412 ;
  assign n25414 = n25409 | n25413 ;
  assign n25415 = n11987 | n25414 ;
  assign n25416 = ( n12310 & n25414 ) | ( n12310 & n25415 ) | ( n25414 & n25415 ) ;
  assign n25417 = x62 & n25416 ;
  assign n25418 = x62 & ~n25417 ;
  assign n25419 = ( n25416 & ~n25417 ) | ( n25416 & n25418 ) | ( ~n25417 & n25418 ) ;
  assign n25420 = ~n25408 & n25419 ;
  assign n25421 = n25408 & ~n25419 ;
  assign n25422 = n25420 | n25421 ;
  assign n25423 = n25356 | n25371 ;
  assign n25424 = ( n25400 & n25422 ) | ( n25400 & ~n25423 ) | ( n25422 & ~n25423 ) ;
  assign n25425 = ( ~n25422 & n25423 ) | ( ~n25422 & n25424 ) | ( n25423 & n25424 ) ;
  assign n25426 = ( ~n25400 & n25424 ) | ( ~n25400 & n25425 ) | ( n25424 & n25425 ) ;
  assign n25427 = ~n25391 & n25426 ;
  assign n25428 = n25391 & ~n25426 ;
  assign n25429 = n25427 | n25428 ;
  assign n25430 = n25381 | n25387 ;
  assign n25431 = ~n25381 & n25388 ;
  assign n25432 = ( n24328 & ~n25430 ) | ( n24328 & n25431 ) | ( ~n25430 & n25431 ) ;
  assign n25433 = n25429 & n25432 ;
  assign n25434 = ~n25429 & n25430 ;
  assign n25435 = n25429 | n25431 ;
  assign n25436 = ( n24328 & ~n25434 ) | ( n24328 & n25435 ) | ( ~n25434 & n25435 ) ;
  assign n25437 = ~n25433 & n25436 ;
  assign n25438 = x127 & ~n10870 ;
  assign n25439 = n11305 & n25438 ;
  assign n25440 = ( x127 & n10879 ) | ( x127 & n25439 ) | ( n10879 & n25439 ) ;
  assign n25441 = ( x126 & n25439 ) | ( x126 & n25440 ) | ( n25439 & n25440 ) ;
  assign n25442 = ( n12685 & n25440 ) | ( n12685 & n25441 ) | ( n25440 & n25441 ) ;
  assign n25443 = x59 & n25442 ;
  assign n25444 = x59 & ~n25443 ;
  assign n25445 = ( n25442 & ~n25443 ) | ( n25442 & n25444 ) | ( ~n25443 & n25444 ) ;
  assign n25446 = x123 & n12808 ;
  assign n25447 = x63 & x122 ;
  assign n25448 = ~n12808 & n25447 ;
  assign n25449 = n25446 | n25448 ;
  assign n25450 = ~n25404 & n25449 ;
  assign n25451 = n25404 & ~n25449 ;
  assign n25452 = n25406 | n25451 ;
  assign n25453 = n25450 | n25452 ;
  assign n25454 = n25407 & ~n25450 ;
  assign n25455 = ( n25419 & ~n25453 ) | ( n25419 & n25454 ) | ( ~n25453 & n25454 ) ;
  assign n25456 = ( n25407 & n25420 ) | ( n25407 & ~n25455 ) | ( n25420 & ~n25455 ) ;
  assign n25457 = n25451 | n25455 ;
  assign n25458 = n25450 | n25457 ;
  assign n25459 = ~n25456 & n25458 ;
  assign n25460 = x126 & n11984 ;
  assign n25461 = x125 & n11979 ;
  assign n25462 = x124 & ~n11978 ;
  assign n25463 = n12430 & n25462 ;
  assign n25464 = n25461 | n25463 ;
  assign n25465 = n25460 | n25464 ;
  assign n25466 = n11987 | n25465 ;
  assign n25467 = ( n12687 & n25465 ) | ( n12687 & n25466 ) | ( n25465 & n25466 ) ;
  assign n25468 = x62 & n25467 ;
  assign n25469 = x62 & ~n25468 ;
  assign n25470 = ( n25467 & ~n25468 ) | ( n25467 & n25469 ) | ( ~n25468 & n25469 ) ;
  assign n25471 = ( n25445 & n25459 ) | ( n25445 & ~n25470 ) | ( n25459 & ~n25470 ) ;
  assign n25472 = ( n25445 & ~n25459 ) | ( n25445 & n25470 ) | ( ~n25459 & n25470 ) ;
  assign n25473 = ( ~n25445 & n25471 ) | ( ~n25445 & n25472 ) | ( n25471 & n25472 ) ;
  assign n25474 = n25425 & ~n25473 ;
  assign n25475 = n25425 & ~n25474 ;
  assign n25476 = n25428 | n25434 ;
  assign n25477 = ~n25428 & n25435 ;
  assign n25478 = ( n24328 & ~n25476 ) | ( n24328 & n25477 ) | ( ~n25476 & n25477 ) ;
  assign n25479 = n25425 | n25473 ;
  assign n25480 = n25478 & n25479 ;
  assign n25481 = ~n25475 & n25480 ;
  assign n25482 = ~n25475 & n25479 ;
  assign n25483 = n25476 & ~n25482 ;
  assign n25484 = n25477 | n25482 ;
  assign n25485 = ( n24328 & ~n25483 ) | ( n24328 & n25484 ) | ( ~n25483 & n25484 ) ;
  assign n25486 = ~n25481 & n25485 ;
  assign n25487 = x127 & n11984 ;
  assign n25488 = x126 & n11979 ;
  assign n25489 = x125 & ~n11978 ;
  assign n25490 = n12430 & n25489 ;
  assign n25491 = n25488 | n25490 ;
  assign n25492 = n25487 | n25491 ;
  assign n25493 = n11987 | n25492 ;
  assign n25494 = ( n12720 & n25492 ) | ( n12720 & n25493 ) | ( n25492 & n25493 ) ;
  assign n25495 = ~x62 & n25494 ;
  assign n25496 = x62 & ~n25494 ;
  assign n25497 = n25495 | n25496 ;
  assign n25498 = x124 & n12808 ;
  assign n25499 = x63 & x123 ;
  assign n25500 = ~n12808 & n25499 ;
  assign n25501 = n25498 | n25500 ;
  assign n25502 = ( x59 & ~n25449 ) | ( x59 & n25501 ) | ( ~n25449 & n25501 ) ;
  assign n25503 = ( ~x59 & n25449 ) | ( ~x59 & n25501 ) | ( n25449 & n25501 ) ;
  assign n25504 = ( ~n25501 & n25502 ) | ( ~n25501 & n25503 ) | ( n25502 & n25503 ) ;
  assign n25505 = ( n25457 & n25497 ) | ( n25457 & ~n25504 ) | ( n25497 & ~n25504 ) ;
  assign n25506 = ( ~n25457 & n25504 ) | ( ~n25457 & n25505 ) | ( n25504 & n25505 ) ;
  assign n25507 = ( ~n25497 & n25505 ) | ( ~n25497 & n25506 ) | ( n25505 & n25506 ) ;
  assign n25508 = n25472 & n25507 ;
  assign n25509 = n25474 | n25483 ;
  assign n25510 = n25472 & ~n25507 ;
  assign n25511 = n25507 | n25510 ;
  assign n25512 = ~n25508 & n25511 ;
  assign n25513 = n25509 & ~n25512 ;
  assign n25514 = ~n25474 & n25484 ;
  assign n25515 = n25512 | n25514 ;
  assign n25516 = ( n24328 & ~n25513 ) | ( n24328 & n25515 ) | ( ~n25513 & n25515 ) ;
  assign n25517 = ( n24328 & ~n25509 ) | ( n24328 & n25514 ) | ( ~n25509 & n25514 ) ;
  assign n25518 = ( n25472 & n25507 ) | ( n25472 & n25517 ) | ( n25507 & n25517 ) ;
  assign n25519 = ( n25508 & n25516 ) | ( n25508 & ~n25518 ) | ( n25516 & ~n25518 ) ;
  assign n25520 = x125 & n12808 ;
  assign n25521 = x63 & x124 ;
  assign n25522 = ~n12808 & n25521 ;
  assign n25523 = n25520 | n25522 ;
  assign n25524 = n25503 & ~n25523 ;
  assign n25525 = ~n25503 & n25523 ;
  assign n25526 = n25524 | n25525 ;
  assign n25527 = x127 & n11979 ;
  assign n25528 = x126 & ~n11978 ;
  assign n25529 = n12430 & n25528 ;
  assign n25530 = n25527 | n25529 ;
  assign n25531 = n11987 | n25530 ;
  assign n25532 = ( n13461 & n25530 ) | ( n13461 & n25531 ) | ( n25530 & n25531 ) ;
  assign n25533 = x62 & n25532 ;
  assign n25534 = x62 & ~n25533 ;
  assign n25535 = ( n25532 & ~n25533 ) | ( n25532 & n25534 ) | ( ~n25533 & n25534 ) ;
  assign n25536 = ~n25526 & n25535 ;
  assign n25537 = n25526 & ~n25535 ;
  assign n25538 = n25536 | n25537 ;
  assign n25539 = n25505 & ~n25538 ;
  assign n25540 = n25505 & ~n25539 ;
  assign n25541 = n25538 | n25539 ;
  assign n25542 = ~n25540 & n25541 ;
  assign n25543 = n25510 | n25513 ;
  assign n25544 = ~n25542 & n25543 ;
  assign n25545 = ~n25510 & n25515 ;
  assign n25546 = n25542 | n25545 ;
  assign n25547 = ( n24328 & ~n25544 ) | ( n24328 & n25546 ) | ( ~n25544 & n25546 ) ;
  assign n25548 = ( n24328 & ~n25543 ) | ( n24328 & n25545 ) | ( ~n25543 & n25545 ) ;
  assign n25549 = n25547 & ~n25548 ;
  assign n25550 = ( ~n25542 & n25547 ) | ( ~n25542 & n25549 ) | ( n25547 & n25549 ) ;
  assign n25551 = n25524 | n25536 ;
  assign n25552 = x126 & n12808 ;
  assign n25553 = x63 & x125 ;
  assign n25554 = ~n12808 & n25553 ;
  assign n25555 = n25552 | n25554 ;
  assign n25556 = ~n25523 & n25555 ;
  assign n25557 = n25523 & ~n25555 ;
  assign n25558 = n25556 | n25557 ;
  assign n25559 = x127 & ~n11978 ;
  assign n25560 = n12430 & n25559 ;
  assign n25561 = ( x127 & n11987 ) | ( x127 & n25560 ) | ( n11987 & n25560 ) ;
  assign n25562 = ( x126 & n25560 ) | ( x126 & n25561 ) | ( n25560 & n25561 ) ;
  assign n25563 = ( n12685 & n25561 ) | ( n12685 & n25562 ) | ( n25561 & n25562 ) ;
  assign n25564 = x62 & n25563 ;
  assign n25565 = x62 & ~n25564 ;
  assign n25566 = ( n25563 & ~n25564 ) | ( n25563 & n25565 ) | ( ~n25564 & n25565 ) ;
  assign n25567 = ~n25558 & n25566 ;
  assign n25568 = n25558 & ~n25566 ;
  assign n25569 = n25567 | n25568 ;
  assign n25570 = n25551 & ~n25569 ;
  assign n25571 = n25551 & ~n25570 ;
  assign n25572 = n25539 | n25544 ;
  assign n25573 = ~n25539 & n25546 ;
  assign n25574 = ( n24328 & ~n25572 ) | ( n24328 & n25573 ) | ( ~n25572 & n25573 ) ;
  assign n25575 = n25551 | n25569 ;
  assign n25576 = n25574 & n25575 ;
  assign n25577 = ~n25571 & n25576 ;
  assign n25578 = ~n25571 & n25575 ;
  assign n25579 = n25572 & ~n25578 ;
  assign n25580 = n25573 | n25578 ;
  assign n25581 = ( n24328 & ~n25579 ) | ( n24328 & n25580 ) | ( ~n25579 & n25580 ) ;
  assign n25582 = ~n25577 & n25581 ;
  assign n25583 = x127 & n12808 ;
  assign n25584 = x63 & x126 ;
  assign n25585 = ~n12808 & n25584 ;
  assign n25586 = n25583 | n25585 ;
  assign n25587 = ~x62 & n25586 ;
  assign n25588 = x62 & ~n25586 ;
  assign n25589 = n25587 | n25588 ;
  assign n25590 = n25523 & ~n25589 ;
  assign n25591 = ~n25523 & n25589 ;
  assign n25592 = n25590 | n25591 ;
  assign n25593 = ( n25556 & n25567 ) | ( n25556 & ~n25592 ) | ( n25567 & ~n25592 ) ;
  assign n25594 = ( n25556 & ~n25557 ) | ( n25556 & n25566 ) | ( ~n25557 & n25566 ) ;
  assign n25595 = n25592 & ~n25594 ;
  assign n25596 = n25593 | n25595 ;
  assign n25597 = n25570 | n25579 ;
  assign n25598 = ~n25570 & n25580 ;
  assign n25599 = ( n24328 & ~n25597 ) | ( n24328 & n25598 ) | ( ~n25597 & n25598 ) ;
  assign n25600 = n25596 & n25599 ;
  assign n25601 = ~n25596 & n25597 ;
  assign n25602 = n25596 | n25598 ;
  assign n25603 = ( n24328 & ~n25601 ) | ( n24328 & n25602 ) | ( ~n25601 & n25602 ) ;
  assign n25604 = ~n25600 & n25603 ;
  assign n25605 = n25587 | n25590 ;
  assign n25606 = x63 & x127 ;
  assign n25607 = ~n12808 & n25606 ;
  assign n25608 = ~n25593 & n25603 ;
  assign n25609 = ( n25605 & ~n25607 ) | ( n25605 & n25608 ) | ( ~n25607 & n25608 ) ;
  assign n25610 = ( n25607 & ~n25608 ) | ( n25607 & n25609 ) | ( ~n25608 & n25609 ) ;
  assign n25611 = ( ~n25605 & n25609 ) | ( ~n25605 & n25610 ) | ( n25609 & n25610 ) ;
  assign y0 = n129 ;
  assign y1 = n150 ;
  assign y2 = n168 ;
  assign y3 = n197 ;
  assign y4 = n241 ;
  assign y5 = n283 ;
  assign y6 = n327 ;
  assign y7 = n393 ;
  assign y8 = n454 ;
  assign y9 = n518 ;
  assign y10 = n597 ;
  assign y11 = n675 ;
  assign y12 = n760 ;
  assign y13 = n857 ;
  assign y14 = n950 ;
  assign y15 = n1048 ;
  assign y16 = n1164 ;
  assign y17 = n1275 ;
  assign y18 = n1390 ;
  assign y19 = n1529 ;
  assign y20 = n1653 ;
  assign y21 = n1784 ;
  assign y22 = n1939 ;
  assign y23 = n2086 ;
  assign y24 = n2233 ;
  assign y25 = n2399 ;
  assign y26 = n2560 ;
  assign y27 = n2731 ;
  assign y28 = n2921 ;
  assign y29 = n3104 ;
  assign y30 = n3283 ;
  assign y31 = n3498 ;
  assign y32 = n3696 ;
  assign y33 = n3892 ;
  assign y34 = n4123 ;
  assign y35 = n4339 ;
  assign y36 = n4551 ;
  assign y37 = n4800 ;
  assign y38 = n5044 ;
  assign y39 = n5283 ;
  assign y40 = n5551 ;
  assign y41 = n5806 ;
  assign y42 = n6057 ;
  assign y43 = n6347 ;
  assign y44 = n6625 ;
  assign y45 = n6902 ;
  assign y46 = n7208 ;
  assign y47 = n7511 ;
  assign y48 = n7799 ;
  assign y49 = n8130 ;
  assign y50 = n8456 ;
  assign y51 = n8767 ;
  assign y52 = n9107 ;
  assign y53 = n9442 ;
  assign y54 = n9778 ;
  assign y55 = n10127 ;
  assign y56 = n10479 ;
  assign y57 = n10830 ;
  assign y58 = n11207 ;
  assign y59 = n11571 ;
  assign y60 = n11938 ;
  assign y61 = n12333 ;
  assign y62 = n12708 ;
  assign y63 = n13085 ;
  assign y64 = n13474 ;
  assign y65 = n13861 ;
  assign y66 = n14205 ;
  assign y67 = n14546 ;
  assign y68 = n14889 ;
  assign y69 = n15243 ;
  assign y70 = n15563 ;
  assign y71 = n15897 ;
  assign y72 = n16224 ;
  assign y73 = n16557 ;
  assign y74 = n16883 ;
  assign y75 = n17198 ;
  assign y76 = n17509 ;
  assign y77 = n17809 ;
  assign y78 = n18112 ;
  assign y79 = n18391 ;
  assign y80 = n18685 ;
  assign y81 = n18977 ;
  assign y82 = n19246 ;
  assign y83 = n19515 ;
  assign y84 = n19785 ;
  assign y85 = n20040 ;
  assign y86 = n20276 ;
  assign y87 = n20516 ;
  assign y88 = n20749 ;
  assign y89 = n20983 ;
  assign y90 = n21216 ;
  assign y91 = n21423 ;
  assign y92 = n21633 ;
  assign y93 = n21850 ;
  assign y94 = n22047 ;
  assign y95 = n22244 ;
  assign y96 = n22448 ;
  assign y97 = n22629 ;
  assign y98 = n22806 ;
  assign y99 = n22989 ;
  assign y100 = n23163 ;
  assign y101 = n23329 ;
  assign y102 = n23485 ;
  assign y103 = n23639 ;
  assign y104 = n23790 ;
  assign y105 = n23934 ;
  assign y106 = n24073 ;
  assign y107 = n24205 ;
  assign y108 = n24329 ;
  assign y109 = n24444 ;
  assign y110 = n24559 ;
  assign y111 = n24668 ;
  assign y112 = n24766 ;
  assign y113 = n24867 ;
  assign y114 = n24966 ;
  assign y115 = n25047 ;
  assign y116 = n25131 ;
  assign y117 = n25199 ;
  assign y118 = n25265 ;
  assign y119 = n25328 ;
  assign y120 = n25390 ;
  assign y121 = n25437 ;
  assign y122 = n25486 ;
  assign y123 = n25519 ;
  assign y124 = n25550 ;
  assign y125 = n25582 ;
  assign y126 = n25604 ;
  assign y127 = n25611 ;
endmodule
