module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 ;
  assign n11 = x3 | x5 ;
  assign n12 = ~x1 & x9 ;
  assign n13 = ~x0 & x9 ;
  assign n14 = x1 & ~n13 ;
  assign n15 = n12 | n14 ;
  assign n16 = n11 | n15 ;
  assign n17 = x0 & ~x9 ;
  assign n18 = x1 | n17 ;
  assign n19 = x1 & ~x9 ;
  assign n20 = x7 | n19 ;
  assign n21 = n18 & ~n20 ;
  assign n22 = n16 & ~n21 ;
  assign n23 = x2 | n22 ;
  assign n24 = x2 | x5 ;
  assign n25 = x1 & x2 ;
  assign n26 = ( ~x0 & n24 ) | ( ~x0 & n25 ) | ( n24 & n25 ) ;
  assign n27 = ~x9 & n26 ;
  assign n28 = x2 | x3 ;
  assign n29 = x9 & n28 ;
  assign n30 = x0 & x3 ;
  assign n31 = n29 | n30 ;
  assign n32 = ~x1 & n31 ;
  assign n33 = x1 & ~x3 ;
  assign n34 = n32 | n33 ;
  assign n35 = n27 | n34 ;
  assign n36 = ~x7 & n35 ;
  assign n37 = n23 & ~n36 ;
  assign n38 = x8 | n37 ;
  assign n39 = x7 & x8 ;
  assign n40 = ~x5 & n39 ;
  assign n41 = ~x7 & x9 ;
  assign n42 = n40 | n41 ;
  assign n43 = x1 & n42 ;
  assign n44 = x1 & ~x7 ;
  assign n45 = x5 | x9 ;
  assign n46 = n44 | n45 ;
  assign n47 = ~n43 & n46 ;
  assign n48 = x0 & ~x2 ;
  assign n49 = ~n47 & n48 ;
  assign n50 = x2 & ~x9 ;
  assign n51 = x0 | x1 ;
  assign n52 = n50 & ~n51 ;
  assign n53 = n40 & n52 ;
  assign n54 = n49 | n53 ;
  assign n55 = ~x3 & n54 ;
  assign n56 = n38 & ~n55 ;
  assign n57 = x6 | n56 ;
  assign n58 = x0 | x2 ;
  assign n59 = n12 & ~n58 ;
  assign n60 = x5 | n59 ;
  assign n61 = x0 | x9 ;
  assign n62 = x0 & x9 ;
  assign n63 = n61 & ~n62 ;
  assign n64 = x1 & ~n63 ;
  assign n65 = x2 & n64 ;
  assign n66 = x5 & n65 ;
  assign n67 = ( x6 & n60 ) | ( x6 & n66 ) | ( n60 & n66 ) ;
  assign n68 = x8 & n67 ;
  assign n69 = x1 | n13 ;
  assign n70 = ~x8 & n69 ;
  assign n71 = ~x1 & x2 ;
  assign n72 = n17 & n71 ;
  assign n73 = n70 | n72 ;
  assign n74 = ~x5 & n73 ;
  assign n75 = n68 | n74 ;
  assign n76 = x3 & n75 ;
  assign n77 = x2 | n17 ;
  assign n78 = x6 & n77 ;
  assign n79 = ~n28 & n64 ;
  assign n80 = n78 | n79 ;
  assign n81 = x5 & n80 ;
  assign n82 = x2 & x9 ;
  assign n83 = ~x2 & n19 ;
  assign n84 = n82 | n83 ;
  assign n85 = x0 | x3 ;
  assign n86 = n84 & ~n85 ;
  assign n87 = x6 & n86 ;
  assign n88 = n81 | n87 ;
  assign n89 = x8 & n88 ;
  assign n90 = x2 & ~x3 ;
  assign n91 = n12 & n90 ;
  assign n92 = x1 & ~x8 ;
  assign n93 = n91 | n92 ;
  assign n94 = ~x0 & n93 ;
  assign n95 = x1 | x9 ;
  assign n96 = ~x2 & x6 ;
  assign n97 = x3 & ~n96 ;
  assign n98 = n95 | n97 ;
  assign n99 = ~n82 & n98 ;
  assign n100 = x8 | n99 ;
  assign n101 = ~n94 & n100 ;
  assign n102 = x5 | n101 ;
  assign n103 = x0 | n28 ;
  assign n104 = x8 | n95 ;
  assign n105 = n103 | n104 ;
  assign n106 = n102 & n105 ;
  assign n107 = ~n89 & n106 ;
  assign n108 = ~n76 & n107 ;
  assign n109 = x7 | n108 ;
  assign n110 = n57 & n109 ;
  assign n111 = x4 | n110 ;
  assign n112 = x4 & x8 ;
  assign n113 = x6 & n112 ;
  assign n114 = ~x6 & x9 ;
  assign n115 = x6 | x8 ;
  assign n116 = ( ~n113 & n114 ) | ( ~n113 & n115 ) | ( n114 & n115 ) ;
  assign n117 = x5 & ~n116 ;
  assign n118 = x6 & ~x9 ;
  assign n119 = x4 & x9 ;
  assign n120 = n118 | n119 ;
  assign n121 = x5 & x6 ;
  assign n122 = n120 & ~n121 ;
  assign n123 = ~x8 & n122 ;
  assign n124 = n117 | n123 ;
  assign n125 = ~x7 & n124 ;
  assign n126 = x1 | x3 ;
  assign n127 = ( n58 & n125 ) | ( n58 & ~n126 ) | ( n125 & ~n126 ) ;
  assign n128 = ~n58 & n127 ;
  assign n129 = n111 & ~n128 ;
  assign n130 = x3 & n25 ;
  assign n131 = ( x5 & n28 ) | ( x5 & n130 ) | ( n28 & n130 ) ;
  assign n132 = x3 & ~x8 ;
  assign n133 = x1 | x2 ;
  assign n134 = n132 & ~n133 ;
  assign n135 = x1 & x5 ;
  assign n136 = x0 & n135 ;
  assign n137 = ( x0 & n134 ) | ( x0 & n136 ) | ( n134 & n136 ) ;
  assign n138 = n131 | n137 ;
  assign n139 = x5 & ~x8 ;
  assign n140 = n130 & n139 ;
  assign n141 = x6 | n140 ;
  assign n142 = ( n138 & n140 ) | ( n138 & n141 ) | ( n140 & n141 ) ;
  assign n143 = ( x4 & x9 ) | ( x4 & ~n142 ) | ( x9 & ~n142 ) ;
  assign n144 = ~x0 & x5 ;
  assign n145 = ~x2 & x8 ;
  assign n146 = x0 & ~x5 ;
  assign n147 = ( x0 & n145 ) | ( x0 & n146 ) | ( n145 & n146 ) ;
  assign n148 = ( x1 & n144 ) | ( x1 & n147 ) | ( n144 & n147 ) ;
  assign n149 = x3 & x8 ;
  assign n150 = n58 | n149 ;
  assign n151 = ( ~x0 & n148 ) | ( ~x0 & n150 ) | ( n148 & n150 ) ;
  assign n152 = ~x5 & x8 ;
  assign n153 = x3 | x8 ;
  assign n154 = ~n152 & n153 ;
  assign n155 = x0 & n154 ;
  assign n156 = x2 | x8 ;
  assign n157 = x5 & ~n156 ;
  assign n158 = ~x1 & n157 ;
  assign n159 = ( ~x1 & n155 ) | ( ~x1 & n158 ) | ( n155 & n158 ) ;
  assign n160 = n151 | n159 ;
  assign n161 = ~x6 & n160 ;
  assign n162 = x2 & x6 ;
  assign n163 = ~x1 & n162 ;
  assign n164 = ~x2 & x3 ;
  assign n165 = x1 | x8 ;
  assign n166 = x3 & n165 ;
  assign n167 = ( n163 & n164 ) | ( n163 & n166 ) | ( n164 & n166 ) ;
  assign n168 = x1 | x6 ;
  assign n169 = x0 & x1 ;
  assign n170 = n168 & ~n169 ;
  assign n171 = ~x0 & x8 ;
  assign n172 = x2 | n171 ;
  assign n173 = n170 & ~n172 ;
  assign n174 = n167 | n173 ;
  assign n175 = ~x5 & n174 ;
  assign n176 = ( ~x4 & x9 ) | ( ~x4 & n175 ) | ( x9 & n175 ) ;
  assign n177 = x4 & ~x9 ;
  assign n178 = ( n161 & n176 ) | ( n161 & ~n177 ) | ( n176 & ~n177 ) ;
  assign n179 = ~n143 & n178 ;
  assign n180 = x6 & x9 ;
  assign n181 = n152 | n180 ;
  assign n182 = ~x0 & n181 ;
  assign n183 = x8 & n180 ;
  assign n184 = x8 | n45 ;
  assign n185 = ~n183 & n184 ;
  assign n186 = ~n182 & n185 ;
  assign n187 = x2 & ~n186 ;
  assign n188 = x0 & x8 ;
  assign n189 = n82 & n188 ;
  assign n190 = n61 | n156 ;
  assign n191 = ~n189 & n190 ;
  assign n192 = x5 & ~n191 ;
  assign n193 = ~x4 & n192 ;
  assign n194 = ( ~x4 & n187 ) | ( ~x4 & n193 ) | ( n187 & n193 ) ;
  assign n195 = n112 | n139 ;
  assign n196 = x6 & ~n119 ;
  assign n197 = ( n119 & n195 ) | ( n119 & ~n196 ) | ( n195 & ~n196 ) ;
  assign n198 = n58 | n114 ;
  assign n199 = n197 & ~n198 ;
  assign n200 = ~x1 & n199 ;
  assign n201 = ( ~x1 & n194 ) | ( ~x1 & n200 ) | ( n194 & n200 ) ;
  assign n202 = ~x0 & x6 ;
  assign n203 = x2 | n202 ;
  assign n204 = n115 & ~n152 ;
  assign n205 = ( n115 & ~n203 ) | ( n115 & n204 ) | ( ~n203 & n204 ) ;
  assign n206 = x9 | n205 ;
  assign n207 = x6 & x8 ;
  assign n208 = x0 & ~n207 ;
  assign n209 = n181 & n208 ;
  assign n210 = ~x8 & x9 ;
  assign n211 = n144 & n210 ;
  assign n212 = ~x2 & n211 ;
  assign n213 = ( ~x2 & n209 ) | ( ~x2 & n212 ) | ( n209 & n212 ) ;
  assign n214 = n206 & ~n213 ;
  assign n215 = ~x6 & x8 ;
  assign n216 = n50 & n215 ;
  assign n217 = x1 | n216 ;
  assign n218 = ~x4 & n217 ;
  assign n219 = ~x4 & n216 ;
  assign n220 = ( ~n214 & n218 ) | ( ~n214 & n219 ) | ( n218 & n219 ) ;
  assign n221 = ~x3 & n220 ;
  assign n222 = ( ~x3 & n201 ) | ( ~x3 & n221 ) | ( n201 & n221 ) ;
  assign n223 = n179 | n222 ;
  assign n224 = ~x7 & n223 ;
  assign n225 = x6 | n11 ;
  assign n226 = n77 | n169 ;
  assign n227 = x2 & n51 ;
  assign n228 = x8 | n227 ;
  assign n229 = n226 & ~n228 ;
  assign n230 = n19 & n145 ;
  assign n231 = x7 & n230 ;
  assign n232 = n52 | n231 ;
  assign n233 = x7 | n52 ;
  assign n234 = ( n229 & n232 ) | ( n229 & n233 ) | ( n232 & n233 ) ;
  assign n235 = ~x4 & n234 ;
  assign n236 = x7 & ~n235 ;
  assign n237 = ( n223 & n235 ) | ( n223 & ~n236 ) | ( n235 & ~n236 ) ;
  assign n238 = ( n224 & ~n225 ) | ( n224 & n237 ) | ( ~n225 & n237 ) ;
  assign n239 = ~x1 & x3 ;
  assign n240 = x5 & ~n239 ;
  assign n241 = x8 | x9 ;
  assign n242 = x2 | n241 ;
  assign n243 = n240 | n242 ;
  assign n244 = ~x1 & x8 ;
  assign n245 = n29 & n244 ;
  assign n246 = n243 & ~n245 ;
  assign n247 = x0 & ~n246 ;
  assign n248 = x8 & n62 ;
  assign n249 = x5 & ~n241 ;
  assign n250 = ( x5 & n248 ) | ( x5 & n249 ) | ( n248 & n249 ) ;
  assign n251 = ~x5 & n82 ;
  assign n252 = x1 & n251 ;
  assign n253 = ( x1 & n250 ) | ( x1 & n252 ) | ( n250 & n252 ) ;
  assign n254 = x8 & ~x9 ;
  assign n255 = n210 | n254 ;
  assign n256 = ( n90 & ~n95 ) | ( n90 & n255 ) | ( ~n95 & n255 ) ;
  assign n257 = n90 & n256 ;
  assign n258 = ( ~x3 & n253 ) | ( ~x3 & n257 ) | ( n253 & n257 ) ;
  assign n259 = n247 | n258 ;
  assign n260 = ~x6 & n259 ;
  assign n261 = x8 & ~n50 ;
  assign n262 = x2 & ~n241 ;
  assign n263 = n261 | n262 ;
  assign n264 = x1 & x9 ;
  assign n265 = x2 & n264 ;
  assign n266 = x6 & n244 ;
  assign n267 = ( x6 & n265 ) | ( x6 & n266 ) | ( n265 & n266 ) ;
  assign n268 = n263 | n267 ;
  assign n269 = x3 & n268 ;
  assign n270 = n95 & ~n264 ;
  assign n271 = n153 | n270 ;
  assign n272 = x6 & ~n12 ;
  assign n273 = x8 & ~n19 ;
  assign n274 = ~n272 & n273 ;
  assign n275 = ( ~x8 & n271 ) | ( ~x8 & n274 ) | ( n271 & n274 ) ;
  assign n276 = x2 | n275 ;
  assign n277 = ~n269 & n276 ;
  assign n278 = n146 & ~n277 ;
  assign n279 = n260 | n278 ;
  assign n280 = ~x4 & n279 ;
  assign n281 = n115 & ~n254 ;
  assign n282 = ~x5 & n281 ;
  assign n283 = ~x3 & x4 ;
  assign n284 = ~x2 & n283 ;
  assign n285 = ~x1 & n284 ;
  assign n286 = ~n282 & n285 ;
  assign n287 = x2 & ~n215 ;
  assign n288 = ( ~x1 & n71 ) | ( ~x1 & n149 ) | ( n71 & n149 ) ;
  assign n289 = n287 | n288 ;
  assign n290 = x5 & n289 ;
  assign n291 = x6 & ~x8 ;
  assign n292 = ~x3 & x9 ;
  assign n293 = x1 & n292 ;
  assign n294 = n291 & n293 ;
  assign n295 = x1 & n207 ;
  assign n296 = ( x6 & x9 ) | ( x6 & ~n295 ) | ( x9 & ~n295 ) ;
  assign n297 = ~x2 & n296 ;
  assign n298 = ~x1 & n210 ;
  assign n299 = x3 & n298 ;
  assign n300 = ( x3 & n297 ) | ( x3 & n299 ) | ( n297 & n299 ) ;
  assign n301 = n294 | n300 ;
  assign n302 = n290 | n301 ;
  assign n303 = n33 | n210 ;
  assign n304 = x6 | n292 ;
  assign n305 = n303 & ~n304 ;
  assign n306 = x2 & ~x5 ;
  assign n307 = ~x3 & x8 ;
  assign n308 = ( x8 & n306 ) | ( x8 & n307 ) | ( n306 & n307 ) ;
  assign n309 = x3 & ~n145 ;
  assign n310 = x5 & ~n309 ;
  assign n311 = n308 | n310 ;
  assign n312 = x1 & n311 ;
  assign n313 = ~x5 & x6 ;
  assign n314 = ~x8 & n313 ;
  assign n315 = ~n126 & n314 ;
  assign n316 = ~x9 & n315 ;
  assign n317 = ( ~x9 & n312 ) | ( ~x9 & n316 ) | ( n312 & n316 ) ;
  assign n318 = n305 | n317 ;
  assign n319 = n302 | n318 ;
  assign n320 = x4 | n286 ;
  assign n321 = n319 & ~n320 ;
  assign n322 = ( ~x0 & n286 ) | ( ~x0 & n321 ) | ( n286 & n321 ) ;
  assign n323 = ~x7 & n322 ;
  assign n324 = ( ~x7 & n280 ) | ( ~x7 & n323 ) | ( n280 & n323 ) ;
  assign n325 = n39 & n62 ;
  assign n326 = x1 & ~n61 ;
  assign n327 = ( x1 & n325 ) | ( x1 & n326 ) | ( n325 & n326 ) ;
  assign n328 = n17 & ~n165 ;
  assign n329 = ~x4 & n328 ;
  assign n330 = ( ~x4 & n327 ) | ( ~x4 & n329 ) | ( n327 & n329 ) ;
  assign n331 = x5 | x6 ;
  assign n332 = n28 | n331 ;
  assign n333 = n330 & ~n332 ;
  assign n334 = n324 | n333 ;
  assign n335 = x3 & ~n114 ;
  assign n336 = n162 | n335 ;
  assign n337 = ~x4 & n336 ;
  assign n338 = x8 & x9 ;
  assign n339 = ~n331 & n338 ;
  assign n340 = n121 | n339 ;
  assign n341 = n284 & n340 ;
  assign n342 = n337 | n341 ;
  assign n343 = ~x1 & n342 ;
  assign n344 = x5 & x8 ;
  assign n345 = n114 & n344 ;
  assign n346 = n184 & ~n345 ;
  assign n347 = x2 & ~n346 ;
  assign n348 = x3 & x5 ;
  assign n349 = ~n215 & n348 ;
  assign n350 = ( x3 & n314 ) | ( x3 & ~n349 ) | ( n314 & ~n349 ) ;
  assign n351 = n347 | n350 ;
  assign n352 = x1 & n351 ;
  assign n353 = x2 & n313 ;
  assign n354 = n352 | n353 ;
  assign n355 = ~x4 & n354 ;
  assign n356 = n343 | n355 ;
  assign n357 = ~x0 & n356 ;
  assign n358 = ( x3 & n11 ) | ( x3 & n210 ) | ( n11 & n210 ) ;
  assign n359 = ~x2 & n358 ;
  assign n360 = x6 | n132 ;
  assign n361 = x3 & ~x5 ;
  assign n362 = n360 & ~n361 ;
  assign n363 = n359 | n362 ;
  assign n364 = ( x2 & ~x9 ) | ( x2 & n344 ) | ( ~x9 & n344 ) ;
  assign n365 = ( x2 & x9 ) | ( x2 & n154 ) | ( x9 & n154 ) ;
  assign n366 = n364 & ~n365 ;
  assign n367 = n363 | n366 ;
  assign n368 = x1 & n367 ;
  assign n369 = ~x3 & n313 ;
  assign n370 = n157 & ~n168 ;
  assign n371 = n369 | n370 ;
  assign n372 = ~x9 & n371 ;
  assign n373 = n368 | n372 ;
  assign n374 = x0 & n373 ;
  assign n375 = n28 & n313 ;
  assign n376 = x3 & ~x6 ;
  assign n377 = x2 & n376 ;
  assign n378 = n375 | n377 ;
  assign n379 = x9 & n378 ;
  assign n380 = ~x9 & n313 ;
  assign n381 = n376 | n380 ;
  assign n382 = ~x8 & n381 ;
  assign n383 = n379 | n382 ;
  assign n384 = ~x1 & n383 ;
  assign n385 = n45 & n115 ;
  assign n386 = x2 | n385 ;
  assign n387 = x5 & x9 ;
  assign n388 = x6 | n387 ;
  assign n389 = n264 | n344 ;
  assign n390 = ~n388 & n389 ;
  assign n391 = n386 & ~n390 ;
  assign n392 = x3 & ~n391 ;
  assign n393 = x1 & n254 ;
  assign n394 = n313 & n393 ;
  assign n395 = n392 | n394 ;
  assign n396 = n384 | n395 ;
  assign n397 = n374 | n396 ;
  assign n398 = ~x4 & n397 ;
  assign n399 = n357 | n398 ;
  assign n400 = ~x7 & n399 ;
  assign n401 = x3 & ~x4 ;
  assign n402 = x0 | n133 ;
  assign n403 = ( x3 & x4 ) | ( x3 & n402 ) | ( x4 & n402 ) ;
  assign n404 = x4 | n227 ;
  assign n405 = ( n401 & ~n403 ) | ( n401 & n404 ) | ( ~n403 & n404 ) ;
  assign n406 = ~x7 & n405 ;
  assign n407 = n121 & n406 ;
  assign n408 = ~n51 & n284 ;
  assign n409 = n401 & n402 ;
  assign n410 = n408 | n409 ;
  assign n411 = ~x7 & n410 ;
  assign n412 = n121 & n411 ;
  assign n413 = ~x1 & x4 ;
  assign n414 = n121 | n413 ;
  assign n415 = ( ~n103 & n121 ) | ( ~n103 & n414 ) | ( n121 & n414 ) ;
  assign n416 = ~x7 & n415 ;
  assign n417 = x0 | x8 ;
  assign n418 = ~n146 & n417 ;
  assign n419 = n19 & n418 ;
  assign n420 = x0 & n207 ;
  assign n421 = ~x2 & n92 ;
  assign n422 = ( ~x2 & n420 ) | ( ~x2 & n421 ) | ( n420 & n421 ) ;
  assign n423 = ~x8 & n169 ;
  assign n424 = x9 & n423 ;
  assign n425 = ( x9 & n422 ) | ( x9 & n424 ) | ( n422 & n424 ) ;
  assign n426 = n419 | n425 ;
  assign n427 = x2 & n19 ;
  assign n428 = x0 & n264 ;
  assign n429 = ( x0 & ~n104 ) | ( x0 & n428 ) | ( ~n104 & n428 ) ;
  assign n430 = n427 | n429 ;
  assign n431 = x0 | x6 ;
  assign n432 = n165 & ~n431 ;
  assign n433 = n270 & n432 ;
  assign n434 = ~x5 & n433 ;
  assign n435 = ( ~x5 & n430 ) | ( ~x5 & n434 ) | ( n430 & n434 ) ;
  assign n436 = n426 | n435 ;
  assign n437 = x3 & n436 ;
  assign n438 = x2 & x8 ;
  assign n439 = n13 & n438 ;
  assign n440 = ~x8 & n431 ;
  assign n441 = ~x9 & n146 ;
  assign n442 = ( ~x9 & n440 ) | ( ~x9 & n441 ) | ( n440 & n441 ) ;
  assign n443 = x2 & ~n439 ;
  assign n444 = ( n439 & n442 ) | ( n439 & ~n443 ) | ( n442 & ~n443 ) ;
  assign n445 = ~x1 & n444 ;
  assign n446 = ~x2 & x5 ;
  assign n447 = ~n63 & n446 ;
  assign n448 = x6 | n306 ;
  assign n449 = n13 & n448 ;
  assign n450 = n447 | n449 ;
  assign n451 = ~x8 & n450 ;
  assign n452 = x2 & n241 ;
  assign n453 = n248 | n452 ;
  assign n454 = x6 & n453 ;
  assign n455 = x1 & n454 ;
  assign n456 = ( x1 & n451 ) | ( x1 & n455 ) | ( n451 & n455 ) ;
  assign n457 = n445 | n456 ;
  assign n458 = n437 | n457 ;
  assign n459 = ~x7 & n458 ;
  assign n460 = x3 | x4 ;
  assign n461 = x5 & n264 ;
  assign n462 = x0 & n461 ;
  assign n463 = x6 | x9 ;
  assign n464 = x1 | x5 ;
  assign n465 = ( x2 & n463 ) | ( x2 & n464 ) | ( n463 & n464 ) ;
  assign n466 = n463 | n465 ;
  assign n467 = ( x0 & n462 ) | ( x0 & ~n466 ) | ( n462 & ~n466 ) ;
  assign n468 = ~x0 & x2 ;
  assign n469 = n45 & n468 ;
  assign n470 = x8 & n469 ;
  assign n471 = ( x8 & n467 ) | ( x8 & n470 ) | ( n467 & n470 ) ;
  assign n472 = x2 & n13 ;
  assign n473 = n104 & ~n472 ;
  assign n474 = x5 & ~n473 ;
  assign n475 = n241 & ~n338 ;
  assign n476 = x6 & ~n475 ;
  assign n477 = ~x2 & x9 ;
  assign n478 = n50 | n477 ;
  assign n479 = n476 & ~n478 ;
  assign n480 = n474 | n479 ;
  assign n481 = n471 | n480 ;
  assign n482 = ~x7 & n481 ;
  assign n483 = n188 & n264 ;
  assign n484 = x7 & ~n241 ;
  assign n485 = ( x7 & n483 ) | ( x7 & n484 ) | ( n483 & n484 ) ;
  assign n486 = ~x2 & n485 ;
  assign n487 = ~x0 & n83 ;
  assign n488 = x7 & n254 ;
  assign n489 = ( ~x8 & n71 ) | ( ~x8 & n488 ) | ( n71 & n488 ) ;
  assign n490 = ( ~x0 & n487 ) | ( ~x0 & n489 ) | ( n487 & n489 ) ;
  assign n491 = n486 | n490 ;
  assign n492 = ~n331 & n491 ;
  assign n493 = ( ~n460 & n482 ) | ( ~n460 & n492 ) | ( n482 & n492 ) ;
  assign n494 = ~n460 & n493 ;
  assign n495 = ( ~x4 & n459 ) | ( ~x4 & n494 ) | ( n459 & n494 ) ;
  assign n496 = n416 | n495 ;
  assign n497 = x3 & ~n338 ;
  assign n498 = ~x6 & n188 ;
  assign n499 = ( ~x6 & n497 ) | ( ~x6 & n498 ) | ( n497 & n498 ) ;
  assign n500 = ~x3 & n338 ;
  assign n501 = x2 & n500 ;
  assign n502 = ( x2 & n499 ) | ( x2 & n501 ) | ( n499 & n501 ) ;
  assign n503 = x6 | n241 ;
  assign n504 = x3 | n503 ;
  assign n505 = ~n502 & n504 ;
  assign n506 = ( x6 & x8 ) | ( x6 & x9 ) | ( x8 & x9 ) ;
  assign n507 = n171 & n376 ;
  assign n508 = x9 & ~n507 ;
  assign n509 = ( n210 & n506 ) | ( n210 & ~n508 ) | ( n506 & ~n508 ) ;
  assign n510 = ( n48 & n180 ) | ( n48 & n307 ) | ( n180 & n307 ) ;
  assign n511 = n48 & n510 ;
  assign n512 = ( ~x2 & n509 ) | ( ~x2 & n511 ) | ( n509 & n511 ) ;
  assign n513 = n505 & ~n512 ;
  assign n514 = ~x9 & n291 ;
  assign n515 = n164 & n514 ;
  assign n516 = ( x1 & ~n513 ) | ( x1 & n515 ) | ( ~n513 & n515 ) ;
  assign n517 = n61 & ~n210 ;
  assign n518 = x2 | x6 ;
  assign n519 = n517 | n518 ;
  assign n520 = n202 & ~n475 ;
  assign n521 = n519 & ~n520 ;
  assign n522 = x3 & ~n521 ;
  assign n523 = x0 | n156 ;
  assign n524 = ~n420 & n523 ;
  assign n525 = x9 | n524 ;
  assign n526 = ~x6 & n153 ;
  assign n527 = n452 & ~n526 ;
  assign n528 = n525 & ~n527 ;
  assign n529 = ~n522 & n528 ;
  assign n530 = ( x1 & ~n515 ) | ( x1 & n529 ) | ( ~n515 & n529 ) ;
  assign n531 = ~n516 & n530 ;
  assign n532 = x5 | n531 ;
  assign n533 = x5 & ~x9 ;
  assign n534 = n164 & n533 ;
  assign n535 = n50 | n348 ;
  assign n536 = ~x0 & n535 ;
  assign n537 = x3 & n446 ;
  assign n538 = ~x8 & n537 ;
  assign n539 = ( ~x8 & n536 ) | ( ~x8 & n538 ) | ( n536 & n538 ) ;
  assign n540 = n534 | n539 ;
  assign n541 = n82 & n139 ;
  assign n542 = ~x3 & n541 ;
  assign n543 = ( x0 & x8 ) | ( x0 & n533 ) | ( x8 & n533 ) ;
  assign n544 = ( ~x0 & x8 ) | ( ~x0 & n478 ) | ( x8 & n478 ) ;
  assign n545 = n543 & n544 ;
  assign n546 = ( ~x3 & n542 ) | ( ~x3 & n545 ) | ( n542 & n545 ) ;
  assign n547 = n540 | n546 ;
  assign n548 = x1 & n547 ;
  assign n549 = x2 & x3 ;
  assign n550 = x8 & n387 ;
  assign n551 = n549 & n550 ;
  assign n552 = x2 | n30 ;
  assign n553 = ~n475 & n552 ;
  assign n554 = x5 & n549 ;
  assign n555 = ( x5 & n553 ) | ( x5 & n554 ) | ( n553 & n554 ) ;
  assign n556 = n30 & n262 ;
  assign n557 = ~x1 & n556 ;
  assign n558 = ( ~x1 & n555 ) | ( ~x1 & n557 ) | ( n555 & n557 ) ;
  assign n559 = n551 | n558 ;
  assign n560 = ~x6 & n559 ;
  assign n561 = ( ~x6 & n548 ) | ( ~x6 & n560 ) | ( n548 & n560 ) ;
  assign n562 = ~x7 & n561 ;
  assign n563 = ( x7 & n532 ) | ( x7 & ~n562 ) | ( n532 & ~n562 ) ;
  assign n564 = n24 | n85 ;
  assign n565 = x4 & ~x7 ;
  assign n566 = ~n168 & n565 ;
  assign n567 = ~n564 & n566 ;
  assign n568 = x4 & ~n567 ;
  assign n569 = ~x9 & n39 ;
  assign n570 = n48 & n569 ;
  assign n571 = n255 & n468 ;
  assign n572 = n570 | n571 ;
  assign n573 = n11 | n168 ;
  assign n574 = n572 & ~n573 ;
  assign n575 = ( n567 & ~n568 ) | ( n567 & n574 ) | ( ~n568 & n574 ) ;
  assign n576 = ( n563 & n568 ) | ( n563 & ~n575 ) | ( n568 & ~n575 ) ;
  assign n577 = ~n11 & n565 ;
  assign n578 = ~n402 & n577 ;
  assign n579 = n156 & ~n438 ;
  assign n580 = x0 | n579 ;
  assign n581 = x0 & n145 ;
  assign n582 = ~x9 & n581 ;
  assign n583 = ( x9 & n580 ) | ( x9 & ~n582 ) | ( n580 & ~n582 ) ;
  assign n584 = n264 & ~n523 ;
  assign n585 = x1 & ~n584 ;
  assign n586 = n82 & ~n417 ;
  assign n587 = ( n584 & ~n585 ) | ( n584 & n586 ) | ( ~n585 & n586 ) ;
  assign n588 = ( n583 & n585 ) | ( n583 & ~n587 ) | ( n585 & ~n587 ) ;
  assign n589 = n225 | n588 ;
  assign n590 = ~x2 & n85 ;
  assign n591 = n135 | n361 ;
  assign n592 = n590 & ~n591 ;
  assign n593 = ~n126 & n146 ;
  assign n594 = x8 & n593 ;
  assign n595 = ( x8 & n592 ) | ( x8 & n594 ) | ( n592 & n594 ) ;
  assign n596 = x5 | n171 ;
  assign n597 = n25 & ~n348 ;
  assign n598 = n596 & n597 ;
  assign n599 = ~x9 & n598 ;
  assign n600 = ( ~x9 & n595 ) | ( ~x9 & n599 ) | ( n595 & n599 ) ;
  assign n601 = ( x3 & ~x8 ) | ( x3 & n549 ) | ( ~x8 & n549 ) ;
  assign n602 = ( n306 & n348 ) | ( n306 & ~n601 ) | ( n348 & ~n601 ) ;
  assign n603 = x1 & n602 ;
  assign n604 = ~n144 & n239 ;
  assign n605 = n145 & n604 ;
  assign n606 = x9 & n605 ;
  assign n607 = ( x9 & n603 ) | ( x9 & n606 ) | ( n603 & n606 ) ;
  assign n608 = n600 | n607 ;
  assign n609 = n95 & ~n292 ;
  assign n610 = ~n591 & n609 ;
  assign n611 = ~x2 & n610 ;
  assign n612 = n90 & ~n464 ;
  assign n613 = ( n90 & ~n270 ) | ( n90 & n612 ) | ( ~n270 & n612 ) ;
  assign n614 = n611 | n613 ;
  assign n615 = ~n133 & n533 ;
  assign n616 = ( n293 & ~n417 ) | ( n293 & n615 ) | ( ~n417 & n615 ) ;
  assign n617 = ~n417 & n616 ;
  assign n618 = ( ~x8 & n614 ) | ( ~x8 & n617 ) | ( n614 & n617 ) ;
  assign n619 = n608 | n618 ;
  assign n620 = ( x2 & n25 ) | ( x2 & ~n241 ) | ( n25 & ~n241 ) ;
  assign n621 = n272 | n620 ;
  assign n622 = x0 & n621 ;
  assign n623 = ( x2 & n92 ) | ( x2 & n162 ) | ( n92 & n162 ) ;
  assign n624 = ( ~x8 & n272 ) | ( ~x8 & n393 ) | ( n272 & n393 ) ;
  assign n625 = n623 | n624 ;
  assign n626 = n622 | n625 ;
  assign n627 = n361 & n626 ;
  assign n628 = x6 & ~n627 ;
  assign n629 = ( n619 & n627 ) | ( n619 & ~n628 ) | ( n627 & ~n628 ) ;
  assign n630 = ~x7 & n589 ;
  assign n631 = n629 & n630 ;
  assign n632 = ( x4 & n589 ) | ( x4 & ~n631 ) | ( n589 & ~n631 ) ;
  assign n633 = ~n578 & n632 ;
  assign n634 = n171 | n180 ;
  assign n635 = ( n180 & n388 ) | ( n180 & n634 ) | ( n388 & n634 ) ;
  assign n636 = ( x3 & n331 ) | ( x3 & n460 ) | ( n331 & n460 ) ;
  assign n637 = ~x3 & n636 ;
  assign n638 = ( ~n635 & n636 ) | ( ~n635 & n637 ) | ( n636 & n637 ) ;
  assign n639 = x2 | n638 ;
  assign n640 = ~x3 & n45 ;
  assign n641 = x8 | n387 ;
  assign n642 = ( ~n71 & n640 ) | ( ~n71 & n641 ) | ( n640 & n641 ) ;
  assign n643 = n71 & n642 ;
  assign n644 = ( x1 & n639 ) | ( x1 & ~n643 ) | ( n639 & ~n643 ) ;
  assign n645 = ( x6 & n90 ) | ( x6 & n121 ) | ( n90 & n121 ) ;
  assign n646 = n644 & ~n645 ;
  assign n647 = x7 & ~n90 ;
  assign n648 = ( x6 & n115 ) | ( x6 & n387 ) | ( n115 & n387 ) ;
  assign n649 = ~x3 & n648 ;
  assign n650 = x5 | n338 ;
  assign n651 = n377 & ~n650 ;
  assign n652 = n649 | n651 ;
  assign n653 = x3 & ~n180 ;
  assign n654 = n171 & ~n653 ;
  assign n655 = ~x2 & n640 ;
  assign n656 = ( ~x2 & n654 ) | ( ~x2 & n655 ) | ( n654 & n655 ) ;
  assign n657 = n652 | n656 ;
  assign n658 = x1 & n657 ;
  assign n659 = n647 | n658 ;
  assign n660 = n646 & ~n659 ;
  assign n661 = ~x1 & n241 ;
  assign n662 = x7 | n146 ;
  assign n663 = ( x7 & n377 ) | ( x7 & n662 ) | ( n377 & n662 ) ;
  assign n664 = ~n661 & n663 ;
  assign n665 = x2 | n126 ;
  assign n666 = ~x7 & n665 ;
  assign n667 = x0 & ~n666 ;
  assign n668 = n664 | n667 ;
  assign n669 = x4 & n665 ;
  assign n670 = n668 | n669 ;
  assign n671 = n660 & ~n670 ;
  assign n672 = ( ~x8 & n14 ) | ( ~x8 & n18 ) | ( n14 & n18 ) ;
  assign n673 = n401 & n672 ;
  assign n674 = x2 & n673 ;
  assign n675 = n408 | n674 ;
  assign n676 = ~x7 & n675 ;
  assign n677 = ~n331 & n676 ;
  assign y0 = ~n129 ;
  assign y1 = n238 ;
  assign y2 = n334 ;
  assign y3 = n400 ;
  assign y4 = n407 ;
  assign y5 = n412 ;
  assign y6 = ~n496 ;
  assign y7 = n576 ;
  assign y8 = n633 ;
  assign y9 = n671 ;
  assign y10 = n677 ;
endmodule
