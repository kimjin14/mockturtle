module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 ;
  assign n129 = x126 & x127 ;
  assign n130 = x125 & ~x126 ;
  assign n131 = ( x125 & n129 ) | ( x125 & n130 ) | ( n129 & n130 ) ;
  assign n132 = ~x125 & x127 ;
  assign n133 = x124 & n132 ;
  assign n134 = ( x124 & n131 ) | ( x124 & n133 ) | ( n131 & n133 ) ;
  assign n135 = x124 | x126 ;
  assign n136 = ( x124 & ~n129 ) | ( x124 & n135 ) | ( ~n129 & n135 ) ;
  assign n137 = x123 & ~n136 ;
  assign n138 = ( x123 & n134 ) | ( x123 & n137 ) | ( n134 & n137 ) ;
  assign n139 = ~x123 & n132 ;
  assign n140 = ( ~x123 & n131 ) | ( ~x123 & n139 ) | ( n131 & n139 ) ;
  assign n141 = x122 & n140 ;
  assign n142 = ( x122 & n138 ) | ( x122 & n141 ) | ( n138 & n141 ) ;
  assign n143 = x122 | n136 ;
  assign n144 = ( x122 & ~n134 ) | ( x122 & n143 ) | ( ~n134 & n143 ) ;
  assign n145 = x121 & ~n144 ;
  assign n146 = ( x121 & n142 ) | ( x121 & n145 ) | ( n142 & n145 ) ;
  assign n147 = ~x121 & n140 ;
  assign n148 = ( ~x121 & n138 ) | ( ~x121 & n147 ) | ( n138 & n147 ) ;
  assign n149 = x120 & n148 ;
  assign n150 = ( x120 & n146 ) | ( x120 & n149 ) | ( n146 & n149 ) ;
  assign n151 = x120 | n144 ;
  assign n152 = ( x120 & ~n142 ) | ( x120 & n151 ) | ( ~n142 & n151 ) ;
  assign n153 = x119 & ~n152 ;
  assign n154 = ( x119 & n150 ) | ( x119 & n153 ) | ( n150 & n153 ) ;
  assign n155 = ~x119 & n148 ;
  assign n156 = ( ~x119 & n146 ) | ( ~x119 & n155 ) | ( n146 & n155 ) ;
  assign n157 = x118 & n156 ;
  assign n158 = ( x118 & n154 ) | ( x118 & n157 ) | ( n154 & n157 ) ;
  assign n159 = x118 | n152 ;
  assign n160 = ( x118 & ~n150 ) | ( x118 & n159 ) | ( ~n150 & n159 ) ;
  assign n161 = x117 & ~n160 ;
  assign n162 = ( x117 & n158 ) | ( x117 & n161 ) | ( n158 & n161 ) ;
  assign n163 = ~x117 & n156 ;
  assign n164 = ( ~x117 & n154 ) | ( ~x117 & n163 ) | ( n154 & n163 ) ;
  assign n165 = x116 & n164 ;
  assign n166 = ( x116 & n162 ) | ( x116 & n165 ) | ( n162 & n165 ) ;
  assign n167 = x116 | n160 ;
  assign n168 = ( x116 & ~n158 ) | ( x116 & n167 ) | ( ~n158 & n167 ) ;
  assign n169 = x115 & ~n168 ;
  assign n170 = ( x115 & n166 ) | ( x115 & n169 ) | ( n166 & n169 ) ;
  assign n171 = ~x115 & n164 ;
  assign n172 = ( ~x115 & n162 ) | ( ~x115 & n171 ) | ( n162 & n171 ) ;
  assign n173 = x114 & n172 ;
  assign n174 = ( x114 & n170 ) | ( x114 & n173 ) | ( n170 & n173 ) ;
  assign n175 = x114 | n168 ;
  assign n176 = ( x114 & ~n166 ) | ( x114 & n175 ) | ( ~n166 & n175 ) ;
  assign n177 = x113 & ~n176 ;
  assign n178 = ( x113 & n174 ) | ( x113 & n177 ) | ( n174 & n177 ) ;
  assign n179 = ~x113 & n172 ;
  assign n180 = ( ~x113 & n170 ) | ( ~x113 & n179 ) | ( n170 & n179 ) ;
  assign n181 = x112 & n180 ;
  assign n182 = ( x112 & n178 ) | ( x112 & n181 ) | ( n178 & n181 ) ;
  assign n183 = x112 | n176 ;
  assign n184 = ( x112 & ~n174 ) | ( x112 & n183 ) | ( ~n174 & n183 ) ;
  assign n185 = x111 & ~n184 ;
  assign n186 = ( x111 & n182 ) | ( x111 & n185 ) | ( n182 & n185 ) ;
  assign n187 = ~x111 & n180 ;
  assign n188 = ( ~x111 & n178 ) | ( ~x111 & n187 ) | ( n178 & n187 ) ;
  assign n189 = x110 & n188 ;
  assign n190 = ( x110 & n186 ) | ( x110 & n189 ) | ( n186 & n189 ) ;
  assign n191 = x110 | n184 ;
  assign n192 = ( x110 & ~n182 ) | ( x110 & n191 ) | ( ~n182 & n191 ) ;
  assign n193 = x109 & ~n192 ;
  assign n194 = ( x109 & n190 ) | ( x109 & n193 ) | ( n190 & n193 ) ;
  assign n195 = ~x109 & n188 ;
  assign n196 = ( ~x109 & n186 ) | ( ~x109 & n195 ) | ( n186 & n195 ) ;
  assign n197 = x108 & n196 ;
  assign n198 = ( x108 & n194 ) | ( x108 & n197 ) | ( n194 & n197 ) ;
  assign n199 = x108 | n192 ;
  assign n200 = ( x108 & ~n190 ) | ( x108 & n199 ) | ( ~n190 & n199 ) ;
  assign n201 = x107 & ~n200 ;
  assign n202 = ( x107 & n198 ) | ( x107 & n201 ) | ( n198 & n201 ) ;
  assign n203 = ~x107 & n196 ;
  assign n204 = ( ~x107 & n194 ) | ( ~x107 & n203 ) | ( n194 & n203 ) ;
  assign n205 = x106 & n204 ;
  assign n206 = ( x106 & n202 ) | ( x106 & n205 ) | ( n202 & n205 ) ;
  assign n207 = x106 | n200 ;
  assign n208 = ( x106 & ~n198 ) | ( x106 & n207 ) | ( ~n198 & n207 ) ;
  assign n209 = x105 & ~n208 ;
  assign n210 = ( x105 & n206 ) | ( x105 & n209 ) | ( n206 & n209 ) ;
  assign n211 = ~x105 & n204 ;
  assign n212 = ( ~x105 & n202 ) | ( ~x105 & n211 ) | ( n202 & n211 ) ;
  assign n213 = x104 & n212 ;
  assign n214 = ( x104 & n210 ) | ( x104 & n213 ) | ( n210 & n213 ) ;
  assign n215 = x104 | n208 ;
  assign n216 = ( x104 & ~n206 ) | ( x104 & n215 ) | ( ~n206 & n215 ) ;
  assign n217 = x103 & ~n216 ;
  assign n218 = ( x103 & n214 ) | ( x103 & n217 ) | ( n214 & n217 ) ;
  assign n219 = ~x103 & n212 ;
  assign n220 = ( ~x103 & n210 ) | ( ~x103 & n219 ) | ( n210 & n219 ) ;
  assign n221 = x102 & n220 ;
  assign n222 = ( x102 & n218 ) | ( x102 & n221 ) | ( n218 & n221 ) ;
  assign n223 = x102 | n216 ;
  assign n224 = ( x102 & ~n214 ) | ( x102 & n223 ) | ( ~n214 & n223 ) ;
  assign n225 = x101 & ~n224 ;
  assign n226 = ( x101 & n222 ) | ( x101 & n225 ) | ( n222 & n225 ) ;
  assign n227 = ~x101 & n220 ;
  assign n228 = ( ~x101 & n218 ) | ( ~x101 & n227 ) | ( n218 & n227 ) ;
  assign n229 = x100 & n228 ;
  assign n230 = ( x100 & n226 ) | ( x100 & n229 ) | ( n226 & n229 ) ;
  assign n231 = x100 | n224 ;
  assign n232 = ( x100 & ~n222 ) | ( x100 & n231 ) | ( ~n222 & n231 ) ;
  assign n233 = x99 & ~n232 ;
  assign n234 = ( x99 & n230 ) | ( x99 & n233 ) | ( n230 & n233 ) ;
  assign n235 = ~x99 & n228 ;
  assign n236 = ( ~x99 & n226 ) | ( ~x99 & n235 ) | ( n226 & n235 ) ;
  assign n237 = x98 & n236 ;
  assign n238 = ( x98 & n234 ) | ( x98 & n237 ) | ( n234 & n237 ) ;
  assign n239 = x98 | n232 ;
  assign n240 = ( x98 & ~n230 ) | ( x98 & n239 ) | ( ~n230 & n239 ) ;
  assign n241 = x97 & ~n240 ;
  assign n242 = ( x97 & n238 ) | ( x97 & n241 ) | ( n238 & n241 ) ;
  assign n243 = ~x97 & n236 ;
  assign n244 = ( ~x97 & n234 ) | ( ~x97 & n243 ) | ( n234 & n243 ) ;
  assign n245 = x96 & n244 ;
  assign n246 = ( x96 & n242 ) | ( x96 & n245 ) | ( n242 & n245 ) ;
  assign n247 = x96 | n240 ;
  assign n248 = ( x96 & ~n238 ) | ( x96 & n247 ) | ( ~n238 & n247 ) ;
  assign n249 = x95 & ~n248 ;
  assign n250 = ( x95 & n246 ) | ( x95 & n249 ) | ( n246 & n249 ) ;
  assign n251 = ~x95 & n244 ;
  assign n252 = ( ~x95 & n242 ) | ( ~x95 & n251 ) | ( n242 & n251 ) ;
  assign n253 = x94 & n252 ;
  assign n254 = ( x94 & n250 ) | ( x94 & n253 ) | ( n250 & n253 ) ;
  assign n255 = x94 | n248 ;
  assign n256 = ( x94 & ~n246 ) | ( x94 & n255 ) | ( ~n246 & n255 ) ;
  assign n257 = x93 & ~n256 ;
  assign n258 = ( x93 & n254 ) | ( x93 & n257 ) | ( n254 & n257 ) ;
  assign n259 = ~x93 & n252 ;
  assign n260 = ( ~x93 & n250 ) | ( ~x93 & n259 ) | ( n250 & n259 ) ;
  assign n261 = x92 & n260 ;
  assign n262 = ( x92 & n258 ) | ( x92 & n261 ) | ( n258 & n261 ) ;
  assign n263 = x92 | n256 ;
  assign n264 = ( x92 & ~n254 ) | ( x92 & n263 ) | ( ~n254 & n263 ) ;
  assign n265 = x91 & ~n264 ;
  assign n266 = ( x91 & n262 ) | ( x91 & n265 ) | ( n262 & n265 ) ;
  assign n267 = ~x91 & n260 ;
  assign n268 = ( ~x91 & n258 ) | ( ~x91 & n267 ) | ( n258 & n267 ) ;
  assign n269 = x90 & n268 ;
  assign n270 = ( x90 & n266 ) | ( x90 & n269 ) | ( n266 & n269 ) ;
  assign n271 = x90 | n264 ;
  assign n272 = ( x90 & ~n262 ) | ( x90 & n271 ) | ( ~n262 & n271 ) ;
  assign n273 = x89 & ~n272 ;
  assign n274 = ( x89 & n270 ) | ( x89 & n273 ) | ( n270 & n273 ) ;
  assign n275 = ~x89 & n268 ;
  assign n276 = ( ~x89 & n266 ) | ( ~x89 & n275 ) | ( n266 & n275 ) ;
  assign n277 = x88 & n276 ;
  assign n278 = ( x88 & n274 ) | ( x88 & n277 ) | ( n274 & n277 ) ;
  assign n279 = x88 | n272 ;
  assign n280 = ( x88 & ~n270 ) | ( x88 & n279 ) | ( ~n270 & n279 ) ;
  assign n281 = x87 & ~n280 ;
  assign n282 = ( x87 & n278 ) | ( x87 & n281 ) | ( n278 & n281 ) ;
  assign n283 = ~x87 & n276 ;
  assign n284 = ( ~x87 & n274 ) | ( ~x87 & n283 ) | ( n274 & n283 ) ;
  assign n285 = x86 & n284 ;
  assign n286 = ( x86 & n282 ) | ( x86 & n285 ) | ( n282 & n285 ) ;
  assign n287 = x86 | n280 ;
  assign n288 = ( x86 & ~n278 ) | ( x86 & n287 ) | ( ~n278 & n287 ) ;
  assign n289 = x85 & ~n288 ;
  assign n290 = ( x85 & n286 ) | ( x85 & n289 ) | ( n286 & n289 ) ;
  assign n291 = ~x85 & n284 ;
  assign n292 = ( ~x85 & n282 ) | ( ~x85 & n291 ) | ( n282 & n291 ) ;
  assign n293 = x84 & n292 ;
  assign n294 = ( x84 & n290 ) | ( x84 & n293 ) | ( n290 & n293 ) ;
  assign n295 = x84 | n288 ;
  assign n296 = ( x84 & ~n286 ) | ( x84 & n295 ) | ( ~n286 & n295 ) ;
  assign n297 = x83 & ~n296 ;
  assign n298 = ( x83 & n294 ) | ( x83 & n297 ) | ( n294 & n297 ) ;
  assign n299 = ~x83 & n292 ;
  assign n300 = ( ~x83 & n290 ) | ( ~x83 & n299 ) | ( n290 & n299 ) ;
  assign n301 = x82 & n300 ;
  assign n302 = ( x82 & n298 ) | ( x82 & n301 ) | ( n298 & n301 ) ;
  assign n303 = x82 | n296 ;
  assign n304 = ( x82 & ~n294 ) | ( x82 & n303 ) | ( ~n294 & n303 ) ;
  assign n305 = x81 & ~n304 ;
  assign n306 = ( x81 & n302 ) | ( x81 & n305 ) | ( n302 & n305 ) ;
  assign n307 = ~x81 & n300 ;
  assign n308 = ( ~x81 & n298 ) | ( ~x81 & n307 ) | ( n298 & n307 ) ;
  assign n309 = x80 & n308 ;
  assign n310 = ( x80 & n306 ) | ( x80 & n309 ) | ( n306 & n309 ) ;
  assign n311 = x80 | n304 ;
  assign n312 = ( x80 & ~n302 ) | ( x80 & n311 ) | ( ~n302 & n311 ) ;
  assign n313 = x79 & ~n312 ;
  assign n314 = ( x79 & n310 ) | ( x79 & n313 ) | ( n310 & n313 ) ;
  assign n315 = ~x79 & n308 ;
  assign n316 = ( ~x79 & n306 ) | ( ~x79 & n315 ) | ( n306 & n315 ) ;
  assign n317 = x78 & n316 ;
  assign n318 = ( x78 & n314 ) | ( x78 & n317 ) | ( n314 & n317 ) ;
  assign n319 = x78 | n312 ;
  assign n320 = ( x78 & ~n310 ) | ( x78 & n319 ) | ( ~n310 & n319 ) ;
  assign n321 = x77 & ~n320 ;
  assign n322 = ( x77 & n318 ) | ( x77 & n321 ) | ( n318 & n321 ) ;
  assign n323 = ~x77 & n316 ;
  assign n324 = ( ~x77 & n314 ) | ( ~x77 & n323 ) | ( n314 & n323 ) ;
  assign n325 = x76 & n324 ;
  assign n326 = ( x76 & n322 ) | ( x76 & n325 ) | ( n322 & n325 ) ;
  assign n327 = x76 | n320 ;
  assign n328 = ( x76 & ~n318 ) | ( x76 & n327 ) | ( ~n318 & n327 ) ;
  assign n329 = x75 & ~n328 ;
  assign n330 = ( x75 & n326 ) | ( x75 & n329 ) | ( n326 & n329 ) ;
  assign n331 = ~x75 & n324 ;
  assign n332 = ( ~x75 & n322 ) | ( ~x75 & n331 ) | ( n322 & n331 ) ;
  assign n333 = x74 & n332 ;
  assign n334 = ( x74 & n330 ) | ( x74 & n333 ) | ( n330 & n333 ) ;
  assign n335 = x74 | n328 ;
  assign n336 = ( x74 & ~n326 ) | ( x74 & n335 ) | ( ~n326 & n335 ) ;
  assign n337 = x73 & ~n336 ;
  assign n338 = ( x73 & n334 ) | ( x73 & n337 ) | ( n334 & n337 ) ;
  assign n339 = ~x73 & n332 ;
  assign n340 = ( ~x73 & n330 ) | ( ~x73 & n339 ) | ( n330 & n339 ) ;
  assign n341 = x72 & n340 ;
  assign n342 = ( x72 & n338 ) | ( x72 & n341 ) | ( n338 & n341 ) ;
  assign n343 = x72 | n336 ;
  assign n344 = ( x72 & ~n334 ) | ( x72 & n343 ) | ( ~n334 & n343 ) ;
  assign n345 = x71 & ~n344 ;
  assign n346 = ( x71 & n342 ) | ( x71 & n345 ) | ( n342 & n345 ) ;
  assign n347 = ~x71 & n340 ;
  assign n348 = ( ~x71 & n338 ) | ( ~x71 & n347 ) | ( n338 & n347 ) ;
  assign n349 = x70 & n348 ;
  assign n350 = ( x70 & n346 ) | ( x70 & n349 ) | ( n346 & n349 ) ;
  assign n351 = x70 | n344 ;
  assign n352 = ( x70 & ~n342 ) | ( x70 & n351 ) | ( ~n342 & n351 ) ;
  assign n353 = x69 & ~n352 ;
  assign n354 = ( x69 & n350 ) | ( x69 & n353 ) | ( n350 & n353 ) ;
  assign n355 = ~x69 & n348 ;
  assign n356 = ( ~x69 & n346 ) | ( ~x69 & n355 ) | ( n346 & n355 ) ;
  assign n357 = x68 & n356 ;
  assign n358 = ( x68 & n354 ) | ( x68 & n357 ) | ( n354 & n357 ) ;
  assign n359 = x68 | n352 ;
  assign n360 = ( x68 & ~n350 ) | ( x68 & n359 ) | ( ~n350 & n359 ) ;
  assign n361 = x67 & ~n360 ;
  assign n362 = ( x67 & n358 ) | ( x67 & n361 ) | ( n358 & n361 ) ;
  assign n363 = ~x67 & n356 ;
  assign n364 = ( ~x67 & n354 ) | ( ~x67 & n363 ) | ( n354 & n363 ) ;
  assign n365 = x66 & n364 ;
  assign n366 = ( x66 & n362 ) | ( x66 & n365 ) | ( n362 & n365 ) ;
  assign n367 = x66 | n360 ;
  assign n368 = ( x66 & ~n358 ) | ( x66 & n367 ) | ( ~n358 & n367 ) ;
  assign n369 = x65 & ~n368 ;
  assign n370 = ( x65 & n366 ) | ( x65 & n369 ) | ( n366 & n369 ) ;
  assign n371 = ~x65 & n364 ;
  assign n372 = ( ~x65 & n362 ) | ( ~x65 & n371 ) | ( n362 & n371 ) ;
  assign n373 = x64 & n372 ;
  assign n374 = ( x64 & n370 ) | ( x64 & n373 ) | ( n370 & n373 ) ;
  assign n375 = x64 | n368 ;
  assign n376 = ( x64 & ~n366 ) | ( x64 & n375 ) | ( ~n366 & n375 ) ;
  assign n377 = x63 & ~n376 ;
  assign n378 = ( x63 & n374 ) | ( x63 & n377 ) | ( n374 & n377 ) ;
  assign n379 = ~x63 & n372 ;
  assign n380 = ( ~x63 & n370 ) | ( ~x63 & n379 ) | ( n370 & n379 ) ;
  assign n381 = x62 & n380 ;
  assign n382 = ( x62 & n378 ) | ( x62 & n381 ) | ( n378 & n381 ) ;
  assign n383 = x62 | n376 ;
  assign n384 = ( x62 & ~n374 ) | ( x62 & n383 ) | ( ~n374 & n383 ) ;
  assign n385 = x61 & ~n384 ;
  assign n386 = ( x61 & n382 ) | ( x61 & n385 ) | ( n382 & n385 ) ;
  assign n387 = ~x61 & n380 ;
  assign n388 = ( ~x61 & n378 ) | ( ~x61 & n387 ) | ( n378 & n387 ) ;
  assign n389 = x60 & n388 ;
  assign n390 = ( x60 & n386 ) | ( x60 & n389 ) | ( n386 & n389 ) ;
  assign n391 = x60 | n384 ;
  assign n392 = ( x60 & ~n382 ) | ( x60 & n391 ) | ( ~n382 & n391 ) ;
  assign n393 = x59 & ~n392 ;
  assign n394 = ( x59 & n390 ) | ( x59 & n393 ) | ( n390 & n393 ) ;
  assign n395 = ~x59 & n388 ;
  assign n396 = ( ~x59 & n386 ) | ( ~x59 & n395 ) | ( n386 & n395 ) ;
  assign n397 = x58 & n396 ;
  assign n398 = ( x58 & n394 ) | ( x58 & n397 ) | ( n394 & n397 ) ;
  assign n399 = x58 | n392 ;
  assign n400 = ( x58 & ~n390 ) | ( x58 & n399 ) | ( ~n390 & n399 ) ;
  assign n401 = x57 & ~n400 ;
  assign n402 = ( x57 & n398 ) | ( x57 & n401 ) | ( n398 & n401 ) ;
  assign n403 = ~x57 & n396 ;
  assign n404 = ( ~x57 & n394 ) | ( ~x57 & n403 ) | ( n394 & n403 ) ;
  assign n405 = x56 & n404 ;
  assign n406 = ( x56 & n402 ) | ( x56 & n405 ) | ( n402 & n405 ) ;
  assign n407 = x56 | n400 ;
  assign n408 = ( x56 & ~n398 ) | ( x56 & n407 ) | ( ~n398 & n407 ) ;
  assign n409 = x55 & ~n408 ;
  assign n410 = ( x55 & n406 ) | ( x55 & n409 ) | ( n406 & n409 ) ;
  assign n411 = ~x55 & n404 ;
  assign n412 = ( ~x55 & n402 ) | ( ~x55 & n411 ) | ( n402 & n411 ) ;
  assign n413 = x54 & n412 ;
  assign n414 = ( x54 & n410 ) | ( x54 & n413 ) | ( n410 & n413 ) ;
  assign n415 = x54 | n408 ;
  assign n416 = ( x54 & ~n406 ) | ( x54 & n415 ) | ( ~n406 & n415 ) ;
  assign n417 = x53 & ~n416 ;
  assign n418 = ( x53 & n414 ) | ( x53 & n417 ) | ( n414 & n417 ) ;
  assign n419 = ~x53 & n412 ;
  assign n420 = ( ~x53 & n410 ) | ( ~x53 & n419 ) | ( n410 & n419 ) ;
  assign n421 = x52 & n420 ;
  assign n422 = ( x52 & n418 ) | ( x52 & n421 ) | ( n418 & n421 ) ;
  assign n423 = x52 | n416 ;
  assign n424 = ( x52 & ~n414 ) | ( x52 & n423 ) | ( ~n414 & n423 ) ;
  assign n425 = x51 & ~n424 ;
  assign n426 = ( x51 & n422 ) | ( x51 & n425 ) | ( n422 & n425 ) ;
  assign n427 = ~x51 & n420 ;
  assign n428 = ( ~x51 & n418 ) | ( ~x51 & n427 ) | ( n418 & n427 ) ;
  assign n429 = x50 & n428 ;
  assign n430 = ( x50 & n426 ) | ( x50 & n429 ) | ( n426 & n429 ) ;
  assign n431 = x50 | n424 ;
  assign n432 = ( x50 & ~n422 ) | ( x50 & n431 ) | ( ~n422 & n431 ) ;
  assign n433 = x49 & ~n432 ;
  assign n434 = ( x49 & n430 ) | ( x49 & n433 ) | ( n430 & n433 ) ;
  assign n435 = ~x49 & n428 ;
  assign n436 = ( ~x49 & n426 ) | ( ~x49 & n435 ) | ( n426 & n435 ) ;
  assign n437 = x48 & n436 ;
  assign n438 = ( x48 & n434 ) | ( x48 & n437 ) | ( n434 & n437 ) ;
  assign n439 = x48 | n432 ;
  assign n440 = ( x48 & ~n430 ) | ( x48 & n439 ) | ( ~n430 & n439 ) ;
  assign n441 = x47 & ~n440 ;
  assign n442 = ( x47 & n438 ) | ( x47 & n441 ) | ( n438 & n441 ) ;
  assign n443 = ~x47 & n436 ;
  assign n444 = ( ~x47 & n434 ) | ( ~x47 & n443 ) | ( n434 & n443 ) ;
  assign n445 = x46 & n444 ;
  assign n446 = ( x46 & n442 ) | ( x46 & n445 ) | ( n442 & n445 ) ;
  assign n447 = x46 | n440 ;
  assign n448 = ( x46 & ~n438 ) | ( x46 & n447 ) | ( ~n438 & n447 ) ;
  assign n449 = x45 & ~n448 ;
  assign n450 = ( x45 & n446 ) | ( x45 & n449 ) | ( n446 & n449 ) ;
  assign n451 = ~x45 & n444 ;
  assign n452 = ( ~x45 & n442 ) | ( ~x45 & n451 ) | ( n442 & n451 ) ;
  assign n453 = x44 & n452 ;
  assign n454 = ( x44 & n450 ) | ( x44 & n453 ) | ( n450 & n453 ) ;
  assign n455 = x44 | n448 ;
  assign n456 = ( x44 & ~n446 ) | ( x44 & n455 ) | ( ~n446 & n455 ) ;
  assign n457 = x43 & ~n456 ;
  assign n458 = ( x43 & n454 ) | ( x43 & n457 ) | ( n454 & n457 ) ;
  assign n459 = ~x43 & n452 ;
  assign n460 = ( ~x43 & n450 ) | ( ~x43 & n459 ) | ( n450 & n459 ) ;
  assign n461 = x42 & n460 ;
  assign n462 = ( x42 & n458 ) | ( x42 & n461 ) | ( n458 & n461 ) ;
  assign n463 = x42 | n456 ;
  assign n464 = ( x42 & ~n454 ) | ( x42 & n463 ) | ( ~n454 & n463 ) ;
  assign n465 = x41 & ~n464 ;
  assign n466 = ( x41 & n462 ) | ( x41 & n465 ) | ( n462 & n465 ) ;
  assign n467 = ~x41 & n460 ;
  assign n468 = ( ~x41 & n458 ) | ( ~x41 & n467 ) | ( n458 & n467 ) ;
  assign n469 = x40 & n468 ;
  assign n470 = ( x40 & n466 ) | ( x40 & n469 ) | ( n466 & n469 ) ;
  assign n471 = x40 | n464 ;
  assign n472 = ( x40 & ~n462 ) | ( x40 & n471 ) | ( ~n462 & n471 ) ;
  assign n473 = x39 & ~n472 ;
  assign n474 = ( x39 & n470 ) | ( x39 & n473 ) | ( n470 & n473 ) ;
  assign n475 = ~x39 & n468 ;
  assign n476 = ( ~x39 & n466 ) | ( ~x39 & n475 ) | ( n466 & n475 ) ;
  assign n477 = x38 & n476 ;
  assign n478 = ( x38 & n474 ) | ( x38 & n477 ) | ( n474 & n477 ) ;
  assign n479 = x38 | n472 ;
  assign n480 = ( x38 & ~n470 ) | ( x38 & n479 ) | ( ~n470 & n479 ) ;
  assign n481 = x37 & ~n480 ;
  assign n482 = ( x37 & n478 ) | ( x37 & n481 ) | ( n478 & n481 ) ;
  assign n483 = ~x37 & n476 ;
  assign n484 = ( ~x37 & n474 ) | ( ~x37 & n483 ) | ( n474 & n483 ) ;
  assign n485 = x36 & n484 ;
  assign n486 = ( x36 & n482 ) | ( x36 & n485 ) | ( n482 & n485 ) ;
  assign n487 = x36 | n480 ;
  assign n488 = ( x36 & ~n478 ) | ( x36 & n487 ) | ( ~n478 & n487 ) ;
  assign n489 = x35 & ~n488 ;
  assign n490 = ( x35 & n486 ) | ( x35 & n489 ) | ( n486 & n489 ) ;
  assign n491 = ~x35 & n484 ;
  assign n492 = ( ~x35 & n482 ) | ( ~x35 & n491 ) | ( n482 & n491 ) ;
  assign n493 = x34 & n492 ;
  assign n494 = ( x34 & n490 ) | ( x34 & n493 ) | ( n490 & n493 ) ;
  assign n495 = x34 | n488 ;
  assign n496 = ( x34 & ~n486 ) | ( x34 & n495 ) | ( ~n486 & n495 ) ;
  assign n497 = x33 & ~n496 ;
  assign n498 = ( x33 & n494 ) | ( x33 & n497 ) | ( n494 & n497 ) ;
  assign n499 = ~x33 & n492 ;
  assign n500 = ( ~x33 & n490 ) | ( ~x33 & n499 ) | ( n490 & n499 ) ;
  assign n501 = x32 & n500 ;
  assign n502 = ( x32 & n498 ) | ( x32 & n501 ) | ( n498 & n501 ) ;
  assign n503 = x32 | n496 ;
  assign n504 = ( x32 & ~n494 ) | ( x32 & n503 ) | ( ~n494 & n503 ) ;
  assign n505 = x31 & ~n504 ;
  assign n506 = ( x31 & n502 ) | ( x31 & n505 ) | ( n502 & n505 ) ;
  assign n507 = ~x31 & n500 ;
  assign n508 = ( ~x31 & n498 ) | ( ~x31 & n507 ) | ( n498 & n507 ) ;
  assign n509 = x30 & n508 ;
  assign n510 = ( x30 & n506 ) | ( x30 & n509 ) | ( n506 & n509 ) ;
  assign n511 = x30 | n504 ;
  assign n512 = ( x30 & ~n502 ) | ( x30 & n511 ) | ( ~n502 & n511 ) ;
  assign n513 = x29 & ~n512 ;
  assign n514 = ( x29 & n510 ) | ( x29 & n513 ) | ( n510 & n513 ) ;
  assign n515 = ~x29 & n508 ;
  assign n516 = ( ~x29 & n506 ) | ( ~x29 & n515 ) | ( n506 & n515 ) ;
  assign n517 = x28 & n516 ;
  assign n518 = ( x28 & n514 ) | ( x28 & n517 ) | ( n514 & n517 ) ;
  assign n519 = x28 | n512 ;
  assign n520 = ( x28 & ~n510 ) | ( x28 & n519 ) | ( ~n510 & n519 ) ;
  assign n521 = x27 & ~n520 ;
  assign n522 = ( x27 & n518 ) | ( x27 & n521 ) | ( n518 & n521 ) ;
  assign n523 = ~x27 & n516 ;
  assign n524 = ( ~x27 & n514 ) | ( ~x27 & n523 ) | ( n514 & n523 ) ;
  assign n525 = x26 & n524 ;
  assign n526 = ( x26 & n522 ) | ( x26 & n525 ) | ( n522 & n525 ) ;
  assign n527 = x26 | n520 ;
  assign n528 = ( x26 & ~n518 ) | ( x26 & n527 ) | ( ~n518 & n527 ) ;
  assign n529 = x25 & ~n528 ;
  assign n530 = ( x25 & n526 ) | ( x25 & n529 ) | ( n526 & n529 ) ;
  assign n531 = ~x25 & n524 ;
  assign n532 = ( ~x25 & n522 ) | ( ~x25 & n531 ) | ( n522 & n531 ) ;
  assign n533 = x24 & n532 ;
  assign n534 = ( x24 & n530 ) | ( x24 & n533 ) | ( n530 & n533 ) ;
  assign n535 = x24 | n528 ;
  assign n536 = ( x24 & ~n526 ) | ( x24 & n535 ) | ( ~n526 & n535 ) ;
  assign n537 = x23 & ~n536 ;
  assign n538 = ( x23 & n534 ) | ( x23 & n537 ) | ( n534 & n537 ) ;
  assign n539 = ~x23 & n532 ;
  assign n540 = ( ~x23 & n530 ) | ( ~x23 & n539 ) | ( n530 & n539 ) ;
  assign n541 = x22 & n540 ;
  assign n542 = ( x22 & n538 ) | ( x22 & n541 ) | ( n538 & n541 ) ;
  assign n543 = x22 | n536 ;
  assign n544 = ( x22 & ~n534 ) | ( x22 & n543 ) | ( ~n534 & n543 ) ;
  assign n545 = x21 & ~n544 ;
  assign n546 = ( x21 & n542 ) | ( x21 & n545 ) | ( n542 & n545 ) ;
  assign n547 = ~x21 & n540 ;
  assign n548 = ( ~x21 & n538 ) | ( ~x21 & n547 ) | ( n538 & n547 ) ;
  assign n549 = x20 & n548 ;
  assign n550 = ( x20 & n546 ) | ( x20 & n549 ) | ( n546 & n549 ) ;
  assign n551 = x20 | n544 ;
  assign n552 = ( x20 & ~n542 ) | ( x20 & n551 ) | ( ~n542 & n551 ) ;
  assign n553 = x19 & ~n552 ;
  assign n554 = ( x19 & n550 ) | ( x19 & n553 ) | ( n550 & n553 ) ;
  assign n555 = ~x19 & n548 ;
  assign n556 = ( ~x19 & n546 ) | ( ~x19 & n555 ) | ( n546 & n555 ) ;
  assign n557 = x18 & n556 ;
  assign n558 = ( x18 & n554 ) | ( x18 & n557 ) | ( n554 & n557 ) ;
  assign n559 = x18 | n552 ;
  assign n560 = ( x18 & ~n550 ) | ( x18 & n559 ) | ( ~n550 & n559 ) ;
  assign n561 = x17 & ~n560 ;
  assign n562 = ( x17 & n558 ) | ( x17 & n561 ) | ( n558 & n561 ) ;
  assign n563 = ~x17 & n556 ;
  assign n564 = ( ~x17 & n554 ) | ( ~x17 & n563 ) | ( n554 & n563 ) ;
  assign n565 = x16 & n564 ;
  assign n566 = ( x16 & n562 ) | ( x16 & n565 ) | ( n562 & n565 ) ;
  assign n567 = x16 | n560 ;
  assign n568 = ( x16 & ~n558 ) | ( x16 & n567 ) | ( ~n558 & n567 ) ;
  assign n569 = x15 & ~n568 ;
  assign n570 = ( x15 & n566 ) | ( x15 & n569 ) | ( n566 & n569 ) ;
  assign n571 = ~x15 & n564 ;
  assign n572 = ( ~x15 & n562 ) | ( ~x15 & n571 ) | ( n562 & n571 ) ;
  assign n573 = x14 & n572 ;
  assign n574 = ( x14 & n570 ) | ( x14 & n573 ) | ( n570 & n573 ) ;
  assign n575 = x14 | n568 ;
  assign n576 = ( x14 & ~n566 ) | ( x14 & n575 ) | ( ~n566 & n575 ) ;
  assign n577 = x13 & ~n576 ;
  assign n578 = ( x13 & n574 ) | ( x13 & n577 ) | ( n574 & n577 ) ;
  assign n579 = ~x13 & n572 ;
  assign n580 = ( ~x13 & n570 ) | ( ~x13 & n579 ) | ( n570 & n579 ) ;
  assign n581 = x12 & n580 ;
  assign n582 = ( x12 & n578 ) | ( x12 & n581 ) | ( n578 & n581 ) ;
  assign n583 = x12 | n576 ;
  assign n584 = ( x12 & ~n574 ) | ( x12 & n583 ) | ( ~n574 & n583 ) ;
  assign n585 = x11 & ~n584 ;
  assign n586 = ( x11 & n582 ) | ( x11 & n585 ) | ( n582 & n585 ) ;
  assign n587 = ~x11 & n580 ;
  assign n588 = ( ~x11 & n578 ) | ( ~x11 & n587 ) | ( n578 & n587 ) ;
  assign n589 = x10 & n588 ;
  assign n590 = ( x10 & n586 ) | ( x10 & n589 ) | ( n586 & n589 ) ;
  assign n591 = x10 | n584 ;
  assign n592 = ( x10 & ~n582 ) | ( x10 & n591 ) | ( ~n582 & n591 ) ;
  assign n593 = x9 & ~n592 ;
  assign n594 = ( x9 & n590 ) | ( x9 & n593 ) | ( n590 & n593 ) ;
  assign n595 = ~x9 & n588 ;
  assign n596 = ( ~x9 & n586 ) | ( ~x9 & n595 ) | ( n586 & n595 ) ;
  assign n597 = x8 & n596 ;
  assign n598 = ( x8 & n594 ) | ( x8 & n597 ) | ( n594 & n597 ) ;
  assign n599 = x8 | n592 ;
  assign n600 = ( x8 & ~n590 ) | ( x8 & n599 ) | ( ~n590 & n599 ) ;
  assign n601 = x7 & ~n600 ;
  assign n602 = ( x7 & n598 ) | ( x7 & n601 ) | ( n598 & n601 ) ;
  assign n603 = ~x7 & n596 ;
  assign n604 = ( ~x7 & n594 ) | ( ~x7 & n603 ) | ( n594 & n603 ) ;
  assign n605 = x6 & n604 ;
  assign n606 = ( x6 & n602 ) | ( x6 & n605 ) | ( n602 & n605 ) ;
  assign n607 = x6 | n600 ;
  assign n608 = ( x6 & ~n598 ) | ( x6 & n607 ) | ( ~n598 & n607 ) ;
  assign n609 = x5 & ~n608 ;
  assign n610 = ( x5 & n606 ) | ( x5 & n609 ) | ( n606 & n609 ) ;
  assign n611 = ~x5 & n604 ;
  assign n612 = ( ~x5 & n602 ) | ( ~x5 & n611 ) | ( n602 & n611 ) ;
  assign n613 = x4 & n612 ;
  assign n614 = ( x4 & n610 ) | ( x4 & n613 ) | ( n610 & n613 ) ;
  assign n615 = x4 | n608 ;
  assign n616 = ( x4 & ~n606 ) | ( x4 & n615 ) | ( ~n606 & n615 ) ;
  assign n617 = x3 & ~n616 ;
  assign n618 = ( x3 & n614 ) | ( x3 & n617 ) | ( n614 & n617 ) ;
  assign n619 = x1 & ~x2 ;
  assign n620 = ~x3 & n612 ;
  assign n621 = ( ~x3 & n610 ) | ( ~x3 & n620 ) | ( n610 & n620 ) ;
  assign n622 = n619 | n621 ;
  assign n623 = n618 | n622 ;
  assign n624 = n616 & n619 ;
  assign n625 = ~n614 & n624 ;
  assign n626 = n623 & ~n625 ;
  assign n627 = x2 | x3 ;
  assign n628 = ~x126 & x127 ;
  assign n629 = x126 | n628 ;
  assign n630 = x124 | x125 ;
  assign n631 = x122 | x123 ;
  assign n632 = ~n630 & n631 ;
  assign n633 = n629 | n632 ;
  assign n634 = x120 & n633 ;
  assign n635 = x121 & ~n631 ;
  assign n636 = n629 | n630 ;
  assign n637 = n635 | n636 ;
  assign n638 = ( x120 & ~n629 ) | ( x120 & n637 ) | ( ~n629 & n637 ) ;
  assign n639 = ~n634 & n638 ;
  assign n640 = x118 | x119 ;
  assign n641 = n639 & n640 ;
  assign n642 = n633 | n640 ;
  assign n643 = ~n641 & n642 ;
  assign n644 = x116 | x117 ;
  assign n645 = n643 & n644 ;
  assign n646 = n639 | n644 ;
  assign n647 = ~n645 & n646 ;
  assign n648 = x114 | x115 ;
  assign n649 = n647 & n648 ;
  assign n650 = n643 | n648 ;
  assign n651 = ~n649 & n650 ;
  assign n652 = x112 | x113 ;
  assign n653 = n651 & n652 ;
  assign n654 = n647 | n652 ;
  assign n655 = ~n653 & n654 ;
  assign n656 = x110 | x111 ;
  assign n657 = n655 & n656 ;
  assign n658 = n651 | n656 ;
  assign n659 = ~n657 & n658 ;
  assign n660 = x108 | x109 ;
  assign n661 = n659 & n660 ;
  assign n662 = n655 | n660 ;
  assign n663 = ~n661 & n662 ;
  assign n664 = x106 | x107 ;
  assign n665 = n663 & n664 ;
  assign n666 = n659 | n664 ;
  assign n667 = ~n665 & n666 ;
  assign n668 = x104 | x105 ;
  assign n669 = n667 & n668 ;
  assign n670 = n663 | n668 ;
  assign n671 = ~n669 & n670 ;
  assign n672 = x102 | x103 ;
  assign n673 = n671 & n672 ;
  assign n674 = n667 | n672 ;
  assign n675 = ~n673 & n674 ;
  assign n676 = x100 | x101 ;
  assign n677 = n675 & n676 ;
  assign n678 = n671 | n676 ;
  assign n679 = ~n677 & n678 ;
  assign n680 = x98 | x99 ;
  assign n681 = n679 & n680 ;
  assign n682 = n675 | n680 ;
  assign n683 = ~n681 & n682 ;
  assign n684 = x96 | x97 ;
  assign n685 = n683 & n684 ;
  assign n686 = n679 | n684 ;
  assign n687 = ~n685 & n686 ;
  assign n688 = x94 | x95 ;
  assign n689 = n687 & n688 ;
  assign n690 = n683 | n688 ;
  assign n691 = ~n689 & n690 ;
  assign n692 = x92 | x93 ;
  assign n693 = n691 & n692 ;
  assign n694 = n687 | n692 ;
  assign n695 = ~n693 & n694 ;
  assign n696 = x90 | x91 ;
  assign n697 = n695 & n696 ;
  assign n698 = n691 | n696 ;
  assign n699 = ~n697 & n698 ;
  assign n700 = x88 | x89 ;
  assign n701 = n699 & n700 ;
  assign n702 = n695 | n700 ;
  assign n703 = ~n701 & n702 ;
  assign n704 = x86 | x87 ;
  assign n705 = n703 & n704 ;
  assign n706 = n699 | n704 ;
  assign n707 = ~n705 & n706 ;
  assign n708 = x84 | x85 ;
  assign n709 = n707 & n708 ;
  assign n710 = n703 | n708 ;
  assign n711 = ~n709 & n710 ;
  assign n712 = x82 | x83 ;
  assign n713 = n711 & n712 ;
  assign n714 = n707 | n712 ;
  assign n715 = ~n713 & n714 ;
  assign n716 = x80 | x81 ;
  assign n717 = n715 & n716 ;
  assign n718 = n711 | n716 ;
  assign n719 = ~n717 & n718 ;
  assign n720 = x78 | x79 ;
  assign n721 = n719 & n720 ;
  assign n722 = n715 | n720 ;
  assign n723 = ~n721 & n722 ;
  assign n724 = x76 | x77 ;
  assign n725 = n723 & n724 ;
  assign n726 = n719 | n724 ;
  assign n727 = ~n725 & n726 ;
  assign n728 = x74 | x75 ;
  assign n729 = n727 & n728 ;
  assign n730 = n723 | n728 ;
  assign n731 = ~n729 & n730 ;
  assign n732 = x72 | x73 ;
  assign n733 = n731 & n732 ;
  assign n734 = n727 | n732 ;
  assign n735 = ~n733 & n734 ;
  assign n736 = x70 | x71 ;
  assign n737 = n735 & n736 ;
  assign n738 = n731 | n736 ;
  assign n739 = ~n737 & n738 ;
  assign n740 = x68 | x69 ;
  assign n741 = n739 & n740 ;
  assign n742 = n735 | n740 ;
  assign n743 = ~n741 & n742 ;
  assign n744 = x66 | x67 ;
  assign n745 = n743 & n744 ;
  assign n746 = n739 | n744 ;
  assign n747 = ~n745 & n746 ;
  assign n748 = x64 | x65 ;
  assign n749 = n747 & n748 ;
  assign n750 = n743 | n748 ;
  assign n751 = ~n749 & n750 ;
  assign n752 = x62 | x63 ;
  assign n753 = n751 & n752 ;
  assign n754 = n747 | n752 ;
  assign n755 = ~n753 & n754 ;
  assign n756 = x60 | x61 ;
  assign n757 = n755 & n756 ;
  assign n758 = n751 | n756 ;
  assign n759 = ~n757 & n758 ;
  assign n760 = x58 | x59 ;
  assign n761 = n759 & n760 ;
  assign n762 = n755 | n760 ;
  assign n763 = ~n761 & n762 ;
  assign n764 = x56 | x57 ;
  assign n765 = n763 & n764 ;
  assign n766 = n759 | n764 ;
  assign n767 = ~n765 & n766 ;
  assign n768 = x54 | x55 ;
  assign n769 = n767 & n768 ;
  assign n770 = n763 | n768 ;
  assign n771 = ~n769 & n770 ;
  assign n772 = x52 | x53 ;
  assign n773 = n771 & n772 ;
  assign n774 = n767 | n772 ;
  assign n775 = ~n773 & n774 ;
  assign n776 = x50 | x51 ;
  assign n777 = n775 & n776 ;
  assign n778 = n771 | n776 ;
  assign n779 = ~n777 & n778 ;
  assign n780 = x48 | x49 ;
  assign n781 = n779 & n780 ;
  assign n782 = n775 | n780 ;
  assign n783 = ~n781 & n782 ;
  assign n784 = x46 | x47 ;
  assign n785 = n783 & n784 ;
  assign n786 = n779 | n784 ;
  assign n787 = ~n785 & n786 ;
  assign n788 = x44 | x45 ;
  assign n789 = n787 & n788 ;
  assign n790 = n783 | n788 ;
  assign n791 = ~n789 & n790 ;
  assign n792 = x42 | x43 ;
  assign n793 = n791 & n792 ;
  assign n794 = n787 | n792 ;
  assign n795 = ~n793 & n794 ;
  assign n796 = x40 | x41 ;
  assign n797 = n795 & n796 ;
  assign n798 = n791 | n796 ;
  assign n799 = ~n797 & n798 ;
  assign n800 = x38 | x39 ;
  assign n801 = n799 & n800 ;
  assign n802 = n795 | n800 ;
  assign n803 = ~n801 & n802 ;
  assign n804 = x36 | x37 ;
  assign n805 = n803 & n804 ;
  assign n806 = n799 | n804 ;
  assign n807 = ~n805 & n806 ;
  assign n808 = x34 | x35 ;
  assign n809 = n807 & n808 ;
  assign n810 = n803 | n808 ;
  assign n811 = ~n809 & n810 ;
  assign n812 = x32 | x33 ;
  assign n813 = n811 & n812 ;
  assign n814 = n807 | n812 ;
  assign n815 = ~n813 & n814 ;
  assign n816 = x30 | x31 ;
  assign n817 = n815 & n816 ;
  assign n818 = n811 | n816 ;
  assign n819 = ~n817 & n818 ;
  assign n820 = x28 | x29 ;
  assign n821 = n819 & n820 ;
  assign n822 = n815 | n820 ;
  assign n823 = ~n821 & n822 ;
  assign n824 = x26 | x27 ;
  assign n825 = n823 & n824 ;
  assign n826 = n819 | n824 ;
  assign n827 = ~n825 & n826 ;
  assign n828 = x24 | x25 ;
  assign n829 = n827 & n828 ;
  assign n830 = n823 | n828 ;
  assign n831 = ~n829 & n830 ;
  assign n832 = x22 | x23 ;
  assign n833 = n831 & n832 ;
  assign n834 = n827 | n832 ;
  assign n835 = ~n833 & n834 ;
  assign n836 = x20 | x21 ;
  assign n837 = n835 & n836 ;
  assign n838 = n831 | n836 ;
  assign n839 = ~n837 & n838 ;
  assign n840 = x18 | x19 ;
  assign n841 = n839 & n840 ;
  assign n842 = n835 | n840 ;
  assign n843 = ~n841 & n842 ;
  assign n844 = x16 | x17 ;
  assign n845 = n843 & n844 ;
  assign n846 = n839 | n844 ;
  assign n847 = ~n845 & n846 ;
  assign n848 = x14 | x15 ;
  assign n849 = n847 & n848 ;
  assign n850 = n843 | n848 ;
  assign n851 = ~n849 & n850 ;
  assign n852 = x12 | x13 ;
  assign n853 = n851 & n852 ;
  assign n854 = n847 | n852 ;
  assign n855 = ~n853 & n854 ;
  assign n856 = x10 | x11 ;
  assign n857 = n855 & n856 ;
  assign n858 = n851 | n856 ;
  assign n859 = ~n857 & n858 ;
  assign n860 = x8 | x9 ;
  assign n861 = n859 & n860 ;
  assign n862 = n855 | n860 ;
  assign n863 = ~n861 & n862 ;
  assign n864 = x4 | x5 ;
  assign n865 = n627 & n864 ;
  assign n866 = ( n627 & ~n863 ) | ( n627 & n865 ) | ( ~n863 & n865 ) ;
  assign n867 = x6 | x7 ;
  assign n868 = n863 & n867 ;
  assign n869 = n859 | n867 ;
  assign n870 = ~n868 & n869 ;
  assign n871 = ( n627 & ~n865 ) | ( n627 & n870 ) | ( ~n865 & n870 ) ;
  assign n872 = ( ~n627 & n866 ) | ( ~n627 & n871 ) | ( n866 & n871 ) ;
  assign n873 = x5 | n867 ;
  assign n874 = x4 | n873 ;
  assign n875 = x109 | n656 ;
  assign n876 = x108 | n875 ;
  assign n877 = x113 | x114 ;
  assign n878 = x112 | n877 ;
  assign n879 = x120 | x121 ;
  assign n880 = n631 | n879 ;
  assign n881 = x117 | n640 ;
  assign n882 = x116 | n881 ;
  assign n883 = x115 & ~n882 ;
  assign n884 = n880 | n883 ;
  assign n885 = ( ~n636 & n878 ) | ( ~n636 & n884 ) | ( n878 & n884 ) ;
  assign n886 = ~n880 & n882 ;
  assign n887 = ( n636 & n878 ) | ( n636 & n886 ) | ( n878 & n886 ) ;
  assign n888 = n885 & ~n887 ;
  assign n889 = n876 & ~n888 ;
  assign n890 = n636 | n886 ;
  assign n891 = ~n876 & n890 ;
  assign n892 = n889 | n891 ;
  assign n893 = x105 | n664 ;
  assign n894 = x104 | n893 ;
  assign n895 = ~n892 & n894 ;
  assign n896 = n888 & ~n894 ;
  assign n897 = n895 | n896 ;
  assign n898 = x101 | n672 ;
  assign n899 = x100 | n898 ;
  assign n900 = ~n897 & n899 ;
  assign n901 = n892 & ~n899 ;
  assign n902 = n900 | n901 ;
  assign n903 = x97 | n680 ;
  assign n904 = x96 | n903 ;
  assign n905 = ~n902 & n904 ;
  assign n906 = n897 & ~n904 ;
  assign n907 = n905 | n906 ;
  assign n908 = x93 | n688 ;
  assign n909 = x92 | n908 ;
  assign n910 = ~n907 & n909 ;
  assign n911 = n902 & ~n909 ;
  assign n912 = n910 | n911 ;
  assign n913 = x89 | n696 ;
  assign n914 = x88 | n913 ;
  assign n915 = ~n912 & n914 ;
  assign n916 = n907 & ~n914 ;
  assign n917 = n915 | n916 ;
  assign n918 = x85 | n704 ;
  assign n919 = x84 | n918 ;
  assign n920 = ~n917 & n919 ;
  assign n921 = n912 & ~n919 ;
  assign n922 = n920 | n921 ;
  assign n923 = x81 | n712 ;
  assign n924 = x80 | n923 ;
  assign n925 = ~n922 & n924 ;
  assign n926 = n917 & ~n924 ;
  assign n927 = n925 | n926 ;
  assign n928 = x77 | n720 ;
  assign n929 = x76 | n928 ;
  assign n930 = ~n927 & n929 ;
  assign n931 = n922 & ~n929 ;
  assign n932 = n930 | n931 ;
  assign n933 = x73 | n728 ;
  assign n934 = x72 | n933 ;
  assign n935 = ~n932 & n934 ;
  assign n936 = n927 & ~n934 ;
  assign n937 = n935 | n936 ;
  assign n938 = x69 | n736 ;
  assign n939 = x68 | n938 ;
  assign n940 = ~n937 & n939 ;
  assign n941 = n932 & ~n939 ;
  assign n942 = n940 | n941 ;
  assign n943 = x65 | n744 ;
  assign n944 = x64 | n943 ;
  assign n945 = ~n942 & n944 ;
  assign n946 = n937 & ~n944 ;
  assign n947 = n945 | n946 ;
  assign n948 = x61 | n752 ;
  assign n949 = x60 | n948 ;
  assign n950 = ~n947 & n949 ;
  assign n951 = n942 & ~n949 ;
  assign n952 = n950 | n951 ;
  assign n953 = x57 | n760 ;
  assign n954 = x56 | n953 ;
  assign n955 = ~n952 & n954 ;
  assign n956 = n947 & ~n954 ;
  assign n957 = n955 | n956 ;
  assign n958 = x53 | n768 ;
  assign n959 = x52 | n958 ;
  assign n960 = ~n957 & n959 ;
  assign n961 = n952 & ~n959 ;
  assign n962 = n960 | n961 ;
  assign n963 = x49 | n776 ;
  assign n964 = x48 | n963 ;
  assign n965 = ~n962 & n964 ;
  assign n966 = n957 & ~n964 ;
  assign n967 = n965 | n966 ;
  assign n968 = x45 | n784 ;
  assign n969 = x44 | n968 ;
  assign n970 = ~n967 & n969 ;
  assign n971 = n962 & ~n969 ;
  assign n972 = n970 | n971 ;
  assign n973 = x41 | n792 ;
  assign n974 = x40 | n973 ;
  assign n975 = ~n972 & n974 ;
  assign n976 = n967 & ~n974 ;
  assign n977 = n975 | n976 ;
  assign n978 = x37 | n800 ;
  assign n979 = x36 | n978 ;
  assign n980 = ~n977 & n979 ;
  assign n981 = n972 & ~n979 ;
  assign n982 = n980 | n981 ;
  assign n983 = x33 | n808 ;
  assign n984 = x32 | n983 ;
  assign n985 = ~n982 & n984 ;
  assign n986 = n977 & ~n984 ;
  assign n987 = n985 | n986 ;
  assign n988 = x29 | n816 ;
  assign n989 = x28 | n988 ;
  assign n990 = ~n987 & n989 ;
  assign n991 = n982 & ~n989 ;
  assign n992 = n990 | n991 ;
  assign n993 = x25 | n824 ;
  assign n994 = x24 | n993 ;
  assign n995 = ~n992 & n994 ;
  assign n996 = n987 & ~n994 ;
  assign n997 = n995 | n996 ;
  assign n998 = x21 | n832 ;
  assign n999 = x20 | n998 ;
  assign n1000 = ~n997 & n999 ;
  assign n1001 = n992 & ~n999 ;
  assign n1002 = n1000 | n1001 ;
  assign n1003 = x17 | n840 ;
  assign n1004 = x16 | n1003 ;
  assign n1005 = ~n1002 & n1004 ;
  assign n1006 = n997 & ~n1004 ;
  assign n1007 = n1005 | n1006 ;
  assign n1008 = x9 | n856 ;
  assign n1009 = x8 | n1008 ;
  assign n1010 = n874 & n1009 ;
  assign n1011 = ( n874 & ~n1007 ) | ( n874 & n1010 ) | ( ~n1007 & n1010 ) ;
  assign n1012 = x13 | n848 ;
  assign n1013 = x12 | n1012 ;
  assign n1014 = ~n1007 & n1013 ;
  assign n1015 = n1002 & ~n1013 ;
  assign n1016 = n1014 | n1015 ;
  assign n1017 = ( n874 & ~n1010 ) | ( n874 & n1016 ) | ( ~n1010 & n1016 ) ;
  assign n1018 = ( ~n874 & n1011 ) | ( ~n874 & n1017 ) | ( n1011 & n1017 ) ;
  assign n1019 = x11 | n1013 ;
  assign n1020 = ( x10 & ~n860 ) | ( x10 & n1019 ) | ( ~n860 & n1019 ) ;
  assign n1021 = n860 | n1020 ;
  assign n1022 = n636 | n880 ;
  assign n1023 = x101 | x102 ;
  assign n1024 = ( x100 & ~n680 ) | ( x100 & n1023 ) | ( ~n680 & n1023 ) ;
  assign n1025 = n680 | n1024 ;
  assign n1026 = x97 | n1025 ;
  assign n1027 = x96 | n1026 ;
  assign n1028 = x107 | n876 ;
  assign n1029 = ( x106 & ~n668 ) | ( x106 & n1028 ) | ( ~n668 & n1028 ) ;
  assign n1030 = n668 | n1029 ;
  assign n1031 = x103 & ~n1030 ;
  assign n1032 = ( n648 & ~n652 ) | ( n648 & n882 ) | ( ~n652 & n882 ) ;
  assign n1033 = n652 | n1032 ;
  assign n1034 = n1031 | n1033 ;
  assign n1035 = ( ~n1022 & n1027 ) | ( ~n1022 & n1034 ) | ( n1027 & n1034 ) ;
  assign n1036 = n1030 & ~n1033 ;
  assign n1037 = ( n1022 & n1027 ) | ( n1022 & n1036 ) | ( n1027 & n1036 ) ;
  assign n1038 = n1035 & ~n1037 ;
  assign n1039 = x91 | n909 ;
  assign n1040 = ( x90 & ~n700 ) | ( x90 & n1039 ) | ( ~n700 & n1039 ) ;
  assign n1041 = n700 | n1040 ;
  assign n1042 = ~n1038 & n1041 ;
  assign n1043 = n1022 | n1036 ;
  assign n1044 = ~n1041 & n1043 ;
  assign n1045 = n1042 | n1044 ;
  assign n1046 = x83 | n919 ;
  assign n1047 = ( x82 & ~n716 ) | ( x82 & n1046 ) | ( ~n716 & n1046 ) ;
  assign n1048 = n716 | n1047 ;
  assign n1049 = ~n1045 & n1048 ;
  assign n1050 = n1038 & ~n1048 ;
  assign n1051 = n1049 | n1050 ;
  assign n1052 = x75 | n929 ;
  assign n1053 = ( x74 & ~n732 ) | ( x74 & n1052 ) | ( ~n732 & n1052 ) ;
  assign n1054 = n732 | n1053 ;
  assign n1055 = ~n1051 & n1054 ;
  assign n1056 = n1045 & ~n1054 ;
  assign n1057 = n1055 | n1056 ;
  assign n1058 = x67 | n939 ;
  assign n1059 = ( x66 & ~n748 ) | ( x66 & n1058 ) | ( ~n748 & n1058 ) ;
  assign n1060 = n748 | n1059 ;
  assign n1061 = ~n1057 & n1060 ;
  assign n1062 = n1051 & ~n1060 ;
  assign n1063 = n1061 | n1062 ;
  assign n1064 = x59 | n949 ;
  assign n1065 = ( x58 & ~n764 ) | ( x58 & n1064 ) | ( ~n764 & n1064 ) ;
  assign n1066 = n764 | n1065 ;
  assign n1067 = ~n1063 & n1066 ;
  assign n1068 = n1057 & ~n1066 ;
  assign n1069 = n1067 | n1068 ;
  assign n1070 = x51 | n959 ;
  assign n1071 = ( x50 & ~n780 ) | ( x50 & n1070 ) | ( ~n780 & n1070 ) ;
  assign n1072 = n780 | n1071 ;
  assign n1073 = ~n1069 & n1072 ;
  assign n1074 = n1063 & ~n1072 ;
  assign n1075 = n1073 | n1074 ;
  assign n1076 = x43 | n969 ;
  assign n1077 = ( x42 & ~n796 ) | ( x42 & n1076 ) | ( ~n796 & n1076 ) ;
  assign n1078 = n796 | n1077 ;
  assign n1079 = ~n1075 & n1078 ;
  assign n1080 = n1069 & ~n1078 ;
  assign n1081 = n1079 | n1080 ;
  assign n1082 = x35 | n979 ;
  assign n1083 = ( x34 & ~n812 ) | ( x34 & n1082 ) | ( ~n812 & n1082 ) ;
  assign n1084 = n812 | n1083 ;
  assign n1085 = ~n1081 & n1084 ;
  assign n1086 = n1075 & ~n1084 ;
  assign n1087 = n1085 | n1086 ;
  assign n1088 = x19 | n999 ;
  assign n1089 = ( x18 & ~n844 ) | ( x18 & n1088 ) | ( ~n844 & n1088 ) ;
  assign n1090 = n844 | n1089 ;
  assign n1091 = n1021 & n1090 ;
  assign n1092 = ( n1021 & ~n1087 ) | ( n1021 & n1091 ) | ( ~n1087 & n1091 ) ;
  assign n1093 = x27 | n989 ;
  assign n1094 = ( x26 & ~n828 ) | ( x26 & n1093 ) | ( ~n828 & n1093 ) ;
  assign n1095 = n828 | n1094 ;
  assign n1096 = ~n1087 & n1095 ;
  assign n1097 = n1081 & ~n1095 ;
  assign n1098 = n1096 | n1097 ;
  assign n1099 = ( n1021 & ~n1091 ) | ( n1021 & n1098 ) | ( ~n1091 & n1098 ) ;
  assign n1100 = ( ~n1021 & n1092 ) | ( ~n1021 & n1099 ) | ( n1092 & n1099 ) ;
  assign n1101 = x23 | n1095 ;
  assign n1102 = ( x22 & ~n836 ) | ( x22 & n1101 ) | ( ~n836 & n1101 ) ;
  assign n1103 = n836 | n1102 ;
  assign n1104 = x19 | n1103 ;
  assign n1105 = ( x18 & ~n844 ) | ( x18 & n1104 ) | ( ~n844 & n1104 ) ;
  assign n1106 = n844 | n1105 ;
  assign n1107 = n1022 | n1033 ;
  assign n1108 = x99 | n899 ;
  assign n1109 = ( x98 & ~n684 ) | ( x98 & n1030 ) | ( ~n684 & n1030 ) ;
  assign n1110 = n684 | n1109 ;
  assign n1111 = n1108 | n1110 ;
  assign n1112 = x87 | n1041 ;
  assign n1113 = ( x86 & ~n708 ) | ( x86 & n1112 ) | ( ~n708 & n1112 ) ;
  assign n1114 = n708 | n1113 ;
  assign n1115 = x83 | n1114 ;
  assign n1116 = ( x82 & ~n716 ) | ( x82 & n1115 ) | ( ~n716 & n1115 ) ;
  assign n1117 = n716 | n1116 ;
  assign n1118 = x79 & ~n1117 ;
  assign n1119 = n1111 | n1118 ;
  assign n1120 = x77 | x78 ;
  assign n1121 = ( x76 & ~n728 ) | ( x76 & n1120 ) | ( ~n728 & n1120 ) ;
  assign n1122 = n728 | n1121 ;
  assign n1123 = x73 | n1122 ;
  assign n1124 = ( x72 & ~n736 ) | ( x72 & n1123 ) | ( ~n736 & n1123 ) ;
  assign n1125 = n736 | n1124 ;
  assign n1126 = x69 | n1125 ;
  assign n1127 = x68 | n1126 ;
  assign n1128 = x67 | n1127 ;
  assign n1129 = ( x66 & ~n748 ) | ( x66 & n1128 ) | ( ~n748 & n1128 ) ;
  assign n1130 = n748 | n1129 ;
  assign n1131 = ( ~n1107 & n1119 ) | ( ~n1107 & n1130 ) | ( n1119 & n1130 ) ;
  assign n1132 = ~n1111 & n1117 ;
  assign n1133 = ( n1107 & n1130 ) | ( n1107 & n1132 ) | ( n1130 & n1132 ) ;
  assign n1134 = n1131 & ~n1133 ;
  assign n1135 = x39 | n1078 ;
  assign n1136 = ( x38 & ~n804 ) | ( x38 & n1135 ) | ( ~n804 & n1135 ) ;
  assign n1137 = n804 | n1136 ;
  assign n1138 = x35 | n1137 ;
  assign n1139 = ( x34 & ~n812 ) | ( x34 & n1138 ) | ( ~n812 & n1138 ) ;
  assign n1140 = n812 | n1139 ;
  assign n1141 = n1106 & n1140 ;
  assign n1142 = ( n1106 & ~n1134 ) | ( n1106 & n1141 ) | ( ~n1134 & n1141 ) ;
  assign n1143 = x55 | n1066 ;
  assign n1144 = ( x54 & ~n772 ) | ( x54 & n1143 ) | ( ~n772 & n1143 ) ;
  assign n1145 = n772 | n1144 ;
  assign n1146 = x51 | n1145 ;
  assign n1147 = ( x50 & ~n780 ) | ( x50 & n1146 ) | ( ~n780 & n1146 ) ;
  assign n1148 = n780 | n1147 ;
  assign n1149 = ~n1134 & n1148 ;
  assign n1150 = n1107 | n1132 ;
  assign n1151 = ~n1148 & n1150 ;
  assign n1152 = n1149 | n1151 ;
  assign n1153 = ( n1106 & ~n1141 ) | ( n1106 & n1152 ) | ( ~n1141 & n1152 ) ;
  assign n1154 = ( ~n1106 & n1142 ) | ( ~n1106 & n1153 ) | ( n1142 & n1153 ) ;
  assign n1155 = n1107 | n1111 ;
  assign n1156 = x71 | n1054 ;
  assign n1157 = ( x70 & ~n740 ) | ( x70 & n1117 ) | ( ~n740 & n1117 ) ;
  assign n1158 = n740 | n1157 ;
  assign n1159 = x67 | n1158 ;
  assign n1160 = x66 | n1159 ;
  assign n1161 = ( ~n748 & n1156 ) | ( ~n748 & n1160 ) | ( n1156 & n1160 ) ;
  assign n1162 = n748 | n1161 ;
  assign n1163 = x47 | n1148 ;
  assign n1164 = ( x46 & ~n788 ) | ( x46 & n1163 ) | ( ~n788 & n1163 ) ;
  assign n1165 = n788 | n1164 ;
  assign n1166 = x43 | n1165 ;
  assign n1167 = ( x42 & ~n796 ) | ( x42 & n1166 ) | ( ~n796 & n1166 ) ;
  assign n1168 = n796 | n1167 ;
  assign n1169 = x39 | n1168 ;
  assign n1170 = ( x38 & ~n804 ) | ( x38 & n1169 ) | ( ~n804 & n1169 ) ;
  assign n1171 = n804 | n1170 ;
  assign n1172 = x35 | n1171 ;
  assign n1173 = ( x34 & ~n812 ) | ( x34 & n1172 ) | ( ~n812 & n1172 ) ;
  assign n1174 = n812 | n1173 ;
  assign n1175 = ~n1162 & n1174 ;
  assign n1176 = n1155 | n1175 ;
  assign n1177 = n1155 | n1162 ;
  assign n1178 = n1106 | n1174 ;
  assign n1179 = n874 | n1178 ;
  assign n1180 = x1 | n1179 ;
  assign n1181 = x0 | n1177 ;
  assign n1182 = ( ~n627 & n1021 ) | ( ~n627 & n1181 ) | ( n1021 & n1181 ) ;
  assign n1183 = n627 | n1182 ;
  assign n1184 = n1180 | n1183 ;
  assign y0 = n626 ;
  assign y1 = n872 ;
  assign y2 = n1018 ;
  assign y3 = n1100 ;
  assign y4 = n1154 ;
  assign y5 = n1176 ;
  assign y6 = n1177 ;
  assign y7 = n1184 ;
endmodule
