module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 ;
  assign n136 = x77 & x128 ;
  assign n137 = x78 & ~x128 ;
  assign n138 = n136 | n137 ;
  assign n139 = x129 & n138 ;
  assign n140 = x80 & ~x128 ;
  assign n141 = x79 & x128 ;
  assign n142 = n140 | n141 ;
  assign n143 = ~x129 & n142 ;
  assign n144 = n139 | n143 ;
  assign n145 = x130 | x131 ;
  assign n146 = n144 & ~n145 ;
  assign n147 = x73 & x128 ;
  assign n148 = x74 & ~x128 ;
  assign n149 = n147 | n148 ;
  assign n150 = x129 & n149 ;
  assign n151 = x76 & ~x128 ;
  assign n152 = x75 & x128 ;
  assign n153 = n151 | n152 ;
  assign n154 = ~x129 & n153 ;
  assign n155 = n150 | n154 ;
  assign n156 = x130 & ~x131 ;
  assign n157 = n155 & n156 ;
  assign n158 = n146 | n157 ;
  assign n159 = x65 & x128 ;
  assign n160 = x66 & ~x128 ;
  assign n161 = n159 | n160 ;
  assign n162 = x129 & n161 ;
  assign n163 = x68 & ~x128 ;
  assign n164 = x67 & x128 ;
  assign n165 = n163 | n164 ;
  assign n166 = ~x129 & n165 ;
  assign n167 = n162 | n166 ;
  assign n168 = x130 & x131 ;
  assign n169 = n167 & n168 ;
  assign n170 = x69 & x128 ;
  assign n171 = x70 & ~x128 ;
  assign n172 = n170 | n171 ;
  assign n173 = x129 & n172 ;
  assign n174 = x72 & ~x128 ;
  assign n175 = x71 & x128 ;
  assign n176 = n174 | n175 ;
  assign n177 = ~x129 & n176 ;
  assign n178 = n173 | n177 ;
  assign n179 = ~x130 & x131 ;
  assign n180 = n178 & n179 ;
  assign n181 = n169 | n180 ;
  assign n182 = n158 | n181 ;
  assign n183 = x132 & x133 ;
  assign n184 = n182 & n183 ;
  assign n185 = x93 & x128 ;
  assign n186 = x94 & ~x128 ;
  assign n187 = n185 | n186 ;
  assign n188 = x129 & n187 ;
  assign n189 = x96 & ~x128 ;
  assign n190 = x95 & x128 ;
  assign n191 = n189 | n190 ;
  assign n192 = ~x129 & n191 ;
  assign n193 = n188 | n192 ;
  assign n194 = ~n145 & n193 ;
  assign n195 = x89 & x128 ;
  assign n196 = x90 & ~x128 ;
  assign n197 = n195 | n196 ;
  assign n198 = x129 & n197 ;
  assign n199 = x92 & ~x128 ;
  assign n200 = x91 & x128 ;
  assign n201 = n199 | n200 ;
  assign n202 = ~x129 & n201 ;
  assign n203 = n198 | n202 ;
  assign n204 = n156 & n203 ;
  assign n205 = n194 | n204 ;
  assign n206 = x81 & x128 ;
  assign n207 = x82 & ~x128 ;
  assign n208 = n206 | n207 ;
  assign n209 = x129 & n208 ;
  assign n210 = x84 & ~x128 ;
  assign n211 = x83 & x128 ;
  assign n212 = n210 | n211 ;
  assign n213 = ~x129 & n212 ;
  assign n214 = n209 | n213 ;
  assign n215 = n168 & n214 ;
  assign n216 = x85 & x128 ;
  assign n217 = x86 & ~x128 ;
  assign n218 = n216 | n217 ;
  assign n219 = x129 & n218 ;
  assign n220 = x88 & ~x128 ;
  assign n221 = x87 & x128 ;
  assign n222 = n220 | n221 ;
  assign n223 = ~x129 & n222 ;
  assign n224 = n219 | n223 ;
  assign n225 = n179 & n224 ;
  assign n226 = n215 | n225 ;
  assign n227 = n205 | n226 ;
  assign n228 = ~x132 & x133 ;
  assign n229 = n227 & n228 ;
  assign n230 = n184 | n229 ;
  assign n231 = x125 & x128 ;
  assign n232 = x126 & ~x128 ;
  assign n233 = n231 | n232 ;
  assign n234 = x129 & n233 ;
  assign n235 = x0 & ~x128 ;
  assign n236 = x127 & x128 ;
  assign n237 = n235 | n236 ;
  assign n238 = ~x129 & n237 ;
  assign n239 = n234 | n238 ;
  assign n240 = ~n145 & n239 ;
  assign n241 = x121 & x128 ;
  assign n242 = x122 & ~x128 ;
  assign n243 = n241 | n242 ;
  assign n244 = x129 & n243 ;
  assign n245 = x124 & ~x128 ;
  assign n246 = x123 & x128 ;
  assign n247 = n245 | n246 ;
  assign n248 = ~x129 & n247 ;
  assign n249 = n244 | n248 ;
  assign n250 = n156 & n249 ;
  assign n251 = n240 | n250 ;
  assign n252 = x113 & x128 ;
  assign n253 = x114 & ~x128 ;
  assign n254 = n252 | n253 ;
  assign n255 = x129 & n254 ;
  assign n256 = x116 & ~x128 ;
  assign n257 = x115 & x128 ;
  assign n258 = n256 | n257 ;
  assign n259 = ~x129 & n258 ;
  assign n260 = n255 | n259 ;
  assign n261 = n168 & n260 ;
  assign n262 = x117 & x128 ;
  assign n263 = x118 & ~x128 ;
  assign n264 = n262 | n263 ;
  assign n265 = x129 & n264 ;
  assign n266 = x120 & ~x128 ;
  assign n267 = x119 & x128 ;
  assign n268 = n266 | n267 ;
  assign n269 = ~x129 & n268 ;
  assign n270 = n265 | n269 ;
  assign n271 = n179 & n270 ;
  assign n272 = n261 | n271 ;
  assign n273 = n251 | n272 ;
  assign n274 = x132 | x133 ;
  assign n275 = n273 & ~n274 ;
  assign n276 = x109 & x128 ;
  assign n277 = x110 & ~x128 ;
  assign n278 = n276 | n277 ;
  assign n279 = x129 & n278 ;
  assign n280 = x112 & ~x128 ;
  assign n281 = x111 & x128 ;
  assign n282 = n280 | n281 ;
  assign n283 = ~x129 & n282 ;
  assign n284 = n279 | n283 ;
  assign n285 = ~n145 & n284 ;
  assign n286 = x105 & x128 ;
  assign n287 = x106 & ~x128 ;
  assign n288 = n286 | n287 ;
  assign n289 = x129 & n288 ;
  assign n290 = x108 & ~x128 ;
  assign n291 = x107 & x128 ;
  assign n292 = n290 | n291 ;
  assign n293 = ~x129 & n292 ;
  assign n294 = n289 | n293 ;
  assign n295 = n156 & n294 ;
  assign n296 = n285 | n295 ;
  assign n297 = x97 & x128 ;
  assign n298 = x98 & ~x128 ;
  assign n299 = n297 | n298 ;
  assign n300 = x129 & n299 ;
  assign n301 = x100 & ~x128 ;
  assign n302 = x99 & x128 ;
  assign n303 = n301 | n302 ;
  assign n304 = ~x129 & n303 ;
  assign n305 = n300 | n304 ;
  assign n306 = n168 & n305 ;
  assign n307 = x101 & x128 ;
  assign n308 = x102 & ~x128 ;
  assign n309 = n307 | n308 ;
  assign n310 = x129 & n309 ;
  assign n311 = x104 & ~x128 ;
  assign n312 = x103 & x128 ;
  assign n313 = n311 | n312 ;
  assign n314 = ~x129 & n313 ;
  assign n315 = n310 | n314 ;
  assign n316 = n179 & n315 ;
  assign n317 = n306 | n316 ;
  assign n318 = n296 | n317 ;
  assign n319 = x132 & ~x133 ;
  assign n320 = n318 & n319 ;
  assign n321 = n275 | n320 ;
  assign n322 = n230 | n321 ;
  assign n323 = ~x134 & n322 ;
  assign n324 = x13 & x128 ;
  assign n325 = x14 & ~x128 ;
  assign n326 = n324 | n325 ;
  assign n327 = x129 & n326 ;
  assign n328 = x16 & ~x128 ;
  assign n329 = x15 & x128 ;
  assign n330 = n328 | n329 ;
  assign n331 = ~x129 & n330 ;
  assign n332 = n327 | n331 ;
  assign n333 = ~n145 & n332 ;
  assign n334 = x9 & x128 ;
  assign n335 = x10 & ~x128 ;
  assign n336 = n334 | n335 ;
  assign n337 = x129 & n336 ;
  assign n338 = x12 & ~x128 ;
  assign n339 = x11 & x128 ;
  assign n340 = n338 | n339 ;
  assign n341 = ~x129 & n340 ;
  assign n342 = n337 | n341 ;
  assign n343 = n156 & n342 ;
  assign n344 = n333 | n343 ;
  assign n345 = x1 & x128 ;
  assign n346 = x2 & ~x128 ;
  assign n347 = n345 | n346 ;
  assign n348 = x129 & n347 ;
  assign n349 = x4 & ~x128 ;
  assign n350 = x3 & x128 ;
  assign n351 = n349 | n350 ;
  assign n352 = ~x129 & n351 ;
  assign n353 = n348 | n352 ;
  assign n354 = n168 & n353 ;
  assign n355 = x5 & x128 ;
  assign n356 = x6 & ~x128 ;
  assign n357 = n355 | n356 ;
  assign n358 = x129 & n357 ;
  assign n359 = x8 & ~x128 ;
  assign n360 = x7 & x128 ;
  assign n361 = n359 | n360 ;
  assign n362 = ~x129 & n361 ;
  assign n363 = n358 | n362 ;
  assign n364 = n179 & n363 ;
  assign n365 = n354 | n364 ;
  assign n366 = n344 | n365 ;
  assign n367 = n183 & n366 ;
  assign n368 = x29 & x128 ;
  assign n369 = x30 & ~x128 ;
  assign n370 = n368 | n369 ;
  assign n371 = x129 & n370 ;
  assign n372 = x32 & ~x128 ;
  assign n373 = x31 & x128 ;
  assign n374 = n372 | n373 ;
  assign n375 = ~x129 & n374 ;
  assign n376 = n371 | n375 ;
  assign n377 = ~n145 & n376 ;
  assign n378 = x25 & x128 ;
  assign n379 = x26 & ~x128 ;
  assign n380 = n378 | n379 ;
  assign n381 = x129 & n380 ;
  assign n382 = x28 & ~x128 ;
  assign n383 = x27 & x128 ;
  assign n384 = n382 | n383 ;
  assign n385 = ~x129 & n384 ;
  assign n386 = n381 | n385 ;
  assign n387 = n156 & n386 ;
  assign n388 = n377 | n387 ;
  assign n389 = x17 & x128 ;
  assign n390 = x18 & ~x128 ;
  assign n391 = n389 | n390 ;
  assign n392 = x129 & n391 ;
  assign n393 = x20 & ~x128 ;
  assign n394 = x19 & x128 ;
  assign n395 = n393 | n394 ;
  assign n396 = ~x129 & n395 ;
  assign n397 = n392 | n396 ;
  assign n398 = n168 & n397 ;
  assign n399 = x21 & x128 ;
  assign n400 = x22 & ~x128 ;
  assign n401 = n399 | n400 ;
  assign n402 = x129 & n401 ;
  assign n403 = x24 & ~x128 ;
  assign n404 = x23 & x128 ;
  assign n405 = n403 | n404 ;
  assign n406 = ~x129 & n405 ;
  assign n407 = n402 | n406 ;
  assign n408 = n179 & n407 ;
  assign n409 = n398 | n408 ;
  assign n410 = n388 | n409 ;
  assign n411 = n228 & n410 ;
  assign n412 = n367 | n411 ;
  assign n413 = x61 & x128 ;
  assign n414 = x62 & ~x128 ;
  assign n415 = n413 | n414 ;
  assign n416 = x129 & n415 ;
  assign n417 = x64 & ~x128 ;
  assign n418 = x63 & x128 ;
  assign n419 = n417 | n418 ;
  assign n420 = ~x129 & n419 ;
  assign n421 = n416 | n420 ;
  assign n422 = ~n145 & n421 ;
  assign n423 = x57 & x128 ;
  assign n424 = x58 & ~x128 ;
  assign n425 = n423 | n424 ;
  assign n426 = x129 & n425 ;
  assign n427 = x60 & ~x128 ;
  assign n428 = x59 & x128 ;
  assign n429 = n427 | n428 ;
  assign n430 = ~x129 & n429 ;
  assign n431 = n426 | n430 ;
  assign n432 = n156 & n431 ;
  assign n433 = n422 | n432 ;
  assign n434 = x49 & x128 ;
  assign n435 = x50 & ~x128 ;
  assign n436 = n434 | n435 ;
  assign n437 = x129 & n436 ;
  assign n438 = x52 & ~x128 ;
  assign n439 = x51 & x128 ;
  assign n440 = n438 | n439 ;
  assign n441 = ~x129 & n440 ;
  assign n442 = n437 | n441 ;
  assign n443 = n168 & n442 ;
  assign n444 = x53 & x128 ;
  assign n445 = x54 & ~x128 ;
  assign n446 = n444 | n445 ;
  assign n447 = x129 & n446 ;
  assign n448 = x56 & ~x128 ;
  assign n449 = x55 & x128 ;
  assign n450 = n448 | n449 ;
  assign n451 = ~x129 & n450 ;
  assign n452 = n447 | n451 ;
  assign n453 = n179 & n452 ;
  assign n454 = n443 | n453 ;
  assign n455 = n433 | n454 ;
  assign n456 = ~n274 & n455 ;
  assign n457 = x33 & x128 ;
  assign n458 = x34 & ~x128 ;
  assign n459 = n457 | n458 ;
  assign n460 = x129 & n459 ;
  assign n461 = x36 & ~x128 ;
  assign n462 = x35 & x128 ;
  assign n463 = n461 | n462 ;
  assign n464 = ~x129 & n463 ;
  assign n465 = n460 | n464 ;
  assign n466 = n168 & n465 ;
  assign n467 = x40 & ~x128 ;
  assign n468 = ~x129 & n467 ;
  assign n469 = x37 & x128 ;
  assign n470 = x129 & n469 ;
  assign n471 = n468 | n470 ;
  assign n472 = x38 & ~x128 ;
  assign n473 = ( x129 & n471 ) | ( x129 & n472 ) | ( n471 & n472 ) ;
  assign n474 = x39 & x128 ;
  assign n475 = ( ~x129 & n471 ) | ( ~x129 & n474 ) | ( n471 & n474 ) ;
  assign n476 = n473 | n475 ;
  assign n477 = n179 & n476 ;
  assign n478 = n466 | n477 ;
  assign n479 = x45 & x128 ;
  assign n480 = x46 & ~x128 ;
  assign n481 = n479 | n480 ;
  assign n482 = x129 & n481 ;
  assign n483 = x48 & ~x128 ;
  assign n484 = x47 & x128 ;
  assign n485 = n483 | n484 ;
  assign n486 = ~x129 & n485 ;
  assign n487 = n482 | n486 ;
  assign n488 = ~n145 & n487 ;
  assign n489 = x41 & x128 ;
  assign n490 = x42 & ~x128 ;
  assign n491 = n489 | n490 ;
  assign n492 = x129 & n491 ;
  assign n493 = x44 & ~x128 ;
  assign n494 = x43 & x128 ;
  assign n495 = n493 | n494 ;
  assign n496 = ~x129 & n495 ;
  assign n497 = n492 | n496 ;
  assign n498 = n156 & n497 ;
  assign n499 = n488 | n498 ;
  assign n500 = n319 & n499 ;
  assign n501 = ( n319 & n478 ) | ( n319 & n500 ) | ( n478 & n500 ) ;
  assign n502 = n456 | n501 ;
  assign n503 = n412 | n502 ;
  assign n504 = x134 & n503 ;
  assign n505 = n323 | n504 ;
  assign n506 = x81 & ~x128 ;
  assign n507 = ~x129 & n506 ;
  assign n508 = x78 & x128 ;
  assign n509 = x129 & n508 ;
  assign n510 = n507 | n509 ;
  assign n511 = x79 & ~x128 ;
  assign n512 = ( x129 & n510 ) | ( x129 & n511 ) | ( n510 & n511 ) ;
  assign n513 = x80 & x128 ;
  assign n514 = ( ~x129 & n510 ) | ( ~x129 & n513 ) | ( n510 & n513 ) ;
  assign n515 = n512 | n514 ;
  assign n516 = ~n145 & n515 ;
  assign n517 = x77 & ~x128 ;
  assign n518 = ~x129 & n517 ;
  assign n519 = x74 & x128 ;
  assign n520 = x129 & n519 ;
  assign n521 = n518 | n520 ;
  assign n522 = x75 & ~x128 ;
  assign n523 = ( x129 & n521 ) | ( x129 & n522 ) | ( n521 & n522 ) ;
  assign n524 = x76 & x128 ;
  assign n525 = ( ~x129 & n521 ) | ( ~x129 & n524 ) | ( n521 & n524 ) ;
  assign n526 = n523 | n525 ;
  assign n527 = n156 & n526 ;
  assign n528 = n516 | n527 ;
  assign n529 = x69 & ~x128 ;
  assign n530 = ~x129 & n529 ;
  assign n531 = x66 & x128 ;
  assign n532 = x129 & n531 ;
  assign n533 = n530 | n532 ;
  assign n534 = x67 & ~x128 ;
  assign n535 = ( x129 & n533 ) | ( x129 & n534 ) | ( n533 & n534 ) ;
  assign n536 = x68 & x128 ;
  assign n537 = ( ~x129 & n533 ) | ( ~x129 & n536 ) | ( n533 & n536 ) ;
  assign n538 = n535 | n537 ;
  assign n539 = n168 & n538 ;
  assign n540 = x73 & ~x128 ;
  assign n541 = ~x129 & n540 ;
  assign n542 = x70 & x128 ;
  assign n543 = x129 & n542 ;
  assign n544 = n541 | n543 ;
  assign n545 = x71 & ~x128 ;
  assign n546 = ( x129 & n544 ) | ( x129 & n545 ) | ( n544 & n545 ) ;
  assign n547 = x72 & x128 ;
  assign n548 = ( ~x129 & n544 ) | ( ~x129 & n547 ) | ( n544 & n547 ) ;
  assign n549 = n546 | n548 ;
  assign n550 = n179 & n549 ;
  assign n551 = n539 | n550 ;
  assign n552 = n528 | n551 ;
  assign n553 = n183 & n552 ;
  assign n554 = x97 & ~x128 ;
  assign n555 = ~x129 & n554 ;
  assign n556 = x94 & x128 ;
  assign n557 = x129 & n556 ;
  assign n558 = n555 | n557 ;
  assign n559 = x95 & ~x128 ;
  assign n560 = ( x129 & n558 ) | ( x129 & n559 ) | ( n558 & n559 ) ;
  assign n561 = x96 & x128 ;
  assign n562 = ( ~x129 & n558 ) | ( ~x129 & n561 ) | ( n558 & n561 ) ;
  assign n563 = n560 | n562 ;
  assign n564 = ~n145 & n563 ;
  assign n565 = x93 & ~x128 ;
  assign n566 = ~x129 & n565 ;
  assign n567 = x90 & x128 ;
  assign n568 = x129 & n567 ;
  assign n569 = n566 | n568 ;
  assign n570 = x91 & ~x128 ;
  assign n571 = ( x129 & n569 ) | ( x129 & n570 ) | ( n569 & n570 ) ;
  assign n572 = x92 & x128 ;
  assign n573 = ( ~x129 & n569 ) | ( ~x129 & n572 ) | ( n569 & n572 ) ;
  assign n574 = n571 | n573 ;
  assign n575 = n156 & n574 ;
  assign n576 = n564 | n575 ;
  assign n577 = x85 & ~x128 ;
  assign n578 = ~x129 & n577 ;
  assign n579 = x82 & x128 ;
  assign n580 = x129 & n579 ;
  assign n581 = n578 | n580 ;
  assign n582 = x83 & ~x128 ;
  assign n583 = ( x129 & n581 ) | ( x129 & n582 ) | ( n581 & n582 ) ;
  assign n584 = x84 & x128 ;
  assign n585 = ( ~x129 & n581 ) | ( ~x129 & n584 ) | ( n581 & n584 ) ;
  assign n586 = n583 | n585 ;
  assign n587 = n168 & n586 ;
  assign n588 = x89 & ~x128 ;
  assign n589 = ~x129 & n588 ;
  assign n590 = x86 & x128 ;
  assign n591 = x129 & n590 ;
  assign n592 = n589 | n591 ;
  assign n593 = x87 & ~x128 ;
  assign n594 = ( x129 & n592 ) | ( x129 & n593 ) | ( n592 & n593 ) ;
  assign n595 = x88 & x128 ;
  assign n596 = ( ~x129 & n592 ) | ( ~x129 & n595 ) | ( n592 & n595 ) ;
  assign n597 = n594 | n596 ;
  assign n598 = n179 & n597 ;
  assign n599 = n587 | n598 ;
  assign n600 = n576 | n599 ;
  assign n601 = n228 & n600 ;
  assign n602 = n553 | n601 ;
  assign n603 = x1 & ~x128 ;
  assign n604 = ~x129 & n603 ;
  assign n605 = x126 & x128 ;
  assign n606 = x129 & n605 ;
  assign n607 = n604 | n606 ;
  assign n608 = x127 & ~x128 ;
  assign n609 = ( x129 & n607 ) | ( x129 & n608 ) | ( n607 & n608 ) ;
  assign n610 = x0 & x128 ;
  assign n611 = ( ~x129 & n607 ) | ( ~x129 & n610 ) | ( n607 & n610 ) ;
  assign n612 = n609 | n611 ;
  assign n613 = ~n145 & n612 ;
  assign n614 = x125 & ~x128 ;
  assign n615 = ~x129 & n614 ;
  assign n616 = x122 & x128 ;
  assign n617 = x129 & n616 ;
  assign n618 = n615 | n617 ;
  assign n619 = x123 & ~x128 ;
  assign n620 = ( x129 & n618 ) | ( x129 & n619 ) | ( n618 & n619 ) ;
  assign n621 = x124 & x128 ;
  assign n622 = ( ~x129 & n618 ) | ( ~x129 & n621 ) | ( n618 & n621 ) ;
  assign n623 = n620 | n622 ;
  assign n624 = n156 & n623 ;
  assign n625 = n613 | n624 ;
  assign n626 = x117 & ~x128 ;
  assign n627 = ~x129 & n626 ;
  assign n628 = x114 & x128 ;
  assign n629 = x129 & n628 ;
  assign n630 = n627 | n629 ;
  assign n631 = x115 & ~x128 ;
  assign n632 = ( x129 & n630 ) | ( x129 & n631 ) | ( n630 & n631 ) ;
  assign n633 = x116 & x128 ;
  assign n634 = ( ~x129 & n630 ) | ( ~x129 & n633 ) | ( n630 & n633 ) ;
  assign n635 = n632 | n634 ;
  assign n636 = n168 & n635 ;
  assign n637 = x121 & ~x128 ;
  assign n638 = ~x129 & n637 ;
  assign n639 = x118 & x128 ;
  assign n640 = x129 & n639 ;
  assign n641 = n638 | n640 ;
  assign n642 = x119 & ~x128 ;
  assign n643 = ( x129 & n641 ) | ( x129 & n642 ) | ( n641 & n642 ) ;
  assign n644 = x120 & x128 ;
  assign n645 = ( ~x129 & n641 ) | ( ~x129 & n644 ) | ( n641 & n644 ) ;
  assign n646 = n643 | n645 ;
  assign n647 = n179 & n646 ;
  assign n648 = n636 | n647 ;
  assign n649 = n625 | n648 ;
  assign n650 = ~n274 & n649 ;
  assign n651 = x113 & ~x128 ;
  assign n652 = ~x129 & n651 ;
  assign n653 = x110 & x128 ;
  assign n654 = x129 & n653 ;
  assign n655 = n652 | n654 ;
  assign n656 = x111 & ~x128 ;
  assign n657 = ( x129 & n655 ) | ( x129 & n656 ) | ( n655 & n656 ) ;
  assign n658 = x112 & x128 ;
  assign n659 = ( ~x129 & n655 ) | ( ~x129 & n658 ) | ( n655 & n658 ) ;
  assign n660 = n657 | n659 ;
  assign n661 = ~n145 & n660 ;
  assign n662 = x109 & ~x128 ;
  assign n663 = ~x129 & n662 ;
  assign n664 = x106 & x128 ;
  assign n665 = x129 & n664 ;
  assign n666 = n663 | n665 ;
  assign n667 = x107 & ~x128 ;
  assign n668 = ( x129 & n666 ) | ( x129 & n667 ) | ( n666 & n667 ) ;
  assign n669 = x108 & x128 ;
  assign n670 = ( ~x129 & n666 ) | ( ~x129 & n669 ) | ( n666 & n669 ) ;
  assign n671 = n668 | n670 ;
  assign n672 = n156 & n671 ;
  assign n673 = n661 | n672 ;
  assign n674 = x101 & ~x128 ;
  assign n675 = ~x129 & n674 ;
  assign n676 = x98 & x128 ;
  assign n677 = x129 & n676 ;
  assign n678 = n675 | n677 ;
  assign n679 = x99 & ~x128 ;
  assign n680 = ( x129 & n678 ) | ( x129 & n679 ) | ( n678 & n679 ) ;
  assign n681 = x100 & x128 ;
  assign n682 = ( ~x129 & n678 ) | ( ~x129 & n681 ) | ( n678 & n681 ) ;
  assign n683 = n680 | n682 ;
  assign n684 = n168 & n683 ;
  assign n685 = x105 & ~x128 ;
  assign n686 = ~x129 & n685 ;
  assign n687 = x102 & x128 ;
  assign n688 = x129 & n687 ;
  assign n689 = n686 | n688 ;
  assign n690 = x103 & ~x128 ;
  assign n691 = ( x129 & n689 ) | ( x129 & n690 ) | ( n689 & n690 ) ;
  assign n692 = x104 & x128 ;
  assign n693 = ( ~x129 & n689 ) | ( ~x129 & n692 ) | ( n689 & n692 ) ;
  assign n694 = n691 | n693 ;
  assign n695 = n179 & n694 ;
  assign n696 = n684 | n695 ;
  assign n697 = n673 | n696 ;
  assign n698 = n319 & n697 ;
  assign n699 = n650 | n698 ;
  assign n700 = n602 | n699 ;
  assign n701 = ~x134 & n700 ;
  assign n702 = x65 & ~x128 ;
  assign n703 = ~x129 & n702 ;
  assign n704 = x62 & x128 ;
  assign n705 = x129 & n704 ;
  assign n706 = n703 | n705 ;
  assign n707 = x63 & ~x128 ;
  assign n708 = ( x129 & n706 ) | ( x129 & n707 ) | ( n706 & n707 ) ;
  assign n709 = x64 & x128 ;
  assign n710 = ( ~x129 & n706 ) | ( ~x129 & n709 ) | ( n706 & n709 ) ;
  assign n711 = n708 | n710 ;
  assign n712 = ~n145 & n711 ;
  assign n713 = x61 & ~x128 ;
  assign n714 = ~x129 & n713 ;
  assign n715 = x58 & x128 ;
  assign n716 = x129 & n715 ;
  assign n717 = n714 | n716 ;
  assign n718 = x59 & ~x128 ;
  assign n719 = ( x129 & n717 ) | ( x129 & n718 ) | ( n717 & n718 ) ;
  assign n720 = x60 & x128 ;
  assign n721 = ( ~x129 & n717 ) | ( ~x129 & n720 ) | ( n717 & n720 ) ;
  assign n722 = n719 | n721 ;
  assign n723 = n156 & n722 ;
  assign n724 = n712 | n723 ;
  assign n725 = x53 & ~x128 ;
  assign n726 = ~x129 & n725 ;
  assign n727 = x50 & x128 ;
  assign n728 = x129 & n727 ;
  assign n729 = n726 | n728 ;
  assign n730 = x51 & ~x128 ;
  assign n731 = ( x129 & n729 ) | ( x129 & n730 ) | ( n729 & n730 ) ;
  assign n732 = x52 & x128 ;
  assign n733 = ( ~x129 & n729 ) | ( ~x129 & n732 ) | ( n729 & n732 ) ;
  assign n734 = n731 | n733 ;
  assign n735 = n168 & n734 ;
  assign n736 = x57 & ~x128 ;
  assign n737 = ~x129 & n736 ;
  assign n738 = x54 & x128 ;
  assign n739 = x129 & n738 ;
  assign n740 = n737 | n739 ;
  assign n741 = x55 & ~x128 ;
  assign n742 = ( x129 & n740 ) | ( x129 & n741 ) | ( n740 & n741 ) ;
  assign n743 = x56 & x128 ;
  assign n744 = ( ~x129 & n740 ) | ( ~x129 & n743 ) | ( n740 & n743 ) ;
  assign n745 = n742 | n744 ;
  assign n746 = n179 & n745 ;
  assign n747 = n735 | n746 ;
  assign n748 = n724 | n747 ;
  assign n749 = ~n274 & n748 ;
  assign n750 = x17 & ~x128 ;
  assign n751 = ~x129 & n750 ;
  assign n752 = x14 & x128 ;
  assign n753 = x129 & n752 ;
  assign n754 = n751 | n753 ;
  assign n755 = x15 & ~x128 ;
  assign n756 = ( x129 & n754 ) | ( x129 & n755 ) | ( n754 & n755 ) ;
  assign n757 = x16 & x128 ;
  assign n758 = ( ~x129 & n754 ) | ( ~x129 & n757 ) | ( n754 & n757 ) ;
  assign n759 = n756 | n758 ;
  assign n760 = ~n145 & n759 ;
  assign n761 = x13 & ~x128 ;
  assign n762 = ~x129 & n761 ;
  assign n763 = x10 & x128 ;
  assign n764 = x129 & n763 ;
  assign n765 = n762 | n764 ;
  assign n766 = x11 & ~x128 ;
  assign n767 = ( x129 & n765 ) | ( x129 & n766 ) | ( n765 & n766 ) ;
  assign n768 = x12 & x128 ;
  assign n769 = ( ~x129 & n765 ) | ( ~x129 & n768 ) | ( n765 & n768 ) ;
  assign n770 = n767 | n769 ;
  assign n771 = n156 & n770 ;
  assign n772 = n760 | n771 ;
  assign n773 = x5 & ~x128 ;
  assign n774 = ~x129 & n773 ;
  assign n775 = x2 & x128 ;
  assign n776 = x129 & n775 ;
  assign n777 = n774 | n776 ;
  assign n778 = x3 & ~x128 ;
  assign n779 = ( x129 & n777 ) | ( x129 & n778 ) | ( n777 & n778 ) ;
  assign n780 = x4 & x128 ;
  assign n781 = ( ~x129 & n777 ) | ( ~x129 & n780 ) | ( n777 & n780 ) ;
  assign n782 = n779 | n781 ;
  assign n783 = n168 & n782 ;
  assign n784 = x9 & ~x128 ;
  assign n785 = ~x129 & n784 ;
  assign n786 = x6 & x128 ;
  assign n787 = x129 & n786 ;
  assign n788 = n785 | n787 ;
  assign n789 = x7 & ~x128 ;
  assign n790 = ( x129 & n788 ) | ( x129 & n789 ) | ( n788 & n789 ) ;
  assign n791 = x8 & x128 ;
  assign n792 = ( ~x129 & n788 ) | ( ~x129 & n791 ) | ( n788 & n791 ) ;
  assign n793 = n790 | n792 ;
  assign n794 = n179 & n793 ;
  assign n795 = n783 | n794 ;
  assign n796 = n772 | n795 ;
  assign n797 = n183 & n796 ;
  assign n798 = n749 | n797 ;
  assign n799 = x49 & ~x128 ;
  assign n800 = ~x129 & n799 ;
  assign n801 = x46 & x128 ;
  assign n802 = x129 & n801 ;
  assign n803 = n800 | n802 ;
  assign n804 = x47 & ~x128 ;
  assign n805 = ( x129 & n803 ) | ( x129 & n804 ) | ( n803 & n804 ) ;
  assign n806 = x48 & x128 ;
  assign n807 = ( ~x129 & n803 ) | ( ~x129 & n806 ) | ( n803 & n806 ) ;
  assign n808 = n805 | n807 ;
  assign n809 = ~n145 & n808 ;
  assign n810 = x42 & x128 ;
  assign n811 = x43 & ~x128 ;
  assign n812 = n810 | n811 ;
  assign n813 = x129 & n812 ;
  assign n814 = x45 & ~x128 ;
  assign n815 = x44 & x128 ;
  assign n816 = n814 | n815 ;
  assign n817 = ~x129 & n816 ;
  assign n818 = n813 | n817 ;
  assign n819 = n156 & n818 ;
  assign n820 = n809 | n819 ;
  assign n821 = x37 & ~x128 ;
  assign n822 = ~x129 & n821 ;
  assign n823 = x34 & x128 ;
  assign n824 = x129 & n823 ;
  assign n825 = n822 | n824 ;
  assign n826 = x35 & ~x128 ;
  assign n827 = ( x129 & n825 ) | ( x129 & n826 ) | ( n825 & n826 ) ;
  assign n828 = x36 & x128 ;
  assign n829 = ( ~x129 & n825 ) | ( ~x129 & n828 ) | ( n825 & n828 ) ;
  assign n830 = n827 | n829 ;
  assign n831 = n168 & n830 ;
  assign n832 = x41 & ~x128 ;
  assign n833 = x40 & x128 ;
  assign n834 = n832 | n833 ;
  assign n835 = ~x129 & n834 ;
  assign n836 = x39 & ~x128 ;
  assign n837 = x38 & x128 ;
  assign n838 = n836 | n837 ;
  assign n839 = x129 & n838 ;
  assign n840 = n835 | n839 ;
  assign n841 = n179 & n840 ;
  assign n842 = n831 | n841 ;
  assign n843 = n820 | n842 ;
  assign n844 = n319 & n843 ;
  assign n845 = x33 & ~x128 ;
  assign n846 = ~x129 & n845 ;
  assign n847 = x30 & x128 ;
  assign n848 = x129 & n847 ;
  assign n849 = n846 | n848 ;
  assign n850 = x31 & ~x128 ;
  assign n851 = ( x129 & n849 ) | ( x129 & n850 ) | ( n849 & n850 ) ;
  assign n852 = x32 & x128 ;
  assign n853 = ( ~x129 & n849 ) | ( ~x129 & n852 ) | ( n849 & n852 ) ;
  assign n854 = n851 | n853 ;
  assign n855 = ~n145 & n854 ;
  assign n856 = x29 & ~x128 ;
  assign n857 = ~x129 & n856 ;
  assign n858 = x26 & x128 ;
  assign n859 = x129 & n858 ;
  assign n860 = n857 | n859 ;
  assign n861 = x27 & ~x128 ;
  assign n862 = ( x129 & n860 ) | ( x129 & n861 ) | ( n860 & n861 ) ;
  assign n863 = x28 & x128 ;
  assign n864 = ( ~x129 & n860 ) | ( ~x129 & n863 ) | ( n860 & n863 ) ;
  assign n865 = n862 | n864 ;
  assign n866 = n156 & n865 ;
  assign n867 = n855 | n866 ;
  assign n868 = x21 & ~x128 ;
  assign n869 = ~x129 & n868 ;
  assign n870 = x18 & x128 ;
  assign n871 = x129 & n870 ;
  assign n872 = n869 | n871 ;
  assign n873 = x19 & ~x128 ;
  assign n874 = ( x129 & n872 ) | ( x129 & n873 ) | ( n872 & n873 ) ;
  assign n875 = x20 & x128 ;
  assign n876 = ( ~x129 & n872 ) | ( ~x129 & n875 ) | ( n872 & n875 ) ;
  assign n877 = n874 | n876 ;
  assign n878 = n168 & n877 ;
  assign n879 = x25 & ~x128 ;
  assign n880 = ~x129 & n879 ;
  assign n881 = x22 & x128 ;
  assign n882 = x129 & n881 ;
  assign n883 = n880 | n882 ;
  assign n884 = x23 & ~x128 ;
  assign n885 = ( x129 & n883 ) | ( x129 & n884 ) | ( n883 & n884 ) ;
  assign n886 = x24 & x128 ;
  assign n887 = ( ~x129 & n883 ) | ( ~x129 & n886 ) | ( n883 & n886 ) ;
  assign n888 = n885 | n887 ;
  assign n889 = n179 & n888 ;
  assign n890 = n878 | n889 ;
  assign n891 = n867 | n890 ;
  assign n892 = n228 & n891 ;
  assign n893 = n844 | n892 ;
  assign n894 = n798 | n893 ;
  assign n895 = x134 & n894 ;
  assign n896 = n701 | n895 ;
  assign n897 = ~x129 & n208 ;
  assign n898 = x129 & n142 ;
  assign n899 = n897 | n898 ;
  assign n900 = ~n145 & n899 ;
  assign n901 = ~x129 & n138 ;
  assign n902 = x129 & n153 ;
  assign n903 = n901 | n902 ;
  assign n904 = n156 & n903 ;
  assign n905 = n900 | n904 ;
  assign n906 = ~x129 & n172 ;
  assign n907 = x129 & n165 ;
  assign n908 = n906 | n907 ;
  assign n909 = n168 & n908 ;
  assign n910 = ~x129 & n149 ;
  assign n911 = x129 & n176 ;
  assign n912 = n910 | n911 ;
  assign n913 = n179 & n912 ;
  assign n914 = n909 | n913 ;
  assign n915 = n905 | n914 ;
  assign n916 = n183 & n915 ;
  assign n917 = ~x129 & n299 ;
  assign n918 = x129 & n191 ;
  assign n919 = n917 | n918 ;
  assign n920 = ~n145 & n919 ;
  assign n921 = ~x129 & n187 ;
  assign n922 = x129 & n201 ;
  assign n923 = n921 | n922 ;
  assign n924 = n156 & n923 ;
  assign n925 = n920 | n924 ;
  assign n926 = ~x129 & n218 ;
  assign n927 = x129 & n212 ;
  assign n928 = n926 | n927 ;
  assign n929 = n168 & n928 ;
  assign n930 = ~x129 & n197 ;
  assign n931 = x129 & n222 ;
  assign n932 = n930 | n931 ;
  assign n933 = n179 & n932 ;
  assign n934 = n929 | n933 ;
  assign n935 = n925 | n934 ;
  assign n936 = n228 & n935 ;
  assign n937 = n916 | n936 ;
  assign n938 = ~x129 & n347 ;
  assign n939 = x129 & n237 ;
  assign n940 = n938 | n939 ;
  assign n941 = ~n145 & n940 ;
  assign n942 = ~x129 & n233 ;
  assign n943 = x129 & n247 ;
  assign n944 = n942 | n943 ;
  assign n945 = n156 & n944 ;
  assign n946 = n941 | n945 ;
  assign n947 = ~x129 & n264 ;
  assign n948 = x129 & n258 ;
  assign n949 = n947 | n948 ;
  assign n950 = n168 & n949 ;
  assign n951 = ~x129 & n243 ;
  assign n952 = x129 & n268 ;
  assign n953 = n951 | n952 ;
  assign n954 = n179 & n953 ;
  assign n955 = n950 | n954 ;
  assign n956 = n946 | n955 ;
  assign n957 = ~n274 & n956 ;
  assign n958 = ~x129 & n254 ;
  assign n959 = x129 & n282 ;
  assign n960 = n958 | n959 ;
  assign n961 = ~n145 & n960 ;
  assign n962 = ~x129 & n278 ;
  assign n963 = x129 & n292 ;
  assign n964 = n962 | n963 ;
  assign n965 = n156 & n964 ;
  assign n966 = n961 | n965 ;
  assign n967 = ~x129 & n309 ;
  assign n968 = x129 & n303 ;
  assign n969 = n967 | n968 ;
  assign n970 = n168 & n969 ;
  assign n971 = ~x129 & n288 ;
  assign n972 = x129 & n313 ;
  assign n973 = n971 | n972 ;
  assign n974 = n179 & n973 ;
  assign n975 = n970 | n974 ;
  assign n976 = n966 | n975 ;
  assign n977 = n319 & n976 ;
  assign n978 = n957 | n977 ;
  assign n979 = n937 | n978 ;
  assign n980 = ~x134 & n979 ;
  assign n981 = ~x129 & n161 ;
  assign n982 = x129 & n419 ;
  assign n983 = n981 | n982 ;
  assign n984 = ~n145 & n983 ;
  assign n985 = ~x129 & n415 ;
  assign n986 = x129 & n429 ;
  assign n987 = n985 | n986 ;
  assign n988 = n156 & n987 ;
  assign n989 = n984 | n988 ;
  assign n990 = ~x129 & n446 ;
  assign n991 = x129 & n440 ;
  assign n992 = n990 | n991 ;
  assign n993 = n168 & n992 ;
  assign n994 = ~x129 & n425 ;
  assign n995 = x129 & n450 ;
  assign n996 = n994 | n995 ;
  assign n997 = n179 & n996 ;
  assign n998 = n993 | n997 ;
  assign n999 = n989 | n998 ;
  assign n1000 = ~n274 & n999 ;
  assign n1001 = ~x129 & n391 ;
  assign n1002 = x129 & n330 ;
  assign n1003 = n1001 | n1002 ;
  assign n1004 = ~n145 & n1003 ;
  assign n1005 = ~x129 & n326 ;
  assign n1006 = x129 & n340 ;
  assign n1007 = n1005 | n1006 ;
  assign n1008 = n156 & n1007 ;
  assign n1009 = n1004 | n1008 ;
  assign n1010 = ~x129 & n357 ;
  assign n1011 = x129 & n351 ;
  assign n1012 = n1010 | n1011 ;
  assign n1013 = n168 & n1012 ;
  assign n1014 = ~x129 & n336 ;
  assign n1015 = x129 & n361 ;
  assign n1016 = n1014 | n1015 ;
  assign n1017 = n179 & n1016 ;
  assign n1018 = n1013 | n1017 ;
  assign n1019 = n1009 | n1018 ;
  assign n1020 = n183 & n1019 ;
  assign n1021 = n1000 | n1020 ;
  assign n1022 = ~x129 & n436 ;
  assign n1023 = x129 & n485 ;
  assign n1024 = n1022 | n1023 ;
  assign n1025 = ~n145 & n1024 ;
  assign n1026 = x129 & n495 ;
  assign n1027 = ~x129 & n481 ;
  assign n1028 = n1026 | n1027 ;
  assign n1029 = n156 & n1028 ;
  assign n1030 = n1025 | n1029 ;
  assign n1031 = n469 | n472 ;
  assign n1032 = ~x129 & n1031 ;
  assign n1033 = x129 & n463 ;
  assign n1034 = n1032 | n1033 ;
  assign n1035 = n168 & n1034 ;
  assign n1036 = ~x129 & n491 ;
  assign n1037 = n467 | n474 ;
  assign n1038 = x129 & n1037 ;
  assign n1039 = n1036 | n1038 ;
  assign n1040 = n179 & n1039 ;
  assign n1041 = n1035 | n1040 ;
  assign n1042 = n1030 | n1041 ;
  assign n1043 = n319 & n1042 ;
  assign n1044 = ~x129 & n459 ;
  assign n1045 = x129 & n374 ;
  assign n1046 = n1044 | n1045 ;
  assign n1047 = ~n145 & n1046 ;
  assign n1048 = ~x129 & n370 ;
  assign n1049 = x129 & n384 ;
  assign n1050 = n1048 | n1049 ;
  assign n1051 = n156 & n1050 ;
  assign n1052 = n1047 | n1051 ;
  assign n1053 = ~x129 & n401 ;
  assign n1054 = x129 & n395 ;
  assign n1055 = n1053 | n1054 ;
  assign n1056 = n168 & n1055 ;
  assign n1057 = ~x129 & n380 ;
  assign n1058 = x129 & n405 ;
  assign n1059 = n1057 | n1058 ;
  assign n1060 = n179 & n1059 ;
  assign n1061 = n1056 | n1060 ;
  assign n1062 = n1052 | n1061 ;
  assign n1063 = n228 & n1062 ;
  assign n1064 = n1043 | n1063 ;
  assign n1065 = n1021 | n1064 ;
  assign n1066 = x134 & n1065 ;
  assign n1067 = n980 | n1066 ;
  assign n1068 = x129 & n651 ;
  assign n1069 = ~x129 & n628 ;
  assign n1070 = n1068 | n1069 ;
  assign n1071 = ( x129 & n658 ) | ( x129 & n1070 ) | ( n658 & n1070 ) ;
  assign n1072 = ( ~x129 & n631 ) | ( ~x129 & n1070 ) | ( n631 & n1070 ) ;
  assign n1073 = n1071 | n1072 ;
  assign n1074 = ~n145 & n1073 ;
  assign n1075 = x129 & n662 ;
  assign n1076 = ~x129 & n653 ;
  assign n1077 = n1075 | n1076 ;
  assign n1078 = ( x129 & n669 ) | ( x129 & n1077 ) | ( n669 & n1077 ) ;
  assign n1079 = ( ~x129 & n656 ) | ( ~x129 & n1077 ) | ( n656 & n1077 ) ;
  assign n1080 = n1078 | n1079 ;
  assign n1081 = n156 & n1080 ;
  assign n1082 = n1074 | n1081 ;
  assign n1083 = x129 & n674 ;
  assign n1084 = ~x129 & n687 ;
  assign n1085 = n1083 | n1084 ;
  assign n1086 = ( x129 & n681 ) | ( x129 & n1085 ) | ( n681 & n1085 ) ;
  assign n1087 = ( ~x129 & n690 ) | ( ~x129 & n1085 ) | ( n690 & n1085 ) ;
  assign n1088 = n1086 | n1087 ;
  assign n1089 = n168 & n1088 ;
  assign n1090 = x129 & n685 ;
  assign n1091 = ~x129 & n664 ;
  assign n1092 = n1090 | n1091 ;
  assign n1093 = ( x129 & n692 ) | ( x129 & n1092 ) | ( n692 & n1092 ) ;
  assign n1094 = ( ~x129 & n667 ) | ( ~x129 & n1092 ) | ( n667 & n1092 ) ;
  assign n1095 = n1093 | n1094 ;
  assign n1096 = n179 & n1095 ;
  assign n1097 = n1089 | n1096 ;
  assign n1098 = n1082 | n1097 ;
  assign n1099 = n319 & n1098 ;
  assign n1100 = x129 & n554 ;
  assign n1101 = ~x129 & n676 ;
  assign n1102 = n1100 | n1101 ;
  assign n1103 = ( x129 & n561 ) | ( x129 & n1102 ) | ( n561 & n1102 ) ;
  assign n1104 = ( ~x129 & n679 ) | ( ~x129 & n1102 ) | ( n679 & n1102 ) ;
  assign n1105 = n1103 | n1104 ;
  assign n1106 = ~n145 & n1105 ;
  assign n1107 = x129 & n565 ;
  assign n1108 = ~x129 & n556 ;
  assign n1109 = n1107 | n1108 ;
  assign n1110 = ( x129 & n572 ) | ( x129 & n1109 ) | ( n572 & n1109 ) ;
  assign n1111 = ( ~x129 & n559 ) | ( ~x129 & n1109 ) | ( n559 & n1109 ) ;
  assign n1112 = n1110 | n1111 ;
  assign n1113 = n156 & n1112 ;
  assign n1114 = n1106 | n1113 ;
  assign n1115 = x129 & n577 ;
  assign n1116 = ~x129 & n590 ;
  assign n1117 = n1115 | n1116 ;
  assign n1118 = ( x129 & n584 ) | ( x129 & n1117 ) | ( n584 & n1117 ) ;
  assign n1119 = ( ~x129 & n593 ) | ( ~x129 & n1117 ) | ( n593 & n1117 ) ;
  assign n1120 = n1118 | n1119 ;
  assign n1121 = n168 & n1120 ;
  assign n1122 = x129 & n588 ;
  assign n1123 = ~x129 & n567 ;
  assign n1124 = n1122 | n1123 ;
  assign n1125 = ( x129 & n595 ) | ( x129 & n1124 ) | ( n595 & n1124 ) ;
  assign n1126 = ( ~x129 & n570 ) | ( ~x129 & n1124 ) | ( n570 & n1124 ) ;
  assign n1127 = n1125 | n1126 ;
  assign n1128 = n179 & n1127 ;
  assign n1129 = n1121 | n1128 ;
  assign n1130 = n1114 | n1129 ;
  assign n1131 = n228 & n1130 ;
  assign n1132 = n1099 | n1131 ;
  assign n1133 = x129 & n603 ;
  assign n1134 = ~x129 & n775 ;
  assign n1135 = n1133 | n1134 ;
  assign n1136 = ( x129 & n610 ) | ( x129 & n1135 ) | ( n610 & n1135 ) ;
  assign n1137 = ( ~x129 & n778 ) | ( ~x129 & n1135 ) | ( n778 & n1135 ) ;
  assign n1138 = n1136 | n1137 ;
  assign n1139 = ~n145 & n1138 ;
  assign n1140 = x129 & n614 ;
  assign n1141 = ~x129 & n605 ;
  assign n1142 = n1140 | n1141 ;
  assign n1143 = ( x129 & n621 ) | ( x129 & n1142 ) | ( n621 & n1142 ) ;
  assign n1144 = ( ~x129 & n608 ) | ( ~x129 & n1142 ) | ( n608 & n1142 ) ;
  assign n1145 = n1143 | n1144 ;
  assign n1146 = n156 & n1145 ;
  assign n1147 = n1139 | n1146 ;
  assign n1148 = x129 & n626 ;
  assign n1149 = ~x129 & n639 ;
  assign n1150 = n1148 | n1149 ;
  assign n1151 = ( x129 & n633 ) | ( x129 & n1150 ) | ( n633 & n1150 ) ;
  assign n1152 = ( ~x129 & n642 ) | ( ~x129 & n1150 ) | ( n642 & n1150 ) ;
  assign n1153 = n1151 | n1152 ;
  assign n1154 = n168 & n1153 ;
  assign n1155 = x129 & n637 ;
  assign n1156 = ~x129 & n616 ;
  assign n1157 = n1155 | n1156 ;
  assign n1158 = ( x129 & n644 ) | ( x129 & n1157 ) | ( n644 & n1157 ) ;
  assign n1159 = ( ~x129 & n619 ) | ( ~x129 & n1157 ) | ( n619 & n1157 ) ;
  assign n1160 = n1158 | n1159 ;
  assign n1161 = n179 & n1160 ;
  assign n1162 = n1154 | n1161 ;
  assign n1163 = n1147 | n1162 ;
  assign n1164 = ~n274 & n1163 ;
  assign n1165 = x129 & n506 ;
  assign n1166 = ~x129 & n579 ;
  assign n1167 = n1165 | n1166 ;
  assign n1168 = ( x129 & n513 ) | ( x129 & n1167 ) | ( n513 & n1167 ) ;
  assign n1169 = ( ~x129 & n582 ) | ( ~x129 & n1167 ) | ( n582 & n1167 ) ;
  assign n1170 = n1168 | n1169 ;
  assign n1171 = ~n145 & n1170 ;
  assign n1172 = x129 & n517 ;
  assign n1173 = ~x129 & n508 ;
  assign n1174 = n1172 | n1173 ;
  assign n1175 = ( x129 & n524 ) | ( x129 & n1174 ) | ( n524 & n1174 ) ;
  assign n1176 = ( ~x129 & n511 ) | ( ~x129 & n1174 ) | ( n511 & n1174 ) ;
  assign n1177 = n1175 | n1176 ;
  assign n1178 = n156 & n1177 ;
  assign n1179 = n1171 | n1178 ;
  assign n1180 = x129 & n529 ;
  assign n1181 = ~x129 & n542 ;
  assign n1182 = n1180 | n1181 ;
  assign n1183 = ( x129 & n536 ) | ( x129 & n1182 ) | ( n536 & n1182 ) ;
  assign n1184 = ( ~x129 & n545 ) | ( ~x129 & n1182 ) | ( n545 & n1182 ) ;
  assign n1185 = n1183 | n1184 ;
  assign n1186 = n168 & n1185 ;
  assign n1187 = x129 & n540 ;
  assign n1188 = ~x129 & n519 ;
  assign n1189 = n1187 | n1188 ;
  assign n1190 = ( x129 & n547 ) | ( x129 & n1189 ) | ( n547 & n1189 ) ;
  assign n1191 = ( ~x129 & n522 ) | ( ~x129 & n1189 ) | ( n522 & n1189 ) ;
  assign n1192 = n1190 | n1191 ;
  assign n1193 = n179 & n1192 ;
  assign n1194 = n1186 | n1193 ;
  assign n1195 = n1179 | n1194 ;
  assign n1196 = n183 & n1195 ;
  assign n1197 = n1164 | n1196 ;
  assign n1198 = n1132 | n1197 ;
  assign n1199 = ~x134 & n1198 ;
  assign n1200 = x129 & n702 ;
  assign n1201 = ~x129 & n531 ;
  assign n1202 = n1200 | n1201 ;
  assign n1203 = ( x129 & n709 ) | ( x129 & n1202 ) | ( n709 & n1202 ) ;
  assign n1204 = ( ~x129 & n534 ) | ( ~x129 & n1202 ) | ( n534 & n1202 ) ;
  assign n1205 = n1203 | n1204 ;
  assign n1206 = ~n145 & n1205 ;
  assign n1207 = x129 & n713 ;
  assign n1208 = ~x129 & n704 ;
  assign n1209 = n1207 | n1208 ;
  assign n1210 = ( x129 & n720 ) | ( x129 & n1209 ) | ( n720 & n1209 ) ;
  assign n1211 = ( ~x129 & n707 ) | ( ~x129 & n1209 ) | ( n707 & n1209 ) ;
  assign n1212 = n1210 | n1211 ;
  assign n1213 = n156 & n1212 ;
  assign n1214 = n1206 | n1213 ;
  assign n1215 = x129 & n725 ;
  assign n1216 = ~x129 & n738 ;
  assign n1217 = n1215 | n1216 ;
  assign n1218 = ( x129 & n732 ) | ( x129 & n1217 ) | ( n732 & n1217 ) ;
  assign n1219 = ( ~x129 & n741 ) | ( ~x129 & n1217 ) | ( n741 & n1217 ) ;
  assign n1220 = n1218 | n1219 ;
  assign n1221 = n168 & n1220 ;
  assign n1222 = x129 & n736 ;
  assign n1223 = ~x129 & n715 ;
  assign n1224 = n1222 | n1223 ;
  assign n1225 = ( x129 & n743 ) | ( x129 & n1224 ) | ( n743 & n1224 ) ;
  assign n1226 = ( ~x129 & n718 ) | ( ~x129 & n1224 ) | ( n718 & n1224 ) ;
  assign n1227 = n1225 | n1226 ;
  assign n1228 = n179 & n1227 ;
  assign n1229 = n1221 | n1228 ;
  assign n1230 = n1214 | n1229 ;
  assign n1231 = ~n274 & n1230 ;
  assign n1232 = x129 & n799 ;
  assign n1233 = ~x129 & n727 ;
  assign n1234 = n1232 | n1233 ;
  assign n1235 = ( x129 & n806 ) | ( x129 & n1234 ) | ( n806 & n1234 ) ;
  assign n1236 = ( ~x129 & n730 ) | ( ~x129 & n1234 ) | ( n730 & n1234 ) ;
  assign n1237 = n1235 | n1236 ;
  assign n1238 = ~n145 & n1237 ;
  assign n1239 = x129 & n816 ;
  assign n1240 = n801 | n804 ;
  assign n1241 = ~x129 & n1240 ;
  assign n1242 = n1239 | n1241 ;
  assign n1243 = n156 & n1242 ;
  assign n1244 = n1238 | n1243 ;
  assign n1245 = x129 & n821 ;
  assign n1246 = ~x129 & n837 ;
  assign n1247 = n1245 | n1246 ;
  assign n1248 = ( x129 & n828 ) | ( x129 & n1247 ) | ( n828 & n1247 ) ;
  assign n1249 = ( ~x129 & n836 ) | ( ~x129 & n1247 ) | ( n836 & n1247 ) ;
  assign n1250 = n1248 | n1249 ;
  assign n1251 = n168 & n1250 ;
  assign n1252 = x129 & n832 ;
  assign n1253 = ~x129 & n810 ;
  assign n1254 = n1252 | n1253 ;
  assign n1255 = ( x129 & n833 ) | ( x129 & n1254 ) | ( n833 & n1254 ) ;
  assign n1256 = ( ~x129 & n811 ) | ( ~x129 & n1254 ) | ( n811 & n1254 ) ;
  assign n1257 = n1255 | n1256 ;
  assign n1258 = n179 & n1257 ;
  assign n1259 = n1251 | n1258 ;
  assign n1260 = n1244 | n1259 ;
  assign n1261 = n319 & n1260 ;
  assign n1262 = n1231 | n1261 ;
  assign n1263 = x129 & n750 ;
  assign n1264 = ~x129 & n870 ;
  assign n1265 = n1263 | n1264 ;
  assign n1266 = ( x129 & n757 ) | ( x129 & n1265 ) | ( n757 & n1265 ) ;
  assign n1267 = ( ~x129 & n873 ) | ( ~x129 & n1265 ) | ( n873 & n1265 ) ;
  assign n1268 = n1266 | n1267 ;
  assign n1269 = ~n145 & n1268 ;
  assign n1270 = x129 & n761 ;
  assign n1271 = ~x129 & n752 ;
  assign n1272 = n1270 | n1271 ;
  assign n1273 = ( x129 & n768 ) | ( x129 & n1272 ) | ( n768 & n1272 ) ;
  assign n1274 = ( ~x129 & n755 ) | ( ~x129 & n1272 ) | ( n755 & n1272 ) ;
  assign n1275 = n1273 | n1274 ;
  assign n1276 = n156 & n1275 ;
  assign n1277 = n1269 | n1276 ;
  assign n1278 = x129 & n773 ;
  assign n1279 = ~x129 & n786 ;
  assign n1280 = n1278 | n1279 ;
  assign n1281 = ( x129 & n780 ) | ( x129 & n1280 ) | ( n780 & n1280 ) ;
  assign n1282 = ( ~x129 & n789 ) | ( ~x129 & n1280 ) | ( n789 & n1280 ) ;
  assign n1283 = n1281 | n1282 ;
  assign n1284 = n168 & n1283 ;
  assign n1285 = x129 & n784 ;
  assign n1286 = ~x129 & n763 ;
  assign n1287 = n1285 | n1286 ;
  assign n1288 = ( x129 & n791 ) | ( x129 & n1287 ) | ( n791 & n1287 ) ;
  assign n1289 = ( ~x129 & n766 ) | ( ~x129 & n1287 ) | ( n766 & n1287 ) ;
  assign n1290 = n1288 | n1289 ;
  assign n1291 = n179 & n1290 ;
  assign n1292 = n1284 | n1291 ;
  assign n1293 = n1277 | n1292 ;
  assign n1294 = n183 & n1293 ;
  assign n1295 = x129 & n845 ;
  assign n1296 = ~x129 & n823 ;
  assign n1297 = n1295 | n1296 ;
  assign n1298 = ( x129 & n852 ) | ( x129 & n1297 ) | ( n852 & n1297 ) ;
  assign n1299 = ( ~x129 & n826 ) | ( ~x129 & n1297 ) | ( n826 & n1297 ) ;
  assign n1300 = n1298 | n1299 ;
  assign n1301 = ~n145 & n1300 ;
  assign n1302 = x129 & n856 ;
  assign n1303 = ~x129 & n847 ;
  assign n1304 = n1302 | n1303 ;
  assign n1305 = ( x129 & n863 ) | ( x129 & n1304 ) | ( n863 & n1304 ) ;
  assign n1306 = ( ~x129 & n850 ) | ( ~x129 & n1304 ) | ( n850 & n1304 ) ;
  assign n1307 = n1305 | n1306 ;
  assign n1308 = n156 & n1307 ;
  assign n1309 = n1301 | n1308 ;
  assign n1310 = x129 & n868 ;
  assign n1311 = ~x129 & n881 ;
  assign n1312 = n1310 | n1311 ;
  assign n1313 = ( x129 & n875 ) | ( x129 & n1312 ) | ( n875 & n1312 ) ;
  assign n1314 = ( ~x129 & n884 ) | ( ~x129 & n1312 ) | ( n884 & n1312 ) ;
  assign n1315 = n1313 | n1314 ;
  assign n1316 = n168 & n1315 ;
  assign n1317 = x129 & n879 ;
  assign n1318 = ~x129 & n858 ;
  assign n1319 = n1317 | n1318 ;
  assign n1320 = ( x129 & n886 ) | ( x129 & n1319 ) | ( n886 & n1319 ) ;
  assign n1321 = ( ~x129 & n861 ) | ( ~x129 & n1319 ) | ( n861 & n1319 ) ;
  assign n1322 = n1320 | n1321 ;
  assign n1323 = n179 & n1322 ;
  assign n1324 = n1316 | n1323 ;
  assign n1325 = n1309 | n1324 ;
  assign n1326 = n228 & n1325 ;
  assign n1327 = n1294 | n1326 ;
  assign n1328 = n1262 | n1327 ;
  assign n1329 = x134 & n1328 ;
  assign n1330 = n1199 | n1329 ;
  assign n1331 = ~n145 & n214 ;
  assign n1332 = n144 & n156 ;
  assign n1333 = n1331 | n1332 ;
  assign n1334 = n168 & n178 ;
  assign n1335 = n155 & n179 ;
  assign n1336 = n1334 | n1335 ;
  assign n1337 = n1333 | n1336 ;
  assign n1338 = n183 & n1337 ;
  assign n1339 = ~n145 & n305 ;
  assign n1340 = n156 & n193 ;
  assign n1341 = n1339 | n1340 ;
  assign n1342 = n168 & n224 ;
  assign n1343 = n179 & n203 ;
  assign n1344 = n1342 | n1343 ;
  assign n1345 = n1341 | n1344 ;
  assign n1346 = n228 & n1345 ;
  assign n1347 = n1338 | n1346 ;
  assign n1348 = ~n145 & n353 ;
  assign n1349 = n156 & n239 ;
  assign n1350 = n1348 | n1349 ;
  assign n1351 = n168 & n270 ;
  assign n1352 = n179 & n249 ;
  assign n1353 = n1351 | n1352 ;
  assign n1354 = n1350 | n1353 ;
  assign n1355 = ~n274 & n1354 ;
  assign n1356 = ~n145 & n260 ;
  assign n1357 = n156 & n284 ;
  assign n1358 = n1356 | n1357 ;
  assign n1359 = n168 & n315 ;
  assign n1360 = n179 & n294 ;
  assign n1361 = n1359 | n1360 ;
  assign n1362 = n1358 | n1361 ;
  assign n1363 = n319 & n1362 ;
  assign n1364 = n1355 | n1363 ;
  assign n1365 = n1347 | n1364 ;
  assign n1366 = ~x134 & n1365 ;
  assign n1367 = ~n145 & n167 ;
  assign n1368 = n156 & n421 ;
  assign n1369 = n1367 | n1368 ;
  assign n1370 = n168 & n452 ;
  assign n1371 = n179 & n431 ;
  assign n1372 = n1370 | n1371 ;
  assign n1373 = n1369 | n1372 ;
  assign n1374 = ~n274 & n1373 ;
  assign n1375 = n168 & n476 ;
  assign n1376 = n179 & n497 ;
  assign n1377 = n1375 | n1376 ;
  assign n1378 = ~n145 & n442 ;
  assign n1379 = n156 & n487 ;
  assign n1380 = n1378 | n1379 ;
  assign n1381 = n319 & n1380 ;
  assign n1382 = ( n319 & n1377 ) | ( n319 & n1381 ) | ( n1377 & n1381 ) ;
  assign n1383 = n1374 | n1382 ;
  assign n1384 = ~n145 & n465 ;
  assign n1385 = n156 & n376 ;
  assign n1386 = n1384 | n1385 ;
  assign n1387 = n168 & n407 ;
  assign n1388 = n179 & n386 ;
  assign n1389 = n1387 | n1388 ;
  assign n1390 = n1386 | n1389 ;
  assign n1391 = n228 & n1390 ;
  assign n1392 = ~n145 & n397 ;
  assign n1393 = n156 & n332 ;
  assign n1394 = n1392 | n1393 ;
  assign n1395 = n168 & n363 ;
  assign n1396 = n179 & n342 ;
  assign n1397 = n1395 | n1396 ;
  assign n1398 = n1394 | n1397 ;
  assign n1399 = n183 & n1398 ;
  assign n1400 = n1391 | n1399 ;
  assign n1401 = n1383 | n1400 ;
  assign n1402 = x134 & n1401 ;
  assign n1403 = n1366 | n1402 ;
  assign n1404 = ~n145 & n586 ;
  assign n1405 = n156 & n515 ;
  assign n1406 = n1404 | n1405 ;
  assign n1407 = n168 & n549 ;
  assign n1408 = n179 & n526 ;
  assign n1409 = n1407 | n1408 ;
  assign n1410 = n1406 | n1409 ;
  assign n1411 = n183 & n1410 ;
  assign n1412 = ~n145 & n683 ;
  assign n1413 = n156 & n563 ;
  assign n1414 = n1412 | n1413 ;
  assign n1415 = n168 & n597 ;
  assign n1416 = n179 & n574 ;
  assign n1417 = n1415 | n1416 ;
  assign n1418 = n1414 | n1417 ;
  assign n1419 = n228 & n1418 ;
  assign n1420 = n1411 | n1419 ;
  assign n1421 = ~n145 & n782 ;
  assign n1422 = n156 & n612 ;
  assign n1423 = n1421 | n1422 ;
  assign n1424 = n168 & n646 ;
  assign n1425 = n179 & n623 ;
  assign n1426 = n1424 | n1425 ;
  assign n1427 = n1423 | n1426 ;
  assign n1428 = ~n274 & n1427 ;
  assign n1429 = ~n145 & n635 ;
  assign n1430 = n156 & n660 ;
  assign n1431 = n1429 | n1430 ;
  assign n1432 = n168 & n694 ;
  assign n1433 = n179 & n671 ;
  assign n1434 = n1432 | n1433 ;
  assign n1435 = n1431 | n1434 ;
  assign n1436 = n319 & n1435 ;
  assign n1437 = n1428 | n1436 ;
  assign n1438 = n1420 | n1437 ;
  assign n1439 = ~x134 & n1438 ;
  assign n1440 = ~n145 & n538 ;
  assign n1441 = n156 & n711 ;
  assign n1442 = n1440 | n1441 ;
  assign n1443 = n168 & n745 ;
  assign n1444 = n179 & n722 ;
  assign n1445 = n1443 | n1444 ;
  assign n1446 = n1442 | n1445 ;
  assign n1447 = ~n274 & n1446 ;
  assign n1448 = ~n145 & n734 ;
  assign n1449 = n156 & n808 ;
  assign n1450 = n1448 | n1449 ;
  assign n1451 = n168 & n840 ;
  assign n1452 = n179 & n818 ;
  assign n1453 = n1451 | n1452 ;
  assign n1454 = n319 & n1453 ;
  assign n1455 = ( n319 & n1450 ) | ( n319 & n1454 ) | ( n1450 & n1454 ) ;
  assign n1456 = n1447 | n1455 ;
  assign n1457 = ~n145 & n830 ;
  assign n1458 = n156 & n854 ;
  assign n1459 = n1457 | n1458 ;
  assign n1460 = n168 & n888 ;
  assign n1461 = n179 & n865 ;
  assign n1462 = n1460 | n1461 ;
  assign n1463 = n1459 | n1462 ;
  assign n1464 = n228 & n1463 ;
  assign n1465 = ~n145 & n877 ;
  assign n1466 = n156 & n759 ;
  assign n1467 = n1465 | n1466 ;
  assign n1468 = n168 & n793 ;
  assign n1469 = n179 & n770 ;
  assign n1470 = n1468 | n1469 ;
  assign n1471 = n1467 | n1470 ;
  assign n1472 = n183 & n1471 ;
  assign n1473 = n1464 | n1472 ;
  assign n1474 = n1456 | n1473 ;
  assign n1475 = x134 & n1474 ;
  assign n1476 = n1439 | n1475 ;
  assign n1477 = ~n145 & n928 ;
  assign n1478 = n156 & n899 ;
  assign n1479 = n1477 | n1478 ;
  assign n1480 = n168 & n912 ;
  assign n1481 = n179 & n903 ;
  assign n1482 = n1480 | n1481 ;
  assign n1483 = n1479 | n1482 ;
  assign n1484 = n183 & n1483 ;
  assign n1485 = ~n145 & n969 ;
  assign n1486 = n156 & n919 ;
  assign n1487 = n1485 | n1486 ;
  assign n1488 = n168 & n932 ;
  assign n1489 = n179 & n923 ;
  assign n1490 = n1488 | n1489 ;
  assign n1491 = n1487 | n1490 ;
  assign n1492 = n228 & n1491 ;
  assign n1493 = n1484 | n1492 ;
  assign n1494 = ~n145 & n1012 ;
  assign n1495 = n156 & n940 ;
  assign n1496 = n1494 | n1495 ;
  assign n1497 = n168 & n953 ;
  assign n1498 = n179 & n944 ;
  assign n1499 = n1497 | n1498 ;
  assign n1500 = n1496 | n1499 ;
  assign n1501 = ~n274 & n1500 ;
  assign n1502 = ~n145 & n949 ;
  assign n1503 = n156 & n960 ;
  assign n1504 = n1502 | n1503 ;
  assign n1505 = n168 & n973 ;
  assign n1506 = n179 & n964 ;
  assign n1507 = n1505 | n1506 ;
  assign n1508 = n1504 | n1507 ;
  assign n1509 = n319 & n1508 ;
  assign n1510 = n1501 | n1509 ;
  assign n1511 = n1493 | n1510 ;
  assign n1512 = ~x134 & n1511 ;
  assign n1513 = ~n145 & n992 ;
  assign n1514 = n156 & n1024 ;
  assign n1515 = n1513 | n1514 ;
  assign n1516 = n168 & n1039 ;
  assign n1517 = n179 & n1028 ;
  assign n1518 = n1516 | n1517 ;
  assign n1519 = n1515 | n1518 ;
  assign n1520 = n319 & n1519 ;
  assign n1521 = ~n145 & n908 ;
  assign n1522 = n156 & n983 ;
  assign n1523 = n1521 | n1522 ;
  assign n1524 = n168 & n996 ;
  assign n1525 = n179 & n987 ;
  assign n1526 = n1524 | n1525 ;
  assign n1527 = n1523 | n1526 ;
  assign n1528 = ~n274 & n1527 ;
  assign n1529 = n1520 | n1528 ;
  assign n1530 = ~n145 & n1034 ;
  assign n1531 = n156 & n1046 ;
  assign n1532 = n1530 | n1531 ;
  assign n1533 = n168 & n1059 ;
  assign n1534 = n179 & n1050 ;
  assign n1535 = n1533 | n1534 ;
  assign n1536 = n1532 | n1535 ;
  assign n1537 = n228 & n1536 ;
  assign n1538 = ~n145 & n1055 ;
  assign n1539 = n156 & n1003 ;
  assign n1540 = n1538 | n1539 ;
  assign n1541 = n168 & n1016 ;
  assign n1542 = n179 & n1007 ;
  assign n1543 = n1541 | n1542 ;
  assign n1544 = n1540 | n1543 ;
  assign n1545 = n183 & n1544 ;
  assign n1546 = n1537 | n1545 ;
  assign n1547 = n1529 | n1546 ;
  assign n1548 = x134 & n1547 ;
  assign n1549 = n1512 | n1548 ;
  assign n1550 = ~n145 & n1120 ;
  assign n1551 = n156 & n1170 ;
  assign n1552 = n1550 | n1551 ;
  assign n1553 = n168 & n1192 ;
  assign n1554 = n179 & n1177 ;
  assign n1555 = n1553 | n1554 ;
  assign n1556 = n1552 | n1555 ;
  assign n1557 = n183 & n1556 ;
  assign n1558 = ~n145 & n1088 ;
  assign n1559 = n156 & n1105 ;
  assign n1560 = n1558 | n1559 ;
  assign n1561 = n168 & n1127 ;
  assign n1562 = n179 & n1112 ;
  assign n1563 = n1561 | n1562 ;
  assign n1564 = n1560 | n1563 ;
  assign n1565 = n228 & n1564 ;
  assign n1566 = n1557 | n1565 ;
  assign n1567 = ~n145 & n1283 ;
  assign n1568 = n156 & n1138 ;
  assign n1569 = n1567 | n1568 ;
  assign n1570 = n168 & n1160 ;
  assign n1571 = n179 & n1145 ;
  assign n1572 = n1570 | n1571 ;
  assign n1573 = n1569 | n1572 ;
  assign n1574 = ~n274 & n1573 ;
  assign n1575 = ~n145 & n1153 ;
  assign n1576 = n156 & n1073 ;
  assign n1577 = n1575 | n1576 ;
  assign n1578 = n168 & n1095 ;
  assign n1579 = n179 & n1080 ;
  assign n1580 = n1578 | n1579 ;
  assign n1581 = n1577 | n1580 ;
  assign n1582 = n319 & n1581 ;
  assign n1583 = n1574 | n1582 ;
  assign n1584 = n1566 | n1583 ;
  assign n1585 = ~x134 & n1584 ;
  assign n1586 = n156 & n1237 ;
  assign n1587 = n179 & n1242 ;
  assign n1588 = n1586 | n1587 ;
  assign n1589 = n168 & n1257 ;
  assign n1590 = ~n145 & n1220 ;
  assign n1591 = n1589 | n1590 ;
  assign n1592 = n1588 | n1591 ;
  assign n1593 = n319 & n1592 ;
  assign n1594 = ~n145 & n1185 ;
  assign n1595 = n156 & n1205 ;
  assign n1596 = n1594 | n1595 ;
  assign n1597 = n168 & n1227 ;
  assign n1598 = n179 & n1212 ;
  assign n1599 = n1597 | n1598 ;
  assign n1600 = n1596 | n1599 ;
  assign n1601 = ~n274 & n1600 ;
  assign n1602 = n1593 | n1601 ;
  assign n1603 = ~n145 & n1250 ;
  assign n1604 = n156 & n1300 ;
  assign n1605 = n1603 | n1604 ;
  assign n1606 = n168 & n1322 ;
  assign n1607 = n179 & n1307 ;
  assign n1608 = n1606 | n1607 ;
  assign n1609 = n1605 | n1608 ;
  assign n1610 = n228 & n1609 ;
  assign n1611 = ~n145 & n1315 ;
  assign n1612 = n156 & n1268 ;
  assign n1613 = n1611 | n1612 ;
  assign n1614 = n168 & n1290 ;
  assign n1615 = n179 & n1275 ;
  assign n1616 = n1614 | n1615 ;
  assign n1617 = n1613 | n1616 ;
  assign n1618 = n183 & n1617 ;
  assign n1619 = n1610 | n1618 ;
  assign n1620 = n1602 | n1619 ;
  assign n1621 = x134 & n1620 ;
  assign n1622 = n1585 | n1621 ;
  assign n1623 = ~n145 & n224 ;
  assign n1624 = n156 & n214 ;
  assign n1625 = n1623 | n1624 ;
  assign n1626 = n155 & n168 ;
  assign n1627 = n144 & n179 ;
  assign n1628 = n1626 | n1627 ;
  assign n1629 = n1625 | n1628 ;
  assign n1630 = n183 & n1629 ;
  assign n1631 = ~n145 & n315 ;
  assign n1632 = n156 & n305 ;
  assign n1633 = n1631 | n1632 ;
  assign n1634 = n168 & n203 ;
  assign n1635 = n179 & n193 ;
  assign n1636 = n1634 | n1635 ;
  assign n1637 = n1633 | n1636 ;
  assign n1638 = n228 & n1637 ;
  assign n1639 = n1630 | n1638 ;
  assign n1640 = ~n145 & n363 ;
  assign n1641 = n156 & n353 ;
  assign n1642 = n1640 | n1641 ;
  assign n1643 = n168 & n249 ;
  assign n1644 = n179 & n239 ;
  assign n1645 = n1643 | n1644 ;
  assign n1646 = n1642 | n1645 ;
  assign n1647 = ~n274 & n1646 ;
  assign n1648 = ~n145 & n270 ;
  assign n1649 = n156 & n260 ;
  assign n1650 = n1648 | n1649 ;
  assign n1651 = n168 & n294 ;
  assign n1652 = n179 & n284 ;
  assign n1653 = n1651 | n1652 ;
  assign n1654 = n1650 | n1653 ;
  assign n1655 = n319 & n1654 ;
  assign n1656 = n1647 | n1655 ;
  assign n1657 = n1639 | n1656 ;
  assign n1658 = ~x134 & n1657 ;
  assign n1659 = ~n145 & n452 ;
  assign n1660 = n156 & n442 ;
  assign n1661 = n1659 | n1660 ;
  assign n1662 = n168 & n497 ;
  assign n1663 = n179 & n487 ;
  assign n1664 = n1662 | n1663 ;
  assign n1665 = n1661 | n1664 ;
  assign n1666 = n319 & n1665 ;
  assign n1667 = ~n145 & n178 ;
  assign n1668 = n156 & n167 ;
  assign n1669 = n1667 | n1668 ;
  assign n1670 = n168 & n431 ;
  assign n1671 = n179 & n421 ;
  assign n1672 = n1670 | n1671 ;
  assign n1673 = n1669 | n1672 ;
  assign n1674 = ~n274 & n1673 ;
  assign n1675 = n1666 | n1674 ;
  assign n1676 = ~n145 & n407 ;
  assign n1677 = n156 & n397 ;
  assign n1678 = n1676 | n1677 ;
  assign n1679 = n168 & n342 ;
  assign n1680 = n179 & n332 ;
  assign n1681 = n1679 | n1680 ;
  assign n1682 = n1678 | n1681 ;
  assign n1683 = n183 & n1682 ;
  assign n1684 = ~n145 & n476 ;
  assign n1685 = n156 & n465 ;
  assign n1686 = n1684 | n1685 ;
  assign n1687 = n168 & n386 ;
  assign n1688 = n179 & n376 ;
  assign n1689 = n1687 | n1688 ;
  assign n1690 = n228 & n1689 ;
  assign n1691 = ( n228 & n1686 ) | ( n228 & n1690 ) | ( n1686 & n1690 ) ;
  assign n1692 = n1683 | n1691 ;
  assign n1693 = n1675 | n1692 ;
  assign n1694 = x134 & n1693 ;
  assign n1695 = n1658 | n1694 ;
  assign n1696 = ~n145 & n597 ;
  assign n1697 = n156 & n586 ;
  assign n1698 = n1696 | n1697 ;
  assign n1699 = n168 & n526 ;
  assign n1700 = n179 & n515 ;
  assign n1701 = n1699 | n1700 ;
  assign n1702 = n1698 | n1701 ;
  assign n1703 = n183 & n1702 ;
  assign n1704 = ~n145 & n694 ;
  assign n1705 = n156 & n683 ;
  assign n1706 = n1704 | n1705 ;
  assign n1707 = n168 & n574 ;
  assign n1708 = n179 & n563 ;
  assign n1709 = n1707 | n1708 ;
  assign n1710 = n1706 | n1709 ;
  assign n1711 = n228 & n1710 ;
  assign n1712 = n1703 | n1711 ;
  assign n1713 = ~n145 & n793 ;
  assign n1714 = n156 & n782 ;
  assign n1715 = n1713 | n1714 ;
  assign n1716 = n168 & n623 ;
  assign n1717 = n179 & n612 ;
  assign n1718 = n1716 | n1717 ;
  assign n1719 = n1715 | n1718 ;
  assign n1720 = ~n274 & n1719 ;
  assign n1721 = ~n145 & n646 ;
  assign n1722 = n156 & n635 ;
  assign n1723 = n1721 | n1722 ;
  assign n1724 = n168 & n671 ;
  assign n1725 = n179 & n660 ;
  assign n1726 = n1724 | n1725 ;
  assign n1727 = n1723 | n1726 ;
  assign n1728 = n319 & n1727 ;
  assign n1729 = n1720 | n1728 ;
  assign n1730 = n1712 | n1729 ;
  assign n1731 = ~x134 & n1730 ;
  assign n1732 = ~n145 & n745 ;
  assign n1733 = n156 & n734 ;
  assign n1734 = n1732 | n1733 ;
  assign n1735 = n168 & n818 ;
  assign n1736 = n179 & n808 ;
  assign n1737 = n1735 | n1736 ;
  assign n1738 = n1734 | n1737 ;
  assign n1739 = n319 & n1738 ;
  assign n1740 = ~n145 & n549 ;
  assign n1741 = n156 & n538 ;
  assign n1742 = n1740 | n1741 ;
  assign n1743 = n168 & n722 ;
  assign n1744 = n179 & n711 ;
  assign n1745 = n1743 | n1744 ;
  assign n1746 = n1742 | n1745 ;
  assign n1747 = ~n274 & n1746 ;
  assign n1748 = n1739 | n1747 ;
  assign n1749 = ~n145 & n840 ;
  assign n1750 = n156 & n830 ;
  assign n1751 = n1749 | n1750 ;
  assign n1752 = n168 & n865 ;
  assign n1753 = n179 & n854 ;
  assign n1754 = n1752 | n1753 ;
  assign n1755 = n1751 | n1754 ;
  assign n1756 = n228 & n1755 ;
  assign n1757 = ~n145 & n888 ;
  assign n1758 = n156 & n877 ;
  assign n1759 = n1757 | n1758 ;
  assign n1760 = n168 & n770 ;
  assign n1761 = n179 & n759 ;
  assign n1762 = n1760 | n1761 ;
  assign n1763 = n1759 | n1762 ;
  assign n1764 = n183 & n1763 ;
  assign n1765 = n1756 | n1764 ;
  assign n1766 = n1748 | n1765 ;
  assign n1767 = x134 & n1766 ;
  assign n1768 = n1731 | n1767 ;
  assign n1769 = ~n145 & n932 ;
  assign n1770 = n156 & n928 ;
  assign n1771 = n1769 | n1770 ;
  assign n1772 = n168 & n903 ;
  assign n1773 = n179 & n899 ;
  assign n1774 = n1772 | n1773 ;
  assign n1775 = n1771 | n1774 ;
  assign n1776 = n183 & n1775 ;
  assign n1777 = ~n145 & n973 ;
  assign n1778 = n156 & n969 ;
  assign n1779 = n1777 | n1778 ;
  assign n1780 = n168 & n923 ;
  assign n1781 = n179 & n919 ;
  assign n1782 = n1780 | n1781 ;
  assign n1783 = n1779 | n1782 ;
  assign n1784 = n228 & n1783 ;
  assign n1785 = n1776 | n1784 ;
  assign n1786 = ~n145 & n1016 ;
  assign n1787 = n156 & n1012 ;
  assign n1788 = n1786 | n1787 ;
  assign n1789 = n168 & n944 ;
  assign n1790 = n179 & n940 ;
  assign n1791 = n1789 | n1790 ;
  assign n1792 = n1788 | n1791 ;
  assign n1793 = ~n274 & n1792 ;
  assign n1794 = ~n145 & n953 ;
  assign n1795 = n156 & n949 ;
  assign n1796 = n1794 | n1795 ;
  assign n1797 = n168 & n964 ;
  assign n1798 = n179 & n960 ;
  assign n1799 = n1797 | n1798 ;
  assign n1800 = n1796 | n1799 ;
  assign n1801 = n319 & n1800 ;
  assign n1802 = n1793 | n1801 ;
  assign n1803 = n1785 | n1802 ;
  assign n1804 = ~x134 & n1803 ;
  assign n1805 = ~n145 & n996 ;
  assign n1806 = n156 & n992 ;
  assign n1807 = n1805 | n1806 ;
  assign n1808 = n168 & n1028 ;
  assign n1809 = n179 & n1024 ;
  assign n1810 = n1808 | n1809 ;
  assign n1811 = n1807 | n1810 ;
  assign n1812 = n319 & n1811 ;
  assign n1813 = ~n145 & n912 ;
  assign n1814 = n156 & n908 ;
  assign n1815 = n1813 | n1814 ;
  assign n1816 = n168 & n987 ;
  assign n1817 = n179 & n983 ;
  assign n1818 = n1816 | n1817 ;
  assign n1819 = n1815 | n1818 ;
  assign n1820 = ~n274 & n1819 ;
  assign n1821 = n1812 | n1820 ;
  assign n1822 = ~n145 & n1039 ;
  assign n1823 = n156 & n1034 ;
  assign n1824 = n1822 | n1823 ;
  assign n1825 = n168 & n1050 ;
  assign n1826 = n179 & n1046 ;
  assign n1827 = n1825 | n1826 ;
  assign n1828 = n1824 | n1827 ;
  assign n1829 = n228 & n1828 ;
  assign n1830 = ~n145 & n1059 ;
  assign n1831 = n156 & n1055 ;
  assign n1832 = n1830 | n1831 ;
  assign n1833 = n168 & n1007 ;
  assign n1834 = n179 & n1003 ;
  assign n1835 = n1833 | n1834 ;
  assign n1836 = n1832 | n1835 ;
  assign n1837 = n183 & n1836 ;
  assign n1838 = n1829 | n1837 ;
  assign n1839 = n1821 | n1838 ;
  assign n1840 = x134 & n1839 ;
  assign n1841 = n1804 | n1840 ;
  assign n1842 = ~n145 & n1127 ;
  assign n1843 = n156 & n1120 ;
  assign n1844 = n1842 | n1843 ;
  assign n1845 = n168 & n1177 ;
  assign n1846 = n179 & n1170 ;
  assign n1847 = n1845 | n1846 ;
  assign n1848 = n1844 | n1847 ;
  assign n1849 = n183 & n1848 ;
  assign n1850 = ~n145 & n1095 ;
  assign n1851 = n156 & n1088 ;
  assign n1852 = n1850 | n1851 ;
  assign n1853 = n168 & n1112 ;
  assign n1854 = n179 & n1105 ;
  assign n1855 = n1853 | n1854 ;
  assign n1856 = n1852 | n1855 ;
  assign n1857 = n228 & n1856 ;
  assign n1858 = n1849 | n1857 ;
  assign n1859 = ~n145 & n1290 ;
  assign n1860 = n156 & n1283 ;
  assign n1861 = n1859 | n1860 ;
  assign n1862 = n168 & n1145 ;
  assign n1863 = n179 & n1138 ;
  assign n1864 = n1862 | n1863 ;
  assign n1865 = n1861 | n1864 ;
  assign n1866 = ~n274 & n1865 ;
  assign n1867 = ~n145 & n1160 ;
  assign n1868 = n156 & n1153 ;
  assign n1869 = n1867 | n1868 ;
  assign n1870 = n168 & n1080 ;
  assign n1871 = n179 & n1073 ;
  assign n1872 = n1870 | n1871 ;
  assign n1873 = n1869 | n1872 ;
  assign n1874 = n319 & n1873 ;
  assign n1875 = n1866 | n1874 ;
  assign n1876 = n1858 | n1875 ;
  assign n1877 = ~x134 & n1876 ;
  assign n1878 = ~n145 & n1227 ;
  assign n1879 = n179 & n1237 ;
  assign n1880 = n1878 | n1879 ;
  assign n1881 = n168 & n1242 ;
  assign n1882 = n156 & n1220 ;
  assign n1883 = n1881 | n1882 ;
  assign n1884 = n1880 | n1883 ;
  assign n1885 = n319 & n1884 ;
  assign n1886 = ~n145 & n1192 ;
  assign n1887 = n156 & n1185 ;
  assign n1888 = n1886 | n1887 ;
  assign n1889 = n168 & n1212 ;
  assign n1890 = n179 & n1205 ;
  assign n1891 = n1889 | n1890 ;
  assign n1892 = n1888 | n1891 ;
  assign n1893 = ~n274 & n1892 ;
  assign n1894 = n1885 | n1893 ;
  assign n1895 = ~n145 & n1257 ;
  assign n1896 = n156 & n1250 ;
  assign n1897 = n1895 | n1896 ;
  assign n1898 = n168 & n1307 ;
  assign n1899 = n179 & n1300 ;
  assign n1900 = n1898 | n1899 ;
  assign n1901 = n1897 | n1900 ;
  assign n1902 = n228 & n1901 ;
  assign n1903 = ~n145 & n1322 ;
  assign n1904 = n156 & n1315 ;
  assign n1905 = n1903 | n1904 ;
  assign n1906 = n168 & n1275 ;
  assign n1907 = n179 & n1268 ;
  assign n1908 = n1906 | n1907 ;
  assign n1909 = n1905 | n1908 ;
  assign n1910 = n183 & n1909 ;
  assign n1911 = n1902 | n1910 ;
  assign n1912 = n1894 | n1911 ;
  assign n1913 = x134 & n1912 ;
  assign n1914 = n1877 | n1913 ;
  assign n1915 = ~n145 & n203 ;
  assign n1916 = n156 & n224 ;
  assign n1917 = n1915 | n1916 ;
  assign n1918 = n144 & n168 ;
  assign n1919 = n179 & n214 ;
  assign n1920 = n1918 | n1919 ;
  assign n1921 = n1917 | n1920 ;
  assign n1922 = n183 & n1921 ;
  assign n1923 = ~n145 & n294 ;
  assign n1924 = n156 & n315 ;
  assign n1925 = n1923 | n1924 ;
  assign n1926 = n168 & n193 ;
  assign n1927 = n179 & n305 ;
  assign n1928 = n1926 | n1927 ;
  assign n1929 = n1925 | n1928 ;
  assign n1930 = n228 & n1929 ;
  assign n1931 = n1922 | n1930 ;
  assign n1932 = ~n145 & n342 ;
  assign n1933 = n156 & n363 ;
  assign n1934 = n1932 | n1933 ;
  assign n1935 = n168 & n239 ;
  assign n1936 = n179 & n353 ;
  assign n1937 = n1935 | n1936 ;
  assign n1938 = n1934 | n1937 ;
  assign n1939 = ~n274 & n1938 ;
  assign n1940 = ~n145 & n249 ;
  assign n1941 = n156 & n270 ;
  assign n1942 = n1940 | n1941 ;
  assign n1943 = n168 & n284 ;
  assign n1944 = n179 & n260 ;
  assign n1945 = n1943 | n1944 ;
  assign n1946 = n1942 | n1945 ;
  assign n1947 = n319 & n1946 ;
  assign n1948 = n1939 | n1947 ;
  assign n1949 = n1931 | n1948 ;
  assign n1950 = ~x134 & n1949 ;
  assign n1951 = ~n145 & n431 ;
  assign n1952 = n156 & n452 ;
  assign n1953 = n1951 | n1952 ;
  assign n1954 = n168 & n487 ;
  assign n1955 = n179 & n442 ;
  assign n1956 = n1954 | n1955 ;
  assign n1957 = n1953 | n1956 ;
  assign n1958 = n319 & n1957 ;
  assign n1959 = ~n145 & n155 ;
  assign n1960 = n156 & n178 ;
  assign n1961 = n1959 | n1960 ;
  assign n1962 = n168 & n421 ;
  assign n1963 = n167 & n179 ;
  assign n1964 = n1962 | n1963 ;
  assign n1965 = n1961 | n1964 ;
  assign n1966 = ~n274 & n1965 ;
  assign n1967 = n1958 | n1966 ;
  assign n1968 = ~n145 & n386 ;
  assign n1969 = n156 & n407 ;
  assign n1970 = n1968 | n1969 ;
  assign n1971 = n168 & n332 ;
  assign n1972 = n179 & n397 ;
  assign n1973 = n1971 | n1972 ;
  assign n1974 = n1970 | n1973 ;
  assign n1975 = n183 & n1974 ;
  assign n1976 = ~n145 & n497 ;
  assign n1977 = n156 & n476 ;
  assign n1978 = n1976 | n1977 ;
  assign n1979 = n168 & n376 ;
  assign n1980 = n179 & n465 ;
  assign n1981 = n1979 | n1980 ;
  assign n1982 = n228 & n1981 ;
  assign n1983 = ( n228 & n1978 ) | ( n228 & n1982 ) | ( n1978 & n1982 ) ;
  assign n1984 = n1975 | n1983 ;
  assign n1985 = n1967 | n1984 ;
  assign n1986 = x134 & n1985 ;
  assign n1987 = n1950 | n1986 ;
  assign n1988 = ~n145 & n574 ;
  assign n1989 = n156 & n597 ;
  assign n1990 = n1988 | n1989 ;
  assign n1991 = n168 & n515 ;
  assign n1992 = n179 & n586 ;
  assign n1993 = n1991 | n1992 ;
  assign n1994 = n1990 | n1993 ;
  assign n1995 = n183 & n1994 ;
  assign n1996 = ~n145 & n671 ;
  assign n1997 = n156 & n694 ;
  assign n1998 = n1996 | n1997 ;
  assign n1999 = n168 & n563 ;
  assign n2000 = n179 & n683 ;
  assign n2001 = n1999 | n2000 ;
  assign n2002 = n1998 | n2001 ;
  assign n2003 = n228 & n2002 ;
  assign n2004 = n1995 | n2003 ;
  assign n2005 = ~n145 & n770 ;
  assign n2006 = n156 & n793 ;
  assign n2007 = n2005 | n2006 ;
  assign n2008 = n168 & n612 ;
  assign n2009 = n179 & n782 ;
  assign n2010 = n2008 | n2009 ;
  assign n2011 = n2007 | n2010 ;
  assign n2012 = ~n274 & n2011 ;
  assign n2013 = ~n145 & n623 ;
  assign n2014 = n156 & n646 ;
  assign n2015 = n2013 | n2014 ;
  assign n2016 = n168 & n660 ;
  assign n2017 = n179 & n635 ;
  assign n2018 = n2016 | n2017 ;
  assign n2019 = n2015 | n2018 ;
  assign n2020 = n319 & n2019 ;
  assign n2021 = n2012 | n2020 ;
  assign n2022 = n2004 | n2021 ;
  assign n2023 = ~x134 & n2022 ;
  assign n2024 = ~n145 & n722 ;
  assign n2025 = n156 & n745 ;
  assign n2026 = n2024 | n2025 ;
  assign n2027 = n168 & n808 ;
  assign n2028 = n179 & n734 ;
  assign n2029 = n2027 | n2028 ;
  assign n2030 = n2026 | n2029 ;
  assign n2031 = n319 & n2030 ;
  assign n2032 = ~n145 & n526 ;
  assign n2033 = n156 & n549 ;
  assign n2034 = n2032 | n2033 ;
  assign n2035 = n168 & n711 ;
  assign n2036 = n179 & n538 ;
  assign n2037 = n2035 | n2036 ;
  assign n2038 = n2034 | n2037 ;
  assign n2039 = ~n274 & n2038 ;
  assign n2040 = n2031 | n2039 ;
  assign n2041 = ~n145 & n865 ;
  assign n2042 = n156 & n888 ;
  assign n2043 = n2041 | n2042 ;
  assign n2044 = n168 & n759 ;
  assign n2045 = n179 & n877 ;
  assign n2046 = n2044 | n2045 ;
  assign n2047 = n2043 | n2046 ;
  assign n2048 = n183 & n2047 ;
  assign n2049 = n168 & n854 ;
  assign n2050 = n179 & n830 ;
  assign n2051 = n2049 | n2050 ;
  assign n2052 = ~n145 & n818 ;
  assign n2053 = n156 & n840 ;
  assign n2054 = n2052 | n2053 ;
  assign n2055 = n228 & n2054 ;
  assign n2056 = ( n228 & n2051 ) | ( n228 & n2055 ) | ( n2051 & n2055 ) ;
  assign n2057 = n2048 | n2056 ;
  assign n2058 = n2040 | n2057 ;
  assign n2059 = x134 & n2058 ;
  assign n2060 = n2023 | n2059 ;
  assign n2061 = ~n145 & n923 ;
  assign n2062 = n156 & n932 ;
  assign n2063 = n2061 | n2062 ;
  assign n2064 = n168 & n899 ;
  assign n2065 = n179 & n928 ;
  assign n2066 = n2064 | n2065 ;
  assign n2067 = n2063 | n2066 ;
  assign n2068 = n183 & n2067 ;
  assign n2069 = ~n145 & n964 ;
  assign n2070 = n156 & n973 ;
  assign n2071 = n2069 | n2070 ;
  assign n2072 = n168 & n919 ;
  assign n2073 = n179 & n969 ;
  assign n2074 = n2072 | n2073 ;
  assign n2075 = n2071 | n2074 ;
  assign n2076 = n228 & n2075 ;
  assign n2077 = n2068 | n2076 ;
  assign n2078 = ~n145 & n1007 ;
  assign n2079 = n156 & n1016 ;
  assign n2080 = n2078 | n2079 ;
  assign n2081 = n168 & n940 ;
  assign n2082 = n179 & n1012 ;
  assign n2083 = n2081 | n2082 ;
  assign n2084 = n2080 | n2083 ;
  assign n2085 = ~n274 & n2084 ;
  assign n2086 = ~n145 & n944 ;
  assign n2087 = n156 & n953 ;
  assign n2088 = n2086 | n2087 ;
  assign n2089 = n168 & n960 ;
  assign n2090 = n179 & n949 ;
  assign n2091 = n2089 | n2090 ;
  assign n2092 = n2088 | n2091 ;
  assign n2093 = n319 & n2092 ;
  assign n2094 = n2085 | n2093 ;
  assign n2095 = n2077 | n2094 ;
  assign n2096 = ~x134 & n2095 ;
  assign n2097 = ~n145 & n987 ;
  assign n2098 = n156 & n996 ;
  assign n2099 = n2097 | n2098 ;
  assign n2100 = n168 & n1024 ;
  assign n2101 = n179 & n992 ;
  assign n2102 = n2100 | n2101 ;
  assign n2103 = n2099 | n2102 ;
  assign n2104 = n319 & n2103 ;
  assign n2105 = ~n145 & n903 ;
  assign n2106 = n156 & n912 ;
  assign n2107 = n2105 | n2106 ;
  assign n2108 = n168 & n983 ;
  assign n2109 = n179 & n908 ;
  assign n2110 = n2108 | n2109 ;
  assign n2111 = n2107 | n2110 ;
  assign n2112 = ~n274 & n2111 ;
  assign n2113 = n2104 | n2112 ;
  assign n2114 = ~n145 & n1028 ;
  assign n2115 = n156 & n1039 ;
  assign n2116 = n2114 | n2115 ;
  assign n2117 = n168 & n1046 ;
  assign n2118 = n179 & n1034 ;
  assign n2119 = n2117 | n2118 ;
  assign n2120 = n2116 | n2119 ;
  assign n2121 = n228 & n2120 ;
  assign n2122 = ~n145 & n1050 ;
  assign n2123 = n156 & n1059 ;
  assign n2124 = n2122 | n2123 ;
  assign n2125 = n168 & n1003 ;
  assign n2126 = n179 & n1055 ;
  assign n2127 = n2125 | n2126 ;
  assign n2128 = n2124 | n2127 ;
  assign n2129 = n183 & n2128 ;
  assign n2130 = n2121 | n2129 ;
  assign n2131 = n2113 | n2130 ;
  assign n2132 = x134 & n2131 ;
  assign n2133 = n2096 | n2132 ;
  assign n2134 = ~n145 & n1112 ;
  assign n2135 = n156 & n1127 ;
  assign n2136 = n2134 | n2135 ;
  assign n2137 = n168 & n1170 ;
  assign n2138 = n179 & n1120 ;
  assign n2139 = n2137 | n2138 ;
  assign n2140 = n2136 | n2139 ;
  assign n2141 = n183 & n2140 ;
  assign n2142 = ~n145 & n1080 ;
  assign n2143 = n156 & n1095 ;
  assign n2144 = n2142 | n2143 ;
  assign n2145 = n168 & n1105 ;
  assign n2146 = n179 & n1088 ;
  assign n2147 = n2145 | n2146 ;
  assign n2148 = n2144 | n2147 ;
  assign n2149 = n228 & n2148 ;
  assign n2150 = n2141 | n2149 ;
  assign n2151 = ~n145 & n1275 ;
  assign n2152 = n156 & n1290 ;
  assign n2153 = n2151 | n2152 ;
  assign n2154 = n168 & n1138 ;
  assign n2155 = n179 & n1283 ;
  assign n2156 = n2154 | n2155 ;
  assign n2157 = n2153 | n2156 ;
  assign n2158 = ~n274 & n2157 ;
  assign n2159 = ~n145 & n1145 ;
  assign n2160 = n156 & n1160 ;
  assign n2161 = n2159 | n2160 ;
  assign n2162 = n168 & n1073 ;
  assign n2163 = n179 & n1153 ;
  assign n2164 = n2162 | n2163 ;
  assign n2165 = n2161 | n2164 ;
  assign n2166 = n319 & n2165 ;
  assign n2167 = n2158 | n2166 ;
  assign n2168 = n2150 | n2167 ;
  assign n2169 = ~x134 & n2168 ;
  assign n2170 = ~n145 & n1212 ;
  assign n2171 = n156 & n1227 ;
  assign n2172 = n2170 | n2171 ;
  assign n2173 = n168 & n1237 ;
  assign n2174 = n179 & n1220 ;
  assign n2175 = n2173 | n2174 ;
  assign n2176 = n2172 | n2175 ;
  assign n2177 = n319 & n2176 ;
  assign n2178 = ~n145 & n1177 ;
  assign n2179 = n156 & n1192 ;
  assign n2180 = n2178 | n2179 ;
  assign n2181 = n168 & n1205 ;
  assign n2182 = n179 & n1185 ;
  assign n2183 = n2181 | n2182 ;
  assign n2184 = n2180 | n2183 ;
  assign n2185 = ~n274 & n2184 ;
  assign n2186 = n2177 | n2185 ;
  assign n2187 = ~n145 & n1242 ;
  assign n2188 = n156 & n1257 ;
  assign n2189 = n2187 | n2188 ;
  assign n2190 = n168 & n1300 ;
  assign n2191 = n179 & n1250 ;
  assign n2192 = n2190 | n2191 ;
  assign n2193 = n2189 | n2192 ;
  assign n2194 = n228 & n2193 ;
  assign n2195 = ~n145 & n1307 ;
  assign n2196 = n156 & n1322 ;
  assign n2197 = n2195 | n2196 ;
  assign n2198 = n168 & n1268 ;
  assign n2199 = n179 & n1315 ;
  assign n2200 = n2198 | n2199 ;
  assign n2201 = n2197 | n2200 ;
  assign n2202 = n183 & n2201 ;
  assign n2203 = n2194 | n2202 ;
  assign n2204 = n2186 | n2203 ;
  assign n2205 = x134 & n2204 ;
  assign n2206 = n2169 | n2205 ;
  assign n2207 = n183 & n227 ;
  assign n2208 = n228 & n318 ;
  assign n2209 = n2207 | n2208 ;
  assign n2210 = ~n274 & n366 ;
  assign n2211 = n273 & n319 ;
  assign n2212 = n2210 | n2211 ;
  assign n2213 = n2209 | n2212 ;
  assign n2214 = ~x134 & n2213 ;
  assign n2215 = n182 & ~n274 ;
  assign n2216 = n183 & n410 ;
  assign n2217 = n2215 | n2216 ;
  assign n2218 = n319 & n455 ;
  assign n2219 = n228 & n499 ;
  assign n2220 = ( n228 & n478 ) | ( n228 & n2219 ) | ( n478 & n2219 ) ;
  assign n2221 = n2218 | n2220 ;
  assign n2222 = n2217 | n2221 ;
  assign n2223 = x134 & n2222 ;
  assign n2224 = n2214 | n2223 ;
  assign n2225 = n183 & n600 ;
  assign n2226 = n228 & n697 ;
  assign n2227 = n2225 | n2226 ;
  assign n2228 = ~n274 & n796 ;
  assign n2229 = n319 & n649 ;
  assign n2230 = n2228 | n2229 ;
  assign n2231 = n2227 | n2230 ;
  assign n2232 = ~x134 & n2231 ;
  assign n2233 = n319 & n748 ;
  assign n2234 = ~n274 & n552 ;
  assign n2235 = n2233 | n2234 ;
  assign n2236 = n228 & n843 ;
  assign n2237 = n183 & n891 ;
  assign n2238 = n2236 | n2237 ;
  assign n2239 = n2235 | n2238 ;
  assign n2240 = x134 & n2239 ;
  assign n2241 = n2232 | n2240 ;
  assign n2242 = n183 & n935 ;
  assign n2243 = n228 & n976 ;
  assign n2244 = n2242 | n2243 ;
  assign n2245 = ~n274 & n1019 ;
  assign n2246 = n319 & n956 ;
  assign n2247 = n2245 | n2246 ;
  assign n2248 = n2244 | n2247 ;
  assign n2249 = ~x134 & n2248 ;
  assign n2250 = n319 & n999 ;
  assign n2251 = ~n274 & n915 ;
  assign n2252 = n2250 | n2251 ;
  assign n2253 = n228 & n1042 ;
  assign n2254 = n183 & n1062 ;
  assign n2255 = n2253 | n2254 ;
  assign n2256 = n2252 | n2255 ;
  assign n2257 = x134 & n2256 ;
  assign n2258 = n2249 | n2257 ;
  assign n2259 = n228 & n1098 ;
  assign n2260 = n183 & n1130 ;
  assign n2261 = n2259 | n2260 ;
  assign n2262 = n319 & n1163 ;
  assign n2263 = ~n274 & n1293 ;
  assign n2264 = n2262 | n2263 ;
  assign n2265 = n2261 | n2264 ;
  assign n2266 = ~x134 & n2265 ;
  assign n2267 = n319 & n1230 ;
  assign n2268 = ~n274 & n1195 ;
  assign n2269 = n2267 | n2268 ;
  assign n2270 = n183 & n1325 ;
  assign n2271 = n228 & n1260 ;
  assign n2272 = n2270 | n2271 ;
  assign n2273 = n2269 | n2272 ;
  assign n2274 = x134 & n2273 ;
  assign n2275 = n2266 | n2274 ;
  assign n2276 = n183 & n1345 ;
  assign n2277 = n228 & n1362 ;
  assign n2278 = n2276 | n2277 ;
  assign n2279 = ~n274 & n1398 ;
  assign n2280 = n319 & n1354 ;
  assign n2281 = n2279 | n2280 ;
  assign n2282 = n2278 | n2281 ;
  assign n2283 = ~x134 & n2282 ;
  assign n2284 = ~n274 & n1337 ;
  assign n2285 = n228 & n1380 ;
  assign n2286 = ( n228 & n1377 ) | ( n228 & n2285 ) | ( n1377 & n2285 ) ;
  assign n2287 = n2284 | n2286 ;
  assign n2288 = n183 & n1390 ;
  assign n2289 = n319 & n1373 ;
  assign n2290 = n2288 | n2289 ;
  assign n2291 = n2287 | n2290 ;
  assign n2292 = x134 & n2291 ;
  assign n2293 = n2283 | n2292 ;
  assign n2294 = n183 & n1418 ;
  assign n2295 = n228 & n1435 ;
  assign n2296 = n2294 | n2295 ;
  assign n2297 = ~n274 & n1471 ;
  assign n2298 = n319 & n1427 ;
  assign n2299 = n2297 | n2298 ;
  assign n2300 = n2296 | n2299 ;
  assign n2301 = ~x134 & n2300 ;
  assign n2302 = ~n274 & n1410 ;
  assign n2303 = n228 & n1453 ;
  assign n2304 = ( n228 & n1450 ) | ( n228 & n2303 ) | ( n1450 & n2303 ) ;
  assign n2305 = n2302 | n2304 ;
  assign n2306 = n183 & n1463 ;
  assign n2307 = n319 & n1446 ;
  assign n2308 = n2306 | n2307 ;
  assign n2309 = n2305 | n2308 ;
  assign n2310 = x134 & n2309 ;
  assign n2311 = n2301 | n2310 ;
  assign n2312 = n183 & n1491 ;
  assign n2313 = n228 & n1508 ;
  assign n2314 = n2312 | n2313 ;
  assign n2315 = ~n274 & n1544 ;
  assign n2316 = n319 & n1500 ;
  assign n2317 = n2315 | n2316 ;
  assign n2318 = n2314 | n2317 ;
  assign n2319 = ~x134 & n2318 ;
  assign n2320 = ~n274 & n1483 ;
  assign n2321 = n228 & n1519 ;
  assign n2322 = n2320 | n2321 ;
  assign n2323 = n183 & n1536 ;
  assign n2324 = n319 & n1527 ;
  assign n2325 = n2323 | n2324 ;
  assign n2326 = n2322 | n2325 ;
  assign n2327 = x134 & n2326 ;
  assign n2328 = n2319 | n2327 ;
  assign n2329 = n183 & n1564 ;
  assign n2330 = ~n274 & n1617 ;
  assign n2331 = n2329 | n2330 ;
  assign n2332 = n319 & n1573 ;
  assign n2333 = n228 & n1581 ;
  assign n2334 = n2332 | n2333 ;
  assign n2335 = n2331 | n2334 ;
  assign n2336 = ~x134 & n2335 ;
  assign n2337 = n228 & n1592 ;
  assign n2338 = n319 & n1600 ;
  assign n2339 = n2337 | n2338 ;
  assign n2340 = n183 & n1609 ;
  assign n2341 = ~n274 & n1556 ;
  assign n2342 = n2340 | n2341 ;
  assign n2343 = n2339 | n2342 ;
  assign n2344 = x134 & n2343 ;
  assign n2345 = n2336 | n2344 ;
  assign n2346 = n183 & n1637 ;
  assign n2347 = ~n274 & n1682 ;
  assign n2348 = n2346 | n2347 ;
  assign n2349 = n319 & n1646 ;
  assign n2350 = n228 & n1654 ;
  assign n2351 = n2349 | n2350 ;
  assign n2352 = n2348 | n2351 ;
  assign n2353 = ~x134 & n2352 ;
  assign n2354 = n228 & n1665 ;
  assign n2355 = n319 & n1673 ;
  assign n2356 = n2354 | n2355 ;
  assign n2357 = ~n274 & n1629 ;
  assign n2358 = n183 & n1689 ;
  assign n2359 = ( n183 & n1686 ) | ( n183 & n2358 ) | ( n1686 & n2358 ) ;
  assign n2360 = n2357 | n2359 ;
  assign n2361 = n2356 | n2360 ;
  assign n2362 = x134 & n2361 ;
  assign n2363 = n2353 | n2362 ;
  assign n2364 = n183 & n1710 ;
  assign n2365 = ~n274 & n1763 ;
  assign n2366 = n2364 | n2365 ;
  assign n2367 = n319 & n1719 ;
  assign n2368 = n228 & n1727 ;
  assign n2369 = n2367 | n2368 ;
  assign n2370 = n2366 | n2369 ;
  assign n2371 = ~x134 & n2370 ;
  assign n2372 = n228 & n1738 ;
  assign n2373 = n319 & n1746 ;
  assign n2374 = n2372 | n2373 ;
  assign n2375 = n183 & n1755 ;
  assign n2376 = ~n274 & n1702 ;
  assign n2377 = n2375 | n2376 ;
  assign n2378 = n2374 | n2377 ;
  assign n2379 = x134 & n2378 ;
  assign n2380 = n2371 | n2379 ;
  assign n2381 = n183 & n1783 ;
  assign n2382 = n228 & n1800 ;
  assign n2383 = n2381 | n2382 ;
  assign n2384 = ~n274 & n1836 ;
  assign n2385 = n319 & n1792 ;
  assign n2386 = n2384 | n2385 ;
  assign n2387 = n2383 | n2386 ;
  assign n2388 = ~x134 & n2387 ;
  assign n2389 = n228 & n1811 ;
  assign n2390 = n319 & n1819 ;
  assign n2391 = n2389 | n2390 ;
  assign n2392 = n183 & n1828 ;
  assign n2393 = ~n274 & n1775 ;
  assign n2394 = n2392 | n2393 ;
  assign n2395 = n2391 | n2394 ;
  assign n2396 = x134 & n2395 ;
  assign n2397 = n2388 | n2396 ;
  assign n2398 = n183 & n1856 ;
  assign n2399 = n228 & n1873 ;
  assign n2400 = n2398 | n2399 ;
  assign n2401 = ~n274 & n1909 ;
  assign n2402 = n319 & n1865 ;
  assign n2403 = n2401 | n2402 ;
  assign n2404 = n2400 | n2403 ;
  assign n2405 = ~x134 & n2404 ;
  assign n2406 = n228 & n1884 ;
  assign n2407 = n319 & n1892 ;
  assign n2408 = n2406 | n2407 ;
  assign n2409 = n183 & n1901 ;
  assign n2410 = ~n274 & n1848 ;
  assign n2411 = n2409 | n2410 ;
  assign n2412 = n2408 | n2411 ;
  assign n2413 = x134 & n2412 ;
  assign n2414 = n2405 | n2413 ;
  assign n2415 = n183 & n1929 ;
  assign n2416 = n228 & n1946 ;
  assign n2417 = n2415 | n2416 ;
  assign n2418 = ~n274 & n1974 ;
  assign n2419 = n319 & n1938 ;
  assign n2420 = n2418 | n2419 ;
  assign n2421 = n2417 | n2420 ;
  assign n2422 = ~x134 & n2421 ;
  assign n2423 = n228 & n1957 ;
  assign n2424 = n319 & n1965 ;
  assign n2425 = n2423 | n2424 ;
  assign n2426 = ~n274 & n1921 ;
  assign n2427 = n183 & n1981 ;
  assign n2428 = ( n183 & n1978 ) | ( n183 & n2427 ) | ( n1978 & n2427 ) ;
  assign n2429 = n2426 | n2428 ;
  assign n2430 = n2425 | n2429 ;
  assign n2431 = x134 & n2430 ;
  assign n2432 = n2422 | n2431 ;
  assign n2433 = n183 & n2002 ;
  assign n2434 = n228 & n2019 ;
  assign n2435 = n2433 | n2434 ;
  assign n2436 = ~n274 & n2047 ;
  assign n2437 = n319 & n2011 ;
  assign n2438 = n2436 | n2437 ;
  assign n2439 = n2435 | n2438 ;
  assign n2440 = ~x134 & n2439 ;
  assign n2441 = n228 & n2030 ;
  assign n2442 = n319 & n2038 ;
  assign n2443 = n2441 | n2442 ;
  assign n2444 = ~n274 & n1994 ;
  assign n2445 = n183 & n2054 ;
  assign n2446 = ( n183 & n2051 ) | ( n183 & n2445 ) | ( n2051 & n2445 ) ;
  assign n2447 = n2444 | n2446 ;
  assign n2448 = n2443 | n2447 ;
  assign n2449 = x134 & n2448 ;
  assign n2450 = n2440 | n2449 ;
  assign n2451 = n183 & n2075 ;
  assign n2452 = n228 & n2092 ;
  assign n2453 = n2451 | n2452 ;
  assign n2454 = ~n274 & n2128 ;
  assign n2455 = n319 & n2084 ;
  assign n2456 = n2454 | n2455 ;
  assign n2457 = n2453 | n2456 ;
  assign n2458 = ~x134 & n2457 ;
  assign n2459 = n228 & n2103 ;
  assign n2460 = n319 & n2111 ;
  assign n2461 = n2459 | n2460 ;
  assign n2462 = n183 & n2120 ;
  assign n2463 = ~n274 & n2067 ;
  assign n2464 = n2462 | n2463 ;
  assign n2465 = n2461 | n2464 ;
  assign n2466 = x134 & n2465 ;
  assign n2467 = n2458 | n2466 ;
  assign n2468 = n183 & n2148 ;
  assign n2469 = n228 & n2165 ;
  assign n2470 = n2468 | n2469 ;
  assign n2471 = ~n274 & n2201 ;
  assign n2472 = n319 & n2157 ;
  assign n2473 = n2471 | n2472 ;
  assign n2474 = n2470 | n2473 ;
  assign n2475 = ~x134 & n2474 ;
  assign n2476 = n228 & n2176 ;
  assign n2477 = n319 & n2184 ;
  assign n2478 = n2476 | n2477 ;
  assign n2479 = n183 & n2193 ;
  assign n2480 = ~n274 & n2140 ;
  assign n2481 = n2479 | n2480 ;
  assign n2482 = n2478 | n2481 ;
  assign n2483 = x134 & n2482 ;
  assign n2484 = n2475 | n2483 ;
  assign n2485 = n183 & n318 ;
  assign n2486 = n228 & n273 ;
  assign n2487 = n2485 | n2486 ;
  assign n2488 = ~n274 & n410 ;
  assign n2489 = n319 & n366 ;
  assign n2490 = n2488 | n2489 ;
  assign n2491 = n2487 | n2490 ;
  assign n2492 = ~x134 & n2491 ;
  assign n2493 = n182 & n319 ;
  assign n2494 = n227 & ~n274 ;
  assign n2495 = n2493 | n2494 ;
  assign n2496 = n228 & n455 ;
  assign n2497 = n183 & n499 ;
  assign n2498 = ( n183 & n478 ) | ( n183 & n2497 ) | ( n478 & n2497 ) ;
  assign n2499 = n2496 | n2498 ;
  assign n2500 = n2495 | n2499 ;
  assign n2501 = x134 & n2500 ;
  assign n2502 = n2492 | n2501 ;
  assign n2503 = n183 & n697 ;
  assign n2504 = n228 & n649 ;
  assign n2505 = n2503 | n2504 ;
  assign n2506 = ~n274 & n891 ;
  assign n2507 = n319 & n796 ;
  assign n2508 = n2506 | n2507 ;
  assign n2509 = n2505 | n2508 ;
  assign n2510 = ~x134 & n2509 ;
  assign n2511 = n228 & n748 ;
  assign n2512 = n319 & n552 ;
  assign n2513 = n2511 | n2512 ;
  assign n2514 = n183 & n843 ;
  assign n2515 = ~n274 & n600 ;
  assign n2516 = n2514 | n2515 ;
  assign n2517 = n2513 | n2516 ;
  assign n2518 = x134 & n2517 ;
  assign n2519 = n2510 | n2518 ;
  assign n2520 = n183 & n976 ;
  assign n2521 = n228 & n956 ;
  assign n2522 = n2520 | n2521 ;
  assign n2523 = ~n274 & n1062 ;
  assign n2524 = n319 & n1019 ;
  assign n2525 = n2523 | n2524 ;
  assign n2526 = n2522 | n2525 ;
  assign n2527 = ~x134 & n2526 ;
  assign n2528 = n228 & n999 ;
  assign n2529 = n319 & n915 ;
  assign n2530 = n2528 | n2529 ;
  assign n2531 = n183 & n1042 ;
  assign n2532 = ~n274 & n935 ;
  assign n2533 = n2531 | n2532 ;
  assign n2534 = n2530 | n2533 ;
  assign n2535 = x134 & n2534 ;
  assign n2536 = n2527 | n2535 ;
  assign n2537 = n183 & n1098 ;
  assign n2538 = ~n274 & n1325 ;
  assign n2539 = n2537 | n2538 ;
  assign n2540 = n228 & n1163 ;
  assign n2541 = n319 & n1293 ;
  assign n2542 = n2540 | n2541 ;
  assign n2543 = n2539 | n2542 ;
  assign n2544 = ~x134 & n2543 ;
  assign n2545 = n228 & n1230 ;
  assign n2546 = ~n274 & n1130 ;
  assign n2547 = n2545 | n2546 ;
  assign n2548 = n183 & n1260 ;
  assign n2549 = n319 & n1195 ;
  assign n2550 = n2548 | n2549 ;
  assign n2551 = n2547 | n2550 ;
  assign n2552 = x134 & n2551 ;
  assign n2553 = n2544 | n2552 ;
  assign n2554 = n183 & n1362 ;
  assign n2555 = n228 & n1354 ;
  assign n2556 = n2554 | n2555 ;
  assign n2557 = ~n274 & n1390 ;
  assign n2558 = n319 & n1398 ;
  assign n2559 = n2557 | n2558 ;
  assign n2560 = n2556 | n2559 ;
  assign n2561 = ~x134 & n2560 ;
  assign n2562 = n319 & n1337 ;
  assign n2563 = ~n274 & n1345 ;
  assign n2564 = n2562 | n2563 ;
  assign n2565 = n228 & n1373 ;
  assign n2566 = n183 & n1380 ;
  assign n2567 = ( n183 & n1377 ) | ( n183 & n2566 ) | ( n1377 & n2566 ) ;
  assign n2568 = n2565 | n2567 ;
  assign n2569 = n2564 | n2568 ;
  assign n2570 = x134 & n2569 ;
  assign n2571 = n2561 | n2570 ;
  assign n2572 = n183 & n1435 ;
  assign n2573 = n228 & n1427 ;
  assign n2574 = n2572 | n2573 ;
  assign n2575 = ~n274 & n1463 ;
  assign n2576 = n319 & n1471 ;
  assign n2577 = n2575 | n2576 ;
  assign n2578 = n2574 | n2577 ;
  assign n2579 = ~x134 & n2578 ;
  assign n2580 = n319 & n1410 ;
  assign n2581 = ~n274 & n1418 ;
  assign n2582 = n2580 | n2581 ;
  assign n2583 = n228 & n1446 ;
  assign n2584 = n183 & n1453 ;
  assign n2585 = ( n183 & n1450 ) | ( n183 & n2584 ) | ( n1450 & n2584 ) ;
  assign n2586 = n2583 | n2585 ;
  assign n2587 = n2582 | n2586 ;
  assign n2588 = x134 & n2587 ;
  assign n2589 = n2579 | n2588 ;
  assign n2590 = n183 & n1508 ;
  assign n2591 = n228 & n1500 ;
  assign n2592 = n2590 | n2591 ;
  assign n2593 = ~n274 & n1536 ;
  assign n2594 = n319 & n1544 ;
  assign n2595 = n2593 | n2594 ;
  assign n2596 = n2592 | n2595 ;
  assign n2597 = ~x134 & n2596 ;
  assign n2598 = n319 & n1483 ;
  assign n2599 = ~n274 & n1491 ;
  assign n2600 = n2598 | n2599 ;
  assign n2601 = n228 & n1527 ;
  assign n2602 = n183 & n1519 ;
  assign n2603 = n2601 | n2602 ;
  assign n2604 = n2600 | n2603 ;
  assign n2605 = x134 & n2604 ;
  assign n2606 = n2597 | n2605 ;
  assign n2607 = n319 & n1617 ;
  assign n2608 = ~n274 & n1609 ;
  assign n2609 = n2607 | n2608 ;
  assign n2610 = n228 & n1573 ;
  assign n2611 = n183 & n1581 ;
  assign n2612 = n2610 | n2611 ;
  assign n2613 = n2609 | n2612 ;
  assign n2614 = ~x134 & n2613 ;
  assign n2615 = n183 & n1592 ;
  assign n2616 = n228 & n1600 ;
  assign n2617 = n2615 | n2616 ;
  assign n2618 = ~n274 & n1564 ;
  assign n2619 = n319 & n1556 ;
  assign n2620 = n2618 | n2619 ;
  assign n2621 = n2617 | n2620 ;
  assign n2622 = x134 & n2621 ;
  assign n2623 = n2614 | n2622 ;
  assign n2624 = n319 & n1682 ;
  assign n2625 = ~n274 & n1689 ;
  assign n2626 = ( ~n274 & n1686 ) | ( ~n274 & n2625 ) | ( n1686 & n2625 ) ;
  assign n2627 = n2624 | n2626 ;
  assign n2628 = n228 & n1646 ;
  assign n2629 = n183 & n1654 ;
  assign n2630 = n2628 | n2629 ;
  assign n2631 = n2627 | n2630 ;
  assign n2632 = ~x134 & n2631 ;
  assign n2633 = n183 & n1665 ;
  assign n2634 = n228 & n1673 ;
  assign n2635 = n2633 | n2634 ;
  assign n2636 = ~n274 & n1637 ;
  assign n2637 = n319 & n1629 ;
  assign n2638 = n2636 | n2637 ;
  assign n2639 = n2635 | n2638 ;
  assign n2640 = x134 & n2639 ;
  assign n2641 = n2632 | n2640 ;
  assign n2642 = n319 & n1763 ;
  assign n2643 = ~n274 & n1755 ;
  assign n2644 = n2642 | n2643 ;
  assign n2645 = n228 & n1719 ;
  assign n2646 = n183 & n1727 ;
  assign n2647 = n2645 | n2646 ;
  assign n2648 = n2644 | n2647 ;
  assign n2649 = ~x134 & n2648 ;
  assign n2650 = n183 & n1738 ;
  assign n2651 = n228 & n1746 ;
  assign n2652 = n2650 | n2651 ;
  assign n2653 = ~n274 & n1710 ;
  assign n2654 = n319 & n1702 ;
  assign n2655 = n2653 | n2654 ;
  assign n2656 = n2652 | n2655 ;
  assign n2657 = x134 & n2656 ;
  assign n2658 = n2649 | n2657 ;
  assign n2659 = n183 & n1800 ;
  assign n2660 = n228 & n1792 ;
  assign n2661 = n2659 | n2660 ;
  assign n2662 = ~n274 & n1828 ;
  assign n2663 = n319 & n1836 ;
  assign n2664 = n2662 | n2663 ;
  assign n2665 = n2661 | n2664 ;
  assign n2666 = ~x134 & n2665 ;
  assign n2667 = n183 & n1811 ;
  assign n2668 = n228 & n1819 ;
  assign n2669 = n2667 | n2668 ;
  assign n2670 = ~n274 & n1783 ;
  assign n2671 = n319 & n1775 ;
  assign n2672 = n2670 | n2671 ;
  assign n2673 = n2669 | n2672 ;
  assign n2674 = x134 & n2673 ;
  assign n2675 = n2666 | n2674 ;
  assign n2676 = n183 & n1873 ;
  assign n2677 = n228 & n1865 ;
  assign n2678 = n2676 | n2677 ;
  assign n2679 = ~n274 & n1901 ;
  assign n2680 = n319 & n1909 ;
  assign n2681 = n2679 | n2680 ;
  assign n2682 = n2678 | n2681 ;
  assign n2683 = ~x134 & n2682 ;
  assign n2684 = n183 & n1884 ;
  assign n2685 = n228 & n1892 ;
  assign n2686 = n2684 | n2685 ;
  assign n2687 = ~n274 & n1856 ;
  assign n2688 = n319 & n1848 ;
  assign n2689 = n2687 | n2688 ;
  assign n2690 = n2686 | n2689 ;
  assign n2691 = x134 & n2690 ;
  assign n2692 = n2683 | n2691 ;
  assign n2693 = n183 & n1946 ;
  assign n2694 = n228 & n1938 ;
  assign n2695 = n2693 | n2694 ;
  assign n2696 = n319 & n1974 ;
  assign n2697 = ~n274 & n1981 ;
  assign n2698 = ( ~n274 & n1978 ) | ( ~n274 & n2697 ) | ( n1978 & n2697 ) ;
  assign n2699 = n2696 | n2698 ;
  assign n2700 = n2695 | n2699 ;
  assign n2701 = ~x134 & n2700 ;
  assign n2702 = n183 & n1957 ;
  assign n2703 = n228 & n1965 ;
  assign n2704 = n2702 | n2703 ;
  assign n2705 = ~n274 & n1929 ;
  assign n2706 = n319 & n1921 ;
  assign n2707 = n2705 | n2706 ;
  assign n2708 = n2704 | n2707 ;
  assign n2709 = x134 & n2708 ;
  assign n2710 = n2701 | n2709 ;
  assign n2711 = n183 & n2019 ;
  assign n2712 = n228 & n2011 ;
  assign n2713 = n2711 | n2712 ;
  assign n2714 = n319 & n2047 ;
  assign n2715 = ~n274 & n2054 ;
  assign n2716 = ( ~n274 & n2051 ) | ( ~n274 & n2715 ) | ( n2051 & n2715 ) ;
  assign n2717 = n2714 | n2716 ;
  assign n2718 = n2713 | n2717 ;
  assign n2719 = ~x134 & n2718 ;
  assign n2720 = n183 & n2030 ;
  assign n2721 = n228 & n2038 ;
  assign n2722 = n2720 | n2721 ;
  assign n2723 = ~n274 & n2002 ;
  assign n2724 = n319 & n1994 ;
  assign n2725 = n2723 | n2724 ;
  assign n2726 = n2722 | n2725 ;
  assign n2727 = x134 & n2726 ;
  assign n2728 = n2719 | n2727 ;
  assign n2729 = n183 & n2092 ;
  assign n2730 = n228 & n2084 ;
  assign n2731 = n2729 | n2730 ;
  assign n2732 = ~n274 & n2120 ;
  assign n2733 = n319 & n2128 ;
  assign n2734 = n2732 | n2733 ;
  assign n2735 = n2731 | n2734 ;
  assign n2736 = ~x134 & n2735 ;
  assign n2737 = n183 & n2103 ;
  assign n2738 = n228 & n2111 ;
  assign n2739 = n2737 | n2738 ;
  assign n2740 = ~n274 & n2075 ;
  assign n2741 = n319 & n2067 ;
  assign n2742 = n2740 | n2741 ;
  assign n2743 = n2739 | n2742 ;
  assign n2744 = x134 & n2743 ;
  assign n2745 = n2736 | n2744 ;
  assign n2746 = n183 & n2165 ;
  assign n2747 = n228 & n2157 ;
  assign n2748 = n2746 | n2747 ;
  assign n2749 = ~n274 & n2193 ;
  assign n2750 = n319 & n2201 ;
  assign n2751 = n2749 | n2750 ;
  assign n2752 = n2748 | n2751 ;
  assign n2753 = ~x134 & n2752 ;
  assign n2754 = n183 & n2176 ;
  assign n2755 = n228 & n2184 ;
  assign n2756 = n2754 | n2755 ;
  assign n2757 = ~n274 & n2148 ;
  assign n2758 = n319 & n2140 ;
  assign n2759 = n2757 | n2758 ;
  assign n2760 = n2756 | n2759 ;
  assign n2761 = x134 & n2760 ;
  assign n2762 = n2753 | n2761 ;
  assign n2763 = n183 & n273 ;
  assign n2764 = n228 & n366 ;
  assign n2765 = n2763 | n2764 ;
  assign n2766 = n319 & n410 ;
  assign n2767 = ~n274 & n499 ;
  assign n2768 = ( ~n274 & n478 ) | ( ~n274 & n2767 ) | ( n478 & n2767 ) ;
  assign n2769 = n2766 | n2768 ;
  assign n2770 = n2765 | n2769 ;
  assign n2771 = ~x134 & n2770 ;
  assign n2772 = n182 & n228 ;
  assign n2773 = n227 & n319 ;
  assign n2774 = n2772 | n2773 ;
  assign n2775 = n183 & n455 ;
  assign n2776 = ~n274 & n318 ;
  assign n2777 = n2775 | n2776 ;
  assign n2778 = n2774 | n2777 ;
  assign n2779 = x134 & n2778 ;
  assign n2780 = n2771 | n2779 ;
  assign n2781 = n183 & n649 ;
  assign n2782 = n228 & n796 ;
  assign n2783 = n2781 | n2782 ;
  assign n2784 = ~n274 & n843 ;
  assign n2785 = n319 & n891 ;
  assign n2786 = n2784 | n2785 ;
  assign n2787 = n2783 | n2786 ;
  assign n2788 = ~x134 & n2787 ;
  assign n2789 = n183 & n748 ;
  assign n2790 = n228 & n552 ;
  assign n2791 = n2789 | n2790 ;
  assign n2792 = ~n274 & n697 ;
  assign n2793 = n319 & n600 ;
  assign n2794 = n2792 | n2793 ;
  assign n2795 = n2791 | n2794 ;
  assign n2796 = x134 & n2795 ;
  assign n2797 = n2788 | n2796 ;
  assign n2798 = n183 & n956 ;
  assign n2799 = n228 & n1019 ;
  assign n2800 = n2798 | n2799 ;
  assign n2801 = ~n274 & n1042 ;
  assign n2802 = n319 & n1062 ;
  assign n2803 = n2801 | n2802 ;
  assign n2804 = n2800 | n2803 ;
  assign n2805 = ~x134 & n2804 ;
  assign n2806 = n183 & n999 ;
  assign n2807 = n228 & n915 ;
  assign n2808 = n2806 | n2807 ;
  assign n2809 = ~n274 & n976 ;
  assign n2810 = n319 & n935 ;
  assign n2811 = n2809 | n2810 ;
  assign n2812 = n2808 | n2811 ;
  assign n2813 = x134 & n2812 ;
  assign n2814 = n2805 | n2813 ;
  assign n2815 = ~n274 & n1260 ;
  assign n2816 = n319 & n1325 ;
  assign n2817 = n2815 | n2816 ;
  assign n2818 = n183 & n1163 ;
  assign n2819 = n228 & n1293 ;
  assign n2820 = n2818 | n2819 ;
  assign n2821 = n2817 | n2820 ;
  assign n2822 = ~x134 & n2821 ;
  assign n2823 = n183 & n1230 ;
  assign n2824 = ~n274 & n1098 ;
  assign n2825 = n2823 | n2824 ;
  assign n2826 = n228 & n1195 ;
  assign n2827 = n319 & n1130 ;
  assign n2828 = n2826 | n2827 ;
  assign n2829 = n2825 | n2828 ;
  assign n2830 = x134 & n2829 ;
  assign n2831 = n2822 | n2830 ;
  assign n2832 = n183 & n1354 ;
  assign n2833 = ~n274 & n1380 ;
  assign n2834 = ( ~n274 & n1377 ) | ( ~n274 & n2833 ) | ( n1377 & n2833 ) ;
  assign n2835 = n2832 | n2834 ;
  assign n2836 = n319 & n1390 ;
  assign n2837 = n228 & n1398 ;
  assign n2838 = n2836 | n2837 ;
  assign n2839 = n2835 | n2838 ;
  assign n2840 = ~x134 & n2839 ;
  assign n2841 = n228 & n1337 ;
  assign n2842 = n319 & n1345 ;
  assign n2843 = n2841 | n2842 ;
  assign n2844 = ~n274 & n1362 ;
  assign n2845 = n183 & n1373 ;
  assign n2846 = n2844 | n2845 ;
  assign n2847 = n2843 | n2846 ;
  assign n2848 = x134 & n2847 ;
  assign n2849 = n2840 | n2848 ;
  assign n2850 = n183 & n1427 ;
  assign n2851 = ~n274 & n1453 ;
  assign n2852 = ( ~n274 & n1450 ) | ( ~n274 & n2851 ) | ( n1450 & n2851 ) ;
  assign n2853 = n2850 | n2852 ;
  assign n2854 = n319 & n1463 ;
  assign n2855 = n228 & n1471 ;
  assign n2856 = n2854 | n2855 ;
  assign n2857 = n2853 | n2856 ;
  assign n2858 = ~x134 & n2857 ;
  assign n2859 = n228 & n1410 ;
  assign n2860 = n319 & n1418 ;
  assign n2861 = n2859 | n2860 ;
  assign n2862 = ~n274 & n1435 ;
  assign n2863 = n183 & n1446 ;
  assign n2864 = n2862 | n2863 ;
  assign n2865 = n2861 | n2864 ;
  assign n2866 = x134 & n2865 ;
  assign n2867 = n2858 | n2866 ;
  assign n2868 = ~n274 & n1519 ;
  assign n2869 = n183 & n1500 ;
  assign n2870 = n2868 | n2869 ;
  assign n2871 = n319 & n1536 ;
  assign n2872 = n228 & n1544 ;
  assign n2873 = n2871 | n2872 ;
  assign n2874 = n2870 | n2873 ;
  assign n2875 = ~x134 & n2874 ;
  assign n2876 = n228 & n1483 ;
  assign n2877 = n319 & n1491 ;
  assign n2878 = n2876 | n2877 ;
  assign n2879 = ~n274 & n1508 ;
  assign n2880 = n183 & n1527 ;
  assign n2881 = n2879 | n2880 ;
  assign n2882 = n2878 | n2881 ;
  assign n2883 = x134 & n2882 ;
  assign n2884 = n2875 | n2883 ;
  assign n2885 = ~n274 & n1592 ;
  assign n2886 = n228 & n1617 ;
  assign n2887 = n2885 | n2886 ;
  assign n2888 = n183 & n1573 ;
  assign n2889 = n319 & n1609 ;
  assign n2890 = n2888 | n2889 ;
  assign n2891 = n2887 | n2890 ;
  assign n2892 = ~x134 & n2891 ;
  assign n2893 = n183 & n1600 ;
  assign n2894 = n228 & n1556 ;
  assign n2895 = n2893 | n2894 ;
  assign n2896 = ~n274 & n1581 ;
  assign n2897 = n319 & n1564 ;
  assign n2898 = n2896 | n2897 ;
  assign n2899 = n2895 | n2898 ;
  assign n2900 = x134 & n2899 ;
  assign n2901 = n2892 | n2900 ;
  assign n2902 = ~n274 & n1665 ;
  assign n2903 = n228 & n1682 ;
  assign n2904 = n2902 | n2903 ;
  assign n2905 = n183 & n1646 ;
  assign n2906 = n319 & n1689 ;
  assign n2907 = ( n319 & n1686 ) | ( n319 & n2906 ) | ( n1686 & n2906 ) ;
  assign n2908 = n2905 | n2907 ;
  assign n2909 = n2904 | n2908 ;
  assign n2910 = ~x134 & n2909 ;
  assign n2911 = n183 & n1673 ;
  assign n2912 = n228 & n1629 ;
  assign n2913 = n2911 | n2912 ;
  assign n2914 = ~n274 & n1654 ;
  assign n2915 = n319 & n1637 ;
  assign n2916 = n2914 | n2915 ;
  assign n2917 = n2913 | n2916 ;
  assign n2918 = x134 & n2917 ;
  assign n2919 = n2910 | n2918 ;
  assign n2920 = ~n274 & n1738 ;
  assign n2921 = n228 & n1763 ;
  assign n2922 = n2920 | n2921 ;
  assign n2923 = n183 & n1719 ;
  assign n2924 = n319 & n1755 ;
  assign n2925 = n2923 | n2924 ;
  assign n2926 = n2922 | n2925 ;
  assign n2927 = ~x134 & n2926 ;
  assign n2928 = n183 & n1746 ;
  assign n2929 = n228 & n1702 ;
  assign n2930 = n2928 | n2929 ;
  assign n2931 = ~n274 & n1727 ;
  assign n2932 = n319 & n1710 ;
  assign n2933 = n2931 | n2932 ;
  assign n2934 = n2930 | n2933 ;
  assign n2935 = x134 & n2934 ;
  assign n2936 = n2927 | n2935 ;
  assign n2937 = ~n274 & n1811 ;
  assign n2938 = n183 & n1792 ;
  assign n2939 = n2937 | n2938 ;
  assign n2940 = n319 & n1828 ;
  assign n2941 = n228 & n1836 ;
  assign n2942 = n2940 | n2941 ;
  assign n2943 = n2939 | n2942 ;
  assign n2944 = ~x134 & n2943 ;
  assign n2945 = n183 & n1819 ;
  assign n2946 = n228 & n1775 ;
  assign n2947 = n2945 | n2946 ;
  assign n2948 = ~n274 & n1800 ;
  assign n2949 = n319 & n1783 ;
  assign n2950 = n2948 | n2949 ;
  assign n2951 = n2947 | n2950 ;
  assign n2952 = x134 & n2951 ;
  assign n2953 = n2944 | n2952 ;
  assign n2954 = ~n274 & n1884 ;
  assign n2955 = n183 & n1865 ;
  assign n2956 = n2954 | n2955 ;
  assign n2957 = n319 & n1901 ;
  assign n2958 = n228 & n1909 ;
  assign n2959 = n2957 | n2958 ;
  assign n2960 = n2956 | n2959 ;
  assign n2961 = ~x134 & n2960 ;
  assign n2962 = n183 & n1892 ;
  assign n2963 = n228 & n1848 ;
  assign n2964 = n2962 | n2963 ;
  assign n2965 = ~n274 & n1873 ;
  assign n2966 = n319 & n1856 ;
  assign n2967 = n2965 | n2966 ;
  assign n2968 = n2964 | n2967 ;
  assign n2969 = x134 & n2968 ;
  assign n2970 = n2961 | n2969 ;
  assign n2971 = ~n274 & n1957 ;
  assign n2972 = n183 & n1938 ;
  assign n2973 = n2971 | n2972 ;
  assign n2974 = n228 & n1974 ;
  assign n2975 = n319 & n1981 ;
  assign n2976 = ( n319 & n1978 ) | ( n319 & n2975 ) | ( n1978 & n2975 ) ;
  assign n2977 = n2974 | n2976 ;
  assign n2978 = n2973 | n2977 ;
  assign n2979 = ~x134 & n2978 ;
  assign n2980 = n183 & n1965 ;
  assign n2981 = n228 & n1921 ;
  assign n2982 = n2980 | n2981 ;
  assign n2983 = ~n274 & n1946 ;
  assign n2984 = n319 & n1929 ;
  assign n2985 = n2983 | n2984 ;
  assign n2986 = n2982 | n2985 ;
  assign n2987 = x134 & n2986 ;
  assign n2988 = n2979 | n2987 ;
  assign n2989 = ~n274 & n2030 ;
  assign n2990 = n183 & n2011 ;
  assign n2991 = n2989 | n2990 ;
  assign n2992 = n228 & n2047 ;
  assign n2993 = n319 & n2054 ;
  assign n2994 = ( n319 & n2051 ) | ( n319 & n2993 ) | ( n2051 & n2993 ) ;
  assign n2995 = n2992 | n2994 ;
  assign n2996 = n2991 | n2995 ;
  assign n2997 = ~x134 & n2996 ;
  assign n2998 = n183 & n2038 ;
  assign n2999 = n228 & n1994 ;
  assign n3000 = n2998 | n2999 ;
  assign n3001 = ~n274 & n2019 ;
  assign n3002 = n319 & n2002 ;
  assign n3003 = n3001 | n3002 ;
  assign n3004 = n3000 | n3003 ;
  assign n3005 = x134 & n3004 ;
  assign n3006 = n2997 | n3005 ;
  assign n3007 = ~n274 & n2103 ;
  assign n3008 = n183 & n2084 ;
  assign n3009 = n3007 | n3008 ;
  assign n3010 = n319 & n2120 ;
  assign n3011 = n228 & n2128 ;
  assign n3012 = n3010 | n3011 ;
  assign n3013 = n3009 | n3012 ;
  assign n3014 = ~x134 & n3013 ;
  assign n3015 = n183 & n2111 ;
  assign n3016 = n228 & n2067 ;
  assign n3017 = n3015 | n3016 ;
  assign n3018 = ~n274 & n2092 ;
  assign n3019 = n319 & n2075 ;
  assign n3020 = n3018 | n3019 ;
  assign n3021 = n3017 | n3020 ;
  assign n3022 = x134 & n3021 ;
  assign n3023 = n3014 | n3022 ;
  assign n3024 = ~n274 & n2176 ;
  assign n3025 = n183 & n2157 ;
  assign n3026 = n3024 | n3025 ;
  assign n3027 = n319 & n2193 ;
  assign n3028 = n228 & n2201 ;
  assign n3029 = n3027 | n3028 ;
  assign n3030 = n3026 | n3029 ;
  assign n3031 = ~x134 & n3030 ;
  assign n3032 = n183 & n2184 ;
  assign n3033 = n228 & n2140 ;
  assign n3034 = n3032 | n3033 ;
  assign n3035 = ~n274 & n2165 ;
  assign n3036 = n319 & n2148 ;
  assign n3037 = n3035 | n3036 ;
  assign n3038 = n3034 | n3037 ;
  assign n3039 = x134 & n3038 ;
  assign n3040 = n3031 | n3039 ;
  assign n3041 = ~x134 & n503 ;
  assign n3042 = x134 & n322 ;
  assign n3043 = n3041 | n3042 ;
  assign n3044 = ~x134 & n894 ;
  assign n3045 = x134 & n700 ;
  assign n3046 = n3044 | n3045 ;
  assign n3047 = ~x134 & n1065 ;
  assign n3048 = x134 & n979 ;
  assign n3049 = n3047 | n3048 ;
  assign n3050 = ~x134 & n1328 ;
  assign n3051 = x134 & n1198 ;
  assign n3052 = n3050 | n3051 ;
  assign n3053 = ~x134 & n1401 ;
  assign n3054 = x134 & n1365 ;
  assign n3055 = n3053 | n3054 ;
  assign n3056 = ~x134 & n1474 ;
  assign n3057 = x134 & n1438 ;
  assign n3058 = n3056 | n3057 ;
  assign n3059 = ~x134 & n1547 ;
  assign n3060 = x134 & n1511 ;
  assign n3061 = n3059 | n3060 ;
  assign n3062 = ~x134 & n1620 ;
  assign n3063 = x134 & n1584 ;
  assign n3064 = n3062 | n3063 ;
  assign n3065 = ~x134 & n1693 ;
  assign n3066 = x134 & n1657 ;
  assign n3067 = n3065 | n3066 ;
  assign n3068 = ~x134 & n1766 ;
  assign n3069 = x134 & n1730 ;
  assign n3070 = n3068 | n3069 ;
  assign n3071 = ~x134 & n1839 ;
  assign n3072 = x134 & n1803 ;
  assign n3073 = n3071 | n3072 ;
  assign n3074 = ~x134 & n1912 ;
  assign n3075 = x134 & n1876 ;
  assign n3076 = n3074 | n3075 ;
  assign n3077 = ~x134 & n1985 ;
  assign n3078 = x134 & n1949 ;
  assign n3079 = n3077 | n3078 ;
  assign n3080 = ~x134 & n2058 ;
  assign n3081 = x134 & n2022 ;
  assign n3082 = n3080 | n3081 ;
  assign n3083 = ~x134 & n2131 ;
  assign n3084 = x134 & n2095 ;
  assign n3085 = n3083 | n3084 ;
  assign n3086 = ~x134 & n2204 ;
  assign n3087 = x134 & n2168 ;
  assign n3088 = n3086 | n3087 ;
  assign n3089 = ~x134 & n2222 ;
  assign n3090 = x134 & n2213 ;
  assign n3091 = n3089 | n3090 ;
  assign n3092 = ~x134 & n2239 ;
  assign n3093 = x134 & n2231 ;
  assign n3094 = n3092 | n3093 ;
  assign n3095 = ~x134 & n2256 ;
  assign n3096 = x134 & n2248 ;
  assign n3097 = n3095 | n3096 ;
  assign n3098 = ~x134 & n2273 ;
  assign n3099 = x134 & n2265 ;
  assign n3100 = n3098 | n3099 ;
  assign n3101 = ~x134 & n2291 ;
  assign n3102 = x134 & n2282 ;
  assign n3103 = n3101 | n3102 ;
  assign n3104 = ~x134 & n2309 ;
  assign n3105 = x134 & n2300 ;
  assign n3106 = n3104 | n3105 ;
  assign n3107 = ~x134 & n2326 ;
  assign n3108 = x134 & n2318 ;
  assign n3109 = n3107 | n3108 ;
  assign n3110 = ~x134 & n2343 ;
  assign n3111 = x134 & n2335 ;
  assign n3112 = n3110 | n3111 ;
  assign n3113 = ~x134 & n2361 ;
  assign n3114 = x134 & n2352 ;
  assign n3115 = n3113 | n3114 ;
  assign n3116 = ~x134 & n2378 ;
  assign n3117 = x134 & n2370 ;
  assign n3118 = n3116 | n3117 ;
  assign n3119 = ~x134 & n2395 ;
  assign n3120 = x134 & n2387 ;
  assign n3121 = n3119 | n3120 ;
  assign n3122 = ~x134 & n2412 ;
  assign n3123 = x134 & n2404 ;
  assign n3124 = n3122 | n3123 ;
  assign n3125 = ~x134 & n2430 ;
  assign n3126 = x134 & n2421 ;
  assign n3127 = n3125 | n3126 ;
  assign n3128 = ~x134 & n2448 ;
  assign n3129 = x134 & n2439 ;
  assign n3130 = n3128 | n3129 ;
  assign n3131 = ~x134 & n2465 ;
  assign n3132 = x134 & n2457 ;
  assign n3133 = n3131 | n3132 ;
  assign n3134 = ~x134 & n2482 ;
  assign n3135 = x134 & n2474 ;
  assign n3136 = n3134 | n3135 ;
  assign n3137 = ~x134 & n2500 ;
  assign n3138 = x134 & n2491 ;
  assign n3139 = n3137 | n3138 ;
  assign n3140 = ~x134 & n2517 ;
  assign n3141 = x134 & n2509 ;
  assign n3142 = n3140 | n3141 ;
  assign n3143 = ~x134 & n2534 ;
  assign n3144 = x134 & n2526 ;
  assign n3145 = n3143 | n3144 ;
  assign n3146 = ~x134 & n2551 ;
  assign n3147 = x134 & n2543 ;
  assign n3148 = n3146 | n3147 ;
  assign n3149 = ~x134 & n2569 ;
  assign n3150 = x134 & n2560 ;
  assign n3151 = n3149 | n3150 ;
  assign n3152 = ~x134 & n2587 ;
  assign n3153 = x134 & n2578 ;
  assign n3154 = n3152 | n3153 ;
  assign n3155 = ~x134 & n2604 ;
  assign n3156 = x134 & n2596 ;
  assign n3157 = n3155 | n3156 ;
  assign n3158 = ~x134 & n2621 ;
  assign n3159 = x134 & n2613 ;
  assign n3160 = n3158 | n3159 ;
  assign n3161 = ~x134 & n2639 ;
  assign n3162 = x134 & n2631 ;
  assign n3163 = n3161 | n3162 ;
  assign n3164 = ~x134 & n2656 ;
  assign n3165 = x134 & n2648 ;
  assign n3166 = n3164 | n3165 ;
  assign n3167 = ~x134 & n2673 ;
  assign n3168 = x134 & n2665 ;
  assign n3169 = n3167 | n3168 ;
  assign n3170 = ~x134 & n2690 ;
  assign n3171 = x134 & n2682 ;
  assign n3172 = n3170 | n3171 ;
  assign n3173 = ~x134 & n2708 ;
  assign n3174 = x134 & n2700 ;
  assign n3175 = n3173 | n3174 ;
  assign n3176 = ~x134 & n2726 ;
  assign n3177 = x134 & n2718 ;
  assign n3178 = n3176 | n3177 ;
  assign n3179 = ~x134 & n2743 ;
  assign n3180 = x134 & n2735 ;
  assign n3181 = n3179 | n3180 ;
  assign n3182 = ~x134 & n2760 ;
  assign n3183 = x134 & n2752 ;
  assign n3184 = n3182 | n3183 ;
  assign n3185 = ~x134 & n2778 ;
  assign n3186 = x134 & n2770 ;
  assign n3187 = n3185 | n3186 ;
  assign n3188 = ~x134 & n2795 ;
  assign n3189 = x134 & n2787 ;
  assign n3190 = n3188 | n3189 ;
  assign n3191 = ~x134 & n2812 ;
  assign n3192 = x134 & n2804 ;
  assign n3193 = n3191 | n3192 ;
  assign n3194 = ~x134 & n2829 ;
  assign n3195 = x134 & n2821 ;
  assign n3196 = n3194 | n3195 ;
  assign n3197 = ~x134 & n2847 ;
  assign n3198 = x134 & n2839 ;
  assign n3199 = n3197 | n3198 ;
  assign n3200 = ~x134 & n2865 ;
  assign n3201 = x134 & n2857 ;
  assign n3202 = n3200 | n3201 ;
  assign n3203 = ~x134 & n2882 ;
  assign n3204 = x134 & n2874 ;
  assign n3205 = n3203 | n3204 ;
  assign n3206 = ~x134 & n2899 ;
  assign n3207 = x134 & n2891 ;
  assign n3208 = n3206 | n3207 ;
  assign n3209 = ~x134 & n2917 ;
  assign n3210 = x134 & n2909 ;
  assign n3211 = n3209 | n3210 ;
  assign n3212 = ~x134 & n2934 ;
  assign n3213 = x134 & n2926 ;
  assign n3214 = n3212 | n3213 ;
  assign n3215 = ~x134 & n2951 ;
  assign n3216 = x134 & n2943 ;
  assign n3217 = n3215 | n3216 ;
  assign n3218 = ~x134 & n2968 ;
  assign n3219 = x134 & n2960 ;
  assign n3220 = n3218 | n3219 ;
  assign n3221 = ~x134 & n2986 ;
  assign n3222 = x134 & n2978 ;
  assign n3223 = n3221 | n3222 ;
  assign n3224 = ~x134 & n3004 ;
  assign n3225 = x134 & n2996 ;
  assign n3226 = n3224 | n3225 ;
  assign n3227 = ~x134 & n3021 ;
  assign n3228 = x134 & n3013 ;
  assign n3229 = n3227 | n3228 ;
  assign n3230 = ~x134 & n3038 ;
  assign n3231 = x134 & n3030 ;
  assign n3232 = n3230 | n3231 ;
  assign y0 = n505 ;
  assign y1 = n896 ;
  assign y2 = n1067 ;
  assign y3 = n1330 ;
  assign y4 = n1403 ;
  assign y5 = n1476 ;
  assign y6 = n1549 ;
  assign y7 = n1622 ;
  assign y8 = n1695 ;
  assign y9 = n1768 ;
  assign y10 = n1841 ;
  assign y11 = n1914 ;
  assign y12 = n1987 ;
  assign y13 = n2060 ;
  assign y14 = n2133 ;
  assign y15 = n2206 ;
  assign y16 = n2224 ;
  assign y17 = n2241 ;
  assign y18 = n2258 ;
  assign y19 = n2275 ;
  assign y20 = n2293 ;
  assign y21 = n2311 ;
  assign y22 = n2328 ;
  assign y23 = n2345 ;
  assign y24 = n2363 ;
  assign y25 = n2380 ;
  assign y26 = n2397 ;
  assign y27 = n2414 ;
  assign y28 = n2432 ;
  assign y29 = n2450 ;
  assign y30 = n2467 ;
  assign y31 = n2484 ;
  assign y32 = n2502 ;
  assign y33 = n2519 ;
  assign y34 = n2536 ;
  assign y35 = n2553 ;
  assign y36 = n2571 ;
  assign y37 = n2589 ;
  assign y38 = n2606 ;
  assign y39 = n2623 ;
  assign y40 = n2641 ;
  assign y41 = n2658 ;
  assign y42 = n2675 ;
  assign y43 = n2692 ;
  assign y44 = n2710 ;
  assign y45 = n2728 ;
  assign y46 = n2745 ;
  assign y47 = n2762 ;
  assign y48 = n2780 ;
  assign y49 = n2797 ;
  assign y50 = n2814 ;
  assign y51 = n2831 ;
  assign y52 = n2849 ;
  assign y53 = n2867 ;
  assign y54 = n2884 ;
  assign y55 = n2901 ;
  assign y56 = n2919 ;
  assign y57 = n2936 ;
  assign y58 = n2953 ;
  assign y59 = n2970 ;
  assign y60 = n2988 ;
  assign y61 = n3006 ;
  assign y62 = n3023 ;
  assign y63 = n3040 ;
  assign y64 = n3043 ;
  assign y65 = n3046 ;
  assign y66 = n3049 ;
  assign y67 = n3052 ;
  assign y68 = n3055 ;
  assign y69 = n3058 ;
  assign y70 = n3061 ;
  assign y71 = n3064 ;
  assign y72 = n3067 ;
  assign y73 = n3070 ;
  assign y74 = n3073 ;
  assign y75 = n3076 ;
  assign y76 = n3079 ;
  assign y77 = n3082 ;
  assign y78 = n3085 ;
  assign y79 = n3088 ;
  assign y80 = n3091 ;
  assign y81 = n3094 ;
  assign y82 = n3097 ;
  assign y83 = n3100 ;
  assign y84 = n3103 ;
  assign y85 = n3106 ;
  assign y86 = n3109 ;
  assign y87 = n3112 ;
  assign y88 = n3115 ;
  assign y89 = n3118 ;
  assign y90 = n3121 ;
  assign y91 = n3124 ;
  assign y92 = n3127 ;
  assign y93 = n3130 ;
  assign y94 = n3133 ;
  assign y95 = n3136 ;
  assign y96 = n3139 ;
  assign y97 = n3142 ;
  assign y98 = n3145 ;
  assign y99 = n3148 ;
  assign y100 = n3151 ;
  assign y101 = n3154 ;
  assign y102 = n3157 ;
  assign y103 = n3160 ;
  assign y104 = n3163 ;
  assign y105 = n3166 ;
  assign y106 = n3169 ;
  assign y107 = n3172 ;
  assign y108 = n3175 ;
  assign y109 = n3178 ;
  assign y110 = n3181 ;
  assign y111 = n3184 ;
  assign y112 = n3187 ;
  assign y113 = n3190 ;
  assign y114 = n3193 ;
  assign y115 = n3196 ;
  assign y116 = n3199 ;
  assign y117 = n3202 ;
  assign y118 = n3205 ;
  assign y119 = n3208 ;
  assign y120 = n3211 ;
  assign y121 = n3214 ;
  assign y122 = n3217 ;
  assign y123 = n3220 ;
  assign y124 = n3223 ;
  assign y125 = n3226 ;
  assign y126 = n3229 ;
  assign y127 = n3232 ;
endmodule
