module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 ;
  wire n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 ;
  assign n148 = x13 | x14 ;
  assign n149 = x6 | x7 ;
  assign n150 = n148 | n149 ;
  assign n151 = x17 | x21 ;
  assign n152 = x8 | x12 ;
  assign n153 = n151 | n152 ;
  assign n154 = n150 | n153 ;
  assign n155 = x18 | x19 ;
  assign n156 = x4 | x16 ;
  assign n157 = n155 | n156 ;
  assign n158 = x5 | x22 ;
  assign n159 = x9 | x11 ;
  assign n160 = n158 | n159 ;
  assign n161 = n157 | n160 ;
  assign n162 = n154 | n161 ;
  assign n163 = x0 | x54 ;
  assign n164 = ( x0 & n162 ) | ( x0 & n163 ) | ( n162 & n163 ) ;
  assign n165 = ~x54 & n164 ;
  assign n166 = ~n158 & n159 ;
  assign n167 = ~x56 & n166 ;
  assign n168 = x54 & n167 ;
  assign n169 = n164 & ~n168 ;
  assign n170 = ~x56 & n158 ;
  assign n171 = x6 | x12 ;
  assign n172 = x17 | n157 ;
  assign n173 = n171 | n172 ;
  assign n174 = x8 | x21 ;
  assign n175 = x7 | n174 ;
  assign n176 = x10 & ~n148 ;
  assign n177 = ~n175 & n176 ;
  assign n178 = ~x13 & x14 ;
  assign n179 = ~n175 & n178 ;
  assign n180 = x14 & ~n179 ;
  assign n181 = x8 & x21 ;
  assign n182 = ( x7 & n174 ) | ( x7 & ~n181 ) | ( n174 & ~n181 ) ;
  assign n183 = ( x7 & x13 ) | ( x7 & n174 ) | ( x13 & n174 ) ;
  assign n184 = x13 & ~n182 ;
  assign n185 = ( n182 & ~n183 ) | ( n182 & n184 ) | ( ~n183 & n184 ) ;
  assign n186 = ( n179 & ~n180 ) | ( n179 & n185 ) | ( ~n180 & n185 ) ;
  assign n187 = ~n177 & n186 ;
  assign n188 = ~x10 & n187 ;
  assign n189 = ( ~n158 & n177 ) | ( ~n158 & n188 ) | ( n177 & n188 ) ;
  assign n190 = ~n170 & n189 ;
  assign n191 = ~n173 & n190 ;
  assign n192 = ( ~n159 & n170 ) | ( ~n159 & n191 ) | ( n170 & n191 ) ;
  assign n193 = ( n165 & n169 ) | ( n165 & ~n192 ) | ( n169 & ~n192 ) ;
  assign n194 = x129 | n193 ;
  assign n195 = x3 | n194 ;
  assign n196 = x11 | x12 ;
  assign n197 = n174 | n196 ;
  assign n198 = n157 | n197 ;
  assign n199 = x10 | x22 ;
  assign n200 = x7 | x13 ;
  assign n201 = x5 | x6 ;
  assign n202 = n200 | n201 ;
  assign n203 = x14 | n202 ;
  assign n204 = n199 | n203 ;
  assign n205 = n198 | n204 ;
  assign n206 = ~x17 & x54 ;
  assign n207 = n205 & n206 ;
  assign n208 = x1 | n207 ;
  assign n209 = ~x14 & x54 ;
  assign n210 = x8 | x11 ;
  assign n211 = n151 | n210 ;
  assign n212 = x6 & x12 ;
  assign n213 = ( x5 & n171 ) | ( x5 & ~n212 ) | ( n171 & ~n212 ) ;
  assign n214 = ( x5 & x7 ) | ( x5 & n171 ) | ( x7 & n171 ) ;
  assign n215 = x7 & ~n213 ;
  assign n216 = ( n213 & ~n214 ) | ( n213 & n215 ) | ( ~n214 & n215 ) ;
  assign n217 = ~x13 & n216 ;
  assign n218 = ~x7 & x13 ;
  assign n219 = x5 | n171 ;
  assign n220 = n218 & ~n219 ;
  assign n221 = n217 | n220 ;
  assign n222 = ( x9 & ~n157 ) | ( x9 & n221 ) | ( ~n157 & n221 ) ;
  assign n223 = n200 | n219 ;
  assign n224 = ( x9 & n157 ) | ( x9 & n223 ) | ( n157 & n223 ) ;
  assign n225 = n222 & ~n224 ;
  assign n226 = ~n211 & n225 ;
  assign n227 = n209 & n226 ;
  assign n228 = ~n199 & n227 ;
  assign n229 = n208 & ~n228 ;
  assign n230 = x129 | n229 ;
  assign n231 = x3 | n230 ;
  assign n232 = x122 & x127 ;
  assign n233 = x45 | x48 ;
  assign n234 = x43 | x47 ;
  assign n235 = n233 | n234 ;
  assign n236 = x15 | x20 ;
  assign n237 = x24 | x49 ;
  assign n238 = n236 | n237 ;
  assign n239 = n235 | n238 ;
  assign n240 = x41 | x46 ;
  assign n241 = x38 | x50 ;
  assign n242 = n240 | n241 ;
  assign n243 = x42 | x44 ;
  assign n244 = x40 | n243 ;
  assign n245 = x2 | n244 ;
  assign n246 = n242 | n245 ;
  assign n247 = n239 | n246 ;
  assign n248 = x82 & n247 ;
  assign n249 = n232 | n248 ;
  assign n250 = x65 | n249 ;
  assign n251 = x24 | x45 ;
  assign n252 = x47 | x48 ;
  assign n253 = n251 | n252 ;
  assign n254 = x49 | n236 ;
  assign n255 = n253 | n254 ;
  assign n256 = x38 | x40 ;
  assign n257 = n243 | n256 ;
  assign n258 = x46 | x50 ;
  assign n259 = x41 | n258 ;
  assign n260 = n257 | n259 ;
  assign n261 = x43 | n260 ;
  assign n262 = n255 | n261 ;
  assign n263 = x82 & n262 ;
  assign n264 = ~x82 & n232 ;
  assign n265 = n263 | n264 ;
  assign n266 = x2 & n265 ;
  assign n267 = n250 & ~n266 ;
  assign n268 = x129 | n267 ;
  assign n269 = x9 | x14 ;
  assign n270 = n199 | n269 ;
  assign n271 = n202 | n270 ;
  assign n272 = x8 | x17 ;
  assign n273 = n196 | n272 ;
  assign n274 = x21 | n157 ;
  assign n275 = n273 | n274 ;
  assign n276 = n271 | n275 ;
  assign n277 = x61 | x118 ;
  assign n278 = n276 & ~n277 ;
  assign n279 = x0 & ~x123 ;
  assign n280 = ~x113 & n279 ;
  assign n281 = n278 | n280 ;
  assign n282 = ~x129 & n281 ;
  assign n283 = x10 & ~x22 ;
  assign n284 = ~n269 & n283 ;
  assign n285 = ~n223 & n284 ;
  assign n286 = x54 & ~n157 ;
  assign n287 = ~n211 & n286 ;
  assign n288 = n285 & n287 ;
  assign n289 = x4 & ~x54 ;
  assign n290 = n288 | n289 ;
  assign n291 = ~x129 & n290 ;
  assign n292 = ~x3 & n291 ;
  assign n293 = x5 & ~x54 ;
  assign n294 = x7 | n171 ;
  assign n295 = x25 | x29 ;
  assign n296 = x28 & ~n295 ;
  assign n297 = ~n294 & n296 ;
  assign n298 = x13 | n270 ;
  assign n299 = n297 & ~n298 ;
  assign n300 = x59 | n211 ;
  assign n301 = ~x16 & x54 ;
  assign n302 = x4 | x19 ;
  assign n303 = x18 | n302 ;
  assign n304 = x5 | n303 ;
  assign n305 = n301 & ~n304 ;
  assign n306 = ~n300 & n305 ;
  assign n307 = n299 & n306 ;
  assign n308 = n293 | n307 ;
  assign n309 = ~x129 & n308 ;
  assign n310 = ~x3 & n309 ;
  assign n311 = x6 & ~x54 ;
  assign n312 = x5 | x7 ;
  assign n313 = x25 & ~x29 ;
  assign n314 = ~x28 & n313 ;
  assign n315 = ~x12 & n314 ;
  assign n316 = ~n312 & n315 ;
  assign n317 = ~n298 & n316 ;
  assign n318 = x6 | n303 ;
  assign n319 = n301 & ~n318 ;
  assign n320 = ~n300 & n319 ;
  assign n321 = n317 & n320 ;
  assign n322 = n311 | n321 ;
  assign n323 = ~x129 & n322 ;
  assign n324 = ~x3 & n323 ;
  assign n325 = x7 & ~x54 ;
  assign n326 = x18 | x21 ;
  assign n327 = x8 & ~x17 ;
  assign n328 = ~n326 & n327 ;
  assign n329 = x7 | n302 ;
  assign n330 = n301 & ~n329 ;
  assign n331 = n328 & n330 ;
  assign n332 = x6 | n196 ;
  assign n333 = x5 | n332 ;
  assign n334 = n298 | n333 ;
  assign n335 = n331 & ~n334 ;
  assign n336 = n325 | n335 ;
  assign n337 = ~x129 & n336 ;
  assign n338 = ~x3 & n337 ;
  assign n339 = x8 & ~x54 ;
  assign n340 = n223 | n270 ;
  assign n341 = x17 | x18 ;
  assign n342 = ~x11 & x21 ;
  assign n343 = ~n341 & n342 ;
  assign n344 = x8 | n302 ;
  assign n345 = n301 & ~n344 ;
  assign n346 = n343 & n345 ;
  assign n347 = ~n340 & n346 ;
  assign n348 = n339 | n347 ;
  assign n349 = ~x129 & n348 ;
  assign n350 = ~x3 & n349 ;
  assign n351 = x9 & ~x54 ;
  assign n352 = n148 | n199 ;
  assign n353 = x11 & ~n312 ;
  assign n354 = ~n171 & n353 ;
  assign n355 = ~n352 & n354 ;
  assign n356 = n272 | n326 ;
  assign n357 = x9 | n302 ;
  assign n358 = n301 & ~n357 ;
  assign n359 = ~n356 & n358 ;
  assign n360 = n355 & n359 ;
  assign n361 = n351 | n360 ;
  assign n362 = ~x129 & n361 ;
  assign n363 = ~x3 & n362 ;
  assign n364 = x10 & ~x54 ;
  assign n365 = x10 | n302 ;
  assign n366 = n301 & ~n365 ;
  assign n367 = ~n356 & n366 ;
  assign n368 = n312 | n332 ;
  assign n369 = x9 | x22 ;
  assign n370 = n178 & ~n369 ;
  assign n371 = ~n368 & n370 ;
  assign n372 = n367 & n371 ;
  assign n373 = n364 | n372 ;
  assign n374 = ~x129 & n373 ;
  assign n375 = ~x3 & n374 ;
  assign n376 = x11 & ~x54 ;
  assign n377 = x11 | n302 ;
  assign n378 = n301 & ~n377 ;
  assign n379 = ~n356 & n378 ;
  assign n380 = ~x10 & x22 ;
  assign n381 = ~n269 & n380 ;
  assign n382 = ~n223 & n381 ;
  assign n383 = n379 & n382 ;
  assign n384 = n376 | n383 ;
  assign n385 = ~x129 & n384 ;
  assign n386 = ~x3 & n385 ;
  assign n387 = x12 & ~x54 ;
  assign n388 = x12 | n302 ;
  assign n389 = n301 & ~n388 ;
  assign n390 = x8 | n151 ;
  assign n391 = x18 & ~n390 ;
  assign n392 = n389 & n391 ;
  assign n393 = x11 | n271 ;
  assign n394 = n392 & ~n393 ;
  assign n395 = n387 | n394 ;
  assign n396 = ~x129 & n395 ;
  assign n397 = ~x3 & n396 ;
  assign n398 = x13 & ~x54 ;
  assign n399 = x13 | n303 ;
  assign n400 = n301 & ~n399 ;
  assign n401 = ~n300 & n400 ;
  assign n402 = ~x25 & x29 ;
  assign n403 = ~x28 & n402 ;
  assign n404 = ~n219 & n403 ;
  assign n405 = x7 | n270 ;
  assign n406 = n404 & ~n405 ;
  assign n407 = n401 & n406 ;
  assign n408 = n398 | n407 ;
  assign n409 = ~x129 & n408 ;
  assign n410 = ~x3 & n409 ;
  assign n411 = x14 & ~x54 ;
  assign n412 = ~x16 & n209 ;
  assign n413 = ~n302 & n412 ;
  assign n414 = ~n356 & n413 ;
  assign n415 = ~x9 & x13 ;
  assign n416 = ~n199 & n415 ;
  assign n417 = ~n368 & n416 ;
  assign n418 = n414 & n417 ;
  assign n419 = n411 | n418 ;
  assign n420 = ~x129 & n419 ;
  assign n421 = ~x3 & n420 ;
  assign n422 = x41 | x43 ;
  assign n423 = n252 | n422 ;
  assign n424 = x45 | n237 ;
  assign n425 = n423 | n424 ;
  assign n426 = x46 | n241 ;
  assign n427 = n244 | n426 ;
  assign n428 = x15 | n427 ;
  assign n429 = n425 | n428 ;
  assign n430 = x82 & n429 ;
  assign n431 = n232 | n430 ;
  assign n432 = x70 | n431 ;
  assign n433 = x48 | n234 ;
  assign n434 = n424 | n433 ;
  assign n435 = n260 | n434 ;
  assign n436 = x15 & n435 ;
  assign n437 = x45 | n252 ;
  assign n438 = x2 | x20 ;
  assign n439 = ~x15 & n438 ;
  assign n440 = ~n261 & n439 ;
  assign n441 = ~n237 & n440 ;
  assign n442 = ~n437 & n441 ;
  assign n443 = n436 | n442 ;
  assign n444 = x82 & n443 ;
  assign n445 = x15 & n264 ;
  assign n446 = n444 | n445 ;
  assign n447 = n432 & ~n446 ;
  assign n448 = x129 | n447 ;
  assign n449 = x16 & ~x54 ;
  assign n450 = x6 & ~x12 ;
  assign n451 = ~x5 & n450 ;
  assign n452 = ~n200 & n451 ;
  assign n453 = ~n270 & n452 ;
  assign n454 = n287 & n453 ;
  assign n455 = n449 | n454 ;
  assign n456 = ~x129 & n455 ;
  assign n457 = ~x3 & n456 ;
  assign n458 = x17 & ~x54 ;
  assign n459 = x7 | n201 ;
  assign n460 = x25 | x28 ;
  assign n461 = x12 | n460 ;
  assign n462 = n459 | n461 ;
  assign n463 = n298 | n462 ;
  assign n464 = ~x16 & n206 ;
  assign n465 = ~n303 & n464 ;
  assign n466 = x11 | n174 ;
  assign n467 = ~x29 & x59 ;
  assign n468 = ~n466 & n467 ;
  assign n469 = n465 & n468 ;
  assign n470 = ~n463 & n469 ;
  assign n471 = n458 | n470 ;
  assign n472 = ~x129 & n471 ;
  assign n473 = ~x3 & n472 ;
  assign n474 = x18 & ~x54 ;
  assign n475 = x16 & x54 ;
  assign n476 = ~n303 & n475 ;
  assign n477 = ~n211 & n476 ;
  assign n478 = ~n340 & n477 ;
  assign n479 = n474 | n478 ;
  assign n480 = ~x129 & n479 ;
  assign n481 = ~x3 & n480 ;
  assign n482 = x19 & ~x54 ;
  assign n483 = x17 & ~n466 ;
  assign n484 = x4 | n155 ;
  assign n485 = n301 & ~n484 ;
  assign n486 = n483 & n485 ;
  assign n487 = ~n340 & n486 ;
  assign n488 = n482 | n487 ;
  assign n489 = ~x129 & n488 ;
  assign n490 = ~x3 & n489 ;
  assign n491 = n234 | n240 ;
  assign n492 = x24 | n233 ;
  assign n493 = n491 | n492 ;
  assign n494 = x40 | x42 ;
  assign n495 = n241 | n494 ;
  assign n496 = x44 | n254 ;
  assign n497 = n495 | n496 ;
  assign n498 = n493 | n497 ;
  assign n499 = x82 & n498 ;
  assign n500 = n232 | n499 ;
  assign n501 = x71 | n500 ;
  assign n502 = x50 | n256 ;
  assign n503 = x15 | x49 ;
  assign n504 = n243 | n503 ;
  assign n505 = n502 | n504 ;
  assign n506 = n493 | n505 ;
  assign n507 = x20 & n506 ;
  assign n508 = x2 & ~n498 ;
  assign n509 = n507 | n508 ;
  assign n510 = x82 & n509 ;
  assign n511 = x20 & n264 ;
  assign n512 = n510 | n511 ;
  assign n513 = n501 & ~n512 ;
  assign n514 = x129 | n513 ;
  assign n515 = x21 & ~x54 ;
  assign n516 = n210 | n341 ;
  assign n517 = ~x21 & x54 ;
  assign n518 = x19 & n517 ;
  assign n519 = ~n156 & n518 ;
  assign n520 = ~n516 & n519 ;
  assign n521 = ~n340 & n520 ;
  assign n522 = n515 | n521 ;
  assign n523 = ~x129 & n522 ;
  assign n524 = ~x3 & n523 ;
  assign n525 = x22 & ~x54 ;
  assign n526 = x22 | n302 ;
  assign n527 = n301 & ~n526 ;
  assign n528 = ~n356 & n527 ;
  assign n529 = x9 | x10 ;
  assign n530 = n148 | n529 ;
  assign n531 = x5 & ~x7 ;
  assign n532 = ~n332 & n531 ;
  assign n533 = ~n530 & n532 ;
  assign n534 = n528 & n533 ;
  assign n535 = n525 | n534 ;
  assign n536 = ~x129 & n535 ;
  assign n537 = ~x3 & n536 ;
  assign n538 = ~x23 & x55 ;
  assign n539 = x129 | n538 ;
  assign n540 = x61 & ~n539 ;
  assign n541 = x47 | n422 ;
  assign n542 = n233 | n541 ;
  assign n543 = n427 | n542 ;
  assign n544 = x82 & n543 ;
  assign n545 = n438 | n503 ;
  assign n546 = x82 & n545 ;
  assign n547 = n232 & ~n546 ;
  assign n548 = n544 | n547 ;
  assign n549 = ~x24 & n548 ;
  assign n550 = x2 | x45 ;
  assign n551 = n252 | n550 ;
  assign n552 = n254 | n551 ;
  assign n553 = n261 | n552 ;
  assign n554 = x82 & n553 ;
  assign n555 = n232 | n554 ;
  assign n556 = x63 & ~n555 ;
  assign n557 = x43 | n240 ;
  assign n558 = n437 | n557 ;
  assign n559 = x24 & x82 ;
  assign n560 = ~n243 & n559 ;
  assign n561 = ~n502 & n560 ;
  assign n562 = ~n558 & n561 ;
  assign n563 = x129 | n562 ;
  assign n564 = n556 | n563 ;
  assign n565 = n549 | n564 ;
  assign n566 = x25 & ~x116 ;
  assign n567 = x26 & n566 ;
  assign n568 = x51 | x52 ;
  assign n569 = x39 | n568 ;
  assign n570 = n567 | n569 ;
  assign n571 = x26 & x116 ;
  assign n572 = x95 | x100 ;
  assign n573 = x97 & ~x110 ;
  assign n574 = ( ~x110 & n572 ) | ( ~x110 & n573 ) | ( n572 & n573 ) ;
  assign n575 = x25 & ~n574 ;
  assign n576 = n571 | n575 ;
  assign n577 = ( n567 & n570 ) | ( n567 & n576 ) | ( n570 & n576 ) ;
  assign n578 = ~x85 & n577 ;
  assign n579 = x26 | x27 ;
  assign n580 = x85 | x110 ;
  assign n581 = x96 | n580 ;
  assign n582 = x85 & x116 ;
  assign n583 = x100 & n582 ;
  assign n584 = ( x100 & ~n581 ) | ( x100 & n583 ) | ( ~n581 & n583 ) ;
  assign n585 = x85 & n566 ;
  assign n586 = ( ~n579 & n584 ) | ( ~n579 & n585 ) | ( n584 & n585 ) ;
  assign n587 = ~n579 & n586 ;
  assign n588 = ( ~x27 & n578 ) | ( ~x27 & n587 ) | ( n578 & n587 ) ;
  assign n589 = ~n569 & n575 ;
  assign n590 = x26 | x85 ;
  assign n591 = x39 | x52 ;
  assign n592 = ~x51 & x116 ;
  assign n593 = ~n591 & n592 ;
  assign n594 = x27 & n566 ;
  assign n595 = ( x27 & n593 ) | ( x27 & n594 ) | ( n593 & n594 ) ;
  assign n596 = ~n590 & n595 ;
  assign n597 = ( n589 & ~n590 ) | ( n589 & n596 ) | ( ~n590 & n596 ) ;
  assign n598 = ~x53 & n597 ;
  assign n599 = ( ~x53 & n588 ) | ( ~x53 & n598 ) | ( n588 & n598 ) ;
  assign n600 = x25 & ~x26 ;
  assign n601 = ~x116 & n600 ;
  assign n602 = x27 | x85 ;
  assign n603 = ~x53 & x58 ;
  assign n604 = ~n602 & n603 ;
  assign n605 = n601 & n604 ;
  assign n606 = x53 & ~x85 ;
  assign n607 = ~x27 & n606 ;
  assign n608 = n601 & n607 ;
  assign n609 = x58 & ~n605 ;
  assign n610 = ( n605 & n608 ) | ( n605 & ~n609 ) | ( n608 & ~n609 ) ;
  assign n611 = ~x129 & n610 ;
  assign n612 = x129 | n609 ;
  assign n613 = ( n599 & n611 ) | ( n599 & ~n612 ) | ( n611 & ~n612 ) ;
  assign n614 = ~x3 & n613 ;
  assign n615 = x85 & ~x116 ;
  assign n616 = x110 | n615 ;
  assign n617 = n571 | n616 ;
  assign n618 = x96 | n617 ;
  assign n619 = ~x26 & n582 ;
  assign n620 = n618 & ~n619 ;
  assign n621 = x100 & ~n620 ;
  assign n622 = x85 | n593 ;
  assign n623 = x26 & ~n622 ;
  assign n624 = n621 | n623 ;
  assign n625 = ~x129 & n624 ;
  assign n626 = ~x3 & n625 ;
  assign n627 = x27 | x53 ;
  assign n628 = x58 | n627 ;
  assign n629 = n626 & ~n628 ;
  assign n630 = x95 & ~x96 ;
  assign n631 = x27 & x116 ;
  assign n632 = n616 | n631 ;
  assign n633 = n630 & ~n632 ;
  assign n634 = ~x27 & n582 ;
  assign n635 = n633 | n634 ;
  assign n636 = ~x100 & n635 ;
  assign n637 = x27 & ~n622 ;
  assign n638 = n636 | n637 ;
  assign n639 = ~x129 & n638 ;
  assign n640 = ~x3 & n639 ;
  assign n641 = x53 | x58 ;
  assign n642 = x26 | n641 ;
  assign n643 = n640 & ~n642 ;
  assign n644 = ~x26 & x39 ;
  assign n645 = ( ~x26 & n568 ) | ( ~x26 & n644 ) | ( n568 & n644 ) ;
  assign n646 = x27 | x51 ;
  assign n647 = n591 | n646 ;
  assign n648 = ~n645 & n647 ;
  assign n649 = n574 | n648 ;
  assign n650 = x26 & ~x27 ;
  assign n651 = ~x26 & x27 ;
  assign n652 = n650 | n651 ;
  assign n653 = ~x116 & n652 ;
  assign n654 = x28 & n653 ;
  assign n655 = ( x28 & ~n649 ) | ( x28 & n654 ) | ( ~n649 & n654 ) ;
  assign n656 = x26 | x100 ;
  assign n657 = x110 | n656 ;
  assign n658 = n630 & ~n657 ;
  assign n659 = x51 | n591 ;
  assign n660 = n571 & ~n659 ;
  assign n661 = n658 | n660 ;
  assign n662 = n631 & n645 ;
  assign n663 = x27 & ~n662 ;
  assign n664 = ( n661 & n662 ) | ( n661 & ~n663 ) | ( n662 & ~n663 ) ;
  assign n665 = n655 | n664 ;
  assign n666 = ~x26 & n606 ;
  assign n667 = x28 & ~x116 ;
  assign n668 = ~x27 & n667 ;
  assign n669 = n666 & n668 ;
  assign n670 = ( ~x85 & x100 ) | ( ~x85 & x116 ) | ( x100 & x116 ) ;
  assign n671 = ( x28 & x85 ) | ( x28 & x116 ) | ( x85 & x116 ) ;
  assign n672 = ~n670 & n671 ;
  assign n673 = ~n579 & n672 ;
  assign n674 = x85 & ~n673 ;
  assign n675 = x53 | n674 ;
  assign n676 = ~n669 & n675 ;
  assign n677 = ~x53 & n673 ;
  assign n678 = n669 | n677 ;
  assign n679 = ( n665 & ~n676 ) | ( n665 & n678 ) | ( ~n676 & n678 ) ;
  assign n680 = ~n590 & n603 ;
  assign n681 = n668 & n680 ;
  assign n682 = x58 & ~n681 ;
  assign n683 = x129 | n682 ;
  assign n684 = x3 | n683 ;
  assign n685 = ~x129 & n681 ;
  assign n686 = ~x3 & n685 ;
  assign n687 = ( n679 & ~n684 ) | ( n679 & n686 ) | ( ~n684 & n686 ) ;
  assign n688 = x29 & ~x116 ;
  assign n689 = ~x58 & x85 ;
  assign n690 = ~n627 & n689 ;
  assign n691 = n688 & n690 ;
  assign n692 = ~x26 & n691 ;
  assign n693 = n602 | n641 ;
  assign n694 = x26 & n688 ;
  assign n695 = ~n693 & n694 ;
  assign n696 = n692 | n695 ;
  assign n697 = x26 & ~n695 ;
  assign n698 = ~x96 & n573 ;
  assign n699 = x97 | n572 ;
  assign n700 = x29 & ~n699 ;
  assign n701 = ( ~n572 & n698 ) | ( ~n572 & n700 ) | ( n698 & n700 ) ;
  assign n702 = x29 & x110 ;
  assign n703 = ~x58 & n702 ;
  assign n704 = ( ~x58 & n701 ) | ( ~x58 & n703 ) | ( n701 & n703 ) ;
  assign n705 = x97 & x116 ;
  assign n706 = ( n603 & n688 ) | ( n603 & n705 ) | ( n688 & n705 ) ;
  assign n707 = n603 & n706 ;
  assign n708 = ( ~x53 & n704 ) | ( ~x53 & n707 ) | ( n704 & n707 ) ;
  assign n709 = x27 & n688 ;
  assign n710 = ~n641 & n709 ;
  assign n711 = x27 & ~n710 ;
  assign n712 = x53 & ~x58 ;
  assign n713 = n688 & n712 ;
  assign n714 = ( n710 & ~n711 ) | ( n710 & n713 ) | ( ~n711 & n713 ) ;
  assign n715 = ( n708 & ~n711 ) | ( n708 & n714 ) | ( ~n711 & n714 ) ;
  assign n716 = ~x85 & n715 ;
  assign n717 = ( n696 & ~n697 ) | ( n696 & n716 ) | ( ~n697 & n716 ) ;
  assign n718 = ~x129 & n717 ;
  assign n719 = ~x3 & n718 ;
  assign n720 = x88 & x106 ;
  assign n721 = ( ~x60 & x106 ) | ( ~x60 & x109 ) | ( x106 & x109 ) ;
  assign n722 = ( x30 & ~x106 ) | ( x30 & x109 ) | ( ~x106 & x109 ) ;
  assign n723 = ~n721 & n722 ;
  assign n724 = n720 | n723 ;
  assign n725 = ~x129 & n724 ;
  assign n726 = x89 & x106 ;
  assign n727 = ( ~x30 & x106 ) | ( ~x30 & x109 ) | ( x106 & x109 ) ;
  assign n728 = ( x31 & ~x106 ) | ( x31 & x109 ) | ( ~x106 & x109 ) ;
  assign n729 = ~n727 & n728 ;
  assign n730 = n726 | n729 ;
  assign n731 = ~x129 & n730 ;
  assign n732 = x99 & x106 ;
  assign n733 = ( ~x31 & x106 ) | ( ~x31 & x109 ) | ( x106 & x109 ) ;
  assign n734 = ( x32 & ~x106 ) | ( x32 & x109 ) | ( ~x106 & x109 ) ;
  assign n735 = ~n733 & n734 ;
  assign n736 = n732 | n735 ;
  assign n737 = ~x129 & n736 ;
  assign n738 = x90 & x106 ;
  assign n739 = ( ~x32 & x106 ) | ( ~x32 & x109 ) | ( x106 & x109 ) ;
  assign n740 = ( x33 & ~x106 ) | ( x33 & x109 ) | ( ~x106 & x109 ) ;
  assign n741 = ~n739 & n740 ;
  assign n742 = n738 | n741 ;
  assign n743 = ~x129 & n742 ;
  assign n744 = x91 & x106 ;
  assign n745 = ( ~x33 & x106 ) | ( ~x33 & x109 ) | ( x106 & x109 ) ;
  assign n746 = ( x34 & ~x106 ) | ( x34 & x109 ) | ( ~x106 & x109 ) ;
  assign n747 = ~n745 & n746 ;
  assign n748 = n744 | n747 ;
  assign n749 = ~x129 & n748 ;
  assign n750 = x92 & x106 ;
  assign n751 = ( ~x34 & x106 ) | ( ~x34 & x109 ) | ( x106 & x109 ) ;
  assign n752 = ( x35 & ~x106 ) | ( x35 & x109 ) | ( ~x106 & x109 ) ;
  assign n753 = ~n751 & n752 ;
  assign n754 = n750 | n753 ;
  assign n755 = ~x129 & n754 ;
  assign n756 = x98 & x106 ;
  assign n757 = ( ~x35 & x106 ) | ( ~x35 & x109 ) | ( x106 & x109 ) ;
  assign n758 = ( x36 & ~x106 ) | ( x36 & x109 ) | ( ~x106 & x109 ) ;
  assign n759 = ~n757 & n758 ;
  assign n760 = n756 | n759 ;
  assign n761 = ~x129 & n760 ;
  assign n762 = x93 & x106 ;
  assign n763 = ( ~x36 & x106 ) | ( ~x36 & x109 ) | ( x106 & x109 ) ;
  assign n764 = ( x37 & ~x106 ) | ( x37 & x109 ) | ( ~x106 & x109 ) ;
  assign n765 = ~n763 & n764 ;
  assign n766 = n762 | n765 ;
  assign n767 = ~x129 & n766 ;
  assign n768 = x82 & n244 ;
  assign n769 = n259 | n433 ;
  assign n770 = n238 | n550 ;
  assign n771 = n769 | n770 ;
  assign n772 = x82 & n771 ;
  assign n773 = n232 & ~n772 ;
  assign n774 = n768 | n773 ;
  assign n775 = ~x38 & n774 ;
  assign n776 = x2 | x48 ;
  assign n777 = n251 | n776 ;
  assign n778 = n254 | n777 ;
  assign n779 = x50 | n244 ;
  assign n780 = n491 | n779 ;
  assign n781 = n778 | n780 ;
  assign n782 = x82 & n781 ;
  assign n783 = n232 | n782 ;
  assign n784 = x74 & ~n783 ;
  assign n785 = ~x44 & x82 ;
  assign n786 = x38 & ~n494 ;
  assign n787 = n785 & n786 ;
  assign n788 = x129 | n787 ;
  assign n789 = n784 | n788 ;
  assign n790 = n775 | n789 ;
  assign n791 = ~x51 & x109 ;
  assign n792 = ~n591 & n791 ;
  assign n793 = x106 | n792 ;
  assign n794 = x109 & ~n568 ;
  assign n795 = x39 & ~n794 ;
  assign n796 = n793 | n795 ;
  assign n797 = ~x129 & n796 ;
  assign n798 = x82 & n243 ;
  assign n799 = n433 | n770 ;
  assign n800 = n242 | n799 ;
  assign n801 = x82 & n800 ;
  assign n802 = n232 & ~n801 ;
  assign n803 = n798 | n802 ;
  assign n804 = ~x40 & n803 ;
  assign n805 = n241 | n243 ;
  assign n806 = n491 | n805 ;
  assign n807 = n778 | n806 ;
  assign n808 = x82 & n807 ;
  assign n809 = n232 | n808 ;
  assign n810 = x73 & ~n809 ;
  assign n811 = x40 & x82 ;
  assign n812 = ~n243 & n811 ;
  assign n813 = x129 | n812 ;
  assign n814 = n810 | n813 ;
  assign n815 = n804 | n814 ;
  assign n816 = x82 & n427 ;
  assign n817 = x82 & n799 ;
  assign n818 = n232 & ~n817 ;
  assign n819 = n816 | n818 ;
  assign n820 = ~x41 & n819 ;
  assign n821 = x82 & n257 ;
  assign n822 = n234 | n258 ;
  assign n823 = n778 | n822 ;
  assign n824 = ( x82 & n821 ) | ( x82 & n823 ) | ( n821 & n823 ) ;
  assign n825 = n232 | n824 ;
  assign n826 = x76 & ~n825 ;
  assign n827 = n256 | n258 ;
  assign n828 = x41 & x82 ;
  assign n829 = ~n243 & n828 ;
  assign n830 = ~n827 & n829 ;
  assign n831 = x129 | n830 ;
  assign n832 = n826 | n831 ;
  assign n833 = n820 | n832 ;
  assign n834 = x44 & x82 ;
  assign n835 = n541 | n827 ;
  assign n836 = n778 | n835 ;
  assign n837 = x82 & n836 ;
  assign n838 = n232 & ~n837 ;
  assign n839 = n834 | n838 ;
  assign n840 = ~x42 & n839 ;
  assign n841 = x44 | n502 ;
  assign n842 = n491 | n841 ;
  assign n843 = n778 | n842 ;
  assign n844 = x82 & n843 ;
  assign n845 = n232 | n844 ;
  assign n846 = x72 & ~n845 ;
  assign n847 = x42 & n785 ;
  assign n848 = x129 | n847 ;
  assign n849 = n846 | n848 ;
  assign n850 = n840 | n849 ;
  assign n851 = x82 & n260 ;
  assign n852 = n238 | n551 ;
  assign n853 = x82 & n852 ;
  assign n854 = n232 & ~n853 ;
  assign n855 = n851 | n854 ;
  assign n856 = ~x43 & n855 ;
  assign n857 = x47 | n778 ;
  assign n858 = ( x82 & n851 ) | ( x82 & n857 ) | ( n851 & n857 ) ;
  assign n859 = n232 | n858 ;
  assign n860 = x77 & ~n859 ;
  assign n861 = x43 & ~n494 ;
  assign n862 = n785 & n861 ;
  assign n863 = ~n242 & n862 ;
  assign n864 = x129 | n863 ;
  assign n865 = n860 | n864 ;
  assign n866 = n856 | n865 ;
  assign n867 = x129 | n834 ;
  assign n868 = n491 | n495 ;
  assign n869 = n778 | n868 ;
  assign n870 = x82 & n869 ;
  assign n871 = ( x44 & n232 ) | ( x44 & n870 ) | ( n232 & n870 ) ;
  assign n872 = ( x67 & n232 ) | ( x67 & ~n870 ) | ( n232 & ~n870 ) ;
  assign n873 = ~n871 & n872 ;
  assign n874 = n867 | n873 ;
  assign n875 = n252 | n557 ;
  assign n876 = n241 | n244 ;
  assign n877 = n875 | n876 ;
  assign n878 = x82 & n877 ;
  assign n879 = x24 | n545 ;
  assign n880 = x82 & n879 ;
  assign n881 = n232 & ~n880 ;
  assign n882 = n878 | n881 ;
  assign n883 = ~x45 & n882 ;
  assign n884 = x2 | n252 ;
  assign n885 = n238 | n884 ;
  assign n886 = n261 | n885 ;
  assign n887 = x82 & n886 ;
  assign n888 = n232 | n887 ;
  assign n889 = x68 & ~n888 ;
  assign n890 = x38 | n494 ;
  assign n891 = x45 & ~n890 ;
  assign n892 = n785 & n891 ;
  assign n893 = ~n769 & n892 ;
  assign n894 = x129 | n893 ;
  assign n895 = n889 | n894 ;
  assign n896 = n883 | n895 ;
  assign n897 = x82 & n876 ;
  assign n898 = n541 | n778 ;
  assign n899 = x82 & n898 ;
  assign n900 = n232 & ~n899 ;
  assign n901 = n897 | n900 ;
  assign n902 = ~x46 & n901 ;
  assign n903 = x50 | n257 ;
  assign n904 = n898 | n903 ;
  assign n905 = x82 & n904 ;
  assign n906 = n232 | n905 ;
  assign n907 = x75 & ~n906 ;
  assign n908 = x46 & x82 ;
  assign n909 = ~n903 & n908 ;
  assign n910 = x129 | n909 ;
  assign n911 = n907 | n910 ;
  assign n912 = n902 | n911 ;
  assign n913 = x82 & n261 ;
  assign n914 = x82 & n778 ;
  assign n915 = n232 & ~n914 ;
  assign n916 = n913 | n915 ;
  assign n917 = ~x47 & n916 ;
  assign n918 = n261 | n778 ;
  assign n919 = x82 & n918 ;
  assign n920 = n232 | n919 ;
  assign n921 = x64 & ~n920 ;
  assign n922 = n422 | n426 ;
  assign n923 = x47 & ~n494 ;
  assign n924 = n785 & n923 ;
  assign n925 = ~n922 & n924 ;
  assign n926 = x129 | n925 ;
  assign n927 = n921 | n926 ;
  assign n928 = n917 | n927 ;
  assign n929 = n491 | n876 ;
  assign n930 = x82 & n929 ;
  assign n931 = x82 & n770 ;
  assign n932 = n232 & ~n931 ;
  assign n933 = n930 | n932 ;
  assign n934 = ~x48 & n933 ;
  assign n935 = x2 | x47 ;
  assign n936 = n251 | n254 ;
  assign n937 = n935 | n936 ;
  assign n938 = ( x82 & n913 ) | ( x82 & n937 ) | ( n913 & n937 ) ;
  assign n939 = n232 | n938 ;
  assign n940 = x62 & ~n939 ;
  assign n941 = n234 | n259 ;
  assign n942 = x48 & ~n890 ;
  assign n943 = n785 & n942 ;
  assign n944 = ~n941 & n943 ;
  assign n945 = x129 | n944 ;
  assign n946 = n940 | n945 ;
  assign n947 = n934 | n946 ;
  assign n948 = n237 | n903 ;
  assign n949 = n558 | n948 ;
  assign n950 = x82 & n949 ;
  assign n951 = n232 | n950 ;
  assign n952 = x69 | n951 ;
  assign n953 = x24 | x42 ;
  assign n954 = n841 | n953 ;
  assign n955 = n558 | n954 ;
  assign n956 = x49 & n955 ;
  assign n957 = x2 | n236 ;
  assign n958 = ~n948 & n957 ;
  assign n959 = ~n491 & n958 ;
  assign n960 = ~n233 & n959 ;
  assign n961 = n956 | n960 ;
  assign n962 = x82 & n961 ;
  assign n963 = x49 & n264 ;
  assign n964 = n962 | n963 ;
  assign n965 = n952 & ~n964 ;
  assign n966 = x129 | n965 ;
  assign n967 = n557 | n884 ;
  assign n968 = n936 | n967 ;
  assign n969 = x82 & n968 ;
  assign n970 = n232 & ~n969 ;
  assign n971 = n821 | n970 ;
  assign n972 = ~x50 & n971 ;
  assign n973 = n491 | n778 ;
  assign n974 = ( x82 & n821 ) | ( x82 & n973 ) | ( n821 & n973 ) ;
  assign n975 = n232 | n974 ;
  assign n976 = x66 & ~n975 ;
  assign n977 = x50 & ~n890 ;
  assign n978 = n785 & n977 ;
  assign n979 = x129 | n978 ;
  assign n980 = n976 | n979 ;
  assign n981 = n972 | n980 ;
  assign n982 = x51 & ~x109 ;
  assign n983 = ( ~x51 & x106 ) | ( ~x51 & x109 ) | ( x106 & x109 ) ;
  assign n984 = ( ~x129 & n982 ) | ( ~x129 & n983 ) | ( n982 & n983 ) ;
  assign n985 = x52 & ~n791 ;
  assign n986 = x106 | n794 ;
  assign n987 = n985 | n986 ;
  assign n988 = ~x129 & n987 ;
  assign n989 = x58 & x116 ;
  assign n990 = x58 | x110 ;
  assign n991 = x96 | n990 ;
  assign n992 = n572 | n991 ;
  assign n993 = ~n989 & n992 ;
  assign n994 = x53 | n993 ;
  assign n995 = x97 & ~n994 ;
  assign n996 = ~x116 & n712 ;
  assign n997 = n995 | n996 ;
  assign n998 = ~x129 & n997 ;
  assign n999 = ~x3 & n998 ;
  assign n1000 = ~n602 & n999 ;
  assign n1001 = ~x26 & n1000 ;
  assign n1002 = n261 | n852 ;
  assign n1003 = x82 & n1002 ;
  assign n1004 = n232 | n1003 ;
  assign n1005 = ~x129 & n1004 ;
  assign n1006 = x123 | x129 ;
  assign n1007 = x114 & ~x122 ;
  assign n1008 = ~n1006 & n1007 ;
  assign n1009 = x58 & ~x116 ;
  assign n1010 = ~x26 & x58 ;
  assign n1011 = x37 & ~x116 ;
  assign n1012 = n1010 | n1011 ;
  assign n1013 = ~n1009 & n1012 ;
  assign n1014 = x26 & ~x58 ;
  assign n1015 = ( x58 & x94 ) | ( x58 & n571 ) | ( x94 & n571 ) ;
  assign n1016 = ( ~x26 & n1014 ) | ( ~x26 & n1015 ) | ( n1014 & n1015 ) ;
  assign n1017 = n1013 | n1016 ;
  assign n1018 = ~x53 & n1017 ;
  assign n1019 = ~x26 & x37 ;
  assign n1020 = ~x58 & n1019 ;
  assign n1021 = n1018 | n1020 ;
  assign n1022 = ~x85 & n1021 ;
  assign n1023 = ~n641 & n1019 ;
  assign n1024 = n1022 | n1023 ;
  assign n1025 = ~x27 & n1024 ;
  assign n1026 = x85 | n641 ;
  assign n1027 = n1019 & ~n1026 ;
  assign n1028 = n1025 | n1027 ;
  assign n1029 = ~x129 & n1028 ;
  assign n1030 = ~x3 & n1029 ;
  assign n1031 = x26 | x53 ;
  assign n1032 = x85 | n1031 ;
  assign n1033 = x116 | n1032 ;
  assign n1034 = ( x26 & x53 ) | ( x26 & x85 ) | ( x53 & x85 ) ;
  assign n1035 = x58 | n1034 ;
  assign n1036 = n1033 & n1035 ;
  assign n1037 = x57 & ~n1036 ;
  assign n1038 = x60 & n989 ;
  assign n1039 = ~n1032 & n1038 ;
  assign n1040 = n1037 | n1039 ;
  assign n1041 = ~x27 & n1040 ;
  assign n1042 = x57 & ~x58 ;
  assign n1043 = ~n1032 & n1042 ;
  assign n1044 = n1041 | n1043 ;
  assign n1045 = ~x129 & n1044 ;
  assign n1046 = ~x3 & n1045 ;
  assign n1047 = ~n579 & n1009 ;
  assign n1048 = x116 & n652 ;
  assign n1049 = ~x58 & n1048 ;
  assign n1050 = ~n659 & n1049 ;
  assign n1051 = n1047 | n1050 ;
  assign n1052 = ~x129 & n1051 ;
  assign n1053 = ~x3 & n1052 ;
  assign n1054 = ~x53 & n1053 ;
  assign n1055 = ~x85 & n1054 ;
  assign n1056 = ( x53 & x58 ) | ( x53 & x116 ) | ( x58 & x116 ) ;
  assign n1057 = n641 & ~n1056 ;
  assign n1058 = ( n574 & n1056 ) | ( n574 & ~n1057 ) | ( n1056 & ~n1057 ) ;
  assign n1059 = x59 & ~n1058 ;
  assign n1060 = x96 & ~n641 ;
  assign n1061 = n574 & n1060 ;
  assign n1062 = ~x85 & n1061 ;
  assign n1063 = ( ~x85 & n1059 ) | ( ~x85 & n1062 ) | ( n1059 & n1062 ) ;
  assign n1064 = x59 & ~x116 ;
  assign n1065 = x27 & ~x85 ;
  assign n1066 = ~n641 & n1065 ;
  assign n1067 = n1064 & n1066 ;
  assign n1068 = x85 & ~n641 ;
  assign n1069 = n1064 & n1068 ;
  assign n1070 = ~x27 & n1069 ;
  assign n1071 = n1067 | n1070 ;
  assign n1072 = x27 & ~n1067 ;
  assign n1073 = ( n1063 & n1071 ) | ( n1063 & ~n1072 ) | ( n1071 & ~n1072 ) ;
  assign n1074 = x26 & n1064 ;
  assign n1075 = ~n693 & n1074 ;
  assign n1076 = x26 & ~n1075 ;
  assign n1077 = x129 | n1076 ;
  assign n1078 = x3 | n1077 ;
  assign n1079 = ~x129 & n1075 ;
  assign n1080 = ~x3 & n1079 ;
  assign n1081 = ( n1073 & ~n1078 ) | ( n1073 & n1080 ) | ( ~n1078 & n1080 ) ;
  assign n1082 = x117 | x122 ;
  assign n1083 = x60 & n1082 ;
  assign n1084 = x123 & ~n1082 ;
  assign n1085 = n1083 | n1084 ;
  assign n1086 = ~x114 & x123 ;
  assign n1087 = ~x122 & n1086 ;
  assign n1088 = ~x129 & n1087 ;
  assign n1089 = x136 & ~x137 ;
  assign n1090 = x132 & x133 ;
  assign n1091 = x131 & n1090 ;
  assign n1092 = ( x138 & n1089 ) | ( x138 & ~n1091 ) | ( n1089 & ~n1091 ) ;
  assign n1093 = n1089 & ~n1092 ;
  assign n1094 = x62 & ~n1093 ;
  assign n1095 = ~x140 & n1089 ;
  assign n1096 = ~x138 & n1091 ;
  assign n1097 = n1095 & n1096 ;
  assign n1098 = n1094 | n1097 ;
  assign n1099 = ~x129 & n1098 ;
  assign n1100 = x63 & ~n1093 ;
  assign n1101 = ~x142 & n1089 ;
  assign n1102 = n1096 & n1101 ;
  assign n1103 = n1100 | n1102 ;
  assign n1104 = ~x129 & n1103 ;
  assign n1105 = x64 & ~n1093 ;
  assign n1106 = ~x139 & n1089 ;
  assign n1107 = n1096 & n1106 ;
  assign n1108 = n1105 | n1107 ;
  assign n1109 = ~x129 & n1108 ;
  assign n1110 = x65 & ~n1093 ;
  assign n1111 = ~x146 & n1089 ;
  assign n1112 = n1096 & n1111 ;
  assign n1113 = n1110 | n1112 ;
  assign n1114 = ~x129 & n1113 ;
  assign n1115 = x136 | x137 ;
  assign n1116 = n1096 & ~n1115 ;
  assign n1117 = ( x129 & x143 ) | ( x129 & n1116 ) | ( x143 & n1116 ) ;
  assign n1118 = ( x66 & ~x129 ) | ( x66 & n1116 ) | ( ~x129 & n1116 ) ;
  assign n1119 = ~n1117 & n1118 ;
  assign n1120 = ( x129 & x139 ) | ( x129 & n1116 ) | ( x139 & n1116 ) ;
  assign n1121 = ( x67 & ~x129 ) | ( x67 & n1116 ) | ( ~x129 & n1116 ) ;
  assign n1122 = ~n1120 & n1121 ;
  assign n1123 = x68 & ~n1093 ;
  assign n1124 = ~x141 & n1089 ;
  assign n1125 = n1096 & n1124 ;
  assign n1126 = n1123 | n1125 ;
  assign n1127 = ~x129 & n1126 ;
  assign n1128 = x69 & ~n1093 ;
  assign n1129 = ~x143 & n1089 ;
  assign n1130 = n1096 & n1129 ;
  assign n1131 = n1128 | n1130 ;
  assign n1132 = ~x129 & n1131 ;
  assign n1133 = x70 & ~n1093 ;
  assign n1134 = ~x144 & n1089 ;
  assign n1135 = n1096 & n1134 ;
  assign n1136 = n1133 | n1135 ;
  assign n1137 = ~x129 & n1136 ;
  assign n1138 = x71 & ~n1093 ;
  assign n1139 = ~x145 & n1089 ;
  assign n1140 = n1096 & n1139 ;
  assign n1141 = n1138 | n1140 ;
  assign n1142 = ~x129 & n1141 ;
  assign n1143 = ( x129 & x140 ) | ( x129 & n1116 ) | ( x140 & n1116 ) ;
  assign n1144 = ( x72 & ~x129 ) | ( x72 & n1116 ) | ( ~x129 & n1116 ) ;
  assign n1145 = ~n1143 & n1144 ;
  assign n1146 = ( x129 & x141 ) | ( x129 & n1116 ) | ( x141 & n1116 ) ;
  assign n1147 = ( x73 & ~x129 ) | ( x73 & n1116 ) | ( ~x129 & n1116 ) ;
  assign n1148 = ~n1146 & n1147 ;
  assign n1149 = ( x129 & x142 ) | ( x129 & n1116 ) | ( x142 & n1116 ) ;
  assign n1150 = ( x74 & ~x129 ) | ( x74 & n1116 ) | ( ~x129 & n1116 ) ;
  assign n1151 = ~n1149 & n1150 ;
  assign n1152 = ( x129 & x144 ) | ( x129 & n1116 ) | ( x144 & n1116 ) ;
  assign n1153 = ( x75 & ~x129 ) | ( x75 & n1116 ) | ( ~x129 & n1116 ) ;
  assign n1154 = ~n1152 & n1153 ;
  assign n1155 = ( x129 & x145 ) | ( x129 & n1116 ) | ( x145 & n1116 ) ;
  assign n1156 = ( x76 & ~x129 ) | ( x76 & n1116 ) | ( ~x129 & n1116 ) ;
  assign n1157 = ~n1155 & n1156 ;
  assign n1158 = ( x129 & x146 ) | ( x129 & n1116 ) | ( x146 & n1116 ) ;
  assign n1159 = ( x77 & ~x129 ) | ( x77 & n1116 ) | ( ~x129 & n1116 ) ;
  assign n1160 = ~n1158 & n1159 ;
  assign n1161 = ~x136 & x137 ;
  assign n1162 = n1096 & n1161 ;
  assign n1163 = ( x129 & ~x142 ) | ( x129 & n1162 ) | ( ~x142 & n1162 ) ;
  assign n1164 = ( x78 & ~x129 ) | ( x78 & n1162 ) | ( ~x129 & n1162 ) ;
  assign n1165 = ~n1163 & n1164 ;
  assign n1166 = ( x129 & ~x143 ) | ( x129 & n1162 ) | ( ~x143 & n1162 ) ;
  assign n1167 = ( x79 & ~x129 ) | ( x79 & n1162 ) | ( ~x129 & n1162 ) ;
  assign n1168 = ~n1166 & n1167 ;
  assign n1169 = ( x129 & ~x144 ) | ( x129 & n1162 ) | ( ~x144 & n1162 ) ;
  assign n1170 = ( x80 & ~x129 ) | ( x80 & n1162 ) | ( ~x129 & n1162 ) ;
  assign n1171 = ~n1169 & n1170 ;
  assign n1172 = ( x129 & ~x145 ) | ( x129 & n1162 ) | ( ~x145 & n1162 ) ;
  assign n1173 = ( x81 & ~x129 ) | ( x81 & n1162 ) | ( ~x129 & n1162 ) ;
  assign n1174 = ~n1172 & n1173 ;
  assign n1175 = ( x129 & ~x146 ) | ( x129 & n1162 ) | ( ~x146 & n1162 ) ;
  assign n1176 = ( x82 & ~x129 ) | ( x82 & n1162 ) | ( ~x129 & n1162 ) ;
  assign n1177 = ~n1175 & n1176 ;
  assign n1178 = ( x89 & x136 ) | ( x89 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1179 = ( ~x62 & x136 ) | ( ~x62 & x138 ) | ( x136 & x138 ) ;
  assign n1180 = n1178 & n1179 ;
  assign n1181 = ( ~x119 & x136 ) | ( ~x119 & x138 ) | ( x136 & x138 ) ;
  assign n1182 = ( x72 & x136 ) | ( x72 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1183 = n1181 | n1182 ;
  assign n1184 = ~n1180 & n1183 ;
  assign n1185 = x137 | n1184 ;
  assign n1186 = x136 & ~x138 ;
  assign n1187 = x31 & n1186 ;
  assign n1188 = ( x115 & x136 ) | ( x115 & x138 ) | ( x136 & x138 ) ;
  assign n1189 = ( x87 & ~x136 ) | ( x87 & x138 ) | ( ~x136 & x138 ) ;
  assign n1190 = ~n1188 & n1189 ;
  assign n1191 = n1187 | n1190 ;
  assign n1192 = x137 & n1191 ;
  assign n1193 = n1185 & ~n1192 ;
  assign n1194 = ( x129 & ~x141 ) | ( x129 & n1162 ) | ( ~x141 & n1162 ) ;
  assign n1195 = ( x84 & ~x129 ) | ( x84 & n1162 ) | ( ~x129 & n1162 ) ;
  assign n1196 = ~n1194 & n1195 ;
  assign n1197 = ( x97 & n572 ) | ( x97 & ~n580 ) | ( n572 & ~n580 ) ;
  assign n1198 = ~n580 & n1197 ;
  assign n1199 = x96 & n1198 ;
  assign n1200 = n615 | n1199 ;
  assign n1201 = ~x129 & n1200 ;
  assign n1202 = ~x3 & n1201 ;
  assign n1203 = ~n628 & n1202 ;
  assign n1204 = ~x26 & n1203 ;
  assign n1205 = ( x129 & ~x139 ) | ( x129 & n1162 ) | ( ~x139 & n1162 ) ;
  assign n1206 = ( x86 & ~x129 ) | ( x86 & n1162 ) | ( ~x129 & n1162 ) ;
  assign n1207 = ~n1205 & n1206 ;
  assign n1208 = ( x129 & ~x140 ) | ( x129 & n1162 ) | ( ~x140 & n1162 ) ;
  assign n1209 = ( x87 & ~x129 ) | ( x87 & n1162 ) | ( ~x129 & n1162 ) ;
  assign n1210 = ~n1208 & n1209 ;
  assign n1211 = x136 & x137 ;
  assign n1212 = n1096 & n1211 ;
  assign n1213 = ( x129 & ~x139 ) | ( x129 & n1212 ) | ( ~x139 & n1212 ) ;
  assign n1214 = ( x88 & ~x129 ) | ( x88 & n1212 ) | ( ~x129 & n1212 ) ;
  assign n1215 = ~n1213 & n1214 ;
  assign n1216 = ( x129 & ~x140 ) | ( x129 & n1212 ) | ( ~x140 & n1212 ) ;
  assign n1217 = ( x89 & ~x129 ) | ( x89 & n1212 ) | ( ~x129 & n1212 ) ;
  assign n1218 = ~n1216 & n1217 ;
  assign n1219 = ( x129 & ~x142 ) | ( x129 & n1212 ) | ( ~x142 & n1212 ) ;
  assign n1220 = ( x90 & ~x129 ) | ( x90 & n1212 ) | ( ~x129 & n1212 ) ;
  assign n1221 = ~n1219 & n1220 ;
  assign n1222 = ( x129 & ~x143 ) | ( x129 & n1212 ) | ( ~x143 & n1212 ) ;
  assign n1223 = ( x91 & ~x129 ) | ( x91 & n1212 ) | ( ~x129 & n1212 ) ;
  assign n1224 = ~n1222 & n1223 ;
  assign n1225 = ( x129 & ~x144 ) | ( x129 & n1212 ) | ( ~x144 & n1212 ) ;
  assign n1226 = ( x92 & ~x129 ) | ( x92 & n1212 ) | ( ~x129 & n1212 ) ;
  assign n1227 = ~n1225 & n1226 ;
  assign n1228 = ( x129 & ~x146 ) | ( x129 & n1212 ) | ( ~x146 & n1212 ) ;
  assign n1229 = ( x93 & ~x129 ) | ( x93 & n1212 ) | ( ~x129 & n1212 ) ;
  assign n1230 = ~n1228 & n1229 ;
  assign n1231 = x138 & n1091 ;
  assign n1232 = x82 & ~n1115 ;
  assign n1233 = n1231 & n1232 ;
  assign n1234 = ( x129 & ~x142 ) | ( x129 & n1233 ) | ( ~x142 & n1233 ) ;
  assign n1235 = ( x94 & ~x129 ) | ( x94 & n1233 ) | ( ~x129 & n1233 ) ;
  assign n1236 = ~n1234 & n1235 ;
  assign n1237 = x3 | n1091 ;
  assign n1238 = x110 | n1237 ;
  assign n1239 = x138 & n1232 ;
  assign n1240 = n1091 & ~n1239 ;
  assign n1241 = n1238 & ~n1240 ;
  assign n1242 = x95 & ~n1241 ;
  assign n1243 = x143 & n1233 ;
  assign n1244 = n1242 | n1243 ;
  assign n1245 = ~x129 & n1244 ;
  assign n1246 = x96 & ~n1241 ;
  assign n1247 = x146 & n1233 ;
  assign n1248 = n1246 | n1247 ;
  assign n1249 = ~x129 & n1248 ;
  assign n1250 = x97 & ~n1241 ;
  assign n1251 = x145 & n1233 ;
  assign n1252 = n1250 | n1251 ;
  assign n1253 = ~x129 & n1252 ;
  assign n1254 = ( x129 & ~x145 ) | ( x129 & n1212 ) | ( ~x145 & n1212 ) ;
  assign n1255 = ( x98 & ~x129 ) | ( x98 & n1212 ) | ( ~x129 & n1212 ) ;
  assign n1256 = ~n1254 & n1255 ;
  assign n1257 = ( x129 & ~x141 ) | ( x129 & n1212 ) | ( ~x141 & n1212 ) ;
  assign n1258 = ( x99 & ~x129 ) | ( x99 & n1212 ) | ( ~x129 & n1212 ) ;
  assign n1259 = ~n1257 & n1258 ;
  assign n1260 = x100 & ~n1241 ;
  assign n1261 = x144 & n1233 ;
  assign n1262 = n1260 | n1261 ;
  assign n1263 = ~x129 & n1262 ;
  assign n1264 = ( ~x124 & x136 ) | ( ~x124 & x138 ) | ( x136 & x138 ) ;
  assign n1265 = ( x77 & x136 ) | ( x77 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1266 = n1264 | n1265 ;
  assign n1267 = ( x93 & x136 ) | ( x93 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1268 = ( ~x65 & x136 ) | ( ~x65 & x138 ) | ( x136 & x138 ) ;
  assign n1269 = n1267 & n1268 ;
  assign n1270 = n1266 & ~n1269 ;
  assign n1271 = x137 | n1270 ;
  assign n1272 = x37 & n1186 ;
  assign n1273 = ( ~x96 & x136 ) | ( ~x96 & x138 ) | ( x136 & x138 ) ;
  assign n1274 = ( x82 & ~x136 ) | ( x82 & x138 ) | ( ~x136 & x138 ) ;
  assign n1275 = ~n1273 & n1274 ;
  assign n1276 = n1272 | n1275 ;
  assign n1277 = x137 & n1276 ;
  assign n1278 = n1271 & ~n1277 ;
  assign n1279 = x91 & n1089 ;
  assign n1280 = x95 & n1161 ;
  assign n1281 = n1279 | n1280 ;
  assign n1282 = x138 & n1281 ;
  assign n1283 = ( x79 & x136 ) | ( x79 & x137 ) | ( x136 & x137 ) ;
  assign n1284 = ( x34 & ~x136 ) | ( x34 & x137 ) | ( ~x136 & x137 ) ;
  assign n1285 = n1283 & n1284 ;
  assign n1286 = ( x69 & x136 ) | ( x69 & x137 ) | ( x136 & x137 ) ;
  assign n1287 = ( x66 & ~x136 ) | ( x66 & x137 ) | ( ~x136 & x137 ) ;
  assign n1288 = n1286 | n1287 ;
  assign n1289 = ~n1285 & n1288 ;
  assign n1290 = x138 | n1289 ;
  assign n1291 = ~n1282 & n1290 ;
  assign n1292 = x90 & n1089 ;
  assign n1293 = x94 & n1161 ;
  assign n1294 = n1292 | n1293 ;
  assign n1295 = x138 & n1294 ;
  assign n1296 = ( x78 & x136 ) | ( x78 & x137 ) | ( x136 & x137 ) ;
  assign n1297 = ( x33 & ~x136 ) | ( x33 & x137 ) | ( ~x136 & x137 ) ;
  assign n1298 = n1296 & n1297 ;
  assign n1299 = ( x63 & x136 ) | ( x63 & x137 ) | ( x136 & x137 ) ;
  assign n1300 = ( x74 & ~x136 ) | ( x74 & x137 ) | ( ~x136 & x137 ) ;
  assign n1301 = n1299 | n1300 ;
  assign n1302 = ~n1298 & n1301 ;
  assign n1303 = x138 | n1302 ;
  assign n1304 = ~n1295 & n1303 ;
  assign n1305 = x99 & n1089 ;
  assign n1306 = ~x112 & n1161 ;
  assign n1307 = n1305 | n1306 ;
  assign n1308 = x138 & n1307 ;
  assign n1309 = ( x68 & x136 ) | ( x68 & x137 ) | ( x136 & x137 ) ;
  assign n1310 = ( x73 & ~x136 ) | ( x73 & x137 ) | ( ~x136 & x137 ) ;
  assign n1311 = n1309 | n1310 ;
  assign n1312 = ( x84 & x136 ) | ( x84 & x137 ) | ( x136 & x137 ) ;
  assign n1313 = ( x32 & ~x136 ) | ( x32 & x137 ) | ( ~x136 & x137 ) ;
  assign n1314 = n1312 & n1313 ;
  assign n1315 = n1311 & ~n1314 ;
  assign n1316 = x138 | n1315 ;
  assign n1317 = ~n1308 & n1316 ;
  assign n1318 = ( x92 & x136 ) | ( x92 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1319 = ( ~x70 & x136 ) | ( ~x70 & x138 ) | ( x136 & x138 ) ;
  assign n1320 = n1318 & n1319 ;
  assign n1321 = ( ~x125 & x136 ) | ( ~x125 & x138 ) | ( x136 & x138 ) ;
  assign n1322 = ( x75 & x136 ) | ( x75 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1323 = n1321 | n1322 ;
  assign n1324 = ~n1320 & n1323 ;
  assign n1325 = x137 | n1324 ;
  assign n1326 = x35 & n1186 ;
  assign n1327 = ( ~x100 & x136 ) | ( ~x100 & x138 ) | ( x136 & x138 ) ;
  assign n1328 = ( x80 & ~x136 ) | ( x80 & x138 ) | ( ~x136 & x138 ) ;
  assign n1329 = ~n1327 & n1328 ;
  assign n1330 = n1326 | n1329 ;
  assign n1331 = x137 & n1330 ;
  assign n1332 = n1325 & ~n1331 ;
  assign n1333 = ~n642 & n1198 ;
  assign n1334 = ~x27 & n1333 ;
  assign n1335 = n582 | n1334 ;
  assign n1336 = ~x129 & n1335 ;
  assign n1337 = ~x3 & n1336 ;
  assign n1338 = ( x98 & x136 ) | ( x98 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1339 = ( ~x71 & x136 ) | ( ~x71 & x138 ) | ( x136 & x138 ) ;
  assign n1340 = n1338 & n1339 ;
  assign n1341 = ( ~x23 & x136 ) | ( ~x23 & x138 ) | ( x136 & x138 ) ;
  assign n1342 = ( x76 & x136 ) | ( x76 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1343 = n1341 | n1342 ;
  assign n1344 = ~n1340 & n1343 ;
  assign n1345 = x137 | n1344 ;
  assign n1346 = x36 & n1186 ;
  assign n1347 = ( ~x97 & x136 ) | ( ~x97 & x138 ) | ( x136 & x138 ) ;
  assign n1348 = ( x81 & ~x136 ) | ( x81 & x138 ) | ( ~x136 & x138 ) ;
  assign n1349 = ~n1347 & n1348 ;
  assign n1350 = n1346 | n1349 ;
  assign n1351 = x137 & n1350 ;
  assign n1352 = n1345 & ~n1351 ;
  assign n1353 = ( x88 & x136 ) | ( x88 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1354 = ( ~x64 & x136 ) | ( ~x64 & x138 ) | ( x136 & x138 ) ;
  assign n1355 = n1353 & n1354 ;
  assign n1356 = ( ~x120 & x136 ) | ( ~x120 & x138 ) | ( x136 & x138 ) ;
  assign n1357 = ( x67 & x136 ) | ( x67 & ~x138 ) | ( x136 & ~x138 ) ;
  assign n1358 = n1356 | n1357 ;
  assign n1359 = ~n1355 & n1358 ;
  assign n1360 = x137 | n1359 ;
  assign n1361 = x30 & n1186 ;
  assign n1362 = ( ~x111 & x136 ) | ( ~x111 & x138 ) | ( x136 & x138 ) ;
  assign n1363 = ( x86 & ~x136 ) | ( x86 & x138 ) | ( ~x136 & x138 ) ;
  assign n1364 = ~n1362 & n1363 ;
  assign n1365 = n1361 | n1364 ;
  assign n1366 = x137 & n1365 ;
  assign n1367 = n1360 & ~n1366 ;
  assign n1368 = n651 & n659 ;
  assign n1369 = n650 | n1368 ;
  assign n1370 = ~x129 & n1369 ;
  assign n1371 = ~x3 & n1370 ;
  assign n1372 = x116 & n1371 ;
  assign n1373 = ~x97 & n603 ;
  assign n1374 = n712 | n1373 ;
  assign n1375 = ~x129 & n1374 ;
  assign n1376 = ~x3 & n1375 ;
  assign n1377 = x116 & n1376 ;
  assign n1378 = x111 & ~n1239 ;
  assign n1379 = ~x136 & x139 ;
  assign n1380 = ~x137 & x138 ;
  assign n1381 = x82 & n1380 ;
  assign n1382 = n1379 & n1381 ;
  assign n1383 = n1378 | n1382 ;
  assign n1384 = n1091 & n1383 ;
  assign n1385 = ~x129 & n1384 ;
  assign n1386 = ~x136 & x141 ;
  assign n1387 = n1381 & n1386 ;
  assign n1388 = x112 | n1239 ;
  assign n1389 = ~n1387 & n1388 ;
  assign n1390 = n1091 & ~n1389 ;
  assign n1391 = ~x129 & n1390 ;
  assign n1392 = ( ~x54 & x113 ) | ( ~x54 & x129 ) | ( x113 & x129 ) ;
  assign n1393 = x11 | x22 ;
  assign n1394 = ( x54 & x129 ) | ( x54 & ~n1393 ) | ( x129 & ~n1393 ) ;
  assign n1395 = n1392 | n1394 ;
  assign n1396 = x3 | n1395 ;
  assign n1397 = ~x136 & x140 ;
  assign n1398 = n1381 & n1397 ;
  assign n1399 = x115 | n1239 ;
  assign n1400 = ~n1398 & n1399 ;
  assign n1401 = n1091 & ~n1400 ;
  assign n1402 = ~x129 & n1401 ;
  assign n1403 = x4 | x12 ;
  assign n1404 = x7 | x9 ;
  assign n1405 = n1403 | n1404 ;
  assign n1406 = ~x129 & n1405 ;
  assign n1407 = ~x3 & n1406 ;
  assign n1408 = x54 & n1407 ;
  assign n1409 = x122 & ~x129 ;
  assign n1410 = ~x54 & x118 ;
  assign n1411 = x54 & ~x59 ;
  assign n1412 = n403 & n1411 ;
  assign n1413 = n1410 | n1412 ;
  assign n1414 = ~x129 & n1413 ;
  assign n1415 = ~x129 & n572 ;
  assign n1416 = x110 | x120 ;
  assign n1417 = x3 | n1416 ;
  assign n1418 = ~x129 & n1417 ;
  assign n1419 = ~x111 & n1418 ;
  assign n1420 = x81 & x120 ;
  assign n1421 = ~x129 & n1420 ;
  assign n1422 = x129 | x134 ;
  assign n1423 = x129 | x135 ;
  assign n1424 = x57 & ~x129 ;
  assign n1425 = ~x96 & x125 ;
  assign n1426 = x3 | n1425 ;
  assign n1427 = ~x129 & n1426 ;
  assign n1428 = ~x126 & n1090 ;
  assign y0 = x108 ;
  assign y1 = x83 ;
  assign y2 = x104 ;
  assign y3 = x103 ;
  assign y4 = x102 ;
  assign y5 = x105 ;
  assign y6 = x107 ;
  assign y7 = x101 ;
  assign y8 = x126 ;
  assign y9 = x121 ;
  assign y10 = x1 ;
  assign y11 = x0 ;
  assign y12 = ~1'b0 ;
  assign y13 = x130 ;
  assign y14 = x128 ;
  assign y15 = n195 ;
  assign y16 = n231 ;
  assign y17 = ~n268 ;
  assign y18 = n282 ;
  assign y19 = n292 ;
  assign y20 = n310 ;
  assign y21 = n324 ;
  assign y22 = n338 ;
  assign y23 = n350 ;
  assign y24 = n363 ;
  assign y25 = n375 ;
  assign y26 = n386 ;
  assign y27 = n397 ;
  assign y28 = n410 ;
  assign y29 = n421 ;
  assign y30 = ~n448 ;
  assign y31 = n457 ;
  assign y32 = n473 ;
  assign y33 = n481 ;
  assign y34 = n490 ;
  assign y35 = ~n514 ;
  assign y36 = n524 ;
  assign y37 = n537 ;
  assign y38 = n540 ;
  assign y39 = ~n565 ;
  assign y40 = n614 ;
  assign y41 = n629 ;
  assign y42 = n643 ;
  assign y43 = n687 ;
  assign y44 = n719 ;
  assign y45 = n725 ;
  assign y46 = n731 ;
  assign y47 = n737 ;
  assign y48 = n743 ;
  assign y49 = n749 ;
  assign y50 = n755 ;
  assign y51 = n761 ;
  assign y52 = n767 ;
  assign y53 = ~n790 ;
  assign y54 = n797 ;
  assign y55 = ~n815 ;
  assign y56 = ~n833 ;
  assign y57 = ~n850 ;
  assign y58 = ~n866 ;
  assign y59 = ~n874 ;
  assign y60 = ~n896 ;
  assign y61 = ~n912 ;
  assign y62 = ~n928 ;
  assign y63 = ~n947 ;
  assign y64 = ~n966 ;
  assign y65 = ~n981 ;
  assign y66 = n984 ;
  assign y67 = n988 ;
  assign y68 = n1001 ;
  assign y69 = ~n1005 ;
  assign y70 = n1008 ;
  assign y71 = n1030 ;
  assign y72 = n1046 ;
  assign y73 = n1055 ;
  assign y74 = n1081 ;
  assign y75 = n1085 ;
  assign y76 = n1088 ;
  assign y77 = ~n1099 ;
  assign y78 = ~n1104 ;
  assign y79 = ~n1109 ;
  assign y80 = ~n1114 ;
  assign y81 = ~n1119 ;
  assign y82 = ~n1122 ;
  assign y83 = ~n1127 ;
  assign y84 = ~n1132 ;
  assign y85 = ~n1137 ;
  assign y86 = ~n1142 ;
  assign y87 = ~n1145 ;
  assign y88 = ~n1148 ;
  assign y89 = ~n1151 ;
  assign y90 = ~n1154 ;
  assign y91 = ~n1157 ;
  assign y92 = ~n1160 ;
  assign y93 = n1165 ;
  assign y94 = n1168 ;
  assign y95 = n1171 ;
  assign y96 = n1174 ;
  assign y97 = n1177 ;
  assign y98 = ~n1193 ;
  assign y99 = n1196 ;
  assign y100 = n1204 ;
  assign y101 = n1207 ;
  assign y102 = n1210 ;
  assign y103 = n1215 ;
  assign y104 = n1218 ;
  assign y105 = n1221 ;
  assign y106 = n1224 ;
  assign y107 = n1227 ;
  assign y108 = n1230 ;
  assign y109 = n1236 ;
  assign y110 = n1245 ;
  assign y111 = n1249 ;
  assign y112 = n1253 ;
  assign y113 = n1256 ;
  assign y114 = n1259 ;
  assign y115 = n1263 ;
  assign y116 = ~n1278 ;
  assign y117 = ~n1291 ;
  assign y118 = ~n1304 ;
  assign y119 = ~n1317 ;
  assign y120 = ~n1332 ;
  assign y121 = n1337 ;
  assign y122 = ~n1352 ;
  assign y123 = ~n1367 ;
  assign y124 = n1372 ;
  assign y125 = n1377 ;
  assign y126 = n1385 ;
  assign y127 = n1391 ;
  assign y128 = ~n1396 ;
  assign y129 = n1006 ;
  assign y130 = n1402 ;
  assign y131 = n1408 ;
  assign y132 = ~n1409 ;
  assign y133 = n1414 ;
  assign y134 = n1415 ;
  assign y135 = n1419 ;
  assign y136 = n1421 ;
  assign y137 = n1422 ;
  assign y138 = n1423 ;
  assign y139 = n1424 ;
  assign y140 = n1427 ;
  assign y141 = n1428 ;
endmodule
